magic
tech EFS8A
magscale 1 2
timestamp 1603297099
<< locali >>
rect 14783 24701 14818 24735
rect 15991 24633 16129 24667
rect 12299 23137 12334 23171
rect 17503 22185 17509 22219
rect 17503 22117 17537 22185
rect 15663 21097 15669 21131
rect 15663 21029 15697 21097
rect 17595 20009 17601 20043
rect 17595 19941 17629 20009
rect 22471 18921 22477 18955
rect 22471 18853 22505 18921
rect 21039 18785 21166 18819
rect 23213 18207 23247 18309
rect 13087 16983 13121 17051
rect 13087 16949 13093 16983
rect 22293 16031 22327 16133
rect 19159 15657 19165 15691
rect 19159 15589 19193 15657
rect 9965 14807 9999 15045
rect 14749 14807 14783 15045
rect 10143 13719 10177 13787
rect 10143 13685 10149 13719
rect 21275 13481 21281 13515
rect 21275 13413 21309 13481
rect 14289 12699 14323 12869
rect 19947 11101 20085 11135
rect 17871 8041 17877 8075
rect 17871 7973 17905 8041
rect 24627 4641 24662 4675
rect 24627 3553 24662 3587
rect 11483 2601 11621 2635
<< viali >>
rect 24660 25313 24694 25347
rect 24731 25109 24765 25143
rect 9965 24905 9999 24939
rect 12909 24905 12943 24939
rect 15209 24905 15243 24939
rect 17325 24905 17359 24939
rect 25145 24905 25179 24939
rect 17003 24837 17037 24871
rect 9572 24701 9606 24735
rect 12516 24701 12550 24735
rect 14749 24701 14783 24735
rect 15920 24701 15954 24735
rect 16313 24701 16347 24735
rect 16932 24701 16966 24735
rect 24660 24701 24694 24735
rect 16129 24633 16163 24667
rect 18153 24633 18187 24667
rect 18245 24633 18279 24667
rect 18797 24633 18831 24667
rect 25513 24633 25547 24667
rect 9643 24565 9677 24599
rect 12587 24565 12621 24599
rect 13737 24565 13771 24599
rect 14887 24565 14921 24599
rect 17877 24565 17911 24599
rect 24731 24565 24765 24599
rect 13001 24361 13035 24395
rect 17003 24361 17037 24395
rect 18153 24361 18187 24395
rect 21097 24361 21131 24395
rect 23857 24361 23891 24395
rect 18889 24293 18923 24327
rect 6444 24225 6478 24259
rect 10584 24225 10618 24259
rect 11564 24225 11598 24259
rect 12817 24225 12851 24259
rect 13988 24225 14022 24259
rect 15853 24225 15887 24259
rect 16900 24225 16934 24259
rect 20913 24225 20947 24259
rect 23673 24225 23707 24259
rect 24844 24225 24878 24259
rect 15301 24157 15335 24191
rect 18797 24157 18831 24191
rect 19073 24157 19107 24191
rect 10655 24089 10689 24123
rect 6515 24021 6549 24055
rect 11667 24021 11701 24055
rect 13737 24021 13771 24055
rect 14059 24021 14093 24055
rect 19809 24021 19843 24055
rect 24915 24021 24949 24055
rect 3709 23817 3743 23851
rect 5825 23817 5859 23851
rect 6469 23817 6503 23851
rect 7849 23817 7883 23851
rect 8953 23817 8987 23851
rect 10425 23817 10459 23851
rect 13553 23817 13587 23851
rect 13921 23817 13955 23851
rect 14289 23817 14323 23851
rect 15853 23817 15887 23851
rect 17417 23817 17451 23851
rect 17877 23817 17911 23851
rect 19165 23817 19199 23851
rect 20913 23817 20947 23851
rect 21465 23817 21499 23851
rect 24869 23817 24903 23851
rect 25421 23817 25455 23851
rect 10057 23749 10091 23783
rect 12817 23749 12851 23783
rect 17049 23749 17083 23783
rect 20361 23749 20395 23783
rect 14933 23681 14967 23715
rect 15577 23681 15611 23715
rect 19809 23681 19843 23715
rect 1444 23613 1478 23647
rect 1869 23613 1903 23647
rect 3300 23613 3334 23647
rect 5432 23613 5466 23647
rect 7456 23613 7490 23647
rect 8560 23613 8594 23647
rect 9572 23613 9606 23647
rect 11069 23613 11103 23647
rect 12633 23613 12667 23647
rect 13185 23613 13219 23647
rect 13737 23613 13771 23647
rect 16773 23613 16807 23647
rect 16865 23613 16899 23647
rect 18245 23613 18279 23647
rect 21281 23613 21315 23647
rect 21833 23613 21867 23647
rect 23489 23613 23523 23647
rect 23765 23613 23799 23647
rect 25237 23613 25271 23647
rect 25789 23613 25823 23647
rect 3387 23545 3421 23579
rect 15025 23545 15059 23579
rect 18889 23545 18923 23579
rect 19533 23545 19567 23579
rect 19901 23545 19935 23579
rect 23121 23545 23155 23579
rect 1547 23477 1581 23511
rect 5503 23477 5537 23511
rect 7527 23477 7561 23511
rect 8631 23477 8665 23511
rect 9643 23477 9677 23511
rect 10793 23477 10827 23511
rect 11529 23477 11563 23511
rect 14749 23477 14783 23511
rect 23949 23477 23983 23511
rect 12403 23273 12437 23307
rect 14841 23273 14875 23307
rect 19257 23273 19291 23307
rect 19901 23273 19935 23307
rect 21051 23273 21085 23307
rect 25375 23273 25409 23307
rect 10885 23205 10919 23239
rect 13461 23205 13495 23239
rect 15485 23205 15519 23239
rect 18889 23205 18923 23239
rect 22293 23205 22327 23239
rect 23857 23205 23891 23239
rect 8344 23137 8378 23171
rect 12265 23137 12299 23171
rect 17176 23137 17210 23171
rect 18245 23137 18279 23171
rect 19717 23137 19751 23171
rect 20948 23137 20982 23171
rect 25304 23137 25338 23171
rect 9689 23069 9723 23103
rect 10793 23069 10827 23103
rect 13369 23069 13403 23103
rect 14013 23069 14047 23103
rect 15393 23069 15427 23103
rect 15669 23069 15703 23103
rect 22201 23069 22235 23103
rect 23765 23069 23799 23103
rect 11345 23001 11379 23035
rect 17279 23001 17313 23035
rect 22753 23001 22787 23035
rect 24317 23001 24351 23035
rect 8447 22933 8481 22967
rect 10609 22933 10643 22967
rect 14381 22933 14415 22967
rect 16497 22933 16531 22967
rect 17601 22933 17635 22967
rect 8309 22729 8343 22763
rect 10149 22729 10183 22763
rect 10609 22729 10643 22763
rect 12587 22729 12621 22763
rect 14933 22729 14967 22763
rect 15669 22729 15703 22763
rect 17417 22729 17451 22763
rect 19073 22729 19107 22763
rect 25789 22729 25823 22763
rect 26157 22729 26191 22763
rect 11345 22661 11379 22695
rect 22661 22661 22695 22695
rect 9229 22593 9263 22627
rect 12909 22593 12943 22627
rect 14013 22593 14047 22627
rect 14289 22593 14323 22627
rect 18153 22593 18187 22627
rect 23121 22593 23155 22627
rect 23765 22593 23799 22627
rect 24041 22593 24075 22627
rect 12484 22525 12518 22559
rect 19533 22525 19567 22559
rect 19717 22525 19751 22559
rect 25304 22525 25338 22559
rect 9321 22457 9355 22491
rect 9873 22457 9907 22491
rect 10793 22457 10827 22491
rect 10885 22457 10919 22491
rect 14105 22457 14139 22491
rect 16497 22457 16531 22491
rect 16589 22457 16623 22491
rect 17141 22457 17175 22491
rect 18245 22457 18279 22491
rect 18797 22457 18831 22491
rect 20913 22457 20947 22491
rect 22109 22457 22143 22491
rect 22201 22457 22235 22491
rect 23857 22457 23891 22491
rect 9045 22389 9079 22423
rect 11713 22389 11747 22423
rect 12265 22389 12299 22423
rect 13277 22389 13311 22423
rect 13829 22389 13863 22423
rect 15301 22389 15335 22423
rect 16313 22389 16347 22423
rect 17877 22389 17911 22423
rect 20085 22389 20119 22423
rect 21465 22389 21499 22423
rect 21925 22389 21959 22423
rect 23397 22389 23431 22423
rect 25375 22389 25409 22423
rect 9229 22185 9263 22219
rect 13829 22185 13863 22219
rect 17509 22185 17543 22219
rect 18061 22185 18095 22219
rect 18337 22185 18371 22219
rect 22477 22185 22511 22219
rect 23765 22185 23799 22219
rect 24041 22185 24075 22219
rect 10333 22117 10367 22151
rect 16313 22117 16347 22151
rect 19441 22117 19475 22151
rect 23397 22117 23431 22151
rect 13461 22049 13495 22083
rect 15945 22049 15979 22083
rect 22753 22049 22787 22083
rect 24660 22049 24694 22083
rect 10241 21981 10275 22015
rect 17141 21981 17175 22015
rect 19349 21981 19383 22015
rect 19993 21981 20027 22015
rect 10793 21913 10827 21947
rect 20361 21913 20395 21947
rect 24731 21913 24765 21947
rect 11161 21845 11195 21879
rect 21833 21845 21867 21879
rect 22201 21845 22235 21879
rect 4813 21641 4847 21675
rect 9045 21641 9079 21675
rect 9689 21641 9723 21675
rect 11069 21641 11103 21675
rect 14381 21641 14415 21675
rect 15945 21641 15979 21675
rect 16221 21641 16255 21675
rect 19349 21641 19383 21675
rect 19901 21641 19935 21675
rect 22661 21641 22695 21675
rect 22937 21641 22971 21675
rect 24777 21641 24811 21675
rect 18889 21573 18923 21607
rect 25789 21573 25823 21607
rect 10057 21505 10091 21539
rect 15393 21505 15427 21539
rect 17141 21505 17175 21539
rect 20085 21505 20119 21539
rect 20545 21505 20579 21539
rect 4420 21437 4454 21471
rect 8493 21437 8527 21471
rect 9229 21437 9263 21471
rect 10149 21437 10183 21471
rect 11345 21437 11379 21471
rect 13461 21437 13495 21471
rect 21741 21437 21775 21471
rect 23489 21437 23523 21471
rect 23765 21437 23799 21471
rect 25304 21437 25338 21471
rect 10511 21369 10545 21403
rect 13369 21369 13403 21403
rect 13823 21369 13857 21403
rect 16497 21369 16531 21403
rect 16589 21369 16623 21403
rect 17509 21369 17543 21403
rect 20177 21369 20211 21403
rect 22062 21369 22096 21403
rect 24409 21369 24443 21403
rect 4491 21301 4525 21335
rect 13001 21301 13035 21335
rect 17785 21301 17819 21335
rect 21649 21301 21683 21335
rect 25375 21301 25409 21335
rect 10609 21097 10643 21131
rect 13645 21097 13679 21131
rect 13921 21097 13955 21131
rect 15669 21097 15703 21131
rect 16221 21097 16255 21131
rect 16497 21097 16531 21131
rect 19717 21097 19751 21131
rect 22477 21097 22511 21131
rect 10051 21029 10085 21063
rect 13087 21029 13121 21063
rect 17233 21029 17267 21063
rect 17785 21029 17819 21063
rect 19159 21029 19193 21063
rect 21878 21029 21912 21063
rect 23489 21029 23523 21063
rect 25053 21029 25087 21063
rect 9689 20893 9723 20927
rect 12725 20893 12759 20927
rect 15301 20893 15335 20927
rect 17141 20893 17175 20927
rect 18797 20893 18831 20927
rect 21557 20893 21591 20927
rect 23397 20893 23431 20927
rect 24961 20893 24995 20927
rect 25237 20893 25271 20927
rect 23949 20825 23983 20859
rect 10885 20757 10919 20791
rect 19993 20757 20027 20791
rect 9781 20553 9815 20587
rect 15209 20553 15243 20587
rect 17233 20553 17267 20587
rect 23121 20553 23155 20587
rect 24961 20553 24995 20587
rect 11805 20485 11839 20519
rect 12265 20485 12299 20519
rect 14197 20485 14231 20519
rect 15577 20485 15611 20519
rect 17601 20485 17635 20519
rect 19349 20485 19383 20519
rect 25789 20485 25823 20519
rect 10885 20417 10919 20451
rect 13461 20417 13495 20451
rect 16589 20417 16623 20451
rect 18797 20417 18831 20451
rect 19901 20417 19935 20451
rect 9413 20349 9447 20383
rect 9873 20349 9907 20383
rect 10333 20349 10367 20383
rect 10609 20349 10643 20383
rect 12725 20349 12759 20383
rect 13277 20349 13311 20383
rect 13829 20349 13863 20383
rect 14289 20349 14323 20383
rect 22604 20349 22638 20383
rect 23673 20349 23707 20383
rect 23765 20349 23799 20383
rect 25304 20349 25338 20383
rect 9045 20281 9079 20315
rect 14651 20281 14685 20315
rect 16313 20281 16347 20315
rect 16405 20281 16439 20315
rect 19993 20281 20027 20315
rect 20545 20281 20579 20315
rect 22385 20281 22419 20315
rect 23489 20281 23523 20315
rect 16129 20213 16163 20247
rect 18705 20213 18739 20247
rect 19625 20213 19659 20247
rect 21649 20213 21683 20247
rect 21925 20213 21959 20247
rect 22707 20213 22741 20247
rect 25375 20213 25409 20247
rect 9781 20009 9815 20043
rect 12817 20009 12851 20043
rect 13553 20009 13587 20043
rect 14381 20009 14415 20043
rect 15393 20009 15427 20043
rect 17601 20009 17635 20043
rect 18153 20009 18187 20043
rect 19533 20009 19567 20043
rect 22753 20009 22787 20043
rect 23305 20009 23339 20043
rect 24961 20009 24995 20043
rect 22195 19941 22229 19975
rect 23949 19941 23983 19975
rect 25329 19941 25363 19975
rect 9781 19873 9815 19907
rect 10149 19873 10183 19907
rect 12817 19873 12851 19907
rect 13093 19873 13127 19907
rect 15301 19873 15335 19907
rect 15761 19873 15795 19907
rect 19349 19873 19383 19907
rect 11253 19805 11287 19839
rect 15117 19805 15151 19839
rect 17233 19805 17267 19839
rect 21833 19805 21867 19839
rect 23857 19805 23891 19839
rect 24225 19805 24259 19839
rect 16313 19669 16347 19703
rect 21373 19669 21407 19703
rect 9781 19465 9815 19499
rect 12725 19465 12759 19499
rect 15301 19465 15335 19499
rect 16129 19465 16163 19499
rect 18981 19465 19015 19499
rect 19349 19465 19383 19499
rect 19625 19465 19659 19499
rect 23121 19465 23155 19499
rect 23489 19397 23523 19431
rect 26065 19397 26099 19431
rect 8677 19329 8711 19363
rect 13645 19329 13679 19363
rect 14565 19329 14599 19363
rect 19901 19329 19935 19363
rect 20545 19329 20579 19363
rect 24317 19329 24351 19363
rect 8284 19261 8318 19295
rect 10701 19261 10735 19295
rect 10885 19261 10919 19295
rect 13829 19261 13863 19295
rect 14381 19261 14415 19295
rect 16313 19261 16347 19295
rect 18061 19261 18095 19295
rect 21281 19261 21315 19295
rect 21373 19261 21407 19295
rect 21833 19261 21867 19295
rect 25580 19261 25614 19295
rect 18382 19193 18416 19227
rect 19993 19193 20027 19227
rect 22109 19193 22143 19227
rect 24041 19193 24075 19227
rect 24133 19193 24167 19227
rect 8355 19125 8389 19159
rect 10149 19125 10183 19159
rect 11253 19125 11287 19159
rect 13093 19125 13127 19159
rect 15025 19125 15059 19159
rect 16865 19125 16899 19159
rect 17325 19125 17359 19159
rect 17877 19125 17911 19159
rect 22385 19125 22419 19159
rect 25651 19125 25685 19159
rect 13921 18921 13955 18955
rect 16313 18921 16347 18955
rect 19901 18921 19935 18955
rect 22477 18921 22511 18955
rect 23029 18921 23063 18955
rect 23949 18921 23983 18955
rect 24777 18921 24811 18955
rect 11345 18853 11379 18887
rect 11897 18853 11931 18887
rect 12909 18853 12943 18887
rect 13461 18853 13495 18887
rect 15485 18853 15519 18887
rect 18981 18853 19015 18887
rect 24317 18853 24351 18887
rect 21005 18785 21039 18819
rect 22109 18785 22143 18819
rect 24593 18785 24627 18819
rect 11253 18717 11287 18751
rect 12817 18717 12851 18751
rect 15393 18717 15427 18751
rect 17785 18717 17819 18751
rect 18889 18717 18923 18751
rect 15945 18649 15979 18683
rect 19441 18649 19475 18683
rect 21235 18649 21269 18683
rect 10333 18581 10367 18615
rect 12541 18581 12575 18615
rect 18245 18581 18279 18615
rect 21833 18581 21867 18615
rect 11529 18377 11563 18411
rect 16129 18377 16163 18411
rect 19809 18377 19843 18411
rect 21833 18377 21867 18411
rect 24685 18377 24719 18411
rect 11897 18309 11931 18343
rect 23213 18309 23247 18343
rect 25421 18309 25455 18343
rect 8861 18241 8895 18275
rect 13277 18241 13311 18275
rect 14197 18241 14231 18275
rect 15485 18241 15519 18275
rect 16313 18241 16347 18275
rect 21373 18241 21407 18275
rect 24225 18241 24259 18275
rect 10333 18173 10367 18207
rect 11253 18173 11287 18207
rect 12633 18173 12667 18207
rect 18337 18173 18371 18207
rect 18981 18173 19015 18207
rect 19441 18173 19475 18207
rect 20545 18173 20579 18207
rect 20913 18173 20947 18207
rect 21097 18173 21131 18207
rect 22604 18173 22638 18207
rect 23029 18173 23063 18207
rect 23213 18173 23247 18207
rect 23489 18173 23523 18207
rect 23673 18173 23707 18207
rect 24133 18173 24167 18207
rect 25237 18173 25271 18207
rect 25789 18173 25823 18207
rect 8677 18105 8711 18139
rect 8953 18105 8987 18139
rect 9505 18105 9539 18139
rect 10654 18105 10688 18139
rect 13369 18105 13403 18139
rect 13921 18105 13955 18139
rect 14841 18105 14875 18139
rect 14933 18105 14967 18139
rect 19165 18105 19199 18139
rect 22707 18105 22741 18139
rect 10149 18037 10183 18071
rect 13093 18037 13127 18071
rect 14657 18037 14691 18071
rect 15761 18037 15795 18071
rect 16957 18037 16991 18071
rect 22201 18037 22235 18071
rect 8861 17833 8895 17867
rect 10609 17833 10643 17867
rect 14841 17833 14875 17867
rect 15761 17833 15795 17867
rect 17969 17833 18003 17867
rect 22017 17833 22051 17867
rect 23029 17833 23063 17867
rect 10010 17765 10044 17799
rect 13823 17765 13857 17799
rect 16773 17765 16807 17799
rect 18981 17765 19015 17799
rect 19073 17765 19107 17799
rect 22430 17765 22464 17799
rect 24041 17765 24075 17799
rect 11529 17697 11563 17731
rect 14381 17697 14415 17731
rect 15393 17697 15427 17731
rect 16865 17697 16899 17731
rect 17325 17697 17359 17731
rect 17693 17697 17727 17731
rect 21164 17697 21198 17731
rect 23673 17697 23707 17731
rect 9689 17629 9723 17663
rect 11437 17629 11471 17663
rect 13461 17629 13495 17663
rect 16405 17629 16439 17663
rect 19441 17629 19475 17663
rect 22109 17629 22143 17663
rect 23949 17629 23983 17663
rect 24225 17629 24259 17663
rect 25421 17629 25455 17663
rect 20729 17561 20763 17595
rect 21649 17561 21683 17595
rect 12725 17493 12759 17527
rect 13277 17493 13311 17527
rect 18245 17493 18279 17527
rect 21235 17493 21269 17527
rect 11529 17289 11563 17323
rect 13645 17289 13679 17323
rect 17141 17289 17175 17323
rect 18981 17289 19015 17323
rect 19257 17289 19291 17323
rect 20361 17289 20395 17323
rect 25421 17289 25455 17323
rect 10885 17221 10919 17255
rect 19625 17221 19659 17255
rect 22707 17221 22741 17255
rect 24777 17221 24811 17255
rect 9413 17153 9447 17187
rect 10333 17153 10367 17187
rect 14841 17153 14875 17187
rect 15577 17153 15611 17187
rect 16957 17153 16991 17187
rect 21557 17153 21591 17187
rect 23121 17153 23155 17187
rect 23765 17153 23799 17187
rect 24041 17153 24075 17187
rect 8585 17085 8619 17119
rect 8953 17085 8987 17119
rect 9229 17085 9263 17119
rect 12725 17085 12759 17119
rect 16037 17085 16071 17119
rect 16865 17085 16899 17119
rect 18061 17085 18095 17119
rect 20821 17085 20855 17119
rect 21281 17085 21315 17119
rect 22636 17085 22670 17119
rect 25237 17085 25271 17119
rect 25789 17085 25823 17119
rect 10425 17017 10459 17051
rect 14565 17017 14599 17051
rect 14657 17017 14691 17051
rect 17877 17017 17911 17051
rect 18423 17017 18457 17051
rect 23857 17017 23891 17051
rect 9781 16949 9815 16983
rect 10149 16949 10183 16983
rect 13093 16949 13127 16983
rect 13921 16949 13955 16983
rect 14381 16949 14415 16983
rect 15853 16949 15887 16983
rect 17417 16949 17451 16983
rect 19809 16949 19843 16983
rect 20729 16949 20763 16983
rect 22201 16949 22235 16983
rect 23489 16949 23523 16983
rect 9505 16745 9539 16779
rect 10149 16745 10183 16779
rect 13277 16745 13311 16779
rect 15117 16745 15151 16779
rect 16773 16745 16807 16779
rect 18705 16745 18739 16779
rect 20085 16745 20119 16779
rect 22661 16745 22695 16779
rect 23581 16745 23615 16779
rect 24317 16745 24351 16779
rect 8769 16677 8803 16711
rect 21649 16677 21683 16711
rect 22109 16677 22143 16711
rect 9873 16609 9907 16643
rect 10425 16609 10459 16643
rect 11529 16609 11563 16643
rect 13093 16609 13127 16643
rect 13461 16609 13495 16643
rect 15301 16609 15335 16643
rect 16497 16609 16531 16643
rect 16957 16609 16991 16643
rect 17325 16609 17359 16643
rect 18705 16609 18739 16643
rect 18889 16609 18923 16643
rect 21189 16609 21223 16643
rect 21373 16609 21407 16643
rect 23949 16609 23983 16643
rect 11437 16541 11471 16575
rect 24869 16541 24903 16575
rect 12725 16473 12759 16507
rect 15485 16473 15519 16507
rect 10977 16405 11011 16439
rect 14197 16405 14231 16439
rect 14473 16405 14507 16439
rect 16129 16405 16163 16439
rect 18061 16405 18095 16439
rect 9045 16201 9079 16235
rect 9413 16201 9447 16235
rect 9781 16201 9815 16235
rect 11529 16201 11563 16235
rect 12265 16201 12299 16235
rect 13553 16201 13587 16235
rect 14381 16201 14415 16235
rect 17141 16201 17175 16235
rect 21097 16201 21131 16235
rect 23397 16201 23431 16235
rect 19165 16133 19199 16167
rect 22293 16133 22327 16167
rect 22385 16133 22419 16167
rect 25605 16133 25639 16167
rect 16957 16065 16991 16099
rect 17417 16065 17451 16099
rect 19533 16065 19567 16099
rect 20085 16065 20119 16099
rect 20545 16065 20579 16099
rect 22109 16065 22143 16099
rect 9873 15997 9907 16031
rect 10425 15997 10459 16031
rect 12541 15997 12575 16031
rect 13001 15997 13035 16031
rect 13921 15997 13955 16031
rect 14197 15997 14231 16031
rect 16037 15997 16071 16031
rect 16865 15997 16899 16031
rect 17877 15997 17911 16031
rect 18337 15997 18371 16031
rect 18521 15997 18555 16031
rect 19809 15997 19843 16031
rect 21624 15997 21658 16031
rect 22293 15997 22327 16031
rect 22604 15997 22638 16031
rect 23949 15997 23983 16031
rect 25421 15997 25455 16031
rect 25973 15997 26007 16031
rect 15853 15929 15887 15963
rect 18797 15929 18831 15963
rect 20177 15929 20211 15963
rect 21373 15929 21407 15963
rect 22707 15929 22741 15963
rect 10149 15861 10183 15895
rect 12633 15861 12667 15895
rect 15301 15861 15335 15895
rect 21695 15861 21729 15895
rect 24133 15861 24167 15895
rect 9873 15657 9907 15691
rect 12633 15657 12667 15691
rect 14197 15657 14231 15691
rect 16221 15657 16255 15691
rect 17233 15657 17267 15691
rect 19165 15657 19199 15691
rect 19993 15657 20027 15691
rect 22109 15657 22143 15691
rect 23397 15657 23431 15691
rect 23949 15657 23983 15691
rect 11253 15589 11287 15623
rect 16497 15589 16531 15623
rect 22798 15589 22832 15623
rect 24409 15589 24443 15623
rect 9689 15521 9723 15555
rect 13553 15521 13587 15555
rect 15669 15521 15703 15555
rect 17049 15521 17083 15555
rect 17509 15521 17543 15555
rect 21097 15521 21131 15555
rect 21373 15521 21407 15555
rect 11161 15453 11195 15487
rect 13921 15453 13955 15487
rect 15485 15453 15519 15487
rect 18797 15453 18831 15487
rect 21649 15453 21683 15487
rect 22477 15453 22511 15487
rect 24317 15453 24351 15487
rect 24593 15453 24627 15487
rect 11713 15385 11747 15419
rect 15853 15385 15887 15419
rect 16957 15385 16991 15419
rect 10241 15317 10275 15351
rect 13001 15317 13035 15351
rect 13461 15317 13495 15351
rect 13691 15317 13725 15351
rect 13829 15317 13863 15351
rect 15025 15317 15059 15351
rect 18061 15317 18095 15351
rect 18429 15317 18463 15351
rect 19717 15317 19751 15351
rect 11437 15113 11471 15147
rect 11805 15113 11839 15147
rect 13921 15113 13955 15147
rect 15485 15113 15519 15147
rect 16773 15113 16807 15147
rect 18337 15113 18371 15147
rect 18705 15113 18739 15147
rect 21005 15113 21039 15147
rect 23397 15113 23431 15147
rect 24041 15113 24075 15147
rect 25237 15113 25271 15147
rect 9965 15045 9999 15079
rect 11161 15045 11195 15079
rect 13001 15045 13035 15079
rect 13737 15045 13771 15079
rect 14749 15045 14783 15079
rect 15301 15045 15335 15079
rect 19165 15045 19199 15079
rect 20545 15045 20579 15079
rect 8585 14977 8619 15011
rect 8953 14909 8987 14943
rect 9229 14909 9263 14943
rect 9413 14841 9447 14875
rect 9781 14841 9815 14875
rect 10241 14977 10275 15011
rect 12449 14977 12483 15011
rect 13608 14977 13642 15011
rect 13829 14977 13863 15011
rect 12265 14909 12299 14943
rect 10562 14841 10596 14875
rect 13461 14841 13495 14875
rect 15172 14977 15206 15011
rect 15393 14977 15427 15011
rect 17417 14977 17451 15011
rect 18429 14977 18463 15011
rect 19993 14977 20027 15011
rect 22109 14977 22143 15011
rect 22385 14977 22419 15011
rect 24317 14977 24351 15011
rect 24777 14977 24811 15011
rect 16589 14909 16623 14943
rect 17049 14909 17083 14943
rect 18208 14909 18242 14943
rect 15025 14841 15059 14875
rect 16037 14841 16071 14875
rect 18061 14841 18095 14875
rect 20085 14841 20119 14875
rect 22201 14841 22235 14875
rect 24409 14841 24443 14875
rect 9965 14773 9999 14807
rect 10057 14773 10091 14807
rect 13369 14773 13403 14807
rect 14565 14773 14599 14807
rect 14749 14773 14783 14807
rect 14841 14773 14875 14807
rect 16497 14773 16531 14807
rect 17785 14773 17819 14807
rect 19717 14773 19751 14807
rect 21281 14773 21315 14807
rect 21925 14773 21959 14807
rect 23029 14773 23063 14807
rect 8769 14569 8803 14603
rect 10241 14569 10275 14603
rect 12909 14569 12943 14603
rect 14473 14569 14507 14603
rect 15025 14569 15059 14603
rect 16405 14569 16439 14603
rect 18521 14569 18555 14603
rect 18889 14569 18923 14603
rect 19533 14569 19567 14603
rect 22477 14569 22511 14603
rect 24317 14569 24351 14603
rect 11253 14501 11287 14535
rect 14105 14501 14139 14535
rect 17877 14501 17911 14535
rect 21465 14501 21499 14535
rect 22017 14501 22051 14535
rect 13277 14433 13311 14467
rect 13369 14433 13403 14467
rect 15393 14433 15427 14467
rect 17141 14433 17175 14467
rect 19533 14433 19567 14467
rect 22937 14433 22971 14467
rect 24593 14433 24627 14467
rect 11161 14365 11195 14399
rect 13737 14365 13771 14399
rect 15301 14365 15335 14399
rect 17509 14365 17543 14399
rect 21373 14365 21407 14399
rect 11713 14297 11747 14331
rect 17049 14297 17083 14331
rect 24777 14297 24811 14331
rect 13507 14229 13541 14263
rect 13645 14229 13679 14263
rect 17279 14229 17313 14263
rect 17417 14229 17451 14263
rect 18153 14229 18187 14263
rect 23305 14229 23339 14263
rect 9321 14025 9355 14059
rect 9689 14025 9723 14059
rect 11161 14025 11195 14059
rect 13626 14025 13660 14059
rect 14841 14025 14875 14059
rect 15853 14025 15887 14059
rect 16681 14025 16715 14059
rect 17417 14025 17451 14059
rect 18337 14025 18371 14059
rect 19533 14025 19567 14059
rect 20545 14025 20579 14059
rect 21925 14025 21959 14059
rect 22937 14025 22971 14059
rect 23397 14025 23431 14059
rect 24685 14025 24719 14059
rect 25421 14025 25455 14059
rect 13001 13957 13035 13991
rect 13369 13957 13403 13991
rect 13737 13957 13771 13991
rect 15209 13957 15243 13991
rect 15577 13957 15611 13991
rect 16543 13957 16577 13991
rect 9781 13889 9815 13923
rect 13829 13889 13863 13923
rect 16773 13889 16807 13923
rect 18208 13889 18242 13923
rect 18429 13889 18463 13923
rect 18797 13889 18831 13923
rect 21005 13889 21039 13923
rect 21373 13889 21407 13923
rect 24041 13889 24075 13923
rect 25789 13889 25823 13923
rect 13461 13821 13495 13855
rect 15393 13821 15427 13855
rect 17141 13821 17175 13855
rect 19073 13821 19107 13855
rect 19625 13821 19659 13855
rect 20085 13821 20119 13855
rect 21833 13821 21867 13855
rect 25237 13821 25271 13855
rect 14197 13753 14231 13787
rect 16405 13753 16439 13787
rect 18061 13753 18095 13787
rect 23765 13753 23799 13787
rect 23857 13753 23891 13787
rect 10149 13685 10183 13719
rect 10701 13685 10735 13719
rect 11437 13685 11471 13719
rect 12265 13685 12299 13719
rect 14565 13685 14599 13719
rect 16221 13685 16255 13719
rect 17877 13685 17911 13719
rect 19809 13685 19843 13719
rect 12633 13481 12667 13515
rect 12909 13481 12943 13515
rect 14105 13481 14139 13515
rect 16497 13481 16531 13515
rect 18061 13481 18095 13515
rect 18521 13481 18555 13515
rect 21281 13481 21315 13515
rect 21833 13481 21867 13515
rect 11069 13413 11103 13447
rect 13461 13413 13495 13447
rect 17049 13413 17083 13447
rect 22753 13413 22787 13447
rect 22845 13413 22879 13447
rect 24409 13413 24443 13447
rect 12449 13345 12483 13379
rect 13369 13345 13403 13379
rect 13608 13345 13642 13379
rect 15301 13345 15335 13379
rect 19257 13345 19291 13379
rect 19717 13345 19751 13379
rect 10977 13277 11011 13311
rect 13829 13277 13863 13311
rect 17417 13277 17451 13311
rect 19993 13277 20027 13311
rect 20913 13277 20947 13311
rect 23029 13277 23063 13311
rect 24317 13277 24351 13311
rect 11529 13209 11563 13243
rect 13737 13209 13771 13243
rect 15025 13209 15059 13243
rect 16865 13209 16899 13243
rect 17325 13209 17359 13243
rect 24869 13209 24903 13243
rect 14657 13141 14691 13175
rect 15485 13141 15519 13175
rect 15853 13141 15887 13175
rect 17214 13141 17248 13175
rect 17693 13141 17727 13175
rect 18797 13141 18831 13175
rect 23765 13141 23799 13175
rect 13277 12937 13311 12971
rect 14730 12937 14764 12971
rect 15577 12937 15611 12971
rect 18199 12937 18233 12971
rect 22385 12937 22419 12971
rect 23121 12937 23155 12971
rect 25145 12937 25179 12971
rect 14289 12869 14323 12903
rect 14841 12869 14875 12903
rect 18337 12869 18371 12903
rect 19809 12869 19843 12903
rect 21925 12869 21959 12903
rect 10885 12801 10919 12835
rect 11897 12801 11931 12835
rect 13369 12801 13403 12835
rect 13148 12733 13182 12767
rect 14105 12733 14139 12767
rect 14933 12801 14967 12835
rect 17141 12801 17175 12835
rect 18429 12801 18463 12835
rect 19257 12801 19291 12835
rect 22753 12801 22787 12835
rect 25237 12801 25271 12835
rect 16497 12733 16531 12767
rect 18061 12733 18095 12767
rect 19625 12733 19659 12767
rect 20085 12733 20119 12767
rect 21005 12733 21039 12767
rect 10241 12665 10275 12699
rect 10333 12665 10367 12699
rect 12173 12665 12207 12699
rect 13001 12665 13035 12699
rect 13737 12665 13771 12699
rect 14289 12665 14323 12699
rect 14565 12665 14599 12699
rect 15301 12665 15335 12699
rect 18797 12665 18831 12699
rect 21326 12665 21360 12699
rect 23765 12665 23799 12699
rect 23857 12665 23891 12699
rect 24409 12665 24443 12699
rect 9965 12597 9999 12631
rect 11161 12597 11195 12631
rect 12909 12597 12943 12631
rect 14473 12597 14507 12631
rect 16221 12597 16255 12631
rect 17417 12597 17451 12631
rect 17785 12597 17819 12631
rect 20545 12597 20579 12631
rect 20821 12597 20855 12631
rect 23489 12597 23523 12631
rect 24685 12597 24719 12631
rect 10149 12393 10183 12427
rect 12357 12393 12391 12427
rect 12725 12393 12759 12427
rect 13093 12393 13127 12427
rect 13369 12393 13403 12427
rect 13645 12393 13679 12427
rect 16405 12393 16439 12427
rect 16773 12393 16807 12427
rect 17049 12393 17083 12427
rect 18613 12393 18647 12427
rect 21097 12393 21131 12427
rect 11161 12325 11195 12359
rect 14013 12325 14047 12359
rect 14749 12325 14783 12359
rect 17233 12325 17267 12359
rect 19993 12325 20027 12359
rect 21465 12325 21499 12359
rect 22062 12325 22096 12359
rect 24409 12325 24443 12359
rect 10517 12257 10551 12291
rect 12173 12257 12207 12291
rect 13185 12257 13219 12291
rect 14197 12257 14231 12291
rect 15301 12257 15335 12291
rect 19257 12257 19291 12291
rect 19717 12257 19751 12291
rect 22661 12257 22695 12291
rect 24225 12257 24259 12291
rect 25237 12257 25271 12291
rect 15669 12189 15703 12223
rect 17601 12189 17635 12223
rect 19165 12189 19199 12223
rect 21741 12189 21775 12223
rect 14381 12121 14415 12155
rect 15466 12121 15500 12155
rect 17509 12121 17543 12155
rect 17877 12121 17911 12155
rect 25421 12121 25455 12155
rect 11529 12053 11563 12087
rect 15025 12053 15059 12087
rect 15577 12053 15611 12087
rect 15945 12053 15979 12087
rect 17371 12053 17405 12087
rect 18245 12053 18279 12087
rect 9689 11849 9723 11883
rect 13921 11849 13955 11883
rect 15669 11849 15703 11883
rect 17785 11849 17819 11883
rect 18889 11849 18923 11883
rect 23811 11849 23845 11883
rect 24225 11849 24259 11883
rect 25513 11849 25547 11883
rect 15393 11781 15427 11815
rect 18245 11781 18279 11815
rect 24823 11781 24857 11815
rect 10333 11713 10367 11747
rect 16405 11713 16439 11747
rect 10517 11645 10551 11679
rect 10885 11645 10919 11679
rect 11069 11645 11103 11679
rect 12633 11645 12667 11679
rect 13277 11645 13311 11679
rect 14289 11645 14323 11679
rect 14565 11645 14599 11679
rect 16497 11645 16531 11679
rect 17417 11645 17451 11679
rect 18061 11645 18095 11679
rect 18521 11645 18555 11679
rect 20085 11645 20119 11679
rect 20545 11645 20579 11679
rect 23740 11645 23774 11679
rect 24501 11645 24535 11679
rect 24752 11645 24786 11679
rect 12449 11577 12483 11611
rect 13001 11577 13035 11611
rect 14749 11577 14783 11611
rect 20821 11577 20855 11611
rect 10057 11509 10091 11543
rect 12265 11509 12299 11543
rect 16313 11509 16347 11543
rect 19257 11509 19291 11543
rect 19901 11509 19935 11543
rect 21741 11509 21775 11543
rect 22109 11509 22143 11543
rect 22569 11509 22603 11543
rect 25237 11509 25271 11543
rect 13185 11305 13219 11339
rect 13553 11305 13587 11339
rect 14473 11305 14507 11339
rect 16957 11305 16991 11339
rect 18843 11305 18877 11339
rect 19349 11305 19383 11339
rect 20361 11305 20395 11339
rect 23673 11305 23707 11339
rect 15025 11237 15059 11271
rect 21649 11237 21683 11271
rect 23074 11237 23108 11271
rect 24685 11237 24719 11271
rect 10333 11169 10367 11203
rect 10977 11169 11011 11203
rect 12449 11169 12483 11203
rect 13737 11169 13771 11203
rect 14013 11169 14047 11203
rect 15485 11169 15519 11203
rect 17141 11169 17175 11203
rect 17693 11169 17727 11203
rect 18740 11169 18774 11203
rect 19876 11169 19910 11203
rect 20913 11169 20947 11203
rect 21373 11169 21407 11203
rect 22753 11169 22787 11203
rect 16497 11101 16531 11135
rect 20085 11101 20119 11135
rect 24593 11101 24627 11135
rect 18521 11033 18555 11067
rect 25145 11033 25179 11067
rect 15577 10965 15611 10999
rect 17233 10965 17267 10999
rect 22017 10965 22051 10999
rect 12725 10761 12759 10795
rect 14197 10761 14231 10795
rect 15577 10761 15611 10795
rect 16865 10761 16899 10795
rect 19809 10761 19843 10795
rect 21281 10761 21315 10795
rect 21649 10761 21683 10795
rect 23305 10761 23339 10795
rect 23949 10761 23983 10795
rect 25513 10761 25547 10795
rect 14473 10693 14507 10727
rect 16681 10693 16715 10727
rect 22937 10693 22971 10727
rect 25145 10693 25179 10727
rect 12909 10625 12943 10659
rect 14657 10625 14691 10659
rect 16773 10625 16807 10659
rect 22661 10625 22695 10659
rect 24593 10625 24627 10659
rect 16552 10557 16586 10591
rect 18337 10557 18371 10591
rect 18705 10557 18739 10591
rect 18889 10557 18923 10591
rect 13230 10489 13264 10523
rect 14978 10489 15012 10523
rect 15945 10489 15979 10523
rect 16405 10489 16439 10523
rect 19165 10489 19199 10523
rect 20361 10489 20395 10523
rect 20453 10489 20487 10523
rect 21005 10489 21039 10523
rect 22017 10489 22051 10523
rect 22109 10489 22143 10523
rect 24685 10489 24719 10523
rect 10241 10421 10275 10455
rect 13829 10421 13863 10455
rect 16221 10421 16255 10455
rect 17417 10421 17451 10455
rect 17785 10421 17819 10455
rect 20085 10421 20119 10455
rect 24409 10421 24443 10455
rect 13001 10217 13035 10251
rect 14749 10217 14783 10251
rect 15117 10217 15151 10251
rect 18429 10217 18463 10251
rect 19717 10217 19751 10251
rect 20361 10217 20395 10251
rect 24409 10217 24443 10251
rect 13277 10149 13311 10183
rect 15485 10149 15519 10183
rect 17785 10149 17819 10183
rect 22569 10149 22603 10183
rect 23121 10149 23155 10183
rect 17233 10081 17267 10115
rect 18705 10081 18739 10115
rect 19165 10081 19199 10115
rect 24225 10081 24259 10115
rect 24961 10081 24995 10115
rect 13185 10013 13219 10047
rect 15393 10013 15427 10047
rect 15669 10013 15703 10047
rect 19441 10013 19475 10047
rect 21373 10013 21407 10047
rect 22477 10013 22511 10047
rect 13737 9945 13771 9979
rect 14197 9877 14231 9911
rect 16405 9877 16439 9911
rect 21925 9877 21959 9911
rect 12173 9673 12207 9707
rect 12909 9673 12943 9707
rect 14841 9673 14875 9707
rect 15945 9673 15979 9707
rect 18337 9673 18371 9707
rect 20361 9673 20395 9707
rect 22753 9673 22787 9707
rect 24041 9673 24075 9707
rect 24777 9673 24811 9707
rect 13277 9537 13311 9571
rect 15669 9537 15703 9571
rect 19165 9537 19199 9571
rect 20913 9537 20947 9571
rect 21833 9469 21867 9503
rect 24593 9469 24627 9503
rect 25145 9469 25179 9503
rect 13461 9401 13495 9435
rect 13553 9401 13587 9435
rect 14105 9401 14139 9435
rect 15025 9401 15059 9435
rect 15117 9401 15151 9435
rect 18613 9401 18647 9435
rect 19486 9401 19520 9435
rect 20729 9401 20763 9435
rect 21234 9401 21268 9435
rect 14473 9333 14507 9367
rect 17141 9333 17175 9367
rect 18981 9333 19015 9367
rect 20085 9333 20119 9367
rect 22477 9333 22511 9367
rect 13461 9129 13495 9163
rect 14933 9129 14967 9163
rect 15301 9129 15335 9163
rect 17509 9129 17543 9163
rect 24133 9129 24167 9163
rect 24777 9129 24811 9163
rect 15761 9061 15795 9095
rect 19993 9061 20027 9095
rect 21373 9061 21407 9095
rect 21925 9061 21959 9095
rect 22753 9061 22787 9095
rect 13277 8993 13311 9027
rect 17233 8993 17267 9027
rect 17417 8993 17451 9027
rect 19349 8993 19383 9027
rect 23029 8993 23063 9027
rect 24593 8993 24627 9027
rect 21281 8925 21315 8959
rect 18153 8789 18187 8823
rect 13185 8585 13219 8619
rect 14105 8585 14139 8619
rect 15025 8585 15059 8619
rect 19349 8585 19383 8619
rect 21281 8585 21315 8619
rect 21649 8585 21683 8619
rect 22707 8585 22741 8619
rect 26157 8585 26191 8619
rect 17693 8517 17727 8551
rect 23029 8517 23063 8551
rect 23857 8517 23891 8551
rect 17325 8449 17359 8483
rect 24133 8449 24167 8483
rect 24409 8449 24443 8483
rect 13921 8381 13955 8415
rect 14381 8381 14415 8415
rect 15209 8381 15243 8415
rect 15669 8381 15703 8415
rect 18153 8381 18187 8415
rect 20085 8381 20119 8415
rect 20269 8381 20303 8415
rect 20729 8381 20763 8415
rect 22636 8381 22670 8415
rect 25672 8381 25706 8415
rect 15945 8313 15979 8347
rect 18797 8313 18831 8347
rect 21005 8313 21039 8347
rect 23397 8313 23431 8347
rect 24225 8313 24259 8347
rect 25053 8245 25087 8279
rect 25743 8245 25777 8279
rect 15485 8041 15519 8075
rect 16957 8041 16991 8075
rect 17877 8041 17911 8075
rect 18429 8041 18463 8075
rect 16082 7973 16116 8007
rect 22062 7973 22096 8007
rect 24225 7973 24259 8007
rect 17509 7905 17543 7939
rect 19257 7905 19291 7939
rect 19717 7905 19751 7939
rect 20269 7905 20303 7939
rect 15761 7837 15795 7871
rect 19993 7837 20027 7871
rect 21741 7837 21775 7871
rect 24133 7837 24167 7871
rect 24409 7837 24443 7871
rect 16681 7701 16715 7735
rect 18705 7701 18739 7735
rect 22661 7701 22695 7735
rect 15853 7497 15887 7531
rect 17509 7497 17543 7531
rect 19441 7497 19475 7531
rect 21189 7497 21223 7531
rect 22661 7497 22695 7531
rect 23489 7497 23523 7531
rect 25743 7497 25777 7531
rect 26157 7497 26191 7531
rect 14749 7429 14783 7463
rect 19165 7429 19199 7463
rect 21557 7429 21591 7463
rect 23949 7429 23983 7463
rect 24685 7429 24719 7463
rect 15577 7361 15611 7395
rect 16497 7361 16531 7395
rect 17141 7361 17175 7395
rect 18153 7361 18187 7395
rect 19993 7361 20027 7395
rect 21741 7361 21775 7395
rect 24133 7361 24167 7395
rect 25421 7361 25455 7395
rect 15117 7293 15151 7327
rect 15301 7293 15335 7327
rect 25672 7293 25706 7327
rect 16589 7225 16623 7259
rect 18245 7225 18279 7259
rect 18797 7225 18831 7259
rect 19717 7225 19751 7259
rect 19809 7225 19843 7259
rect 22062 7225 22096 7259
rect 24225 7225 24259 7259
rect 16313 7157 16347 7191
rect 25053 7157 25087 7191
rect 14933 6953 14967 6987
rect 15761 6953 15795 6987
rect 17417 6953 17451 6987
rect 18613 6953 18647 6987
rect 19395 6953 19429 6987
rect 16773 6885 16807 6919
rect 17785 6885 17819 6919
rect 18337 6885 18371 6919
rect 19717 6885 19751 6919
rect 22109 6885 22143 6919
rect 23305 6885 23339 6919
rect 24317 6885 24351 6919
rect 16681 6817 16715 6851
rect 19292 6817 19326 6851
rect 22661 6817 22695 6851
rect 17693 6749 17727 6783
rect 21741 6749 21775 6783
rect 24225 6749 24259 6783
rect 24501 6749 24535 6783
rect 20085 6613 20119 6647
rect 16129 6409 16163 6443
rect 17693 6409 17727 6443
rect 19257 6409 19291 6443
rect 22661 6409 22695 6443
rect 23397 6409 23431 6443
rect 25375 6409 25409 6443
rect 25789 6409 25823 6443
rect 18153 6273 18187 6307
rect 24409 6273 24443 6307
rect 24685 6273 24719 6307
rect 23765 6205 23799 6239
rect 25304 6205 25338 6239
rect 17325 6069 17359 6103
rect 18199 5865 18233 5899
rect 23489 5865 23523 5899
rect 18128 5729 18162 5763
rect 24660 5729 24694 5763
rect 24731 5593 24765 5627
rect 24225 5525 24259 5559
rect 24685 5321 24719 5355
rect 18337 4981 18371 5015
rect 24731 4709 24765 4743
rect 24593 4641 24627 4675
rect 24685 4233 24719 4267
rect 24731 3621 24765 3655
rect 24593 3553 24627 3587
rect 24685 3145 24719 3179
rect 11621 2601 11655 2635
rect 24731 2601 24765 2635
rect 11412 2465 11446 2499
rect 24660 2465 24694 2499
rect 11897 2397 11931 2431
rect 25145 2261 25179 2295
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 13906 25440 13912 25492
rect 13964 25480 13970 25492
rect 20070 25480 20076 25492
rect 13964 25452 20076 25480
rect 13964 25440 13970 25452
rect 20070 25440 20076 25452
rect 20128 25440 20134 25492
rect 24648 25347 24706 25353
rect 24648 25313 24660 25347
rect 24694 25344 24706 25347
rect 25498 25344 25504 25356
rect 24694 25316 25504 25344
rect 24694 25313 24706 25316
rect 24648 25307 24706 25313
rect 25498 25304 25504 25316
rect 25556 25304 25562 25356
rect 23842 25100 23848 25152
rect 23900 25140 23906 25152
rect 24719 25143 24777 25149
rect 24719 25140 24731 25143
rect 23900 25112 24731 25140
rect 23900 25100 23906 25112
rect 24719 25109 24731 25112
rect 24765 25109 24777 25143
rect 24719 25103 24777 25109
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 9950 24936 9956 24948
rect 9911 24908 9956 24936
rect 9950 24896 9956 24908
rect 10008 24896 10014 24948
rect 12894 24936 12900 24948
rect 12855 24908 12900 24936
rect 12894 24896 12900 24908
rect 12952 24896 12958 24948
rect 14826 24896 14832 24948
rect 14884 24936 14890 24948
rect 15197 24939 15255 24945
rect 15197 24936 15209 24939
rect 14884 24908 15209 24936
rect 14884 24896 14890 24908
rect 15197 24905 15209 24908
rect 15243 24905 15255 24939
rect 17310 24936 17316 24948
rect 17271 24908 17316 24936
rect 15197 24899 15255 24905
rect 17310 24896 17316 24908
rect 17368 24896 17374 24948
rect 25130 24936 25136 24948
rect 25091 24908 25136 24936
rect 25130 24896 25136 24908
rect 25188 24896 25194 24948
rect 16206 24828 16212 24880
rect 16264 24868 16270 24880
rect 16991 24871 17049 24877
rect 16991 24868 17003 24871
rect 16264 24840 17003 24868
rect 16264 24828 16270 24840
rect 16991 24837 17003 24840
rect 17037 24837 17049 24871
rect 16991 24831 17049 24837
rect 9560 24735 9618 24741
rect 9560 24701 9572 24735
rect 9606 24732 9618 24735
rect 9950 24732 9956 24744
rect 9606 24704 9956 24732
rect 9606 24701 9618 24704
rect 9560 24695 9618 24701
rect 9950 24692 9956 24704
rect 10008 24692 10014 24744
rect 12504 24735 12562 24741
rect 12504 24701 12516 24735
rect 12550 24732 12562 24735
rect 12894 24732 12900 24744
rect 12550 24704 12900 24732
rect 12550 24701 12562 24704
rect 12504 24695 12562 24701
rect 12894 24692 12900 24704
rect 12952 24692 12958 24744
rect 14737 24735 14795 24741
rect 14737 24701 14749 24735
rect 14783 24732 14795 24735
rect 14826 24732 14832 24744
rect 14783 24704 14832 24732
rect 14783 24701 14795 24704
rect 14737 24695 14795 24701
rect 14826 24692 14832 24704
rect 14884 24692 14890 24744
rect 15562 24692 15568 24744
rect 15620 24732 15626 24744
rect 15908 24735 15966 24741
rect 15908 24732 15920 24735
rect 15620 24704 15920 24732
rect 15620 24692 15626 24704
rect 15908 24701 15920 24704
rect 15954 24732 15966 24735
rect 16301 24735 16359 24741
rect 16301 24732 16313 24735
rect 15954 24704 16313 24732
rect 15954 24701 15966 24704
rect 15908 24695 15966 24701
rect 16301 24701 16313 24704
rect 16347 24701 16359 24735
rect 16301 24695 16359 24701
rect 16920 24735 16978 24741
rect 16920 24701 16932 24735
rect 16966 24732 16978 24735
rect 17310 24732 17316 24744
rect 16966 24704 17316 24732
rect 16966 24701 16978 24704
rect 16920 24695 16978 24701
rect 17310 24692 17316 24704
rect 17368 24692 17374 24744
rect 24648 24735 24706 24741
rect 24648 24701 24660 24735
rect 24694 24732 24706 24735
rect 25130 24732 25136 24744
rect 24694 24704 25136 24732
rect 24694 24701 24706 24704
rect 24648 24695 24706 24701
rect 25130 24692 25136 24704
rect 25188 24692 25194 24744
rect 16117 24667 16175 24673
rect 16117 24633 16129 24667
rect 16163 24664 16175 24667
rect 17954 24664 17960 24676
rect 16163 24636 17960 24664
rect 16163 24633 16175 24636
rect 16117 24627 16175 24633
rect 17954 24624 17960 24636
rect 18012 24624 18018 24676
rect 18138 24664 18144 24676
rect 18099 24636 18144 24664
rect 18138 24624 18144 24636
rect 18196 24624 18202 24676
rect 18233 24667 18291 24673
rect 18233 24633 18245 24667
rect 18279 24633 18291 24667
rect 18233 24627 18291 24633
rect 18785 24667 18843 24673
rect 18785 24633 18797 24667
rect 18831 24664 18843 24667
rect 20346 24664 20352 24676
rect 18831 24636 20352 24664
rect 18831 24633 18843 24636
rect 18785 24627 18843 24633
rect 9631 24599 9689 24605
rect 9631 24565 9643 24599
rect 9677 24596 9689 24599
rect 11698 24596 11704 24608
rect 9677 24568 11704 24596
rect 9677 24565 9689 24568
rect 9631 24559 9689 24565
rect 11698 24556 11704 24568
rect 11756 24556 11762 24608
rect 12575 24599 12633 24605
rect 12575 24565 12587 24599
rect 12621 24596 12633 24599
rect 13630 24596 13636 24608
rect 12621 24568 13636 24596
rect 12621 24565 12633 24568
rect 12575 24559 12633 24565
rect 13630 24556 13636 24568
rect 13688 24556 13694 24608
rect 13725 24599 13783 24605
rect 13725 24565 13737 24599
rect 13771 24596 13783 24599
rect 14734 24596 14740 24608
rect 13771 24568 14740 24596
rect 13771 24565 13783 24568
rect 13725 24559 13783 24565
rect 14734 24556 14740 24568
rect 14792 24556 14798 24608
rect 14875 24599 14933 24605
rect 14875 24565 14887 24599
rect 14921 24596 14933 24599
rect 15746 24596 15752 24608
rect 14921 24568 15752 24596
rect 14921 24565 14933 24568
rect 14875 24559 14933 24565
rect 15746 24556 15752 24568
rect 15804 24556 15810 24608
rect 17862 24596 17868 24608
rect 17775 24568 17868 24596
rect 17862 24556 17868 24568
rect 17920 24596 17926 24608
rect 18248 24596 18276 24627
rect 20346 24624 20352 24636
rect 20404 24624 20410 24676
rect 25498 24664 25504 24676
rect 25459 24636 25504 24664
rect 25498 24624 25504 24636
rect 25556 24624 25562 24676
rect 17920 24568 18276 24596
rect 17920 24556 17926 24568
rect 22002 24556 22008 24608
rect 22060 24596 22066 24608
rect 24719 24599 24777 24605
rect 24719 24596 24731 24599
rect 22060 24568 24731 24596
rect 22060 24556 22066 24568
rect 24719 24565 24731 24568
rect 24765 24565 24777 24599
rect 24719 24559 24777 24565
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 12989 24395 13047 24401
rect 12989 24361 13001 24395
rect 13035 24392 13047 24395
rect 16991 24395 17049 24401
rect 13035 24364 13814 24392
rect 13035 24361 13047 24364
rect 12989 24355 13047 24361
rect 11790 24324 11796 24336
rect 10587 24296 11796 24324
rect 6432 24259 6490 24265
rect 6432 24225 6444 24259
rect 6478 24256 6490 24259
rect 6638 24256 6644 24268
rect 6478 24228 6644 24256
rect 6478 24225 6490 24228
rect 6432 24219 6490 24225
rect 6638 24216 6644 24228
rect 6696 24216 6702 24268
rect 10410 24216 10416 24268
rect 10468 24256 10474 24268
rect 10587 24265 10615 24296
rect 11790 24284 11796 24296
rect 11848 24284 11854 24336
rect 13786 24324 13814 24364
rect 16991 24361 17003 24395
rect 17037 24392 17049 24395
rect 18138 24392 18144 24404
rect 17037 24364 18144 24392
rect 17037 24361 17049 24364
rect 16991 24355 17049 24361
rect 18138 24352 18144 24364
rect 18196 24352 18202 24404
rect 19058 24392 19064 24404
rect 18708 24364 19064 24392
rect 18708 24324 18736 24364
rect 19058 24352 19064 24364
rect 19116 24352 19122 24404
rect 21085 24395 21143 24401
rect 21085 24361 21097 24395
rect 21131 24392 21143 24395
rect 22186 24392 22192 24404
rect 21131 24364 22192 24392
rect 21131 24361 21143 24364
rect 21085 24355 21143 24361
rect 22186 24352 22192 24364
rect 22244 24352 22250 24404
rect 23845 24395 23903 24401
rect 23845 24361 23857 24395
rect 23891 24392 23903 24395
rect 25314 24392 25320 24404
rect 23891 24364 25320 24392
rect 23891 24361 23903 24364
rect 23845 24355 23903 24361
rect 25314 24352 25320 24364
rect 25372 24352 25378 24404
rect 18874 24324 18880 24336
rect 13786 24296 18736 24324
rect 18835 24296 18880 24324
rect 18874 24284 18880 24296
rect 18932 24284 18938 24336
rect 10572 24259 10630 24265
rect 10572 24256 10584 24259
rect 10468 24228 10584 24256
rect 10468 24216 10474 24228
rect 10572 24225 10584 24228
rect 10618 24225 10630 24259
rect 10572 24219 10630 24225
rect 11330 24216 11336 24268
rect 11388 24256 11394 24268
rect 11552 24259 11610 24265
rect 11552 24256 11564 24259
rect 11388 24228 11564 24256
rect 11388 24216 11394 24228
rect 11552 24225 11564 24228
rect 11598 24225 11610 24259
rect 12802 24256 12808 24268
rect 12715 24228 12808 24256
rect 11552 24219 11610 24225
rect 12802 24216 12808 24228
rect 12860 24256 12866 24268
rect 13538 24256 13544 24268
rect 12860 24228 13544 24256
rect 12860 24216 12866 24228
rect 13538 24216 13544 24228
rect 13596 24216 13602 24268
rect 13976 24259 14034 24265
rect 13976 24225 13988 24259
rect 14022 24256 14034 24259
rect 14182 24256 14188 24268
rect 14022 24228 14188 24256
rect 14022 24225 14034 24228
rect 13976 24219 14034 24225
rect 14182 24216 14188 24228
rect 14240 24216 14246 24268
rect 15838 24256 15844 24268
rect 15799 24228 15844 24256
rect 15838 24216 15844 24228
rect 15896 24216 15902 24268
rect 15930 24216 15936 24268
rect 15988 24256 15994 24268
rect 16888 24259 16946 24265
rect 16888 24256 16900 24259
rect 15988 24228 16900 24256
rect 15988 24216 15994 24228
rect 16888 24225 16900 24228
rect 16934 24256 16946 24259
rect 17402 24256 17408 24268
rect 16934 24228 17408 24256
rect 16934 24225 16946 24228
rect 16888 24219 16946 24225
rect 17402 24216 17408 24228
rect 17460 24216 17466 24268
rect 20898 24256 20904 24268
rect 20859 24228 20904 24256
rect 20898 24216 20904 24228
rect 20956 24216 20962 24268
rect 23658 24256 23664 24268
rect 23619 24228 23664 24256
rect 23658 24216 23664 24228
rect 23716 24216 23722 24268
rect 24854 24265 24860 24268
rect 24832 24259 24860 24265
rect 24832 24256 24844 24259
rect 24767 24228 24844 24256
rect 24832 24225 24844 24228
rect 24912 24256 24918 24268
rect 27338 24256 27344 24268
rect 24912 24228 27344 24256
rect 24832 24219 24860 24225
rect 24854 24216 24860 24219
rect 24912 24216 24918 24228
rect 27338 24216 27344 24228
rect 27396 24216 27402 24268
rect 11698 24148 11704 24200
rect 11756 24188 11762 24200
rect 15286 24188 15292 24200
rect 11756 24160 13814 24188
rect 15247 24160 15292 24188
rect 11756 24148 11762 24160
rect 10643 24123 10701 24129
rect 10643 24089 10655 24123
rect 10689 24120 10701 24123
rect 13446 24120 13452 24132
rect 10689 24092 13452 24120
rect 10689 24089 10701 24092
rect 10643 24083 10701 24089
rect 13446 24080 13452 24092
rect 13504 24080 13510 24132
rect 13786 24120 13814 24160
rect 15286 24148 15292 24160
rect 15344 24148 15350 24200
rect 18782 24188 18788 24200
rect 18743 24160 18788 24188
rect 18782 24148 18788 24160
rect 18840 24148 18846 24200
rect 18966 24148 18972 24200
rect 19024 24188 19030 24200
rect 19061 24191 19119 24197
rect 19061 24188 19073 24191
rect 19024 24160 19073 24188
rect 19024 24148 19030 24160
rect 19061 24157 19073 24160
rect 19107 24157 19119 24191
rect 19061 24151 19119 24157
rect 18322 24120 18328 24132
rect 13786 24092 18328 24120
rect 18322 24080 18328 24092
rect 18380 24080 18386 24132
rect 6503 24055 6561 24061
rect 6503 24021 6515 24055
rect 6549 24052 6561 24055
rect 6822 24052 6828 24064
rect 6549 24024 6828 24052
rect 6549 24021 6561 24024
rect 6503 24015 6561 24021
rect 6822 24012 6828 24024
rect 6880 24012 6886 24064
rect 11655 24055 11713 24061
rect 11655 24021 11667 24055
rect 11701 24052 11713 24055
rect 13722 24052 13728 24064
rect 11701 24024 13728 24052
rect 11701 24021 11713 24024
rect 11655 24015 11713 24021
rect 13722 24012 13728 24024
rect 13780 24012 13786 24064
rect 14047 24055 14105 24061
rect 14047 24021 14059 24055
rect 14093 24052 14105 24055
rect 18506 24052 18512 24064
rect 14093 24024 18512 24052
rect 14093 24021 14105 24024
rect 14047 24015 14105 24021
rect 18506 24012 18512 24024
rect 18564 24012 18570 24064
rect 19794 24052 19800 24064
rect 19755 24024 19800 24052
rect 19794 24012 19800 24024
rect 19852 24012 19858 24064
rect 24118 24012 24124 24064
rect 24176 24052 24182 24064
rect 24903 24055 24961 24061
rect 24903 24052 24915 24055
rect 24176 24024 24915 24052
rect 24176 24012 24182 24024
rect 24903 24021 24915 24024
rect 24949 24021 24961 24055
rect 24903 24015 24961 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 3694 23848 3700 23860
rect 3655 23820 3700 23848
rect 3694 23808 3700 23820
rect 3752 23808 3758 23860
rect 5534 23808 5540 23860
rect 5592 23848 5598 23860
rect 5813 23851 5871 23857
rect 5813 23848 5825 23851
rect 5592 23820 5825 23848
rect 5592 23808 5598 23820
rect 5813 23817 5825 23820
rect 5859 23817 5871 23851
rect 5813 23811 5871 23817
rect 6457 23851 6515 23857
rect 6457 23817 6469 23851
rect 6503 23848 6515 23851
rect 6638 23848 6644 23860
rect 6503 23820 6644 23848
rect 6503 23817 6515 23820
rect 6457 23811 6515 23817
rect 6638 23808 6644 23820
rect 6696 23808 6702 23860
rect 7834 23848 7840 23860
rect 7795 23820 7840 23848
rect 7834 23808 7840 23820
rect 7892 23808 7898 23860
rect 8938 23848 8944 23860
rect 8899 23820 8944 23848
rect 8938 23808 8944 23820
rect 8996 23808 9002 23860
rect 10410 23848 10416 23860
rect 10371 23820 10416 23848
rect 10410 23808 10416 23820
rect 10468 23808 10474 23860
rect 13538 23848 13544 23860
rect 13499 23820 13544 23848
rect 13538 23808 13544 23820
rect 13596 23808 13602 23860
rect 13906 23848 13912 23860
rect 13867 23820 13912 23848
rect 13906 23808 13912 23820
rect 13964 23808 13970 23860
rect 14182 23808 14188 23860
rect 14240 23848 14246 23860
rect 14277 23851 14335 23857
rect 14277 23848 14289 23851
rect 14240 23820 14289 23848
rect 14240 23808 14246 23820
rect 14277 23817 14289 23820
rect 14323 23817 14335 23851
rect 14277 23811 14335 23817
rect 15470 23808 15476 23860
rect 15528 23848 15534 23860
rect 15838 23848 15844 23860
rect 15528 23820 15844 23848
rect 15528 23808 15534 23820
rect 15838 23808 15844 23820
rect 15896 23808 15902 23860
rect 17402 23848 17408 23860
rect 17363 23820 17408 23848
rect 17402 23808 17408 23820
rect 17460 23808 17466 23860
rect 17862 23848 17868 23860
rect 17823 23820 17868 23848
rect 17862 23808 17868 23820
rect 17920 23808 17926 23860
rect 18874 23808 18880 23860
rect 18932 23848 18938 23860
rect 19150 23848 19156 23860
rect 18932 23820 19156 23848
rect 18932 23808 18938 23820
rect 19150 23808 19156 23820
rect 19208 23808 19214 23860
rect 20898 23848 20904 23860
rect 20859 23820 20904 23848
rect 20898 23808 20904 23820
rect 20956 23808 20962 23860
rect 21453 23851 21511 23857
rect 21453 23817 21465 23851
rect 21499 23848 21511 23851
rect 23198 23848 23204 23860
rect 21499 23820 23204 23848
rect 21499 23817 21511 23820
rect 21453 23811 21511 23817
rect 23198 23808 23204 23820
rect 23256 23808 23262 23860
rect 24854 23848 24860 23860
rect 24815 23820 24860 23848
rect 24854 23808 24860 23820
rect 24912 23808 24918 23860
rect 25409 23851 25467 23857
rect 25409 23817 25421 23851
rect 25455 23848 25467 23851
rect 26326 23848 26332 23860
rect 25455 23820 26332 23848
rect 25455 23817 25467 23820
rect 25409 23811 25467 23817
rect 26326 23808 26332 23820
rect 26384 23808 26390 23860
rect 10045 23783 10103 23789
rect 10045 23749 10057 23783
rect 10091 23780 10103 23783
rect 10778 23780 10784 23792
rect 10091 23752 10784 23780
rect 10091 23749 10103 23752
rect 10045 23743 10103 23749
rect 474 23604 480 23656
rect 532 23644 538 23656
rect 1432 23647 1490 23653
rect 1432 23644 1444 23647
rect 532 23616 1444 23644
rect 532 23604 538 23616
rect 1432 23613 1444 23616
rect 1478 23644 1490 23647
rect 1857 23647 1915 23653
rect 1857 23644 1869 23647
rect 1478 23616 1869 23644
rect 1478 23613 1490 23616
rect 1432 23607 1490 23613
rect 1857 23613 1869 23616
rect 1903 23613 1915 23647
rect 1857 23607 1915 23613
rect 3288 23647 3346 23653
rect 3288 23613 3300 23647
rect 3334 23644 3346 23647
rect 3694 23644 3700 23656
rect 3334 23616 3700 23644
rect 3334 23613 3346 23616
rect 3288 23607 3346 23613
rect 3694 23604 3700 23616
rect 3752 23604 3758 23656
rect 5420 23647 5478 23653
rect 5420 23613 5432 23647
rect 5466 23644 5478 23647
rect 5534 23644 5540 23656
rect 5466 23616 5540 23644
rect 5466 23613 5478 23616
rect 5420 23607 5478 23613
rect 5534 23604 5540 23616
rect 5592 23604 5598 23656
rect 7444 23647 7502 23653
rect 7444 23613 7456 23647
rect 7490 23644 7502 23647
rect 7834 23644 7840 23656
rect 7490 23616 7840 23644
rect 7490 23613 7502 23616
rect 7444 23607 7502 23613
rect 7834 23604 7840 23616
rect 7892 23604 7898 23656
rect 8548 23647 8606 23653
rect 8548 23613 8560 23647
rect 8594 23644 8606 23647
rect 8938 23644 8944 23656
rect 8594 23616 8944 23644
rect 8594 23613 8606 23616
rect 8548 23607 8606 23613
rect 8938 23604 8944 23616
rect 8996 23604 9002 23656
rect 9560 23647 9618 23653
rect 9560 23613 9572 23647
rect 9606 23644 9618 23647
rect 10060 23644 10088 23743
rect 10778 23740 10784 23752
rect 10836 23740 10842 23792
rect 12805 23783 12863 23789
rect 12805 23749 12817 23783
rect 12851 23780 12863 23783
rect 17034 23780 17040 23792
rect 12851 23752 16963 23780
rect 16995 23752 17040 23780
rect 12851 23749 12863 23752
rect 12805 23743 12863 23749
rect 14734 23672 14740 23724
rect 14792 23712 14798 23724
rect 14921 23715 14979 23721
rect 14921 23712 14933 23715
rect 14792 23684 14933 23712
rect 14792 23672 14798 23684
rect 14921 23681 14933 23684
rect 14967 23681 14979 23715
rect 15562 23712 15568 23724
rect 15523 23684 15568 23712
rect 14921 23675 14979 23681
rect 15562 23672 15568 23684
rect 15620 23672 15626 23724
rect 16935 23712 16963 23752
rect 17034 23740 17040 23752
rect 17092 23740 17098 23792
rect 20346 23780 20352 23792
rect 20307 23752 20352 23780
rect 20346 23740 20352 23752
rect 20404 23740 20410 23792
rect 18046 23712 18052 23724
rect 16935 23684 18052 23712
rect 18046 23672 18052 23684
rect 18104 23672 18110 23724
rect 19794 23712 19800 23724
rect 19707 23684 19800 23712
rect 19794 23672 19800 23684
rect 19852 23712 19858 23724
rect 21358 23712 21364 23724
rect 19852 23684 21364 23712
rect 19852 23672 19858 23684
rect 21358 23672 21364 23684
rect 21416 23672 21422 23724
rect 11054 23644 11060 23656
rect 9606 23616 10088 23644
rect 11015 23616 11060 23644
rect 9606 23613 9618 23616
rect 9560 23607 9618 23613
rect 11054 23604 11060 23616
rect 11112 23604 11118 23656
rect 12618 23644 12624 23656
rect 12531 23616 12624 23644
rect 12618 23604 12624 23616
rect 12676 23644 12682 23656
rect 13173 23647 13231 23653
rect 13173 23644 13185 23647
rect 12676 23616 13185 23644
rect 12676 23604 12682 23616
rect 13173 23613 13185 23616
rect 13219 23613 13231 23647
rect 13722 23644 13728 23656
rect 13683 23616 13728 23644
rect 13173 23607 13231 23613
rect 13722 23604 13728 23616
rect 13780 23604 13786 23656
rect 16761 23647 16819 23653
rect 16761 23613 16773 23647
rect 16807 23644 16819 23647
rect 16853 23647 16911 23653
rect 16853 23644 16865 23647
rect 16807 23616 16865 23644
rect 16807 23613 16819 23616
rect 16761 23607 16819 23613
rect 16853 23613 16865 23616
rect 16899 23644 16911 23647
rect 17034 23644 17040 23656
rect 16899 23616 17040 23644
rect 16899 23613 16911 23616
rect 16853 23607 16911 23613
rect 17034 23604 17040 23616
rect 17092 23604 17098 23656
rect 17862 23604 17868 23656
rect 17920 23644 17926 23656
rect 18138 23644 18144 23656
rect 17920 23616 18144 23644
rect 17920 23604 17926 23616
rect 18138 23604 18144 23616
rect 18196 23644 18202 23656
rect 18233 23647 18291 23653
rect 18233 23644 18245 23647
rect 18196 23616 18245 23644
rect 18196 23604 18202 23616
rect 18233 23613 18245 23616
rect 18279 23613 18291 23647
rect 21266 23644 21272 23656
rect 21179 23616 21272 23644
rect 18233 23607 18291 23613
rect 21266 23604 21272 23616
rect 21324 23644 21330 23656
rect 21821 23647 21879 23653
rect 21821 23644 21833 23647
rect 21324 23616 21833 23644
rect 21324 23604 21330 23616
rect 21821 23613 21833 23616
rect 21867 23613 21879 23647
rect 21821 23607 21879 23613
rect 22186 23604 22192 23656
rect 22244 23644 22250 23656
rect 23477 23647 23535 23653
rect 23477 23644 23489 23647
rect 22244 23616 23489 23644
rect 22244 23604 22250 23616
rect 23477 23613 23489 23616
rect 23523 23644 23535 23647
rect 23753 23647 23811 23653
rect 23753 23644 23765 23647
rect 23523 23616 23765 23644
rect 23523 23613 23535 23616
rect 23477 23607 23535 23613
rect 23753 23613 23765 23616
rect 23799 23613 23811 23647
rect 25222 23644 25228 23656
rect 25135 23616 25228 23644
rect 23753 23607 23811 23613
rect 25222 23604 25228 23616
rect 25280 23644 25286 23656
rect 25777 23647 25835 23653
rect 25777 23644 25789 23647
rect 25280 23616 25789 23644
rect 25280 23604 25286 23616
rect 25777 23613 25789 23616
rect 25823 23613 25835 23647
rect 25777 23607 25835 23613
rect 3375 23579 3433 23585
rect 3375 23545 3387 23579
rect 3421 23576 3433 23579
rect 15013 23579 15071 23585
rect 3421 23548 4154 23576
rect 3421 23545 3433 23548
rect 3375 23539 3433 23545
rect 1535 23511 1593 23517
rect 1535 23477 1547 23511
rect 1581 23508 1593 23511
rect 1670 23508 1676 23520
rect 1581 23480 1676 23508
rect 1581 23477 1593 23480
rect 1535 23471 1593 23477
rect 1670 23468 1676 23480
rect 1728 23468 1734 23520
rect 4126 23508 4154 23548
rect 15013 23545 15025 23579
rect 15059 23576 15071 23579
rect 15286 23576 15292 23588
rect 15059 23548 15292 23576
rect 15059 23545 15071 23548
rect 15013 23539 15071 23545
rect 5350 23508 5356 23520
rect 4126 23480 5356 23508
rect 5350 23468 5356 23480
rect 5408 23468 5414 23520
rect 5491 23511 5549 23517
rect 5491 23477 5503 23511
rect 5537 23508 5549 23511
rect 7374 23508 7380 23520
rect 5537 23480 7380 23508
rect 5537 23477 5549 23480
rect 5491 23471 5549 23477
rect 7374 23468 7380 23480
rect 7432 23468 7438 23520
rect 7515 23511 7573 23517
rect 7515 23477 7527 23511
rect 7561 23508 7573 23511
rect 7650 23508 7656 23520
rect 7561 23480 7656 23508
rect 7561 23477 7573 23480
rect 7515 23471 7573 23477
rect 7650 23468 7656 23480
rect 7708 23468 7714 23520
rect 8619 23511 8677 23517
rect 8619 23477 8631 23511
rect 8665 23508 8677 23511
rect 8754 23508 8760 23520
rect 8665 23480 8760 23508
rect 8665 23477 8677 23480
rect 8619 23471 8677 23477
rect 8754 23468 8760 23480
rect 8812 23468 8818 23520
rect 9490 23468 9496 23520
rect 9548 23508 9554 23520
rect 9631 23511 9689 23517
rect 9631 23508 9643 23511
rect 9548 23480 9643 23508
rect 9548 23468 9554 23480
rect 9631 23477 9643 23480
rect 9677 23477 9689 23511
rect 10778 23508 10784 23520
rect 10739 23480 10784 23508
rect 9631 23471 9689 23477
rect 10778 23468 10784 23480
rect 10836 23468 10842 23520
rect 11330 23468 11336 23520
rect 11388 23508 11394 23520
rect 11517 23511 11575 23517
rect 11517 23508 11529 23511
rect 11388 23480 11529 23508
rect 11388 23468 11394 23480
rect 11517 23477 11529 23480
rect 11563 23477 11575 23511
rect 11517 23471 11575 23477
rect 14737 23511 14795 23517
rect 14737 23477 14749 23511
rect 14783 23508 14795 23511
rect 15028 23508 15056 23539
rect 15286 23536 15292 23548
rect 15344 23536 15350 23588
rect 18877 23579 18935 23585
rect 18877 23545 18889 23579
rect 18923 23576 18935 23579
rect 19521 23579 19579 23585
rect 19521 23576 19533 23579
rect 18923 23548 19533 23576
rect 18923 23545 18935 23548
rect 18877 23539 18935 23545
rect 19521 23545 19533 23548
rect 19567 23545 19579 23579
rect 19521 23539 19579 23545
rect 19889 23579 19947 23585
rect 19889 23545 19901 23579
rect 19935 23545 19947 23579
rect 19889 23539 19947 23545
rect 23109 23579 23167 23585
rect 23109 23545 23121 23579
rect 23155 23576 23167 23579
rect 23658 23576 23664 23588
rect 23155 23548 23664 23576
rect 23155 23545 23167 23548
rect 23109 23539 23167 23545
rect 14783 23480 15056 23508
rect 19536 23508 19564 23539
rect 19904 23508 19932 23539
rect 23658 23536 23664 23548
rect 23716 23536 23722 23588
rect 23934 23508 23940 23520
rect 19536 23480 19932 23508
rect 23895 23480 23940 23508
rect 14783 23477 14795 23480
rect 14737 23471 14795 23477
rect 23934 23468 23940 23480
rect 23992 23468 23998 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 12391 23307 12449 23313
rect 12391 23273 12403 23307
rect 12437 23304 12449 23307
rect 12618 23304 12624 23316
rect 12437 23276 12624 23304
rect 12437 23273 12449 23276
rect 12391 23267 12449 23273
rect 12618 23264 12624 23276
rect 12676 23264 12682 23316
rect 14734 23264 14740 23316
rect 14792 23304 14798 23316
rect 14829 23307 14887 23313
rect 14829 23304 14841 23307
rect 14792 23276 14841 23304
rect 14792 23264 14798 23276
rect 14829 23273 14841 23276
rect 14875 23273 14887 23307
rect 14829 23267 14887 23273
rect 18782 23264 18788 23316
rect 18840 23304 18846 23316
rect 19245 23307 19303 23313
rect 19245 23304 19257 23307
rect 18840 23276 19257 23304
rect 18840 23264 18846 23276
rect 19245 23273 19257 23276
rect 19291 23304 19303 23307
rect 19889 23307 19947 23313
rect 19291 23276 19472 23304
rect 19291 23273 19303 23276
rect 19245 23267 19303 23273
rect 10594 23196 10600 23248
rect 10652 23236 10658 23248
rect 10778 23236 10784 23248
rect 10652 23208 10784 23236
rect 10652 23196 10658 23208
rect 10778 23196 10784 23208
rect 10836 23236 10842 23248
rect 10873 23239 10931 23245
rect 10873 23236 10885 23239
rect 10836 23208 10885 23236
rect 10836 23196 10842 23208
rect 10873 23205 10885 23208
rect 10919 23205 10931 23239
rect 10873 23199 10931 23205
rect 13170 23196 13176 23248
rect 13228 23236 13234 23248
rect 13449 23239 13507 23245
rect 13449 23236 13461 23239
rect 13228 23208 13461 23236
rect 13228 23196 13234 23208
rect 13449 23205 13461 23208
rect 13495 23205 13507 23239
rect 15470 23236 15476 23248
rect 15431 23208 15476 23236
rect 13449 23199 13507 23205
rect 15470 23196 15476 23208
rect 15528 23196 15534 23248
rect 18877 23239 18935 23245
rect 18877 23205 18889 23239
rect 18923 23236 18935 23239
rect 19150 23236 19156 23248
rect 18923 23208 19156 23236
rect 18923 23205 18935 23208
rect 18877 23199 18935 23205
rect 19150 23196 19156 23208
rect 19208 23196 19214 23248
rect 19444 23236 19472 23276
rect 19889 23273 19901 23307
rect 19935 23304 19947 23307
rect 20806 23304 20812 23316
rect 19935 23276 20812 23304
rect 19935 23273 19947 23276
rect 19889 23267 19947 23273
rect 20806 23264 20812 23276
rect 20864 23264 20870 23316
rect 21039 23307 21097 23313
rect 21039 23273 21051 23307
rect 21085 23304 21097 23307
rect 21266 23304 21272 23316
rect 21085 23276 21272 23304
rect 21085 23273 21097 23276
rect 21039 23267 21097 23273
rect 21266 23264 21272 23276
rect 21324 23264 21330 23316
rect 21358 23264 21364 23316
rect 21416 23304 21422 23316
rect 25363 23307 25421 23313
rect 25363 23304 25375 23307
rect 21416 23276 25375 23304
rect 21416 23264 21422 23276
rect 25363 23273 25375 23276
rect 25409 23273 25421 23307
rect 25363 23267 25421 23273
rect 22002 23236 22008 23248
rect 19444 23208 22008 23236
rect 22002 23196 22008 23208
rect 22060 23196 22066 23248
rect 22186 23196 22192 23248
rect 22244 23236 22250 23248
rect 22281 23239 22339 23245
rect 22281 23236 22293 23239
rect 22244 23208 22293 23236
rect 22244 23196 22250 23208
rect 22281 23205 22293 23208
rect 22327 23205 22339 23239
rect 22281 23199 22339 23205
rect 23750 23196 23756 23248
rect 23808 23236 23814 23248
rect 23845 23239 23903 23245
rect 23845 23236 23857 23239
rect 23808 23208 23857 23236
rect 23808 23196 23814 23208
rect 23845 23205 23857 23208
rect 23891 23236 23903 23239
rect 23934 23236 23940 23248
rect 23891 23208 23940 23236
rect 23891 23205 23903 23208
rect 23845 23199 23903 23205
rect 23934 23196 23940 23208
rect 23992 23196 23998 23248
rect 2498 23128 2504 23180
rect 2556 23168 2562 23180
rect 8294 23168 8300 23180
rect 8352 23177 8358 23180
rect 8352 23171 8390 23177
rect 2556 23140 8300 23168
rect 2556 23128 2562 23140
rect 8294 23128 8300 23140
rect 8378 23137 8390 23171
rect 12250 23168 12256 23180
rect 12211 23140 12256 23168
rect 8352 23131 8390 23137
rect 8352 23128 8358 23131
rect 12250 23128 12256 23140
rect 12308 23128 12314 23180
rect 17164 23171 17222 23177
rect 17164 23168 17176 23171
rect 17144 23137 17176 23168
rect 17210 23137 17222 23171
rect 18230 23168 18236 23180
rect 18191 23140 18236 23168
rect 17144 23131 17222 23137
rect 9677 23103 9735 23109
rect 9677 23069 9689 23103
rect 9723 23100 9735 23103
rect 10134 23100 10140 23112
rect 9723 23072 10140 23100
rect 9723 23069 9735 23072
rect 9677 23063 9735 23069
rect 10134 23060 10140 23072
rect 10192 23100 10198 23112
rect 10781 23103 10839 23109
rect 10781 23100 10793 23103
rect 10192 23072 10793 23100
rect 10192 23060 10198 23072
rect 10781 23069 10793 23072
rect 10827 23069 10839 23103
rect 13354 23100 13360 23112
rect 10781 23063 10839 23069
rect 10888 23072 13360 23100
rect 5350 22992 5356 23044
rect 5408 23032 5414 23044
rect 10888 23032 10916 23072
rect 13354 23060 13360 23072
rect 13412 23060 13418 23112
rect 14001 23103 14059 23109
rect 14001 23069 14013 23103
rect 14047 23100 14059 23103
rect 14274 23100 14280 23112
rect 14047 23072 14280 23100
rect 14047 23069 14059 23072
rect 14001 23063 14059 23069
rect 14274 23060 14280 23072
rect 14332 23100 14338 23112
rect 15378 23100 15384 23112
rect 14332 23072 15384 23100
rect 14332 23060 14338 23072
rect 15378 23060 15384 23072
rect 15436 23060 15442 23112
rect 15562 23060 15568 23112
rect 15620 23100 15626 23112
rect 15657 23103 15715 23109
rect 15657 23100 15669 23103
rect 15620 23072 15669 23100
rect 15620 23060 15626 23072
rect 15657 23069 15669 23072
rect 15703 23069 15715 23103
rect 15657 23063 15715 23069
rect 11330 23032 11336 23044
rect 5408 23004 10916 23032
rect 11291 23004 11336 23032
rect 5408 22992 5414 23004
rect 11330 22992 11336 23004
rect 11388 22992 11394 23044
rect 17144 22976 17172 23131
rect 18230 23128 18236 23140
rect 18288 23128 18294 23180
rect 19702 23168 19708 23180
rect 19663 23140 19708 23168
rect 19702 23128 19708 23140
rect 19760 23128 19766 23180
rect 20806 23128 20812 23180
rect 20864 23168 20870 23180
rect 20936 23171 20994 23177
rect 20936 23168 20948 23171
rect 20864 23140 20948 23168
rect 20864 23128 20870 23140
rect 20936 23137 20948 23140
rect 20982 23137 20994 23171
rect 20936 23131 20994 23137
rect 25292 23171 25350 23177
rect 25292 23137 25304 23171
rect 25338 23168 25350 23171
rect 26142 23168 26148 23180
rect 25338 23140 26148 23168
rect 25338 23137 25350 23140
rect 25292 23131 25350 23137
rect 26142 23128 26148 23140
rect 26200 23128 26206 23180
rect 18506 23060 18512 23112
rect 18564 23100 18570 23112
rect 22189 23103 22247 23109
rect 22189 23100 22201 23103
rect 18564 23072 22201 23100
rect 18564 23060 18570 23072
rect 22189 23069 22201 23072
rect 22235 23100 22247 23103
rect 22462 23100 22468 23112
rect 22235 23072 22468 23100
rect 22235 23069 22247 23072
rect 22189 23063 22247 23069
rect 22462 23060 22468 23072
rect 22520 23060 22526 23112
rect 23753 23103 23811 23109
rect 23753 23069 23765 23103
rect 23799 23100 23811 23103
rect 24026 23100 24032 23112
rect 23799 23072 24032 23100
rect 23799 23069 23811 23072
rect 23753 23063 23811 23069
rect 24026 23060 24032 23072
rect 24084 23060 24090 23112
rect 17267 23035 17325 23041
rect 17267 23001 17279 23035
rect 17313 23032 17325 23035
rect 20898 23032 20904 23044
rect 17313 23004 20904 23032
rect 17313 23001 17325 23004
rect 17267 22995 17325 23001
rect 20898 22992 20904 23004
rect 20956 22992 20962 23044
rect 22741 23035 22799 23041
rect 22741 23001 22753 23035
rect 22787 23032 22799 23035
rect 23934 23032 23940 23044
rect 22787 23004 23940 23032
rect 22787 23001 22799 23004
rect 22741 22995 22799 23001
rect 23934 22992 23940 23004
rect 23992 23032 23998 23044
rect 24305 23035 24363 23041
rect 24305 23032 24317 23035
rect 23992 23004 24317 23032
rect 23992 22992 23998 23004
rect 24305 23001 24317 23004
rect 24351 23001 24363 23035
rect 24305 22995 24363 23001
rect 8435 22967 8493 22973
rect 8435 22933 8447 22967
rect 8481 22964 8493 22967
rect 9214 22964 9220 22976
rect 8481 22936 9220 22964
rect 8481 22933 8493 22936
rect 8435 22927 8493 22933
rect 9214 22924 9220 22936
rect 9272 22924 9278 22976
rect 10597 22967 10655 22973
rect 10597 22933 10609 22967
rect 10643 22964 10655 22967
rect 11054 22964 11060 22976
rect 10643 22936 11060 22964
rect 10643 22933 10655 22936
rect 10597 22927 10655 22933
rect 11054 22924 11060 22936
rect 11112 22924 11118 22976
rect 14366 22964 14372 22976
rect 14327 22936 14372 22964
rect 14366 22924 14372 22936
rect 14424 22924 14430 22976
rect 16482 22964 16488 22976
rect 16443 22936 16488 22964
rect 16482 22924 16488 22936
rect 16540 22924 16546 22976
rect 17126 22924 17132 22976
rect 17184 22964 17190 22976
rect 17589 22967 17647 22973
rect 17589 22964 17601 22967
rect 17184 22936 17601 22964
rect 17184 22924 17190 22936
rect 17589 22933 17601 22936
rect 17635 22933 17647 22967
rect 17589 22927 17647 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 8294 22760 8300 22772
rect 8255 22732 8300 22760
rect 8294 22720 8300 22732
rect 8352 22720 8358 22772
rect 10134 22760 10140 22772
rect 10095 22732 10140 22760
rect 10134 22720 10140 22732
rect 10192 22720 10198 22772
rect 10594 22760 10600 22772
rect 10555 22732 10600 22760
rect 10594 22720 10600 22732
rect 10652 22720 10658 22772
rect 12575 22763 12633 22769
rect 12575 22729 12587 22763
rect 12621 22760 12633 22763
rect 12802 22760 12808 22772
rect 12621 22732 12808 22760
rect 12621 22729 12633 22732
rect 12575 22723 12633 22729
rect 12802 22720 12808 22732
rect 12860 22720 12866 22772
rect 13354 22720 13360 22772
rect 13412 22760 13418 22772
rect 14921 22763 14979 22769
rect 14921 22760 14933 22763
rect 13412 22732 14933 22760
rect 13412 22720 13418 22732
rect 14921 22729 14933 22732
rect 14967 22729 14979 22763
rect 14921 22723 14979 22729
rect 15378 22720 15384 22772
rect 15436 22760 15442 22772
rect 15657 22763 15715 22769
rect 15657 22760 15669 22763
rect 15436 22732 15669 22760
rect 15436 22720 15442 22732
rect 15657 22729 15669 22732
rect 15703 22729 15715 22763
rect 15657 22723 15715 22729
rect 15838 22720 15844 22772
rect 15896 22760 15902 22772
rect 17405 22763 17463 22769
rect 17405 22760 17417 22763
rect 15896 22732 17417 22760
rect 15896 22720 15902 22732
rect 17405 22729 17417 22732
rect 17451 22729 17463 22763
rect 17405 22723 17463 22729
rect 11330 22692 11336 22704
rect 11291 22664 11336 22692
rect 11330 22652 11336 22664
rect 11388 22652 11394 22704
rect 14366 22692 14372 22704
rect 14016 22664 14372 22692
rect 9214 22624 9220 22636
rect 9175 22596 9220 22624
rect 9214 22584 9220 22596
rect 9272 22584 9278 22636
rect 11698 22584 11704 22636
rect 11756 22624 11762 22636
rect 12250 22624 12256 22636
rect 11756 22596 12256 22624
rect 11756 22584 11762 22596
rect 12250 22584 12256 22596
rect 12308 22624 12314 22636
rect 14016 22633 14044 22664
rect 14366 22652 14372 22664
rect 14424 22692 14430 22704
rect 14734 22692 14740 22704
rect 14424 22664 14740 22692
rect 14424 22652 14430 22664
rect 14734 22652 14740 22664
rect 14792 22652 14798 22704
rect 12897 22627 12955 22633
rect 12897 22624 12909 22627
rect 12308 22596 12909 22624
rect 12308 22584 12314 22596
rect 12897 22593 12909 22596
rect 12943 22593 12955 22627
rect 12897 22587 12955 22593
rect 14001 22627 14059 22633
rect 14001 22593 14013 22627
rect 14047 22593 14059 22627
rect 14274 22624 14280 22636
rect 14235 22596 14280 22624
rect 14001 22587 14059 22593
rect 14274 22584 14280 22596
rect 14332 22584 14338 22636
rect 17420 22624 17448 22723
rect 17954 22720 17960 22772
rect 18012 22760 18018 22772
rect 19061 22763 19119 22769
rect 19061 22760 19073 22763
rect 18012 22732 19073 22760
rect 18012 22720 18018 22732
rect 19061 22729 19073 22732
rect 19107 22760 19119 22763
rect 19702 22760 19708 22772
rect 19107 22732 19708 22760
rect 19107 22729 19119 22732
rect 19061 22723 19119 22729
rect 19702 22720 19708 22732
rect 19760 22720 19766 22772
rect 25774 22760 25780 22772
rect 25735 22732 25780 22760
rect 25774 22720 25780 22732
rect 25832 22720 25838 22772
rect 26142 22760 26148 22772
rect 26103 22732 26148 22760
rect 26142 22720 26148 22732
rect 26200 22720 26206 22772
rect 22649 22695 22707 22701
rect 22649 22661 22661 22695
rect 22695 22692 22707 22695
rect 23566 22692 23572 22704
rect 22695 22664 23572 22692
rect 22695 22661 22707 22664
rect 22649 22655 22707 22661
rect 23566 22652 23572 22664
rect 23624 22692 23630 22704
rect 23624 22664 24072 22692
rect 23624 22652 23630 22664
rect 18141 22627 18199 22633
rect 18141 22624 18153 22627
rect 17420 22596 18153 22624
rect 18141 22593 18153 22596
rect 18187 22593 18199 22627
rect 18141 22587 18199 22593
rect 23109 22627 23167 22633
rect 23109 22593 23121 22627
rect 23155 22624 23167 22627
rect 23753 22627 23811 22633
rect 23753 22624 23765 22627
rect 23155 22596 23765 22624
rect 23155 22593 23167 22596
rect 23109 22587 23167 22593
rect 23753 22593 23765 22596
rect 23799 22624 23811 22627
rect 23842 22624 23848 22636
rect 23799 22596 23848 22624
rect 23799 22593 23811 22596
rect 23753 22587 23811 22593
rect 23842 22584 23848 22596
rect 23900 22584 23906 22636
rect 24044 22633 24072 22664
rect 24029 22627 24087 22633
rect 24029 22593 24041 22627
rect 24075 22593 24087 22627
rect 24029 22587 24087 22593
rect 12472 22559 12530 22565
rect 12472 22556 12484 22559
rect 12268 22528 12484 22556
rect 9309 22491 9367 22497
rect 9309 22457 9321 22491
rect 9355 22457 9367 22491
rect 9309 22451 9367 22457
rect 9861 22491 9919 22497
rect 9861 22457 9873 22491
rect 9907 22488 9919 22491
rect 10778 22488 10784 22500
rect 9907 22460 10784 22488
rect 9907 22457 9919 22460
rect 9861 22451 9919 22457
rect 9030 22420 9036 22432
rect 8991 22392 9036 22420
rect 9030 22380 9036 22392
rect 9088 22420 9094 22432
rect 9324 22420 9352 22451
rect 10778 22448 10784 22460
rect 10836 22448 10842 22500
rect 10873 22491 10931 22497
rect 10873 22457 10885 22491
rect 10919 22488 10931 22491
rect 11054 22488 11060 22500
rect 10919 22460 11060 22488
rect 10919 22457 10931 22460
rect 10873 22451 10931 22457
rect 11054 22448 11060 22460
rect 11112 22448 11118 22500
rect 9088 22392 9352 22420
rect 10796 22420 10824 22448
rect 12268 22432 12296 22528
rect 12472 22525 12484 22528
rect 12518 22525 12530 22559
rect 12472 22519 12530 22525
rect 19426 22516 19432 22568
rect 19484 22556 19490 22568
rect 19521 22559 19579 22565
rect 19521 22556 19533 22559
rect 19484 22528 19533 22556
rect 19484 22516 19490 22528
rect 19521 22525 19533 22528
rect 19567 22556 19579 22559
rect 19705 22559 19763 22565
rect 19705 22556 19717 22559
rect 19567 22528 19717 22556
rect 19567 22525 19579 22528
rect 19521 22519 19579 22525
rect 19705 22525 19717 22528
rect 19751 22525 19763 22559
rect 19705 22519 19763 22525
rect 25292 22559 25350 22565
rect 25292 22525 25304 22559
rect 25338 22556 25350 22559
rect 25774 22556 25780 22568
rect 25338 22528 25780 22556
rect 25338 22525 25350 22528
rect 25292 22519 25350 22525
rect 25774 22516 25780 22528
rect 25832 22516 25838 22568
rect 14093 22491 14151 22497
rect 14093 22457 14105 22491
rect 14139 22457 14151 22491
rect 14093 22451 14151 22457
rect 11701 22423 11759 22429
rect 11701 22420 11713 22423
rect 10796 22392 11713 22420
rect 9088 22380 9094 22392
rect 11701 22389 11713 22392
rect 11747 22389 11759 22423
rect 12250 22420 12256 22432
rect 12211 22392 12256 22420
rect 11701 22383 11759 22389
rect 12250 22380 12256 22392
rect 12308 22380 12314 22432
rect 13170 22380 13176 22432
rect 13228 22420 13234 22432
rect 13265 22423 13323 22429
rect 13265 22420 13277 22423
rect 13228 22392 13277 22420
rect 13228 22380 13234 22392
rect 13265 22389 13277 22392
rect 13311 22389 13323 22423
rect 13265 22383 13323 22389
rect 13814 22380 13820 22432
rect 13872 22420 13878 22432
rect 14108 22420 14136 22451
rect 15378 22448 15384 22500
rect 15436 22488 15442 22500
rect 16482 22488 16488 22500
rect 15436 22460 16488 22488
rect 15436 22448 15442 22460
rect 16482 22448 16488 22460
rect 16540 22448 16546 22500
rect 16577 22491 16635 22497
rect 16577 22457 16589 22491
rect 16623 22457 16635 22491
rect 17126 22488 17132 22500
rect 17087 22460 17132 22488
rect 16577 22451 16635 22457
rect 13872 22392 14136 22420
rect 13872 22380 13878 22392
rect 14366 22380 14372 22432
rect 14424 22420 14430 22432
rect 15289 22423 15347 22429
rect 15289 22420 15301 22423
rect 14424 22392 15301 22420
rect 14424 22380 14430 22392
rect 15289 22389 15301 22392
rect 15335 22420 15347 22423
rect 15470 22420 15476 22432
rect 15335 22392 15476 22420
rect 15335 22389 15347 22392
rect 15289 22383 15347 22389
rect 15470 22380 15476 22392
rect 15528 22380 15534 22432
rect 16298 22420 16304 22432
rect 16259 22392 16304 22420
rect 16298 22380 16304 22392
rect 16356 22420 16362 22432
rect 16592 22420 16620 22451
rect 17126 22448 17132 22460
rect 17184 22448 17190 22500
rect 18230 22448 18236 22500
rect 18288 22488 18294 22500
rect 18782 22488 18788 22500
rect 18288 22460 18333 22488
rect 18743 22460 18788 22488
rect 18288 22448 18294 22460
rect 18782 22448 18788 22460
rect 18840 22448 18846 22500
rect 19242 22448 19248 22500
rect 19300 22488 19306 22500
rect 20806 22488 20812 22500
rect 19300 22460 20812 22488
rect 19300 22448 19306 22460
rect 20806 22448 20812 22460
rect 20864 22488 20870 22500
rect 20901 22491 20959 22497
rect 20901 22488 20913 22491
rect 20864 22460 20913 22488
rect 20864 22448 20870 22460
rect 20901 22457 20913 22460
rect 20947 22457 20959 22491
rect 22097 22491 22155 22497
rect 22097 22488 22109 22491
rect 20901 22451 20959 22457
rect 21468 22460 22109 22488
rect 16356 22392 16620 22420
rect 17865 22423 17923 22429
rect 16356 22380 16362 22392
rect 17865 22389 17877 22423
rect 17911 22420 17923 22423
rect 18248 22420 18276 22448
rect 21468 22432 21496 22460
rect 22097 22457 22109 22460
rect 22143 22457 22155 22491
rect 22097 22451 22155 22457
rect 22189 22491 22247 22497
rect 22189 22457 22201 22491
rect 22235 22457 22247 22491
rect 22189 22451 22247 22457
rect 23845 22491 23903 22497
rect 23845 22457 23857 22491
rect 23891 22457 23903 22491
rect 23845 22451 23903 22457
rect 20070 22420 20076 22432
rect 17911 22392 18276 22420
rect 20031 22392 20076 22420
rect 17911 22389 17923 22392
rect 17865 22383 17923 22389
rect 20070 22380 20076 22392
rect 20128 22380 20134 22432
rect 21450 22420 21456 22432
rect 21411 22392 21456 22420
rect 21450 22380 21456 22392
rect 21508 22380 21514 22432
rect 21913 22423 21971 22429
rect 21913 22389 21925 22423
rect 21959 22420 21971 22423
rect 22204 22420 22232 22451
rect 22738 22420 22744 22432
rect 21959 22392 22744 22420
rect 21959 22389 21971 22392
rect 21913 22383 21971 22389
rect 22738 22380 22744 22392
rect 22796 22380 22802 22432
rect 23382 22420 23388 22432
rect 23343 22392 23388 22420
rect 23382 22380 23388 22392
rect 23440 22420 23446 22432
rect 23860 22420 23888 22451
rect 23440 22392 23888 22420
rect 23440 22380 23446 22392
rect 24026 22380 24032 22432
rect 24084 22420 24090 22432
rect 25363 22423 25421 22429
rect 25363 22420 25375 22423
rect 24084 22392 25375 22420
rect 24084 22380 24090 22392
rect 25363 22389 25375 22392
rect 25409 22389 25421 22423
rect 25363 22383 25421 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 9214 22216 9220 22228
rect 9175 22188 9220 22216
rect 9214 22176 9220 22188
rect 9272 22176 9278 22228
rect 13814 22176 13820 22228
rect 13872 22216 13878 22228
rect 17494 22216 17500 22228
rect 13872 22188 13917 22216
rect 17455 22188 17500 22216
rect 13872 22176 13878 22188
rect 17494 22176 17500 22188
rect 17552 22176 17558 22228
rect 18049 22219 18107 22225
rect 18049 22185 18061 22219
rect 18095 22216 18107 22219
rect 18230 22216 18236 22228
rect 18095 22188 18236 22216
rect 18095 22185 18107 22188
rect 18049 22179 18107 22185
rect 18230 22176 18236 22188
rect 18288 22216 18294 22228
rect 18325 22219 18383 22225
rect 18325 22216 18337 22219
rect 18288 22188 18337 22216
rect 18288 22176 18294 22188
rect 18325 22185 18337 22188
rect 18371 22185 18383 22219
rect 22462 22216 22468 22228
rect 22423 22188 22468 22216
rect 18325 22179 18383 22185
rect 22462 22176 22468 22188
rect 22520 22176 22526 22228
rect 23750 22216 23756 22228
rect 23711 22188 23756 22216
rect 23750 22176 23756 22188
rect 23808 22176 23814 22228
rect 24026 22216 24032 22228
rect 23987 22188 24032 22216
rect 24026 22176 24032 22188
rect 24084 22176 24090 22228
rect 9674 22108 9680 22160
rect 9732 22148 9738 22160
rect 10321 22151 10379 22157
rect 10321 22148 10333 22151
rect 9732 22120 10333 22148
rect 9732 22108 9738 22120
rect 10321 22117 10333 22120
rect 10367 22117 10379 22151
rect 16298 22148 16304 22160
rect 16259 22120 16304 22148
rect 10321 22111 10379 22117
rect 16298 22108 16304 22120
rect 16356 22108 16362 22160
rect 19426 22148 19432 22160
rect 19387 22120 19432 22148
rect 19426 22108 19432 22120
rect 19484 22108 19490 22160
rect 23382 22148 23388 22160
rect 23343 22120 23388 22148
rect 23382 22108 23388 22120
rect 23440 22108 23446 22160
rect 13170 22040 13176 22092
rect 13228 22080 13234 22092
rect 13449 22083 13507 22089
rect 13449 22080 13461 22083
rect 13228 22052 13461 22080
rect 13228 22040 13234 22052
rect 13449 22049 13461 22052
rect 13495 22049 13507 22083
rect 15930 22080 15936 22092
rect 15891 22052 15936 22080
rect 13449 22043 13507 22049
rect 15930 22040 15936 22052
rect 15988 22040 15994 22092
rect 22738 22080 22744 22092
rect 22699 22052 22744 22080
rect 22738 22040 22744 22052
rect 22796 22040 22802 22092
rect 24648 22083 24706 22089
rect 24648 22049 24660 22083
rect 24694 22080 24706 22083
rect 24762 22080 24768 22092
rect 24694 22052 24768 22080
rect 24694 22049 24706 22052
rect 24648 22043 24706 22049
rect 24762 22040 24768 22052
rect 24820 22040 24826 22092
rect 9950 21972 9956 22024
rect 10008 22012 10014 22024
rect 10229 22015 10287 22021
rect 10229 22012 10241 22015
rect 10008 21984 10241 22012
rect 10008 21972 10014 21984
rect 10229 21981 10241 21984
rect 10275 21981 10287 22015
rect 10229 21975 10287 21981
rect 17129 22015 17187 22021
rect 17129 21981 17141 22015
rect 17175 22012 17187 22015
rect 17678 22012 17684 22024
rect 17175 21984 17684 22012
rect 17175 21981 17187 21984
rect 17129 21975 17187 21981
rect 17678 21972 17684 21984
rect 17736 21972 17742 22024
rect 18874 21972 18880 22024
rect 18932 22012 18938 22024
rect 19337 22015 19395 22021
rect 19337 22012 19349 22015
rect 18932 21984 19349 22012
rect 18932 21972 18938 21984
rect 19337 21981 19349 21984
rect 19383 21981 19395 22015
rect 19337 21975 19395 21981
rect 19981 22015 20039 22021
rect 19981 21981 19993 22015
rect 20027 22012 20039 22015
rect 20530 22012 20536 22024
rect 20027 21984 20536 22012
rect 20027 21981 20039 21984
rect 19981 21975 20039 21981
rect 20530 21972 20536 21984
rect 20588 21972 20594 22024
rect 10778 21944 10784 21956
rect 10739 21916 10784 21944
rect 10778 21904 10784 21916
rect 10836 21904 10842 21956
rect 20346 21944 20352 21956
rect 20259 21916 20352 21944
rect 20346 21904 20352 21916
rect 20404 21944 20410 21956
rect 24719 21947 24777 21953
rect 24719 21944 24731 21947
rect 20404 21916 24731 21944
rect 20404 21904 20410 21916
rect 24719 21913 24731 21916
rect 24765 21913 24777 21947
rect 24719 21907 24777 21913
rect 11054 21836 11060 21888
rect 11112 21876 11118 21888
rect 11149 21879 11207 21885
rect 11149 21876 11161 21879
rect 11112 21848 11161 21876
rect 11112 21836 11118 21848
rect 11149 21845 11161 21848
rect 11195 21845 11207 21879
rect 21818 21876 21824 21888
rect 21779 21848 21824 21876
rect 11149 21839 11207 21845
rect 21818 21836 21824 21848
rect 21876 21836 21882 21888
rect 22186 21876 22192 21888
rect 22147 21848 22192 21876
rect 22186 21836 22192 21848
rect 22244 21836 22250 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 4798 21672 4804 21684
rect 4759 21644 4804 21672
rect 4798 21632 4804 21644
rect 4856 21632 4862 21684
rect 9033 21675 9091 21681
rect 9033 21641 9045 21675
rect 9079 21672 9091 21675
rect 9674 21672 9680 21684
rect 9079 21644 9680 21672
rect 9079 21641 9091 21644
rect 9033 21635 9091 21641
rect 9674 21632 9680 21644
rect 9732 21632 9738 21684
rect 11054 21672 11060 21684
rect 11015 21644 11060 21672
rect 11054 21632 11060 21644
rect 11112 21632 11118 21684
rect 14366 21672 14372 21684
rect 14327 21644 14372 21672
rect 14366 21632 14372 21644
rect 14424 21632 14430 21684
rect 15930 21672 15936 21684
rect 15891 21644 15936 21672
rect 15930 21632 15936 21644
rect 15988 21672 15994 21684
rect 16209 21675 16267 21681
rect 16209 21672 16221 21675
rect 15988 21644 16221 21672
rect 15988 21632 15994 21644
rect 16209 21641 16221 21644
rect 16255 21641 16267 21675
rect 16209 21635 16267 21641
rect 19337 21675 19395 21681
rect 19337 21641 19349 21675
rect 19383 21672 19395 21675
rect 19426 21672 19432 21684
rect 19383 21644 19432 21672
rect 19383 21641 19395 21644
rect 19337 21635 19395 21641
rect 19426 21632 19432 21644
rect 19484 21632 19490 21684
rect 19889 21675 19947 21681
rect 19889 21641 19901 21675
rect 19935 21672 19947 21675
rect 20070 21672 20076 21684
rect 19935 21644 20076 21672
rect 19935 21641 19947 21644
rect 19889 21635 19947 21641
rect 20070 21632 20076 21644
rect 20128 21632 20134 21684
rect 22186 21632 22192 21684
rect 22244 21672 22250 21684
rect 22649 21675 22707 21681
rect 22649 21672 22661 21675
rect 22244 21644 22661 21672
rect 22244 21632 22250 21644
rect 22649 21641 22661 21644
rect 22695 21641 22707 21675
rect 22649 21635 22707 21641
rect 22738 21632 22744 21684
rect 22796 21672 22802 21684
rect 22925 21675 22983 21681
rect 22925 21672 22937 21675
rect 22796 21644 22937 21672
rect 22796 21632 22802 21644
rect 22925 21641 22937 21644
rect 22971 21641 22983 21675
rect 24762 21672 24768 21684
rect 24723 21644 24768 21672
rect 22925 21635 22983 21641
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 13538 21564 13544 21616
rect 13596 21604 13602 21616
rect 18874 21604 18880 21616
rect 13596 21576 18880 21604
rect 13596 21564 13602 21576
rect 18874 21564 18880 21576
rect 18932 21564 18938 21616
rect 25774 21604 25780 21616
rect 25735 21576 25780 21604
rect 25774 21564 25780 21576
rect 25832 21564 25838 21616
rect 10045 21539 10103 21545
rect 10045 21505 10057 21539
rect 10091 21536 10103 21539
rect 10226 21536 10232 21548
rect 10091 21508 10232 21536
rect 10091 21505 10103 21508
rect 10045 21499 10103 21505
rect 10226 21496 10232 21508
rect 10284 21496 10290 21548
rect 15378 21536 15384 21548
rect 15339 21508 15384 21536
rect 15378 21496 15384 21508
rect 15436 21496 15442 21548
rect 17126 21536 17132 21548
rect 17087 21508 17132 21536
rect 17126 21496 17132 21508
rect 17184 21496 17190 21548
rect 20073 21539 20131 21545
rect 20073 21505 20085 21539
rect 20119 21536 20131 21539
rect 20346 21536 20352 21548
rect 20119 21508 20352 21536
rect 20119 21505 20131 21508
rect 20073 21499 20131 21505
rect 20346 21496 20352 21508
rect 20404 21496 20410 21548
rect 20530 21536 20536 21548
rect 20491 21508 20536 21536
rect 20530 21496 20536 21508
rect 20588 21496 20594 21548
rect 4408 21471 4466 21477
rect 4408 21437 4420 21471
rect 4454 21468 4466 21471
rect 4798 21468 4804 21480
rect 4454 21440 4804 21468
rect 4454 21437 4466 21440
rect 4408 21431 4466 21437
rect 4798 21428 4804 21440
rect 4856 21428 4862 21480
rect 8481 21471 8539 21477
rect 8481 21437 8493 21471
rect 8527 21468 8539 21471
rect 9030 21468 9036 21480
rect 8527 21440 9036 21468
rect 8527 21437 8539 21440
rect 8481 21431 8539 21437
rect 9030 21428 9036 21440
rect 9088 21468 9094 21480
rect 9214 21468 9220 21480
rect 9088 21440 9220 21468
rect 9088 21428 9094 21440
rect 9214 21428 9220 21440
rect 9272 21428 9278 21480
rect 10137 21471 10195 21477
rect 10137 21437 10149 21471
rect 10183 21468 10195 21471
rect 10686 21468 10692 21480
rect 10183 21440 10692 21468
rect 10183 21437 10195 21440
rect 10137 21431 10195 21437
rect 10686 21428 10692 21440
rect 10744 21468 10750 21480
rect 11333 21471 11391 21477
rect 11333 21468 11345 21471
rect 10744 21440 11345 21468
rect 10744 21428 10750 21440
rect 11333 21437 11345 21440
rect 11379 21437 11391 21471
rect 11333 21431 11391 21437
rect 13449 21471 13507 21477
rect 13449 21437 13461 21471
rect 13495 21468 13507 21471
rect 13906 21468 13912 21480
rect 13495 21440 13912 21468
rect 13495 21437 13507 21440
rect 13449 21431 13507 21437
rect 13906 21428 13912 21440
rect 13964 21428 13970 21480
rect 21729 21471 21787 21477
rect 21729 21437 21741 21471
rect 21775 21468 21787 21471
rect 21818 21468 21824 21480
rect 21775 21440 21824 21468
rect 21775 21437 21787 21440
rect 21729 21431 21787 21437
rect 21818 21428 21824 21440
rect 21876 21468 21882 21480
rect 22278 21468 22284 21480
rect 21876 21440 22284 21468
rect 21876 21428 21882 21440
rect 22278 21428 22284 21440
rect 22336 21428 22342 21480
rect 23474 21428 23480 21480
rect 23532 21468 23538 21480
rect 23753 21471 23811 21477
rect 23753 21468 23765 21471
rect 23532 21440 23765 21468
rect 23532 21428 23538 21440
rect 23753 21437 23765 21440
rect 23799 21437 23811 21471
rect 23753 21431 23811 21437
rect 25292 21471 25350 21477
rect 25292 21437 25304 21471
rect 25338 21468 25350 21471
rect 25792 21468 25820 21564
rect 25338 21440 25820 21468
rect 25338 21437 25350 21440
rect 25292 21431 25350 21437
rect 10226 21360 10232 21412
rect 10284 21400 10290 21412
rect 10499 21403 10557 21409
rect 10499 21400 10511 21403
rect 10284 21372 10511 21400
rect 10284 21360 10290 21372
rect 10499 21369 10511 21372
rect 10545 21400 10557 21403
rect 13354 21400 13360 21412
rect 10545 21372 13360 21400
rect 10545 21369 10557 21372
rect 10499 21363 10557 21369
rect 13354 21360 13360 21372
rect 13412 21400 13418 21412
rect 13811 21403 13869 21409
rect 13811 21400 13823 21403
rect 13412 21372 13823 21400
rect 13412 21360 13418 21372
rect 13811 21369 13823 21372
rect 13857 21400 13869 21403
rect 13998 21400 14004 21412
rect 13857 21372 14004 21400
rect 13857 21369 13869 21372
rect 13811 21363 13869 21369
rect 13998 21360 14004 21372
rect 14056 21360 14062 21412
rect 16482 21400 16488 21412
rect 16443 21372 16488 21400
rect 16482 21360 16488 21372
rect 16540 21360 16546 21412
rect 16577 21403 16635 21409
rect 16577 21369 16589 21403
rect 16623 21369 16635 21403
rect 17494 21400 17500 21412
rect 17407 21372 17500 21400
rect 16577 21363 16635 21369
rect 4479 21335 4537 21341
rect 4479 21301 4491 21335
rect 4525 21332 4537 21335
rect 9122 21332 9128 21344
rect 4525 21304 9128 21332
rect 4525 21301 4537 21304
rect 4479 21295 4537 21301
rect 9122 21292 9128 21304
rect 9180 21292 9186 21344
rect 12989 21335 13047 21341
rect 12989 21301 13001 21335
rect 13035 21332 13047 21335
rect 13170 21332 13176 21344
rect 13035 21304 13176 21332
rect 13035 21301 13047 21304
rect 12989 21295 13047 21301
rect 13170 21292 13176 21304
rect 13228 21292 13234 21344
rect 15930 21292 15936 21344
rect 15988 21332 15994 21344
rect 16592 21332 16620 21363
rect 17494 21360 17500 21372
rect 17552 21400 17558 21412
rect 19334 21400 19340 21412
rect 17552 21372 19340 21400
rect 17552 21360 17558 21372
rect 19334 21360 19340 21372
rect 19392 21360 19398 21412
rect 20162 21360 20168 21412
rect 20220 21400 20226 21412
rect 22050 21403 22108 21409
rect 20220 21372 20265 21400
rect 20220 21360 20226 21372
rect 22050 21369 22062 21403
rect 22096 21369 22108 21403
rect 24394 21400 24400 21412
rect 24355 21372 24400 21400
rect 22050 21363 22108 21369
rect 15988 21304 16620 21332
rect 15988 21292 15994 21304
rect 17678 21292 17684 21344
rect 17736 21332 17742 21344
rect 17773 21335 17831 21341
rect 17773 21332 17785 21335
rect 17736 21304 17785 21332
rect 17736 21292 17742 21304
rect 17773 21301 17785 21304
rect 17819 21301 17831 21335
rect 21634 21332 21640 21344
rect 21595 21304 21640 21332
rect 17773 21295 17831 21301
rect 21634 21292 21640 21304
rect 21692 21332 21698 21344
rect 22065 21332 22093 21363
rect 24394 21360 24400 21372
rect 24452 21360 24458 21412
rect 21692 21304 22093 21332
rect 21692 21292 21698 21304
rect 25038 21292 25044 21344
rect 25096 21332 25102 21344
rect 25363 21335 25421 21341
rect 25363 21332 25375 21335
rect 25096 21304 25375 21332
rect 25096 21292 25102 21304
rect 25363 21301 25375 21304
rect 25409 21301 25421 21335
rect 25363 21295 25421 21301
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 9214 21088 9220 21140
rect 9272 21128 9278 21140
rect 10597 21131 10655 21137
rect 10597 21128 10609 21131
rect 9272 21100 10609 21128
rect 9272 21088 9278 21100
rect 10597 21097 10609 21100
rect 10643 21097 10655 21131
rect 10597 21091 10655 21097
rect 13170 21088 13176 21140
rect 13228 21128 13234 21140
rect 13633 21131 13691 21137
rect 13633 21128 13645 21131
rect 13228 21100 13645 21128
rect 13228 21088 13234 21100
rect 13633 21097 13645 21100
rect 13679 21097 13691 21131
rect 13906 21128 13912 21140
rect 13867 21100 13912 21128
rect 13633 21091 13691 21097
rect 13906 21088 13912 21100
rect 13964 21088 13970 21140
rect 15654 21128 15660 21140
rect 15615 21100 15660 21128
rect 15654 21088 15660 21100
rect 15712 21088 15718 21140
rect 15930 21088 15936 21140
rect 15988 21128 15994 21140
rect 16209 21131 16267 21137
rect 16209 21128 16221 21131
rect 15988 21100 16221 21128
rect 15988 21088 15994 21100
rect 16209 21097 16221 21100
rect 16255 21097 16267 21131
rect 16482 21128 16488 21140
rect 16443 21100 16488 21128
rect 16209 21091 16267 21097
rect 16482 21088 16488 21100
rect 16540 21128 16546 21140
rect 16540 21100 17816 21128
rect 16540 21088 16546 21100
rect 10039 21063 10097 21069
rect 10039 21029 10051 21063
rect 10085 21060 10097 21063
rect 10134 21060 10140 21072
rect 10085 21032 10140 21060
rect 10085 21029 10097 21032
rect 10039 21023 10097 21029
rect 10134 21020 10140 21032
rect 10192 21020 10198 21072
rect 13075 21063 13133 21069
rect 13075 21029 13087 21063
rect 13121 21060 13133 21063
rect 13354 21060 13360 21072
rect 13121 21032 13360 21060
rect 13121 21029 13133 21032
rect 13075 21023 13133 21029
rect 13354 21020 13360 21032
rect 13412 21020 13418 21072
rect 17218 21060 17224 21072
rect 17179 21032 17224 21060
rect 17218 21020 17224 21032
rect 17276 21020 17282 21072
rect 17788 21069 17816 21100
rect 19426 21088 19432 21140
rect 19484 21128 19490 21140
rect 19705 21131 19763 21137
rect 19705 21128 19717 21131
rect 19484 21100 19717 21128
rect 19484 21088 19490 21100
rect 19705 21097 19717 21100
rect 19751 21097 19763 21131
rect 19705 21091 19763 21097
rect 22465 21131 22523 21137
rect 22465 21097 22477 21131
rect 22511 21128 22523 21131
rect 22738 21128 22744 21140
rect 22511 21100 22744 21128
rect 22511 21097 22523 21100
rect 22465 21091 22523 21097
rect 22738 21088 22744 21100
rect 22796 21088 22802 21140
rect 17773 21063 17831 21069
rect 17773 21029 17785 21063
rect 17819 21029 17831 21063
rect 17773 21023 17831 21029
rect 19147 21063 19205 21069
rect 19147 21029 19159 21063
rect 19193 21060 19205 21063
rect 19334 21060 19340 21072
rect 19193 21032 19340 21060
rect 19193 21029 19205 21032
rect 19147 21023 19205 21029
rect 19334 21020 19340 21032
rect 19392 21020 19398 21072
rect 21634 21020 21640 21072
rect 21692 21060 21698 21072
rect 21866 21063 21924 21069
rect 21866 21060 21878 21063
rect 21692 21032 21878 21060
rect 21692 21020 21698 21032
rect 21866 21029 21878 21032
rect 21912 21029 21924 21063
rect 21866 21023 21924 21029
rect 23474 21020 23480 21072
rect 23532 21060 23538 21072
rect 23532 21032 23577 21060
rect 23532 21020 23538 21032
rect 24394 21020 24400 21072
rect 24452 21060 24458 21072
rect 24946 21060 24952 21072
rect 24452 21032 24952 21060
rect 24452 21020 24458 21032
rect 24946 21020 24952 21032
rect 25004 21060 25010 21072
rect 25041 21063 25099 21069
rect 25041 21060 25053 21063
rect 25004 21032 25053 21060
rect 25004 21020 25010 21032
rect 25041 21029 25053 21032
rect 25087 21029 25099 21063
rect 25041 21023 25099 21029
rect 9674 20924 9680 20936
rect 9635 20896 9680 20924
rect 9674 20884 9680 20896
rect 9732 20884 9738 20936
rect 12710 20924 12716 20936
rect 12671 20896 12716 20924
rect 12710 20884 12716 20896
rect 12768 20884 12774 20936
rect 15289 20927 15347 20933
rect 15289 20893 15301 20927
rect 15335 20924 15347 20927
rect 15378 20924 15384 20936
rect 15335 20896 15384 20924
rect 15335 20893 15347 20896
rect 15289 20887 15347 20893
rect 15378 20884 15384 20896
rect 15436 20884 15442 20936
rect 17126 20924 17132 20936
rect 17087 20896 17132 20924
rect 17126 20884 17132 20896
rect 17184 20884 17190 20936
rect 18690 20884 18696 20936
rect 18748 20924 18754 20936
rect 18785 20927 18843 20933
rect 18785 20924 18797 20927
rect 18748 20896 18797 20924
rect 18748 20884 18754 20896
rect 18785 20893 18797 20896
rect 18831 20893 18843 20927
rect 18785 20887 18843 20893
rect 21545 20927 21603 20933
rect 21545 20893 21557 20927
rect 21591 20924 21603 20927
rect 21910 20924 21916 20936
rect 21591 20896 21916 20924
rect 21591 20893 21603 20896
rect 21545 20887 21603 20893
rect 21910 20884 21916 20896
rect 21968 20884 21974 20936
rect 23382 20924 23388 20936
rect 23343 20896 23388 20924
rect 23382 20884 23388 20896
rect 23440 20884 23446 20936
rect 24949 20927 25007 20933
rect 24949 20893 24961 20927
rect 24995 20924 25007 20927
rect 25038 20924 25044 20936
rect 24995 20896 25044 20924
rect 24995 20893 25007 20896
rect 24949 20887 25007 20893
rect 25038 20884 25044 20896
rect 25096 20884 25102 20936
rect 25225 20927 25283 20933
rect 25225 20893 25237 20927
rect 25271 20893 25283 20927
rect 25225 20887 25283 20893
rect 23937 20859 23995 20865
rect 23937 20825 23949 20859
rect 23983 20856 23995 20859
rect 24854 20856 24860 20868
rect 23983 20828 24860 20856
rect 23983 20825 23995 20828
rect 23937 20819 23995 20825
rect 24854 20816 24860 20828
rect 24912 20856 24918 20868
rect 25240 20856 25268 20887
rect 24912 20828 25268 20856
rect 24912 20816 24918 20828
rect 9950 20748 9956 20800
rect 10008 20788 10014 20800
rect 10873 20791 10931 20797
rect 10873 20788 10885 20791
rect 10008 20760 10885 20788
rect 10008 20748 10014 20760
rect 10873 20757 10885 20760
rect 10919 20757 10931 20791
rect 19978 20788 19984 20800
rect 19939 20760 19984 20788
rect 10873 20751 10931 20757
rect 19978 20748 19984 20760
rect 20036 20748 20042 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 9769 20587 9827 20593
rect 9769 20553 9781 20587
rect 9815 20584 9827 20587
rect 10134 20584 10140 20596
rect 9815 20556 10140 20584
rect 9815 20553 9827 20556
rect 9769 20547 9827 20553
rect 10134 20544 10140 20556
rect 10192 20544 10198 20596
rect 15197 20587 15255 20593
rect 15197 20553 15209 20587
rect 15243 20584 15255 20587
rect 16298 20584 16304 20596
rect 15243 20556 16304 20584
rect 15243 20553 15255 20556
rect 15197 20547 15255 20553
rect 16298 20544 16304 20556
rect 16356 20584 16362 20596
rect 17218 20584 17224 20596
rect 16356 20556 17224 20584
rect 16356 20544 16362 20556
rect 17218 20544 17224 20556
rect 17276 20544 17282 20596
rect 22738 20544 22744 20596
rect 22796 20584 22802 20596
rect 23109 20587 23167 20593
rect 23109 20584 23121 20587
rect 22796 20556 23121 20584
rect 22796 20544 22802 20556
rect 23109 20553 23121 20556
rect 23155 20584 23167 20587
rect 23474 20584 23480 20596
rect 23155 20556 23480 20584
rect 23155 20553 23167 20556
rect 23109 20547 23167 20553
rect 23474 20544 23480 20556
rect 23532 20544 23538 20596
rect 24946 20584 24952 20596
rect 24907 20556 24952 20584
rect 24946 20544 24952 20556
rect 25004 20544 25010 20596
rect 11793 20519 11851 20525
rect 11793 20516 11805 20519
rect 9600 20488 11805 20516
rect 1486 20340 1492 20392
rect 1544 20380 1550 20392
rect 7374 20380 7380 20392
rect 1544 20352 7380 20380
rect 1544 20340 1550 20352
rect 7374 20340 7380 20352
rect 7432 20340 7438 20392
rect 9401 20383 9459 20389
rect 9401 20349 9413 20383
rect 9447 20380 9459 20383
rect 9600 20380 9628 20488
rect 11793 20485 11805 20488
rect 11839 20485 11851 20519
rect 11793 20479 11851 20485
rect 12253 20519 12311 20525
rect 12253 20485 12265 20519
rect 12299 20516 12311 20519
rect 13998 20516 14004 20528
rect 12299 20488 14004 20516
rect 12299 20485 12311 20488
rect 12253 20479 12311 20485
rect 9674 20408 9680 20460
rect 9732 20448 9738 20460
rect 10873 20451 10931 20457
rect 10873 20448 10885 20451
rect 9732 20420 10885 20448
rect 9732 20408 9738 20420
rect 10873 20417 10885 20420
rect 10919 20417 10931 20451
rect 10873 20411 10931 20417
rect 9858 20380 9864 20392
rect 9447 20352 9864 20380
rect 9447 20349 9459 20352
rect 9401 20343 9459 20349
rect 9858 20340 9864 20352
rect 9916 20340 9922 20392
rect 10134 20340 10140 20392
rect 10192 20380 10198 20392
rect 10321 20383 10379 20389
rect 10321 20380 10333 20383
rect 10192 20352 10333 20380
rect 10192 20340 10198 20352
rect 10321 20349 10333 20352
rect 10367 20349 10379 20383
rect 10321 20343 10379 20349
rect 10597 20383 10655 20389
rect 10597 20349 10609 20383
rect 10643 20380 10655 20383
rect 10686 20380 10692 20392
rect 10643 20352 10692 20380
rect 10643 20349 10655 20352
rect 10597 20343 10655 20349
rect 10686 20340 10692 20352
rect 10744 20340 10750 20392
rect 11808 20380 11836 20479
rect 13998 20476 14004 20488
rect 14056 20516 14062 20528
rect 14185 20519 14243 20525
rect 14185 20516 14197 20519
rect 14056 20488 14197 20516
rect 14056 20476 14062 20488
rect 14185 20485 14197 20488
rect 14231 20516 14243 20519
rect 15565 20519 15623 20525
rect 15565 20516 15577 20519
rect 14231 20488 15577 20516
rect 14231 20485 14243 20488
rect 14185 20479 14243 20485
rect 13449 20451 13507 20457
rect 13449 20417 13461 20451
rect 13495 20448 13507 20451
rect 13906 20448 13912 20460
rect 13495 20420 13912 20448
rect 13495 20417 13507 20420
rect 13449 20411 13507 20417
rect 13906 20408 13912 20420
rect 13964 20408 13970 20460
rect 12713 20383 12771 20389
rect 12713 20380 12725 20383
rect 11808 20352 12725 20380
rect 12713 20349 12725 20352
rect 12759 20380 12771 20383
rect 13078 20380 13084 20392
rect 12759 20352 13084 20380
rect 12759 20349 12771 20352
rect 12713 20343 12771 20349
rect 13078 20340 13084 20352
rect 13136 20340 13142 20392
rect 13265 20383 13323 20389
rect 13265 20349 13277 20383
rect 13311 20380 13323 20383
rect 13814 20380 13820 20392
rect 13311 20352 13820 20380
rect 13311 20349 13323 20352
rect 13265 20343 13323 20349
rect 13814 20340 13820 20352
rect 13872 20380 13878 20392
rect 14274 20380 14280 20392
rect 13872 20352 13965 20380
rect 14235 20352 14280 20380
rect 13872 20340 13878 20352
rect 14274 20340 14280 20352
rect 14332 20340 14338 20392
rect 9033 20315 9091 20321
rect 9033 20281 9045 20315
rect 9079 20312 9091 20315
rect 10152 20312 10180 20340
rect 14654 20321 14682 20488
rect 15565 20485 15577 20488
rect 15611 20516 15623 20519
rect 15654 20516 15660 20528
rect 15611 20488 15660 20516
rect 15611 20485 15623 20488
rect 15565 20479 15623 20485
rect 15654 20476 15660 20488
rect 15712 20516 15718 20528
rect 15712 20488 16712 20516
rect 15712 20476 15718 20488
rect 16482 20408 16488 20460
rect 16540 20448 16546 20460
rect 16577 20451 16635 20457
rect 16577 20448 16589 20451
rect 16540 20420 16589 20448
rect 16540 20408 16546 20420
rect 16577 20417 16589 20420
rect 16623 20417 16635 20451
rect 16684 20448 16712 20488
rect 17126 20476 17132 20528
rect 17184 20516 17190 20528
rect 17589 20519 17647 20525
rect 17589 20516 17601 20519
rect 17184 20488 17601 20516
rect 17184 20476 17190 20488
rect 17589 20485 17601 20488
rect 17635 20485 17647 20519
rect 19334 20516 19340 20528
rect 19247 20488 19340 20516
rect 17589 20479 17647 20485
rect 19334 20476 19340 20488
rect 19392 20516 19398 20528
rect 21634 20516 21640 20528
rect 19392 20488 21640 20516
rect 19392 20476 19398 20488
rect 21634 20476 21640 20488
rect 21692 20476 21698 20528
rect 25774 20516 25780 20528
rect 25735 20488 25780 20516
rect 25774 20476 25780 20488
rect 25832 20476 25838 20528
rect 18785 20451 18843 20457
rect 16684 20420 17172 20448
rect 16577 20411 16635 20417
rect 17144 20380 17172 20420
rect 18785 20417 18797 20451
rect 18831 20448 18843 20451
rect 19889 20451 19947 20457
rect 19889 20448 19901 20451
rect 18831 20420 19901 20448
rect 18831 20417 18843 20420
rect 18785 20411 18843 20417
rect 19889 20417 19901 20420
rect 19935 20448 19947 20451
rect 19978 20448 19984 20460
rect 19935 20420 19984 20448
rect 19935 20417 19947 20420
rect 19889 20411 19947 20417
rect 19978 20408 19984 20420
rect 20036 20408 20042 20460
rect 17586 20380 17592 20392
rect 17144 20352 17592 20380
rect 17586 20340 17592 20352
rect 17644 20340 17650 20392
rect 22592 20383 22650 20389
rect 22592 20380 22604 20383
rect 22388 20352 22604 20380
rect 9079 20284 10180 20312
rect 14639 20315 14697 20321
rect 9079 20281 9091 20284
rect 9033 20275 9091 20281
rect 14639 20281 14651 20315
rect 14685 20281 14697 20315
rect 14639 20275 14697 20281
rect 16022 20272 16028 20324
rect 16080 20312 16086 20324
rect 16301 20315 16359 20321
rect 16301 20312 16313 20315
rect 16080 20284 16313 20312
rect 16080 20272 16086 20284
rect 16301 20281 16313 20284
rect 16347 20281 16359 20315
rect 16301 20275 16359 20281
rect 16393 20315 16451 20321
rect 16393 20281 16405 20315
rect 16439 20281 16451 20315
rect 16393 20275 16451 20281
rect 19981 20315 20039 20321
rect 19981 20281 19993 20315
rect 20027 20281 20039 20315
rect 20530 20312 20536 20324
rect 20491 20284 20536 20312
rect 19981 20275 20039 20281
rect 16114 20244 16120 20256
rect 16075 20216 16120 20244
rect 16114 20204 16120 20216
rect 16172 20244 16178 20256
rect 16408 20244 16436 20275
rect 18690 20244 18696 20256
rect 16172 20216 16436 20244
rect 18651 20216 18696 20244
rect 16172 20204 16178 20216
rect 18690 20204 18696 20216
rect 18748 20204 18754 20256
rect 19518 20204 19524 20256
rect 19576 20244 19582 20256
rect 19613 20247 19671 20253
rect 19613 20244 19625 20247
rect 19576 20216 19625 20244
rect 19576 20204 19582 20216
rect 19613 20213 19625 20216
rect 19659 20244 19671 20247
rect 19996 20244 20024 20275
rect 20530 20272 20536 20284
rect 20588 20312 20594 20324
rect 22388 20321 22416 20352
rect 22592 20349 22604 20352
rect 22638 20349 22650 20383
rect 22592 20343 22650 20349
rect 23382 20340 23388 20392
rect 23440 20380 23446 20392
rect 23661 20383 23719 20389
rect 23661 20380 23673 20383
rect 23440 20352 23673 20380
rect 23440 20340 23446 20352
rect 23661 20349 23673 20352
rect 23707 20349 23719 20383
rect 23661 20343 23719 20349
rect 23753 20383 23811 20389
rect 23753 20349 23765 20383
rect 23799 20349 23811 20383
rect 23753 20343 23811 20349
rect 25292 20383 25350 20389
rect 25292 20349 25304 20383
rect 25338 20380 25350 20383
rect 25792 20380 25820 20476
rect 25338 20352 25820 20380
rect 25338 20349 25350 20352
rect 25292 20343 25350 20349
rect 22373 20315 22431 20321
rect 22373 20312 22385 20315
rect 20588 20284 22385 20312
rect 20588 20272 20594 20284
rect 22373 20281 22385 20284
rect 22419 20281 22431 20315
rect 22373 20275 22431 20281
rect 23477 20315 23535 20321
rect 23477 20281 23489 20315
rect 23523 20312 23535 20315
rect 23768 20312 23796 20343
rect 23934 20312 23940 20324
rect 23523 20284 23940 20312
rect 23523 20281 23535 20284
rect 23477 20275 23535 20281
rect 23934 20272 23940 20284
rect 23992 20272 23998 20324
rect 21634 20244 21640 20256
rect 19659 20216 20024 20244
rect 21595 20216 21640 20244
rect 19659 20213 19671 20216
rect 19613 20207 19671 20213
rect 21634 20204 21640 20216
rect 21692 20204 21698 20256
rect 21910 20244 21916 20256
rect 21871 20216 21916 20244
rect 21910 20204 21916 20216
rect 21968 20204 21974 20256
rect 22695 20247 22753 20253
rect 22695 20213 22707 20247
rect 22741 20244 22753 20247
rect 23106 20244 23112 20256
rect 22741 20216 23112 20244
rect 22741 20213 22753 20216
rect 22695 20207 22753 20213
rect 23106 20204 23112 20216
rect 23164 20204 23170 20256
rect 23750 20204 23756 20256
rect 23808 20244 23814 20256
rect 25363 20247 25421 20253
rect 25363 20244 25375 20247
rect 23808 20216 25375 20244
rect 23808 20204 23814 20216
rect 25363 20213 25375 20216
rect 25409 20213 25421 20247
rect 25363 20207 25421 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 9674 20000 9680 20052
rect 9732 20040 9738 20052
rect 9769 20043 9827 20049
rect 9769 20040 9781 20043
rect 9732 20012 9781 20040
rect 9732 20000 9738 20012
rect 9769 20009 9781 20012
rect 9815 20009 9827 20043
rect 9769 20003 9827 20009
rect 12710 20000 12716 20052
rect 12768 20040 12774 20052
rect 12805 20043 12863 20049
rect 12805 20040 12817 20043
rect 12768 20012 12817 20040
rect 12768 20000 12774 20012
rect 12805 20009 12817 20012
rect 12851 20040 12863 20043
rect 13541 20043 13599 20049
rect 13541 20040 13553 20043
rect 12851 20012 13553 20040
rect 12851 20009 12863 20012
rect 12805 20003 12863 20009
rect 13541 20009 13553 20012
rect 13587 20009 13599 20043
rect 13541 20003 13599 20009
rect 14274 20000 14280 20052
rect 14332 20040 14338 20052
rect 14369 20043 14427 20049
rect 14369 20040 14381 20043
rect 14332 20012 14381 20040
rect 14332 20000 14338 20012
rect 14369 20009 14381 20012
rect 14415 20040 14427 20043
rect 15381 20043 15439 20049
rect 15381 20040 15393 20043
rect 14415 20012 15393 20040
rect 14415 20009 14427 20012
rect 14369 20003 14427 20009
rect 15381 20009 15393 20012
rect 15427 20009 15439 20043
rect 17586 20040 17592 20052
rect 17547 20012 17592 20040
rect 15381 20003 15439 20009
rect 17586 20000 17592 20012
rect 17644 20000 17650 20052
rect 18138 20040 18144 20052
rect 18099 20012 18144 20040
rect 18138 20000 18144 20012
rect 18196 20000 18202 20052
rect 19518 20040 19524 20052
rect 19479 20012 19524 20040
rect 19518 20000 19524 20012
rect 19576 20000 19582 20052
rect 22738 20040 22744 20052
rect 22699 20012 22744 20040
rect 22738 20000 22744 20012
rect 22796 20000 22802 20052
rect 23290 20040 23296 20052
rect 23251 20012 23296 20040
rect 23290 20000 23296 20012
rect 23348 20000 23354 20052
rect 24949 20043 25007 20049
rect 24949 20009 24961 20043
rect 24995 20040 25007 20043
rect 25038 20040 25044 20052
rect 24995 20012 25044 20040
rect 24995 20009 25007 20012
rect 24949 20003 25007 20009
rect 25038 20000 25044 20012
rect 25096 20000 25102 20052
rect 12820 19944 15332 19972
rect 9766 19904 9772 19916
rect 9727 19876 9772 19904
rect 9766 19864 9772 19876
rect 9824 19864 9830 19916
rect 10134 19904 10140 19916
rect 10095 19876 10140 19904
rect 10134 19864 10140 19876
rect 10192 19864 10198 19916
rect 12710 19864 12716 19916
rect 12768 19904 12774 19916
rect 12820 19913 12848 19944
rect 15304 19916 15332 19944
rect 21634 19932 21640 19984
rect 21692 19972 21698 19984
rect 22183 19975 22241 19981
rect 22183 19972 22195 19975
rect 21692 19944 22195 19972
rect 21692 19932 21698 19944
rect 22183 19941 22195 19944
rect 22229 19972 22241 19975
rect 22370 19972 22376 19984
rect 22229 19944 22376 19972
rect 22229 19941 22241 19944
rect 22183 19935 22241 19941
rect 22370 19932 22376 19944
rect 22428 19932 22434 19984
rect 23934 19972 23940 19984
rect 23895 19944 23940 19972
rect 23934 19932 23940 19944
rect 23992 19932 23998 19984
rect 24026 19932 24032 19984
rect 24084 19972 24090 19984
rect 25317 19975 25375 19981
rect 25317 19972 25329 19975
rect 24084 19944 25329 19972
rect 24084 19932 24090 19944
rect 25317 19941 25329 19944
rect 25363 19941 25375 19975
rect 25317 19935 25375 19941
rect 12805 19907 12863 19913
rect 12805 19904 12817 19907
rect 12768 19876 12817 19904
rect 12768 19864 12774 19876
rect 12805 19873 12817 19876
rect 12851 19873 12863 19907
rect 12805 19867 12863 19873
rect 13081 19907 13139 19913
rect 13081 19873 13093 19907
rect 13127 19904 13139 19907
rect 13814 19904 13820 19916
rect 13127 19876 13820 19904
rect 13127 19873 13139 19876
rect 13081 19867 13139 19873
rect 13814 19864 13820 19876
rect 13872 19864 13878 19916
rect 15286 19904 15292 19916
rect 15247 19876 15292 19904
rect 15286 19864 15292 19876
rect 15344 19864 15350 19916
rect 15470 19864 15476 19916
rect 15528 19904 15534 19916
rect 15749 19907 15807 19913
rect 15749 19904 15761 19907
rect 15528 19876 15761 19904
rect 15528 19864 15534 19876
rect 15749 19873 15761 19876
rect 15795 19873 15807 19907
rect 19334 19904 19340 19916
rect 19295 19876 19340 19904
rect 15749 19867 15807 19873
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 11241 19839 11299 19845
rect 11241 19805 11253 19839
rect 11287 19836 11299 19839
rect 11330 19836 11336 19848
rect 11287 19808 11336 19836
rect 11287 19805 11299 19808
rect 11241 19799 11299 19805
rect 11330 19796 11336 19808
rect 11388 19796 11394 19848
rect 14550 19796 14556 19848
rect 14608 19836 14614 19848
rect 15105 19839 15163 19845
rect 15105 19836 15117 19839
rect 14608 19808 15117 19836
rect 14608 19796 14614 19808
rect 15105 19805 15117 19808
rect 15151 19836 15163 19839
rect 15378 19836 15384 19848
rect 15151 19808 15384 19836
rect 15151 19805 15163 19808
rect 15105 19799 15163 19805
rect 15378 19796 15384 19808
rect 15436 19796 15442 19848
rect 16758 19796 16764 19848
rect 16816 19836 16822 19848
rect 17221 19839 17279 19845
rect 17221 19836 17233 19839
rect 16816 19808 17233 19836
rect 16816 19796 16822 19808
rect 17221 19805 17233 19808
rect 17267 19805 17279 19839
rect 17221 19799 17279 19805
rect 21542 19796 21548 19848
rect 21600 19836 21606 19848
rect 21821 19839 21879 19845
rect 21821 19836 21833 19839
rect 21600 19808 21833 19836
rect 21600 19796 21606 19808
rect 21821 19805 21833 19808
rect 21867 19805 21879 19839
rect 23842 19836 23848 19848
rect 23803 19808 23848 19836
rect 21821 19799 21879 19805
rect 23842 19796 23848 19808
rect 23900 19796 23906 19848
rect 24210 19836 24216 19848
rect 24171 19808 24216 19836
rect 24210 19796 24216 19808
rect 24268 19796 24274 19848
rect 16022 19660 16028 19712
rect 16080 19700 16086 19712
rect 16301 19703 16359 19709
rect 16301 19700 16313 19703
rect 16080 19672 16313 19700
rect 16080 19660 16086 19672
rect 16301 19669 16313 19672
rect 16347 19669 16359 19703
rect 16301 19663 16359 19669
rect 20806 19660 20812 19712
rect 20864 19700 20870 19712
rect 21361 19703 21419 19709
rect 21361 19700 21373 19703
rect 20864 19672 21373 19700
rect 20864 19660 20870 19672
rect 21361 19669 21373 19672
rect 21407 19669 21419 19703
rect 21361 19663 21419 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 9030 19456 9036 19508
rect 9088 19496 9094 19508
rect 9766 19496 9772 19508
rect 9088 19468 9772 19496
rect 9088 19456 9094 19468
rect 9766 19456 9772 19468
rect 9824 19496 9830 19508
rect 12342 19496 12348 19508
rect 9824 19468 12348 19496
rect 9824 19456 9830 19468
rect 12342 19456 12348 19468
rect 12400 19496 12406 19508
rect 12710 19496 12716 19508
rect 12400 19468 12716 19496
rect 12400 19456 12406 19468
rect 12710 19456 12716 19468
rect 12768 19456 12774 19508
rect 15286 19496 15292 19508
rect 15247 19468 15292 19496
rect 15286 19456 15292 19468
rect 15344 19456 15350 19508
rect 16114 19496 16120 19508
rect 16075 19468 16120 19496
rect 16114 19456 16120 19468
rect 16172 19456 16178 19508
rect 18969 19499 19027 19505
rect 18969 19465 18981 19499
rect 19015 19496 19027 19499
rect 19334 19496 19340 19508
rect 19015 19468 19340 19496
rect 19015 19465 19027 19468
rect 18969 19459 19027 19465
rect 19334 19456 19340 19468
rect 19392 19496 19398 19508
rect 19613 19499 19671 19505
rect 19613 19496 19625 19499
rect 19392 19468 19625 19496
rect 19392 19456 19398 19468
rect 19613 19465 19625 19468
rect 19659 19496 19671 19499
rect 19978 19496 19984 19508
rect 19659 19468 19984 19496
rect 19659 19465 19671 19468
rect 19613 19459 19671 19465
rect 19978 19456 19984 19468
rect 20036 19456 20042 19508
rect 23014 19456 23020 19508
rect 23072 19496 23078 19508
rect 23109 19499 23167 19505
rect 23109 19496 23121 19499
rect 23072 19468 23121 19496
rect 23072 19456 23078 19468
rect 23109 19465 23121 19468
rect 23155 19496 23167 19499
rect 23934 19496 23940 19508
rect 23155 19468 23940 19496
rect 23155 19465 23167 19468
rect 23109 19459 23167 19465
rect 23934 19456 23940 19468
rect 23992 19456 23998 19508
rect 20438 19428 20444 19440
rect 19904 19400 20444 19428
rect 7374 19320 7380 19372
rect 7432 19360 7438 19372
rect 8665 19363 8723 19369
rect 8665 19360 8677 19363
rect 7432 19332 8677 19360
rect 7432 19320 7438 19332
rect 8287 19301 8315 19332
rect 8665 19329 8677 19332
rect 8711 19329 8723 19363
rect 8665 19323 8723 19329
rect 13078 19320 13084 19372
rect 13136 19360 13142 19372
rect 13633 19363 13691 19369
rect 13633 19360 13645 19363
rect 13136 19332 13645 19360
rect 13136 19320 13142 19332
rect 13633 19329 13645 19332
rect 13679 19329 13691 19363
rect 14550 19360 14556 19372
rect 14511 19332 14556 19360
rect 13633 19323 13691 19329
rect 8272 19295 8330 19301
rect 8272 19261 8284 19295
rect 8318 19261 8330 19295
rect 8272 19255 8330 19261
rect 10689 19295 10747 19301
rect 10689 19261 10701 19295
rect 10735 19292 10747 19295
rect 10870 19292 10876 19304
rect 10735 19264 10876 19292
rect 10735 19261 10747 19264
rect 10689 19255 10747 19261
rect 10870 19252 10876 19264
rect 10928 19252 10934 19304
rect 13648 19292 13676 19323
rect 14550 19320 14556 19332
rect 14608 19320 14614 19372
rect 19904 19369 19932 19400
rect 20438 19388 20444 19400
rect 20496 19388 20502 19440
rect 23477 19431 23535 19437
rect 23477 19397 23489 19431
rect 23523 19428 23535 19431
rect 24026 19428 24032 19440
rect 23523 19400 24032 19428
rect 23523 19397 23535 19400
rect 23477 19391 23535 19397
rect 24026 19388 24032 19400
rect 24084 19388 24090 19440
rect 26050 19428 26056 19440
rect 26011 19400 26056 19428
rect 26050 19388 26056 19400
rect 26108 19388 26114 19440
rect 19889 19363 19947 19369
rect 19889 19329 19901 19363
rect 19935 19329 19947 19363
rect 20530 19360 20536 19372
rect 20491 19332 20536 19360
rect 19889 19323 19947 19329
rect 20530 19320 20536 19332
rect 20588 19320 20594 19372
rect 20990 19320 20996 19372
rect 21048 19360 21054 19372
rect 22002 19360 22008 19372
rect 21048 19332 22008 19360
rect 21048 19320 21054 19332
rect 22002 19320 22008 19332
rect 22060 19360 22066 19372
rect 24210 19360 24216 19372
rect 22060 19332 24216 19360
rect 22060 19320 22066 19332
rect 24210 19320 24216 19332
rect 24268 19360 24274 19372
rect 24305 19363 24363 19369
rect 24305 19360 24317 19363
rect 24268 19332 24317 19360
rect 24268 19320 24274 19332
rect 24305 19329 24317 19332
rect 24351 19329 24363 19363
rect 24305 19323 24363 19329
rect 13817 19295 13875 19301
rect 13817 19292 13829 19295
rect 13648 19264 13829 19292
rect 13817 19261 13829 19264
rect 13863 19261 13875 19295
rect 13817 19255 13875 19261
rect 13906 19252 13912 19304
rect 13964 19292 13970 19304
rect 14369 19295 14427 19301
rect 14369 19292 14381 19295
rect 13964 19264 14381 19292
rect 13964 19252 13970 19264
rect 14369 19261 14381 19264
rect 14415 19292 14427 19295
rect 16298 19292 16304 19304
rect 14415 19264 15056 19292
rect 16259 19264 16304 19292
rect 14415 19261 14427 19264
rect 14369 19255 14427 19261
rect 13188 19196 13860 19224
rect 13188 19168 13216 19196
rect 13832 19168 13860 19196
rect 8343 19159 8401 19165
rect 8343 19125 8355 19159
rect 8389 19156 8401 19159
rect 8846 19156 8852 19168
rect 8389 19128 8852 19156
rect 8389 19125 8401 19128
rect 8343 19119 8401 19125
rect 8846 19116 8852 19128
rect 8904 19116 8910 19168
rect 10134 19156 10140 19168
rect 10047 19128 10140 19156
rect 10134 19116 10140 19128
rect 10192 19156 10198 19168
rect 11054 19156 11060 19168
rect 10192 19128 11060 19156
rect 10192 19116 10198 19128
rect 11054 19116 11060 19128
rect 11112 19116 11118 19168
rect 11238 19156 11244 19168
rect 11199 19128 11244 19156
rect 11238 19116 11244 19128
rect 11296 19116 11302 19168
rect 13081 19159 13139 19165
rect 13081 19125 13093 19159
rect 13127 19156 13139 19159
rect 13170 19156 13176 19168
rect 13127 19128 13176 19156
rect 13127 19125 13139 19128
rect 13081 19119 13139 19125
rect 13170 19116 13176 19128
rect 13228 19116 13234 19168
rect 13814 19116 13820 19168
rect 13872 19116 13878 19168
rect 15028 19165 15056 19264
rect 16298 19252 16304 19264
rect 16356 19252 16362 19304
rect 17954 19252 17960 19304
rect 18012 19292 18018 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 18012 19264 18061 19292
rect 18012 19252 18018 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 21266 19292 21272 19304
rect 21179 19264 21272 19292
rect 18049 19255 18107 19261
rect 21266 19252 21272 19264
rect 21324 19292 21330 19304
rect 21361 19295 21419 19301
rect 21361 19292 21373 19295
rect 21324 19264 21373 19292
rect 21324 19252 21330 19264
rect 21361 19261 21373 19264
rect 21407 19261 21419 19295
rect 21361 19255 21419 19261
rect 21821 19295 21879 19301
rect 21821 19261 21833 19295
rect 21867 19261 21879 19295
rect 21821 19255 21879 19261
rect 25568 19295 25626 19301
rect 25568 19261 25580 19295
rect 25614 19292 25626 19295
rect 26068 19292 26096 19388
rect 25614 19264 26096 19292
rect 25614 19261 25626 19264
rect 25568 19255 25626 19261
rect 18370 19227 18428 19233
rect 18370 19224 18382 19227
rect 18156 19196 18382 19224
rect 18156 19168 18184 19196
rect 18370 19193 18382 19196
rect 18416 19193 18428 19227
rect 18370 19187 18428 19193
rect 19978 19184 19984 19236
rect 20036 19224 20042 19236
rect 20036 19196 20081 19224
rect 20036 19184 20042 19196
rect 20806 19184 20812 19236
rect 20864 19224 20870 19236
rect 21836 19224 21864 19255
rect 22094 19224 22100 19236
rect 20864 19196 21864 19224
rect 22055 19196 22100 19224
rect 20864 19184 20870 19196
rect 22094 19184 22100 19196
rect 22152 19184 22158 19236
rect 24026 19224 24032 19236
rect 23987 19196 24032 19224
rect 24026 19184 24032 19196
rect 24084 19184 24090 19236
rect 24121 19227 24179 19233
rect 24121 19193 24133 19227
rect 24167 19193 24179 19227
rect 24121 19187 24179 19193
rect 15013 19159 15071 19165
rect 15013 19125 15025 19159
rect 15059 19156 15071 19159
rect 15470 19156 15476 19168
rect 15059 19128 15476 19156
rect 15059 19125 15071 19128
rect 15013 19119 15071 19125
rect 15470 19116 15476 19128
rect 15528 19116 15534 19168
rect 16758 19116 16764 19168
rect 16816 19156 16822 19168
rect 16853 19159 16911 19165
rect 16853 19156 16865 19159
rect 16816 19128 16865 19156
rect 16816 19116 16822 19128
rect 16853 19125 16865 19128
rect 16899 19125 16911 19159
rect 16853 19119 16911 19125
rect 17313 19159 17371 19165
rect 17313 19125 17325 19159
rect 17359 19156 17371 19159
rect 17586 19156 17592 19168
rect 17359 19128 17592 19156
rect 17359 19125 17371 19128
rect 17313 19119 17371 19125
rect 17586 19116 17592 19128
rect 17644 19156 17650 19168
rect 17865 19159 17923 19165
rect 17865 19156 17877 19159
rect 17644 19128 17877 19156
rect 17644 19116 17650 19128
rect 17865 19125 17877 19128
rect 17911 19156 17923 19159
rect 18138 19156 18144 19168
rect 17911 19128 18144 19156
rect 17911 19125 17923 19128
rect 17865 19119 17923 19125
rect 18138 19116 18144 19128
rect 18196 19116 18202 19168
rect 22370 19156 22376 19168
rect 22331 19128 22376 19156
rect 22370 19116 22376 19128
rect 22428 19116 22434 19168
rect 22462 19116 22468 19168
rect 22520 19156 22526 19168
rect 23750 19156 23756 19168
rect 22520 19128 23756 19156
rect 22520 19116 22526 19128
rect 23750 19116 23756 19128
rect 23808 19116 23814 19168
rect 23934 19116 23940 19168
rect 23992 19156 23998 19168
rect 24136 19156 24164 19187
rect 23992 19128 24164 19156
rect 23992 19116 23998 19128
rect 25130 19116 25136 19168
rect 25188 19156 25194 19168
rect 25639 19159 25697 19165
rect 25639 19156 25651 19159
rect 25188 19128 25651 19156
rect 25188 19116 25194 19128
rect 25639 19125 25651 19128
rect 25685 19125 25697 19159
rect 25639 19119 25697 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 12250 18952 12256 18964
rect 11900 18924 12256 18952
rect 11238 18844 11244 18896
rect 11296 18884 11302 18896
rect 11900 18893 11928 18924
rect 12250 18912 12256 18924
rect 12308 18952 12314 18964
rect 13906 18952 13912 18964
rect 12308 18924 13492 18952
rect 13867 18924 13912 18952
rect 12308 18912 12314 18924
rect 11333 18887 11391 18893
rect 11333 18884 11345 18887
rect 11296 18856 11345 18884
rect 11296 18844 11302 18856
rect 11333 18853 11345 18856
rect 11379 18853 11391 18887
rect 11333 18847 11391 18853
rect 11885 18887 11943 18893
rect 11885 18853 11897 18887
rect 11931 18853 11943 18887
rect 12894 18884 12900 18896
rect 12855 18856 12900 18884
rect 11885 18847 11943 18853
rect 12894 18844 12900 18856
rect 12952 18844 12958 18896
rect 13464 18893 13492 18924
rect 13906 18912 13912 18924
rect 13964 18912 13970 18964
rect 16298 18952 16304 18964
rect 16259 18924 16304 18952
rect 16298 18912 16304 18924
rect 16356 18912 16362 18964
rect 19889 18955 19947 18961
rect 19889 18921 19901 18955
rect 19935 18952 19947 18955
rect 20438 18952 20444 18964
rect 19935 18924 20444 18952
rect 19935 18921 19947 18924
rect 19889 18915 19947 18921
rect 20438 18912 20444 18924
rect 20496 18912 20502 18964
rect 22370 18912 22376 18964
rect 22428 18952 22434 18964
rect 22465 18955 22523 18961
rect 22465 18952 22477 18955
rect 22428 18924 22477 18952
rect 22428 18912 22434 18924
rect 22465 18921 22477 18924
rect 22511 18921 22523 18955
rect 23014 18952 23020 18964
rect 22975 18924 23020 18952
rect 22465 18915 22523 18921
rect 23014 18912 23020 18924
rect 23072 18912 23078 18964
rect 23382 18912 23388 18964
rect 23440 18952 23446 18964
rect 23934 18952 23940 18964
rect 23440 18924 23940 18952
rect 23440 18912 23446 18924
rect 23934 18912 23940 18924
rect 23992 18912 23998 18964
rect 24765 18955 24823 18961
rect 24765 18921 24777 18955
rect 24811 18952 24823 18955
rect 27614 18952 27620 18964
rect 24811 18924 27620 18952
rect 24811 18921 24823 18924
rect 24765 18915 24823 18921
rect 27614 18912 27620 18924
rect 27672 18912 27678 18964
rect 13449 18887 13507 18893
rect 13449 18853 13461 18887
rect 13495 18853 13507 18887
rect 13449 18847 13507 18853
rect 15473 18887 15531 18893
rect 15473 18853 15485 18887
rect 15519 18884 15531 18887
rect 15746 18884 15752 18896
rect 15519 18856 15752 18884
rect 15519 18853 15531 18856
rect 15473 18847 15531 18853
rect 15746 18844 15752 18856
rect 15804 18844 15810 18896
rect 18966 18884 18972 18896
rect 18927 18856 18972 18884
rect 18966 18844 18972 18856
rect 19024 18844 19030 18896
rect 23842 18844 23848 18896
rect 23900 18884 23906 18896
rect 24305 18887 24363 18893
rect 24305 18884 24317 18887
rect 23900 18856 24317 18884
rect 23900 18844 23906 18856
rect 24305 18853 24317 18856
rect 24351 18853 24363 18887
rect 24305 18847 24363 18853
rect 20990 18816 20996 18828
rect 20951 18788 20996 18816
rect 20990 18776 20996 18788
rect 21048 18776 21054 18828
rect 22094 18816 22100 18828
rect 22055 18788 22100 18816
rect 22094 18776 22100 18788
rect 22152 18776 22158 18828
rect 23106 18776 23112 18828
rect 23164 18816 23170 18828
rect 24581 18819 24639 18825
rect 24581 18816 24593 18819
rect 23164 18788 24593 18816
rect 23164 18776 23170 18788
rect 24581 18785 24593 18788
rect 24627 18816 24639 18819
rect 24670 18816 24676 18828
rect 24627 18788 24676 18816
rect 24627 18785 24639 18788
rect 24581 18779 24639 18785
rect 24670 18776 24676 18788
rect 24728 18776 24734 18828
rect 11241 18751 11299 18757
rect 11241 18717 11253 18751
rect 11287 18748 11299 18751
rect 11330 18748 11336 18760
rect 11287 18720 11336 18748
rect 11287 18717 11299 18720
rect 11241 18711 11299 18717
rect 11330 18708 11336 18720
rect 11388 18708 11394 18760
rect 12805 18751 12863 18757
rect 12805 18748 12817 18751
rect 12544 18720 12817 18748
rect 12544 18624 12572 18720
rect 12805 18717 12817 18720
rect 12851 18717 12863 18751
rect 12805 18711 12863 18717
rect 15381 18751 15439 18757
rect 15381 18717 15393 18751
rect 15427 18748 15439 18751
rect 16114 18748 16120 18760
rect 15427 18720 16120 18748
rect 15427 18717 15439 18720
rect 15381 18711 15439 18717
rect 16114 18708 16120 18720
rect 16172 18708 16178 18760
rect 17770 18748 17776 18760
rect 17731 18720 17776 18748
rect 17770 18708 17776 18720
rect 17828 18708 17834 18760
rect 18874 18748 18880 18760
rect 18835 18720 18880 18748
rect 18874 18708 18880 18720
rect 18932 18708 18938 18760
rect 23474 18708 23480 18760
rect 23532 18748 23538 18760
rect 25222 18748 25228 18760
rect 23532 18720 25228 18748
rect 23532 18708 23538 18720
rect 25222 18708 25228 18720
rect 25280 18708 25286 18760
rect 15930 18680 15936 18692
rect 15891 18652 15936 18680
rect 15930 18640 15936 18652
rect 15988 18680 15994 18692
rect 19242 18680 19248 18692
rect 15988 18652 19248 18680
rect 15988 18640 15994 18652
rect 19242 18640 19248 18652
rect 19300 18640 19306 18692
rect 19426 18680 19432 18692
rect 19387 18652 19432 18680
rect 19426 18640 19432 18652
rect 19484 18640 19490 18692
rect 21223 18683 21281 18689
rect 21223 18649 21235 18683
rect 21269 18680 21281 18683
rect 21269 18652 24691 18680
rect 21269 18649 21281 18652
rect 21223 18643 21281 18649
rect 10134 18572 10140 18624
rect 10192 18612 10198 18624
rect 10321 18615 10379 18621
rect 10321 18612 10333 18615
rect 10192 18584 10333 18612
rect 10192 18572 10198 18584
rect 10321 18581 10333 18584
rect 10367 18581 10379 18615
rect 12526 18612 12532 18624
rect 12487 18584 12532 18612
rect 10321 18575 10379 18581
rect 12526 18572 12532 18584
rect 12584 18572 12590 18624
rect 17954 18572 17960 18624
rect 18012 18612 18018 18624
rect 18233 18615 18291 18621
rect 18233 18612 18245 18615
rect 18012 18584 18245 18612
rect 18012 18572 18018 18584
rect 18233 18581 18245 18584
rect 18279 18581 18291 18615
rect 18233 18575 18291 18581
rect 21542 18572 21548 18624
rect 21600 18612 21606 18624
rect 21821 18615 21879 18621
rect 21821 18612 21833 18615
rect 21600 18584 21833 18612
rect 21600 18572 21606 18584
rect 21821 18581 21833 18584
rect 21867 18581 21879 18615
rect 24663 18612 24691 18652
rect 25222 18612 25228 18624
rect 24663 18584 25228 18612
rect 21821 18575 21879 18581
rect 25222 18572 25228 18584
rect 25280 18572 25286 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 11238 18368 11244 18420
rect 11296 18408 11302 18420
rect 11517 18411 11575 18417
rect 11517 18408 11529 18411
rect 11296 18380 11529 18408
rect 11296 18368 11302 18380
rect 11517 18377 11529 18380
rect 11563 18377 11575 18411
rect 16114 18408 16120 18420
rect 16075 18380 16120 18408
rect 11517 18371 11575 18377
rect 16114 18368 16120 18380
rect 16172 18408 16178 18420
rect 16172 18380 16344 18408
rect 16172 18368 16178 18380
rect 7466 18300 7472 18352
rect 7524 18340 7530 18352
rect 7524 18312 10593 18340
rect 7524 18300 7530 18312
rect 8846 18272 8852 18284
rect 8807 18244 8852 18272
rect 8846 18232 8852 18244
rect 8904 18232 8910 18284
rect 10565 18272 10593 18312
rect 11330 18300 11336 18352
rect 11388 18340 11394 18352
rect 11885 18343 11943 18349
rect 11885 18340 11897 18343
rect 11388 18312 11897 18340
rect 11388 18300 11394 18312
rect 11885 18309 11897 18312
rect 11931 18309 11943 18343
rect 11885 18303 11943 18309
rect 13265 18275 13323 18281
rect 13265 18272 13277 18275
rect 10565 18244 13277 18272
rect 13265 18241 13277 18244
rect 13311 18272 13323 18275
rect 14185 18275 14243 18281
rect 14185 18272 14197 18275
rect 13311 18244 14197 18272
rect 13311 18241 13323 18244
rect 13265 18235 13323 18241
rect 14185 18241 14197 18244
rect 14231 18241 14243 18275
rect 14185 18235 14243 18241
rect 15473 18275 15531 18281
rect 15473 18241 15485 18275
rect 15519 18272 15531 18275
rect 15930 18272 15936 18284
rect 15519 18244 15936 18272
rect 15519 18241 15531 18244
rect 15473 18235 15531 18241
rect 15930 18232 15936 18244
rect 15988 18232 15994 18284
rect 16316 18281 16344 18380
rect 18874 18368 18880 18420
rect 18932 18408 18938 18420
rect 19797 18411 19855 18417
rect 19797 18408 19809 18411
rect 18932 18380 19809 18408
rect 18932 18368 18938 18380
rect 19797 18377 19809 18380
rect 19843 18377 19855 18411
rect 19797 18371 19855 18377
rect 21821 18411 21879 18417
rect 21821 18377 21833 18411
rect 21867 18408 21879 18411
rect 22094 18408 22100 18420
rect 21867 18380 22100 18408
rect 21867 18377 21879 18380
rect 21821 18371 21879 18377
rect 22094 18368 22100 18380
rect 22152 18368 22158 18420
rect 24670 18408 24676 18420
rect 24631 18380 24676 18408
rect 24670 18368 24676 18380
rect 24728 18368 24734 18420
rect 23201 18343 23259 18349
rect 23201 18340 23213 18343
rect 21284 18312 23213 18340
rect 16301 18275 16359 18281
rect 16301 18241 16313 18275
rect 16347 18241 16359 18275
rect 21284 18272 21312 18312
rect 23201 18309 23213 18312
rect 23247 18309 23259 18343
rect 23201 18303 23259 18309
rect 25409 18343 25467 18349
rect 25409 18309 25421 18343
rect 25455 18340 25467 18343
rect 27614 18340 27620 18352
rect 25455 18312 27620 18340
rect 25455 18309 25467 18312
rect 25409 18303 25467 18309
rect 27614 18300 27620 18312
rect 27672 18300 27678 18352
rect 16301 18235 16359 18241
rect 20916 18244 21312 18272
rect 21361 18275 21419 18281
rect 10134 18164 10140 18216
rect 10192 18204 10198 18216
rect 10321 18207 10379 18213
rect 10321 18204 10333 18207
rect 10192 18176 10333 18204
rect 10192 18164 10198 18176
rect 10321 18173 10333 18176
rect 10367 18173 10379 18207
rect 10321 18167 10379 18173
rect 10870 18164 10876 18216
rect 10928 18204 10934 18216
rect 11241 18207 11299 18213
rect 11241 18204 11253 18207
rect 10928 18176 11253 18204
rect 10928 18164 10934 18176
rect 11241 18173 11253 18176
rect 11287 18204 11299 18207
rect 12621 18207 12679 18213
rect 12621 18204 12633 18207
rect 11287 18176 12633 18204
rect 11287 18173 11299 18176
rect 11241 18167 11299 18173
rect 12621 18173 12633 18176
rect 12667 18204 12679 18207
rect 12894 18204 12900 18216
rect 12667 18176 12900 18204
rect 12667 18173 12679 18176
rect 12621 18167 12679 18173
rect 12894 18164 12900 18176
rect 12952 18164 12958 18216
rect 18325 18207 18383 18213
rect 18325 18173 18337 18207
rect 18371 18204 18383 18207
rect 18966 18204 18972 18216
rect 18371 18176 18972 18204
rect 18371 18173 18383 18176
rect 18325 18167 18383 18173
rect 18966 18164 18972 18176
rect 19024 18204 19030 18216
rect 19429 18207 19487 18213
rect 19429 18204 19441 18207
rect 19024 18176 19441 18204
rect 19024 18164 19030 18176
rect 19429 18173 19441 18176
rect 19475 18173 19487 18207
rect 19429 18167 19487 18173
rect 20346 18164 20352 18216
rect 20404 18204 20410 18216
rect 20916 18213 20944 18244
rect 21361 18241 21373 18275
rect 21407 18272 21419 18275
rect 21910 18272 21916 18284
rect 21407 18244 21916 18272
rect 21407 18241 21419 18244
rect 21361 18235 21419 18241
rect 21910 18232 21916 18244
rect 21968 18232 21974 18284
rect 22278 18232 22284 18284
rect 22336 18272 22342 18284
rect 24213 18275 24271 18281
rect 24213 18272 24225 18275
rect 22336 18244 24225 18272
rect 22336 18232 22342 18244
rect 24213 18241 24225 18244
rect 24259 18241 24271 18275
rect 24213 18235 24271 18241
rect 20533 18207 20591 18213
rect 20533 18204 20545 18207
rect 20404 18176 20545 18204
rect 20404 18164 20410 18176
rect 20533 18173 20545 18176
rect 20579 18204 20591 18207
rect 20901 18207 20959 18213
rect 20901 18204 20913 18207
rect 20579 18176 20913 18204
rect 20579 18173 20591 18176
rect 20533 18167 20591 18173
rect 20901 18173 20913 18176
rect 20947 18173 20959 18207
rect 21082 18204 21088 18216
rect 21043 18176 21088 18204
rect 20901 18167 20959 18173
rect 21082 18164 21088 18176
rect 21140 18164 21146 18216
rect 22592 18207 22650 18213
rect 22592 18173 22604 18207
rect 22638 18204 22650 18207
rect 23017 18207 23075 18213
rect 23017 18204 23029 18207
rect 22638 18176 23029 18204
rect 22638 18173 22650 18176
rect 22592 18167 22650 18173
rect 23017 18173 23029 18176
rect 23063 18173 23075 18207
rect 23017 18167 23075 18173
rect 23201 18207 23259 18213
rect 23201 18173 23213 18207
rect 23247 18204 23259 18207
rect 23477 18207 23535 18213
rect 23477 18204 23489 18207
rect 23247 18176 23489 18204
rect 23247 18173 23259 18176
rect 23201 18167 23259 18173
rect 23477 18173 23489 18176
rect 23523 18204 23535 18207
rect 23661 18207 23719 18213
rect 23661 18204 23673 18207
rect 23523 18176 23673 18204
rect 23523 18173 23535 18176
rect 23477 18167 23535 18173
rect 23661 18173 23673 18176
rect 23707 18173 23719 18207
rect 23661 18167 23719 18173
rect 8665 18139 8723 18145
rect 8665 18105 8677 18139
rect 8711 18136 8723 18139
rect 8938 18136 8944 18148
rect 8711 18108 8944 18136
rect 8711 18105 8723 18108
rect 8665 18099 8723 18105
rect 8938 18096 8944 18108
rect 8996 18096 9002 18148
rect 9490 18136 9496 18148
rect 9451 18108 9496 18136
rect 9490 18096 9496 18108
rect 9548 18096 9554 18148
rect 10642 18139 10700 18145
rect 10642 18136 10654 18139
rect 10152 18108 10654 18136
rect 9766 18028 9772 18080
rect 9824 18068 9830 18080
rect 10152 18077 10180 18108
rect 10642 18105 10654 18108
rect 10688 18105 10700 18139
rect 10642 18099 10700 18105
rect 13357 18139 13415 18145
rect 13357 18105 13369 18139
rect 13403 18105 13415 18139
rect 13357 18099 13415 18105
rect 13909 18139 13967 18145
rect 13909 18105 13921 18139
rect 13955 18136 13967 18139
rect 14826 18136 14832 18148
rect 13955 18108 14832 18136
rect 13955 18105 13967 18108
rect 13909 18099 13967 18105
rect 10137 18071 10195 18077
rect 10137 18068 10149 18071
rect 9824 18040 10149 18068
rect 9824 18028 9830 18040
rect 10137 18037 10149 18040
rect 10183 18037 10195 18071
rect 10137 18031 10195 18037
rect 13081 18071 13139 18077
rect 13081 18037 13093 18071
rect 13127 18068 13139 18071
rect 13372 18068 13400 18099
rect 14826 18096 14832 18108
rect 14884 18096 14890 18148
rect 14921 18139 14979 18145
rect 14921 18105 14933 18139
rect 14967 18105 14979 18139
rect 19150 18136 19156 18148
rect 19111 18108 19156 18136
rect 14921 18099 14979 18105
rect 13630 18068 13636 18080
rect 13127 18040 13636 18068
rect 13127 18037 13139 18040
rect 13081 18031 13139 18037
rect 13630 18028 13636 18040
rect 13688 18028 13694 18080
rect 14645 18071 14703 18077
rect 14645 18037 14657 18071
rect 14691 18068 14703 18071
rect 14936 18068 14964 18099
rect 19150 18096 19156 18108
rect 19208 18096 19214 18148
rect 19518 18096 19524 18148
rect 19576 18136 19582 18148
rect 22607 18136 22635 18167
rect 24026 18164 24032 18216
rect 24084 18204 24090 18216
rect 24121 18207 24179 18213
rect 24121 18204 24133 18207
rect 24084 18176 24133 18204
rect 24084 18164 24090 18176
rect 24121 18173 24133 18176
rect 24167 18173 24179 18207
rect 25222 18204 25228 18216
rect 25183 18176 25228 18204
rect 24121 18167 24179 18173
rect 25222 18164 25228 18176
rect 25280 18204 25286 18216
rect 25777 18207 25835 18213
rect 25777 18204 25789 18207
rect 25280 18176 25789 18204
rect 25280 18164 25286 18176
rect 25777 18173 25789 18176
rect 25823 18173 25835 18207
rect 25777 18167 25835 18173
rect 19576 18108 22635 18136
rect 22695 18139 22753 18145
rect 19576 18096 19582 18108
rect 22695 18105 22707 18139
rect 22741 18136 22753 18139
rect 25038 18136 25044 18148
rect 22741 18108 25044 18136
rect 22741 18105 22753 18108
rect 22695 18099 22753 18105
rect 25038 18096 25044 18108
rect 25096 18096 25102 18148
rect 15378 18068 15384 18080
rect 14691 18040 15384 18068
rect 14691 18037 14703 18040
rect 14645 18031 14703 18037
rect 15378 18028 15384 18040
rect 15436 18028 15442 18080
rect 15746 18068 15752 18080
rect 15707 18040 15752 18068
rect 15746 18028 15752 18040
rect 15804 18028 15810 18080
rect 16942 18068 16948 18080
rect 16903 18040 16948 18068
rect 16942 18028 16948 18040
rect 17000 18028 17006 18080
rect 22189 18071 22247 18077
rect 22189 18037 22201 18071
rect 22235 18068 22247 18071
rect 22278 18068 22284 18080
rect 22235 18040 22284 18068
rect 22235 18037 22247 18040
rect 22189 18031 22247 18037
rect 22278 18028 22284 18040
rect 22336 18028 22342 18080
rect 23382 18028 23388 18080
rect 23440 18068 23446 18080
rect 24026 18068 24032 18080
rect 23440 18040 24032 18068
rect 23440 18028 23446 18040
rect 24026 18028 24032 18040
rect 24084 18028 24090 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 8846 17864 8852 17876
rect 8807 17836 8852 17864
rect 8846 17824 8852 17836
rect 8904 17824 8910 17876
rect 8938 17824 8944 17876
rect 8996 17864 9002 17876
rect 10597 17867 10655 17873
rect 10597 17864 10609 17867
rect 8996 17836 10609 17864
rect 8996 17824 9002 17836
rect 10597 17833 10609 17836
rect 10643 17864 10655 17867
rect 14826 17864 14832 17876
rect 10643 17836 11560 17864
rect 14787 17836 14832 17864
rect 10643 17833 10655 17836
rect 10597 17827 10655 17833
rect 9766 17756 9772 17808
rect 9824 17796 9830 17808
rect 9998 17799 10056 17805
rect 9998 17796 10010 17799
rect 9824 17768 10010 17796
rect 9824 17756 9830 17768
rect 9998 17765 10010 17768
rect 10044 17765 10056 17799
rect 9998 17759 10056 17765
rect 11532 17740 11560 17836
rect 14826 17824 14832 17836
rect 14884 17824 14890 17876
rect 15746 17864 15752 17876
rect 15707 17836 15752 17864
rect 15746 17824 15752 17836
rect 15804 17824 15810 17876
rect 17954 17864 17960 17876
rect 17915 17836 17960 17864
rect 17954 17824 17960 17836
rect 18012 17824 18018 17876
rect 22002 17864 22008 17876
rect 21963 17836 22008 17864
rect 22002 17824 22008 17836
rect 22060 17824 22066 17876
rect 23017 17867 23075 17873
rect 23017 17833 23029 17867
rect 23063 17864 23075 17867
rect 23063 17836 24072 17864
rect 23063 17833 23075 17836
rect 23017 17827 23075 17833
rect 13811 17799 13869 17805
rect 13811 17765 13823 17799
rect 13857 17796 13869 17799
rect 13998 17796 14004 17808
rect 13857 17768 14004 17796
rect 13857 17765 13869 17768
rect 13811 17759 13869 17765
rect 13998 17756 14004 17768
rect 14056 17756 14062 17808
rect 16761 17799 16819 17805
rect 16761 17765 16773 17799
rect 16807 17796 16819 17799
rect 16807 17768 17724 17796
rect 16807 17765 16819 17768
rect 16761 17759 16819 17765
rect 11514 17728 11520 17740
rect 11427 17700 11520 17728
rect 11514 17688 11520 17700
rect 11572 17688 11578 17740
rect 14369 17731 14427 17737
rect 14369 17697 14381 17731
rect 14415 17728 14427 17731
rect 15378 17728 15384 17740
rect 14415 17700 15384 17728
rect 14415 17697 14427 17700
rect 14369 17691 14427 17697
rect 15378 17688 15384 17700
rect 15436 17688 15442 17740
rect 16850 17728 16856 17740
rect 16811 17700 16856 17728
rect 16850 17688 16856 17700
rect 16908 17688 16914 17740
rect 16942 17688 16948 17740
rect 17000 17728 17006 17740
rect 17696 17737 17724 17768
rect 17770 17756 17776 17808
rect 17828 17796 17834 17808
rect 18782 17796 18788 17808
rect 17828 17768 18788 17796
rect 17828 17756 17834 17768
rect 18782 17756 18788 17768
rect 18840 17796 18846 17808
rect 18969 17799 19027 17805
rect 18969 17796 18981 17799
rect 18840 17768 18981 17796
rect 18840 17756 18846 17768
rect 18969 17765 18981 17768
rect 19015 17765 19027 17799
rect 18969 17759 19027 17765
rect 19061 17799 19119 17805
rect 19061 17765 19073 17799
rect 19107 17796 19119 17799
rect 19150 17796 19156 17808
rect 19107 17768 19156 17796
rect 19107 17765 19119 17768
rect 19061 17759 19119 17765
rect 19150 17756 19156 17768
rect 19208 17756 19214 17808
rect 20806 17756 20812 17808
rect 20864 17796 20870 17808
rect 20864 17768 22093 17796
rect 20864 17756 20870 17768
rect 17313 17731 17371 17737
rect 17313 17728 17325 17731
rect 17000 17700 17325 17728
rect 17000 17688 17006 17700
rect 17313 17697 17325 17700
rect 17359 17697 17371 17731
rect 17313 17691 17371 17697
rect 17681 17731 17739 17737
rect 17681 17697 17693 17731
rect 17727 17728 17739 17731
rect 17862 17728 17868 17740
rect 17727 17700 17868 17728
rect 17727 17697 17739 17700
rect 17681 17691 17739 17697
rect 17862 17688 17868 17700
rect 17920 17688 17926 17740
rect 21152 17731 21210 17737
rect 21152 17697 21164 17731
rect 21198 17728 21210 17731
rect 22065 17728 22093 17768
rect 22278 17756 22284 17808
rect 22336 17796 22342 17808
rect 24044 17805 24072 17836
rect 22418 17799 22476 17805
rect 22418 17796 22430 17799
rect 22336 17768 22430 17796
rect 22336 17756 22342 17768
rect 22418 17765 22430 17768
rect 22464 17765 22476 17799
rect 22418 17759 22476 17765
rect 24029 17799 24087 17805
rect 24029 17765 24041 17799
rect 24075 17796 24087 17799
rect 24762 17796 24768 17808
rect 24075 17768 24768 17796
rect 24075 17765 24087 17768
rect 24029 17759 24087 17765
rect 24762 17756 24768 17768
rect 24820 17756 24826 17808
rect 23382 17728 23388 17740
rect 21198 17700 21680 17728
rect 22065 17700 23388 17728
rect 21198 17697 21210 17700
rect 21152 17691 21210 17697
rect 9674 17660 9680 17672
rect 9635 17632 9680 17660
rect 9674 17620 9680 17632
rect 9732 17620 9738 17672
rect 10410 17620 10416 17672
rect 10468 17660 10474 17672
rect 11425 17663 11483 17669
rect 11425 17660 11437 17663
rect 10468 17632 11437 17660
rect 10468 17620 10474 17632
rect 11425 17629 11437 17632
rect 11471 17629 11483 17663
rect 13449 17663 13507 17669
rect 13449 17660 13461 17663
rect 11425 17623 11483 17629
rect 13280 17632 13461 17660
rect 13280 17536 13308 17632
rect 13449 17629 13461 17632
rect 13495 17629 13507 17663
rect 13449 17623 13507 17629
rect 16393 17663 16451 17669
rect 16393 17629 16405 17663
rect 16439 17660 16451 17663
rect 16960 17660 16988 17688
rect 19426 17660 19432 17672
rect 16439 17632 16988 17660
rect 19387 17632 19432 17660
rect 16439 17629 16451 17632
rect 16393 17623 16451 17629
rect 19426 17620 19432 17632
rect 19484 17620 19490 17672
rect 20717 17595 20775 17601
rect 20717 17561 20729 17595
rect 20763 17592 20775 17595
rect 21082 17592 21088 17604
rect 20763 17564 21088 17592
rect 20763 17561 20775 17564
rect 20717 17555 20775 17561
rect 21082 17552 21088 17564
rect 21140 17592 21146 17604
rect 21358 17592 21364 17604
rect 21140 17564 21364 17592
rect 21140 17552 21146 17564
rect 21358 17552 21364 17564
rect 21416 17552 21422 17604
rect 21652 17601 21680 17700
rect 23382 17688 23388 17700
rect 23440 17728 23446 17740
rect 23661 17731 23719 17737
rect 23661 17728 23673 17731
rect 23440 17700 23673 17728
rect 23440 17688 23446 17700
rect 23661 17697 23673 17700
rect 23707 17697 23719 17731
rect 23661 17691 23719 17697
rect 22094 17660 22100 17672
rect 22055 17632 22100 17660
rect 22094 17620 22100 17632
rect 22152 17620 22158 17672
rect 23566 17620 23572 17672
rect 23624 17660 23630 17672
rect 23750 17660 23756 17672
rect 23624 17632 23756 17660
rect 23624 17620 23630 17632
rect 23750 17620 23756 17632
rect 23808 17660 23814 17672
rect 23937 17663 23995 17669
rect 23937 17660 23949 17663
rect 23808 17632 23949 17660
rect 23808 17620 23814 17632
rect 23937 17629 23949 17632
rect 23983 17629 23995 17663
rect 23937 17623 23995 17629
rect 24213 17663 24271 17669
rect 24213 17629 24225 17663
rect 24259 17629 24271 17663
rect 24213 17623 24271 17629
rect 21637 17595 21695 17601
rect 21637 17561 21649 17595
rect 21683 17592 21695 17595
rect 24026 17592 24032 17604
rect 21683 17564 24032 17592
rect 21683 17561 21695 17564
rect 21637 17555 21695 17561
rect 24026 17552 24032 17564
rect 24084 17592 24090 17604
rect 24228 17592 24256 17623
rect 24670 17620 24676 17672
rect 24728 17660 24734 17672
rect 25409 17663 25467 17669
rect 25409 17660 25421 17663
rect 24728 17632 25421 17660
rect 24728 17620 24734 17632
rect 25409 17629 25421 17632
rect 25455 17629 25467 17663
rect 25409 17623 25467 17629
rect 24084 17564 24256 17592
rect 24084 17552 24090 17564
rect 12618 17484 12624 17536
rect 12676 17524 12682 17536
rect 12713 17527 12771 17533
rect 12713 17524 12725 17527
rect 12676 17496 12725 17524
rect 12676 17484 12682 17496
rect 12713 17493 12725 17496
rect 12759 17493 12771 17527
rect 13262 17524 13268 17536
rect 13223 17496 13268 17524
rect 12713 17487 12771 17493
rect 13262 17484 13268 17496
rect 13320 17484 13326 17536
rect 18230 17524 18236 17536
rect 18191 17496 18236 17524
rect 18230 17484 18236 17496
rect 18288 17484 18294 17536
rect 21223 17527 21281 17533
rect 21223 17493 21235 17527
rect 21269 17524 21281 17527
rect 21818 17524 21824 17536
rect 21269 17496 21824 17524
rect 21269 17493 21281 17496
rect 21223 17487 21281 17493
rect 21818 17484 21824 17496
rect 21876 17484 21882 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 11514 17320 11520 17332
rect 11475 17292 11520 17320
rect 11514 17280 11520 17292
rect 11572 17280 11578 17332
rect 13630 17320 13636 17332
rect 13591 17292 13636 17320
rect 13630 17280 13636 17292
rect 13688 17280 13694 17332
rect 17129 17323 17187 17329
rect 17129 17289 17141 17323
rect 17175 17320 17187 17323
rect 17678 17320 17684 17332
rect 17175 17292 17684 17320
rect 17175 17289 17187 17292
rect 17129 17283 17187 17289
rect 17678 17280 17684 17292
rect 17736 17280 17742 17332
rect 18966 17320 18972 17332
rect 18927 17292 18972 17320
rect 18966 17280 18972 17292
rect 19024 17280 19030 17332
rect 19150 17280 19156 17332
rect 19208 17320 19214 17332
rect 19245 17323 19303 17329
rect 19245 17320 19257 17323
rect 19208 17292 19257 17320
rect 19208 17280 19214 17292
rect 19245 17289 19257 17292
rect 19291 17289 19303 17323
rect 20346 17320 20352 17332
rect 20307 17292 20352 17320
rect 19245 17283 19303 17289
rect 20346 17280 20352 17292
rect 20404 17280 20410 17332
rect 25222 17320 25228 17332
rect 23446 17292 25228 17320
rect 9490 17212 9496 17264
rect 9548 17252 9554 17264
rect 10873 17255 10931 17261
rect 10873 17252 10885 17255
rect 9548 17224 10885 17252
rect 9548 17212 9554 17224
rect 10873 17221 10885 17224
rect 10919 17252 10931 17255
rect 12526 17252 12532 17264
rect 10919 17224 12532 17252
rect 10919 17221 10931 17224
rect 10873 17215 10931 17221
rect 12526 17212 12532 17224
rect 12584 17212 12590 17264
rect 18782 17212 18788 17264
rect 18840 17252 18846 17264
rect 19613 17255 19671 17261
rect 19613 17252 19625 17255
rect 18840 17224 19625 17252
rect 18840 17212 18846 17224
rect 19613 17221 19625 17224
rect 19659 17221 19671 17255
rect 20364 17252 20392 17280
rect 22695 17255 22753 17261
rect 20364 17224 20484 17252
rect 19613 17215 19671 17221
rect 9401 17187 9459 17193
rect 9401 17153 9413 17187
rect 9447 17184 9459 17187
rect 9674 17184 9680 17196
rect 9447 17156 9680 17184
rect 9447 17153 9459 17156
rect 9401 17147 9459 17153
rect 9674 17144 9680 17156
rect 9732 17144 9738 17196
rect 10321 17187 10379 17193
rect 10321 17153 10333 17187
rect 10367 17184 10379 17187
rect 10962 17184 10968 17196
rect 10367 17156 10968 17184
rect 10367 17153 10379 17156
rect 10321 17147 10379 17153
rect 10962 17144 10968 17156
rect 11020 17144 11026 17196
rect 14826 17184 14832 17196
rect 14787 17156 14832 17184
rect 14826 17144 14832 17156
rect 14884 17144 14890 17196
rect 15565 17187 15623 17193
rect 15565 17153 15577 17187
rect 15611 17184 15623 17187
rect 16942 17184 16948 17196
rect 15611 17156 16804 17184
rect 16903 17156 16948 17184
rect 15611 17153 15623 17156
rect 15565 17147 15623 17153
rect 8573 17119 8631 17125
rect 8573 17085 8585 17119
rect 8619 17116 8631 17119
rect 8941 17119 8999 17125
rect 8941 17116 8953 17119
rect 8619 17088 8953 17116
rect 8619 17085 8631 17088
rect 8573 17079 8631 17085
rect 8941 17085 8953 17088
rect 8987 17116 8999 17119
rect 9030 17116 9036 17128
rect 8987 17088 9036 17116
rect 8987 17085 8999 17088
rect 8941 17079 8999 17085
rect 9030 17076 9036 17088
rect 9088 17076 9094 17128
rect 9214 17116 9220 17128
rect 9175 17088 9220 17116
rect 9214 17076 9220 17088
rect 9272 17076 9278 17128
rect 12618 17076 12624 17128
rect 12676 17116 12682 17128
rect 12713 17119 12771 17125
rect 12713 17116 12725 17119
rect 12676 17088 12725 17116
rect 12676 17076 12682 17088
rect 12713 17085 12725 17088
rect 12759 17085 12771 17119
rect 12713 17079 12771 17085
rect 13630 17076 13636 17128
rect 13688 17116 13694 17128
rect 14182 17116 14188 17128
rect 13688 17088 14188 17116
rect 13688 17076 13694 17088
rect 14182 17076 14188 17088
rect 14240 17076 14246 17128
rect 16025 17119 16083 17125
rect 16025 17116 16037 17119
rect 15856 17088 16037 17116
rect 10410 17008 10416 17060
rect 10468 17048 10474 17060
rect 10468 17020 10513 17048
rect 10468 17008 10474 17020
rect 14274 17008 14280 17060
rect 14332 17048 14338 17060
rect 14553 17051 14611 17057
rect 14553 17048 14565 17051
rect 14332 17020 14565 17048
rect 14332 17008 14338 17020
rect 14553 17017 14565 17020
rect 14599 17017 14611 17051
rect 14553 17011 14611 17017
rect 14645 17051 14703 17057
rect 14645 17017 14657 17051
rect 14691 17017 14703 17051
rect 14645 17011 14703 17017
rect 9766 16980 9772 16992
rect 9727 16952 9772 16980
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 10137 16983 10195 16989
rect 10137 16949 10149 16983
rect 10183 16980 10195 16983
rect 10428 16980 10456 17008
rect 10183 16952 10456 16980
rect 10183 16949 10195 16952
rect 10137 16943 10195 16949
rect 12710 16940 12716 16992
rect 12768 16980 12774 16992
rect 13081 16983 13139 16989
rect 13081 16980 13093 16983
rect 12768 16952 13093 16980
rect 12768 16940 12774 16952
rect 13081 16949 13093 16952
rect 13127 16980 13139 16983
rect 13909 16983 13967 16989
rect 13909 16980 13921 16983
rect 13127 16952 13921 16980
rect 13127 16949 13139 16952
rect 13081 16943 13139 16949
rect 13909 16949 13921 16952
rect 13955 16980 13967 16983
rect 13998 16980 14004 16992
rect 13955 16952 14004 16980
rect 13955 16949 13967 16952
rect 13909 16943 13967 16949
rect 13998 16940 14004 16952
rect 14056 16940 14062 16992
rect 14366 16980 14372 16992
rect 14327 16952 14372 16980
rect 14366 16940 14372 16952
rect 14424 16980 14430 16992
rect 14660 16980 14688 17011
rect 15856 16992 15884 17088
rect 16025 17085 16037 17088
rect 16071 17085 16083 17119
rect 16776 17116 16804 17156
rect 16942 17144 16948 17156
rect 17000 17144 17006 17196
rect 18322 17144 18328 17196
rect 18380 17184 18386 17196
rect 20346 17184 20352 17196
rect 18380 17156 20352 17184
rect 18380 17144 18386 17156
rect 20346 17144 20352 17156
rect 20404 17144 20410 17196
rect 16853 17119 16911 17125
rect 16853 17116 16865 17119
rect 16776 17088 16865 17116
rect 16025 17079 16083 17085
rect 16853 17085 16865 17088
rect 16899 17085 16911 17119
rect 16853 17079 16911 17085
rect 16868 17048 16896 17079
rect 17126 17076 17132 17128
rect 17184 17116 17190 17128
rect 18049 17119 18107 17125
rect 18049 17116 18061 17119
rect 17184 17088 18061 17116
rect 17184 17076 17190 17088
rect 18049 17085 18061 17088
rect 18095 17116 18107 17119
rect 18230 17116 18236 17128
rect 18095 17088 18236 17116
rect 18095 17085 18107 17088
rect 18049 17079 18107 17085
rect 18230 17076 18236 17088
rect 18288 17076 18294 17128
rect 20456 17116 20484 17224
rect 22695 17221 22707 17255
rect 22741 17252 22753 17255
rect 23446 17252 23474 17292
rect 25222 17280 25228 17292
rect 25280 17280 25286 17332
rect 25406 17320 25412 17332
rect 25367 17292 25412 17320
rect 25406 17280 25412 17292
rect 25464 17280 25470 17332
rect 24670 17252 24676 17264
rect 22741 17224 23474 17252
rect 23768 17224 24676 17252
rect 22741 17221 22753 17224
rect 22695 17215 22753 17221
rect 21542 17184 21548 17196
rect 21503 17156 21548 17184
rect 21542 17144 21548 17156
rect 21600 17144 21606 17196
rect 23768 17193 23796 17224
rect 24670 17212 24676 17224
rect 24728 17212 24734 17264
rect 24762 17212 24768 17264
rect 24820 17252 24826 17264
rect 24820 17224 24865 17252
rect 24820 17212 24826 17224
rect 23109 17187 23167 17193
rect 23109 17153 23121 17187
rect 23155 17184 23167 17187
rect 23753 17187 23811 17193
rect 23753 17184 23765 17187
rect 23155 17156 23765 17184
rect 23155 17153 23167 17156
rect 23109 17147 23167 17153
rect 23753 17153 23765 17156
rect 23799 17153 23811 17187
rect 24026 17184 24032 17196
rect 23987 17156 24032 17184
rect 23753 17147 23811 17153
rect 24026 17144 24032 17156
rect 24084 17144 24090 17196
rect 20809 17119 20867 17125
rect 20809 17116 20821 17119
rect 20456 17088 20821 17116
rect 20809 17085 20821 17088
rect 20855 17085 20867 17119
rect 21269 17119 21327 17125
rect 21269 17116 21281 17119
rect 20809 17079 20867 17085
rect 21192 17088 21281 17116
rect 17218 17048 17224 17060
rect 16868 17020 17224 17048
rect 17218 17008 17224 17020
rect 17276 17008 17282 17060
rect 17865 17051 17923 17057
rect 17865 17017 17877 17051
rect 17911 17048 17923 17051
rect 18138 17048 18144 17060
rect 17911 17020 18144 17048
rect 17911 17017 17923 17020
rect 17865 17011 17923 17017
rect 18138 17008 18144 17020
rect 18196 17048 18202 17060
rect 18411 17051 18469 17057
rect 18411 17048 18423 17051
rect 18196 17020 18423 17048
rect 18196 17008 18202 17020
rect 18411 17017 18423 17020
rect 18457 17048 18469 17051
rect 19150 17048 19156 17060
rect 18457 17020 19156 17048
rect 18457 17017 18469 17020
rect 18411 17011 18469 17017
rect 19150 17008 19156 17020
rect 19208 17008 19214 17060
rect 21192 16992 21220 17088
rect 21269 17085 21281 17088
rect 21315 17085 21327 17119
rect 21269 17079 21327 17085
rect 22624 17119 22682 17125
rect 22624 17085 22636 17119
rect 22670 17116 22682 17119
rect 22738 17116 22744 17128
rect 22670 17088 22744 17116
rect 22670 17085 22682 17088
rect 22624 17079 22682 17085
rect 22738 17076 22744 17088
rect 22796 17076 22802 17128
rect 25038 17076 25044 17128
rect 25096 17116 25102 17128
rect 25225 17119 25283 17125
rect 25225 17116 25237 17119
rect 25096 17088 25237 17116
rect 25096 17076 25102 17088
rect 25225 17085 25237 17088
rect 25271 17116 25283 17119
rect 25777 17119 25835 17125
rect 25777 17116 25789 17119
rect 25271 17088 25789 17116
rect 25271 17085 25283 17088
rect 25225 17079 25283 17085
rect 25777 17085 25789 17088
rect 25823 17085 25835 17119
rect 25777 17079 25835 17085
rect 23845 17051 23903 17057
rect 23845 17017 23857 17051
rect 23891 17017 23903 17051
rect 23845 17011 23903 17017
rect 15838 16980 15844 16992
rect 14424 16952 14688 16980
rect 15799 16952 15844 16980
rect 14424 16940 14430 16952
rect 15838 16940 15844 16952
rect 15896 16940 15902 16992
rect 16482 16940 16488 16992
rect 16540 16980 16546 16992
rect 16850 16980 16856 16992
rect 16540 16952 16856 16980
rect 16540 16940 16546 16952
rect 16850 16940 16856 16952
rect 16908 16980 16914 16992
rect 17405 16983 17463 16989
rect 17405 16980 17417 16983
rect 16908 16952 17417 16980
rect 16908 16940 16914 16952
rect 17405 16949 17417 16952
rect 17451 16949 17463 16983
rect 17405 16943 17463 16949
rect 19797 16983 19855 16989
rect 19797 16949 19809 16983
rect 19843 16980 19855 16983
rect 19978 16980 19984 16992
rect 19843 16952 19984 16980
rect 19843 16949 19855 16952
rect 19797 16943 19855 16949
rect 19978 16940 19984 16952
rect 20036 16940 20042 16992
rect 20717 16983 20775 16989
rect 20717 16949 20729 16983
rect 20763 16980 20775 16983
rect 21174 16980 21180 16992
rect 20763 16952 21180 16980
rect 20763 16949 20775 16952
rect 20717 16943 20775 16949
rect 21174 16940 21180 16952
rect 21232 16940 21238 16992
rect 22189 16983 22247 16989
rect 22189 16949 22201 16983
rect 22235 16980 22247 16983
rect 22278 16980 22284 16992
rect 22235 16952 22284 16980
rect 22235 16949 22247 16952
rect 22189 16943 22247 16949
rect 22278 16940 22284 16952
rect 22336 16940 22342 16992
rect 23477 16983 23535 16989
rect 23477 16949 23489 16983
rect 23523 16980 23535 16983
rect 23566 16980 23572 16992
rect 23523 16952 23572 16980
rect 23523 16949 23535 16952
rect 23477 16943 23535 16949
rect 23566 16940 23572 16952
rect 23624 16980 23630 16992
rect 23860 16980 23888 17011
rect 23624 16952 23888 16980
rect 23624 16940 23630 16952
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 9493 16779 9551 16785
rect 9493 16745 9505 16779
rect 9539 16776 9551 16779
rect 9674 16776 9680 16788
rect 9539 16748 9680 16776
rect 9539 16745 9551 16748
rect 9493 16739 9551 16745
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 10134 16776 10140 16788
rect 10095 16748 10140 16776
rect 10134 16736 10140 16748
rect 10192 16736 10198 16788
rect 13262 16776 13268 16788
rect 13223 16748 13268 16776
rect 13262 16736 13268 16748
rect 13320 16736 13326 16788
rect 15105 16779 15163 16785
rect 15105 16745 15117 16779
rect 15151 16776 15163 16779
rect 15378 16776 15384 16788
rect 15151 16748 15384 16776
rect 15151 16745 15163 16748
rect 15105 16739 15163 16745
rect 15378 16736 15384 16748
rect 15436 16736 15442 16788
rect 16758 16776 16764 16788
rect 16719 16748 16764 16776
rect 16758 16736 16764 16748
rect 16816 16736 16822 16788
rect 18690 16776 18696 16788
rect 18651 16748 18696 16776
rect 18690 16736 18696 16748
rect 18748 16736 18754 16788
rect 20070 16776 20076 16788
rect 19983 16748 20076 16776
rect 20070 16736 20076 16748
rect 20128 16776 20134 16788
rect 20622 16776 20628 16788
rect 20128 16748 20628 16776
rect 20128 16736 20134 16748
rect 20622 16736 20628 16748
rect 20680 16736 20686 16788
rect 22649 16779 22707 16785
rect 22649 16745 22661 16779
rect 22695 16776 22707 16779
rect 22738 16776 22744 16788
rect 22695 16748 22744 16776
rect 22695 16745 22707 16748
rect 22649 16739 22707 16745
rect 22738 16736 22744 16748
rect 22796 16736 22802 16788
rect 23566 16776 23572 16788
rect 23527 16748 23572 16776
rect 23566 16736 23572 16748
rect 23624 16736 23630 16788
rect 23750 16736 23756 16788
rect 23808 16776 23814 16788
rect 24305 16779 24363 16785
rect 24305 16776 24317 16779
rect 23808 16748 24317 16776
rect 23808 16736 23814 16748
rect 24305 16745 24317 16748
rect 24351 16745 24363 16779
rect 24305 16739 24363 16745
rect 8757 16711 8815 16717
rect 8757 16677 8769 16711
rect 8803 16708 8815 16711
rect 9214 16708 9220 16720
rect 8803 16680 9220 16708
rect 8803 16677 8815 16680
rect 8757 16671 8815 16677
rect 9214 16668 9220 16680
rect 9272 16708 9278 16720
rect 13906 16708 13912 16720
rect 9272 16680 13912 16708
rect 9272 16668 9278 16680
rect 9858 16640 9864 16652
rect 9819 16612 9864 16640
rect 9858 16600 9864 16612
rect 9916 16600 9922 16652
rect 10428 16649 10456 16680
rect 13906 16668 13912 16680
rect 13964 16668 13970 16720
rect 21266 16708 21272 16720
rect 21192 16680 21272 16708
rect 10413 16643 10471 16649
rect 10413 16609 10425 16643
rect 10459 16609 10471 16643
rect 11514 16640 11520 16652
rect 11475 16612 11520 16640
rect 10413 16603 10471 16609
rect 11514 16600 11520 16612
rect 11572 16600 11578 16652
rect 13078 16640 13084 16652
rect 13039 16612 13084 16640
rect 13078 16600 13084 16612
rect 13136 16600 13142 16652
rect 13446 16640 13452 16652
rect 13407 16612 13452 16640
rect 13446 16600 13452 16612
rect 13504 16600 13510 16652
rect 15286 16640 15292 16652
rect 15247 16612 15292 16640
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 16482 16640 16488 16652
rect 16443 16612 16488 16640
rect 16482 16600 16488 16612
rect 16540 16600 16546 16652
rect 16942 16640 16948 16652
rect 16903 16612 16948 16640
rect 16942 16600 16948 16612
rect 17000 16600 17006 16652
rect 17218 16600 17224 16652
rect 17276 16640 17282 16652
rect 17313 16643 17371 16649
rect 17313 16640 17325 16643
rect 17276 16612 17325 16640
rect 17276 16600 17282 16612
rect 17313 16609 17325 16612
rect 17359 16640 17371 16643
rect 18690 16640 18696 16652
rect 17359 16612 18696 16640
rect 17359 16609 17371 16612
rect 17313 16603 17371 16609
rect 18690 16600 18696 16612
rect 18748 16600 18754 16652
rect 21192 16649 21220 16680
rect 21266 16668 21272 16680
rect 21324 16668 21330 16720
rect 21637 16711 21695 16717
rect 21637 16677 21649 16711
rect 21683 16708 21695 16711
rect 22094 16708 22100 16720
rect 21683 16680 22100 16708
rect 21683 16677 21695 16680
rect 21637 16671 21695 16677
rect 22094 16668 22100 16680
rect 22152 16668 22158 16720
rect 18877 16643 18935 16649
rect 18877 16609 18889 16643
rect 18923 16609 18935 16643
rect 18877 16603 18935 16609
rect 21177 16643 21235 16649
rect 21177 16609 21189 16643
rect 21223 16609 21235 16643
rect 21358 16640 21364 16652
rect 21319 16612 21364 16640
rect 21177 16603 21235 16609
rect 11422 16572 11428 16584
rect 11383 16544 11428 16572
rect 11422 16532 11428 16544
rect 11480 16532 11486 16584
rect 13096 16572 13124 16600
rect 13538 16572 13544 16584
rect 13096 16544 13544 16572
rect 13538 16532 13544 16544
rect 13596 16572 13602 16584
rect 18892 16572 18920 16603
rect 21358 16600 21364 16612
rect 21416 16600 21422 16652
rect 23382 16600 23388 16652
rect 23440 16640 23446 16652
rect 23937 16643 23995 16649
rect 23937 16640 23949 16643
rect 23440 16612 23949 16640
rect 23440 16600 23446 16612
rect 23937 16609 23949 16612
rect 23983 16640 23995 16643
rect 24762 16640 24768 16652
rect 23983 16612 24768 16640
rect 23983 16609 23995 16612
rect 23937 16603 23995 16609
rect 24762 16600 24768 16612
rect 24820 16600 24826 16652
rect 13596 16544 13814 16572
rect 13596 16532 13602 16544
rect 9766 16464 9772 16516
rect 9824 16504 9830 16516
rect 12710 16504 12716 16516
rect 9824 16476 12716 16504
rect 9824 16464 9830 16476
rect 12710 16464 12716 16476
rect 12768 16464 12774 16516
rect 13786 16504 13814 16544
rect 18064 16544 18920 16572
rect 15473 16507 15531 16513
rect 15473 16504 15485 16507
rect 13786 16476 15485 16504
rect 15473 16473 15485 16476
rect 15519 16473 15531 16507
rect 15473 16467 15531 16473
rect 10962 16436 10968 16448
rect 10923 16408 10968 16436
rect 10962 16396 10968 16408
rect 11020 16396 11026 16448
rect 14182 16436 14188 16448
rect 14143 16408 14188 16436
rect 14182 16396 14188 16408
rect 14240 16396 14246 16448
rect 14274 16396 14280 16448
rect 14332 16436 14338 16448
rect 14461 16439 14519 16445
rect 14461 16436 14473 16439
rect 14332 16408 14473 16436
rect 14332 16396 14338 16408
rect 14461 16405 14473 16408
rect 14507 16405 14519 16439
rect 14461 16399 14519 16405
rect 16117 16439 16175 16445
rect 16117 16405 16129 16439
rect 16163 16436 16175 16439
rect 16758 16436 16764 16448
rect 16163 16408 16764 16436
rect 16163 16405 16175 16408
rect 16117 16399 16175 16405
rect 16758 16396 16764 16408
rect 16816 16396 16822 16448
rect 17954 16396 17960 16448
rect 18012 16436 18018 16448
rect 18064 16445 18092 16544
rect 24670 16532 24676 16584
rect 24728 16572 24734 16584
rect 24857 16575 24915 16581
rect 24857 16572 24869 16575
rect 24728 16544 24869 16572
rect 24728 16532 24734 16544
rect 24857 16541 24869 16544
rect 24903 16541 24915 16575
rect 24857 16535 24915 16541
rect 18049 16439 18107 16445
rect 18049 16436 18061 16439
rect 18012 16408 18061 16436
rect 18012 16396 18018 16408
rect 18049 16405 18061 16408
rect 18095 16405 18107 16439
rect 18049 16399 18107 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 9033 16235 9091 16241
rect 9033 16201 9045 16235
rect 9079 16232 9091 16235
rect 9214 16232 9220 16244
rect 9079 16204 9220 16232
rect 9079 16201 9091 16204
rect 9033 16195 9091 16201
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 9401 16235 9459 16241
rect 9401 16201 9413 16235
rect 9447 16232 9459 16235
rect 9769 16235 9827 16241
rect 9769 16232 9781 16235
rect 9447 16204 9781 16232
rect 9447 16201 9459 16204
rect 9401 16195 9459 16201
rect 9769 16201 9781 16204
rect 9815 16232 9827 16235
rect 9858 16232 9864 16244
rect 9815 16204 9864 16232
rect 9815 16201 9827 16204
rect 9769 16195 9827 16201
rect 9858 16192 9864 16204
rect 9916 16192 9922 16244
rect 11514 16232 11520 16244
rect 11475 16204 11520 16232
rect 11514 16192 11520 16204
rect 11572 16192 11578 16244
rect 12253 16235 12311 16241
rect 12253 16201 12265 16235
rect 12299 16232 12311 16235
rect 12342 16232 12348 16244
rect 12299 16204 12348 16232
rect 12299 16201 12311 16204
rect 12253 16195 12311 16201
rect 12342 16192 12348 16204
rect 12400 16192 12406 16244
rect 13538 16232 13544 16244
rect 13499 16204 13544 16232
rect 13538 16192 13544 16204
rect 13596 16192 13602 16244
rect 14366 16232 14372 16244
rect 14327 16204 14372 16232
rect 14366 16192 14372 16204
rect 14424 16192 14430 16244
rect 17126 16192 17132 16244
rect 17184 16232 17190 16244
rect 21085 16235 21143 16241
rect 21085 16232 21097 16235
rect 17184 16204 17229 16232
rect 18432 16204 21097 16232
rect 17184 16192 17190 16204
rect 16942 16096 16948 16108
rect 16903 16068 16948 16096
rect 16942 16056 16948 16068
rect 17000 16096 17006 16108
rect 17405 16099 17463 16105
rect 17405 16096 17417 16099
rect 17000 16068 17417 16096
rect 17000 16056 17006 16068
rect 17405 16065 17417 16068
rect 17451 16065 17463 16099
rect 17405 16059 17463 16065
rect 9858 16028 9864 16040
rect 9819 16000 9864 16028
rect 9858 15988 9864 16000
rect 9916 15988 9922 16040
rect 10413 16031 10471 16037
rect 10413 15997 10425 16031
rect 10459 16028 10471 16031
rect 10686 16028 10692 16040
rect 10459 16000 10692 16028
rect 10459 15997 10471 16000
rect 10413 15991 10471 15997
rect 10686 15988 10692 16000
rect 10744 15988 10750 16040
rect 12342 15988 12348 16040
rect 12400 16028 12406 16040
rect 12529 16031 12587 16037
rect 12529 16028 12541 16031
rect 12400 16000 12541 16028
rect 12400 15988 12406 16000
rect 12529 15997 12541 16000
rect 12575 15997 12587 16031
rect 12986 16028 12992 16040
rect 12947 16000 12992 16028
rect 12529 15991 12587 15997
rect 12986 15988 12992 16000
rect 13044 16028 13050 16040
rect 13446 16028 13452 16040
rect 13044 16000 13452 16028
rect 13044 15988 13050 16000
rect 13446 15988 13452 16000
rect 13504 16028 13510 16040
rect 13909 16031 13967 16037
rect 13909 16028 13921 16031
rect 13504 16000 13921 16028
rect 13504 15988 13510 16000
rect 13909 15997 13921 16000
rect 13955 15997 13967 16031
rect 14182 16028 14188 16040
rect 14143 16000 14188 16028
rect 13909 15991 13967 15997
rect 14182 15988 14188 16000
rect 14240 15988 14246 16040
rect 16025 16031 16083 16037
rect 16025 15997 16037 16031
rect 16071 15997 16083 16031
rect 16025 15991 16083 15997
rect 14642 15920 14648 15972
rect 14700 15960 14706 15972
rect 15838 15960 15844 15972
rect 14700 15932 15844 15960
rect 14700 15920 14706 15932
rect 15838 15920 15844 15932
rect 15896 15960 15902 15972
rect 16040 15960 16068 15991
rect 16758 15988 16764 16040
rect 16816 16028 16822 16040
rect 16853 16031 16911 16037
rect 16853 16028 16865 16031
rect 16816 16000 16865 16028
rect 16816 15988 16822 16000
rect 16853 15997 16865 16000
rect 16899 16028 16911 16031
rect 17862 16028 17868 16040
rect 16899 16000 17868 16028
rect 16899 15997 16911 16000
rect 16853 15991 16911 15997
rect 17862 15988 17868 16000
rect 17920 16028 17926 16040
rect 18325 16031 18383 16037
rect 18325 16028 18337 16031
rect 17920 16000 18337 16028
rect 17920 15988 17926 16000
rect 18325 15997 18337 16000
rect 18371 16028 18383 16031
rect 18432 16028 18460 16204
rect 21085 16201 21097 16204
rect 21131 16232 21143 16235
rect 21266 16232 21272 16244
rect 21131 16204 21272 16232
rect 21131 16201 21143 16204
rect 21085 16195 21143 16201
rect 21266 16192 21272 16204
rect 21324 16192 21330 16244
rect 21818 16192 21824 16244
rect 21876 16232 21882 16244
rect 23382 16232 23388 16244
rect 21876 16204 22829 16232
rect 23343 16204 23388 16232
rect 21876 16192 21882 16204
rect 18690 16124 18696 16176
rect 18748 16164 18754 16176
rect 19153 16167 19211 16173
rect 19153 16164 19165 16167
rect 18748 16136 19165 16164
rect 18748 16124 18754 16136
rect 19153 16133 19165 16136
rect 19199 16164 19211 16167
rect 20254 16164 20260 16176
rect 19199 16136 20260 16164
rect 19199 16133 19211 16136
rect 19153 16127 19211 16133
rect 20254 16124 20260 16136
rect 20312 16124 20318 16176
rect 22281 16167 22339 16173
rect 22281 16164 22293 16167
rect 20548 16136 22293 16164
rect 20548 16108 20576 16136
rect 22281 16133 22293 16136
rect 22327 16164 22339 16167
rect 22373 16167 22431 16173
rect 22373 16164 22385 16167
rect 22327 16136 22385 16164
rect 22327 16133 22339 16136
rect 22281 16127 22339 16133
rect 22373 16133 22385 16136
rect 22419 16133 22431 16167
rect 22373 16127 22431 16133
rect 19521 16099 19579 16105
rect 19521 16096 19533 16099
rect 18524 16068 19533 16096
rect 18524 16037 18552 16068
rect 19521 16065 19533 16068
rect 19567 16065 19579 16099
rect 20070 16096 20076 16108
rect 20031 16068 20076 16096
rect 19521 16059 19579 16065
rect 20070 16056 20076 16068
rect 20128 16056 20134 16108
rect 20530 16096 20536 16108
rect 20491 16068 20536 16096
rect 20530 16056 20536 16068
rect 20588 16056 20594 16108
rect 22097 16099 22155 16105
rect 22097 16096 22109 16099
rect 21627 16068 22109 16096
rect 18371 16000 18460 16028
rect 18509 16031 18567 16037
rect 18371 15997 18383 16000
rect 18325 15991 18383 15997
rect 18509 15997 18521 16031
rect 18555 15997 18567 16031
rect 18509 15991 18567 15997
rect 15896 15932 16068 15960
rect 15896 15920 15902 15932
rect 17954 15920 17960 15972
rect 18012 15960 18018 15972
rect 18524 15960 18552 15991
rect 19426 15988 19432 16040
rect 19484 16028 19490 16040
rect 21627 16037 21655 16068
rect 22097 16065 22109 16068
rect 22143 16096 22155 16099
rect 22801 16096 22829 16204
rect 23382 16192 23388 16204
rect 23440 16192 23446 16244
rect 25593 16167 25651 16173
rect 25593 16133 25605 16167
rect 25639 16164 25651 16167
rect 27614 16164 27620 16176
rect 25639 16136 27620 16164
rect 25639 16133 25651 16136
rect 25593 16127 25651 16133
rect 27614 16124 27620 16136
rect 27672 16124 27678 16176
rect 22143 16068 22738 16096
rect 22801 16068 25452 16096
rect 22143 16065 22155 16068
rect 22097 16059 22155 16065
rect 19797 16031 19855 16037
rect 19797 16028 19809 16031
rect 19484 16000 19809 16028
rect 19484 15988 19490 16000
rect 19797 15997 19809 16000
rect 19843 15997 19855 16031
rect 19797 15991 19855 15997
rect 21612 16031 21670 16037
rect 21612 15997 21624 16031
rect 21658 15997 21670 16031
rect 21612 15991 21670 15997
rect 22281 16031 22339 16037
rect 22281 15997 22293 16031
rect 22327 16028 22339 16031
rect 22592 16031 22650 16037
rect 22592 16028 22604 16031
rect 22327 16000 22604 16028
rect 22327 15997 22339 16000
rect 22281 15991 22339 15997
rect 22592 15997 22604 16000
rect 22638 15997 22650 16031
rect 22710 16028 22738 16068
rect 23934 16028 23940 16040
rect 22710 16000 23796 16028
rect 23895 16000 23940 16028
rect 22592 15991 22650 15997
rect 18012 15932 18552 15960
rect 18785 15963 18843 15969
rect 18012 15920 18018 15932
rect 18785 15929 18797 15963
rect 18831 15960 18843 15963
rect 18874 15960 18880 15972
rect 18831 15932 18880 15960
rect 18831 15929 18843 15932
rect 18785 15923 18843 15929
rect 18874 15920 18880 15932
rect 18932 15920 18938 15972
rect 10134 15892 10140 15904
rect 10095 15864 10140 15892
rect 10134 15852 10140 15864
rect 10192 15852 10198 15904
rect 12618 15892 12624 15904
rect 12579 15864 12624 15892
rect 12618 15852 12624 15864
rect 12676 15852 12682 15904
rect 15286 15892 15292 15904
rect 15247 15864 15292 15892
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 19812 15892 19840 15991
rect 20165 15963 20223 15969
rect 20165 15929 20177 15963
rect 20211 15929 20223 15963
rect 20165 15923 20223 15929
rect 20180 15892 20208 15923
rect 20898 15920 20904 15972
rect 20956 15960 20962 15972
rect 21358 15960 21364 15972
rect 20956 15932 21364 15960
rect 20956 15920 20962 15932
rect 21358 15920 21364 15932
rect 21416 15920 21422 15972
rect 22695 15963 22753 15969
rect 22695 15929 22707 15963
rect 22741 15960 22753 15963
rect 23566 15960 23572 15972
rect 22741 15932 23572 15960
rect 22741 15929 22753 15932
rect 22695 15923 22753 15929
rect 23566 15920 23572 15932
rect 23624 15920 23630 15972
rect 23768 15960 23796 16000
rect 23934 15988 23940 16000
rect 23992 15988 23998 16040
rect 25424 16037 25452 16068
rect 25409 16031 25467 16037
rect 25409 15997 25421 16031
rect 25455 16028 25467 16031
rect 25961 16031 26019 16037
rect 25961 16028 25973 16031
rect 25455 16000 25973 16028
rect 25455 15997 25467 16000
rect 25409 15991 25467 15997
rect 25961 15997 25973 16000
rect 26007 15997 26019 16031
rect 25961 15991 26019 15997
rect 24578 15960 24584 15972
rect 23768 15932 24584 15960
rect 24578 15920 24584 15932
rect 24636 15920 24642 15972
rect 19812 15864 20208 15892
rect 21683 15895 21741 15901
rect 21683 15861 21695 15895
rect 21729 15892 21741 15895
rect 22554 15892 22560 15904
rect 21729 15864 22560 15892
rect 21729 15861 21741 15864
rect 21683 15855 21741 15861
rect 22554 15852 22560 15864
rect 22612 15852 22618 15904
rect 24026 15852 24032 15904
rect 24084 15892 24090 15904
rect 24121 15895 24179 15901
rect 24121 15892 24133 15895
rect 24084 15864 24133 15892
rect 24084 15852 24090 15864
rect 24121 15861 24133 15864
rect 24167 15861 24179 15895
rect 24121 15855 24179 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 9030 15648 9036 15700
rect 9088 15688 9094 15700
rect 9861 15691 9919 15697
rect 9861 15688 9873 15691
rect 9088 15660 9873 15688
rect 9088 15648 9094 15660
rect 9861 15657 9873 15660
rect 9907 15657 9919 15691
rect 9861 15651 9919 15657
rect 12621 15691 12679 15697
rect 12621 15657 12633 15691
rect 12667 15688 12679 15691
rect 12986 15688 12992 15700
rect 12667 15660 12992 15688
rect 12667 15657 12679 15660
rect 12621 15651 12679 15657
rect 12986 15648 12992 15660
rect 13044 15688 13050 15700
rect 14185 15691 14243 15697
rect 14185 15688 14197 15691
rect 13044 15660 14197 15688
rect 13044 15648 13050 15660
rect 14185 15657 14197 15660
rect 14231 15657 14243 15691
rect 14185 15651 14243 15657
rect 16209 15691 16267 15697
rect 16209 15657 16221 15691
rect 16255 15688 16267 15691
rect 16942 15688 16948 15700
rect 16255 15660 16948 15688
rect 16255 15657 16267 15660
rect 16209 15651 16267 15657
rect 16942 15648 16948 15660
rect 17000 15688 17006 15700
rect 17221 15691 17279 15697
rect 17221 15688 17233 15691
rect 17000 15660 17233 15688
rect 17000 15648 17006 15660
rect 17221 15657 17233 15660
rect 17267 15657 17279 15691
rect 19150 15688 19156 15700
rect 19111 15660 19156 15688
rect 17221 15651 17279 15657
rect 19150 15648 19156 15660
rect 19208 15648 19214 15700
rect 19978 15688 19984 15700
rect 19939 15660 19984 15688
rect 19978 15648 19984 15660
rect 20036 15648 20042 15700
rect 22094 15688 22100 15700
rect 22007 15660 22100 15688
rect 22094 15648 22100 15660
rect 22152 15688 22158 15700
rect 22462 15688 22468 15700
rect 22152 15660 22468 15688
rect 22152 15648 22158 15660
rect 22462 15648 22468 15660
rect 22520 15648 22526 15700
rect 23382 15688 23388 15700
rect 23295 15660 23388 15688
rect 23382 15648 23388 15660
rect 23440 15688 23446 15700
rect 23934 15688 23940 15700
rect 23440 15660 23940 15688
rect 23440 15648 23446 15660
rect 23934 15648 23940 15660
rect 23992 15688 23998 15700
rect 23992 15660 24440 15688
rect 23992 15648 23998 15660
rect 11241 15623 11299 15629
rect 11241 15589 11253 15623
rect 11287 15620 11299 15623
rect 11422 15620 11428 15632
rect 11287 15592 11428 15620
rect 11287 15589 11299 15592
rect 11241 15583 11299 15589
rect 11422 15580 11428 15592
rect 11480 15580 11486 15632
rect 16482 15620 16488 15632
rect 13786 15592 16488 15620
rect 9674 15552 9680 15564
rect 9635 15524 9680 15552
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 13541 15555 13599 15561
rect 13541 15552 13553 15555
rect 13004 15524 13553 15552
rect 11149 15487 11207 15493
rect 11149 15453 11161 15487
rect 11195 15484 11207 15487
rect 11790 15484 11796 15496
rect 11195 15456 11796 15484
rect 11195 15453 11207 15456
rect 11149 15447 11207 15453
rect 11790 15444 11796 15456
rect 11848 15444 11854 15496
rect 11698 15416 11704 15428
rect 11659 15388 11704 15416
rect 11698 15376 11704 15388
rect 11756 15376 11762 15428
rect 10042 15308 10048 15360
rect 10100 15348 10106 15360
rect 10229 15351 10287 15357
rect 10229 15348 10241 15351
rect 10100 15320 10241 15348
rect 10100 15308 10106 15320
rect 10229 15317 10241 15320
rect 10275 15348 10287 15351
rect 10686 15348 10692 15360
rect 10275 15320 10692 15348
rect 10275 15317 10287 15320
rect 10229 15311 10287 15317
rect 10686 15308 10692 15320
rect 10744 15348 10750 15360
rect 11606 15348 11612 15360
rect 10744 15320 11612 15348
rect 10744 15308 10750 15320
rect 11606 15308 11612 15320
rect 11664 15308 11670 15360
rect 12894 15308 12900 15360
rect 12952 15348 12958 15360
rect 13004 15357 13032 15524
rect 13541 15521 13553 15524
rect 13587 15552 13599 15555
rect 13786 15552 13814 15592
rect 16482 15580 16488 15592
rect 16540 15580 16546 15632
rect 21266 15620 21272 15632
rect 21100 15592 21272 15620
rect 13587 15524 13814 15552
rect 13587 15521 13599 15524
rect 13541 15515 13599 15521
rect 15378 15512 15384 15564
rect 15436 15552 15442 15564
rect 15657 15555 15715 15561
rect 15657 15552 15669 15555
rect 15436 15524 15669 15552
rect 15436 15512 15442 15524
rect 15657 15521 15669 15524
rect 15703 15521 15715 15555
rect 15657 15515 15715 15521
rect 16942 15512 16948 15564
rect 17000 15552 17006 15564
rect 21100 15561 21128 15592
rect 21266 15580 21272 15592
rect 21324 15580 21330 15632
rect 22278 15580 22284 15632
rect 22336 15620 22342 15632
rect 24412 15629 24440 15660
rect 22786 15623 22844 15629
rect 22786 15620 22798 15623
rect 22336 15592 22798 15620
rect 22336 15580 22342 15592
rect 22786 15589 22798 15592
rect 22832 15589 22844 15623
rect 22786 15583 22844 15589
rect 24397 15623 24455 15629
rect 24397 15589 24409 15623
rect 24443 15589 24455 15623
rect 24397 15583 24455 15589
rect 17037 15555 17095 15561
rect 17037 15552 17049 15555
rect 17000 15524 17049 15552
rect 17000 15512 17006 15524
rect 17037 15521 17049 15524
rect 17083 15552 17095 15555
rect 17497 15555 17555 15561
rect 17497 15552 17509 15555
rect 17083 15524 17509 15552
rect 17083 15521 17095 15524
rect 17037 15515 17095 15521
rect 17497 15521 17509 15524
rect 17543 15521 17555 15555
rect 17497 15515 17555 15521
rect 21085 15555 21143 15561
rect 21085 15521 21097 15555
rect 21131 15521 21143 15555
rect 21085 15515 21143 15521
rect 21174 15512 21180 15564
rect 21232 15552 21238 15564
rect 21361 15555 21419 15561
rect 21361 15552 21373 15555
rect 21232 15524 21373 15552
rect 21232 15512 21238 15524
rect 21361 15521 21373 15524
rect 21407 15521 21419 15555
rect 21361 15515 21419 15521
rect 13078 15444 13084 15496
rect 13136 15484 13142 15496
rect 13909 15487 13967 15493
rect 13909 15484 13921 15487
rect 13136 15456 13921 15484
rect 13136 15444 13142 15456
rect 13909 15453 13921 15456
rect 13955 15484 13967 15487
rect 15473 15487 15531 15493
rect 15473 15484 15485 15487
rect 13955 15456 15485 15484
rect 13955 15453 13967 15456
rect 13909 15447 13967 15453
rect 15473 15453 15485 15456
rect 15519 15484 15531 15487
rect 15562 15484 15568 15496
rect 15519 15456 15568 15484
rect 15519 15453 15531 15456
rect 15473 15447 15531 15453
rect 15562 15444 15568 15456
rect 15620 15444 15626 15496
rect 18785 15487 18843 15493
rect 18785 15453 18797 15487
rect 18831 15484 18843 15487
rect 18874 15484 18880 15496
rect 18831 15456 18880 15484
rect 18831 15453 18843 15456
rect 18785 15447 18843 15453
rect 18874 15444 18880 15456
rect 18932 15444 18938 15496
rect 21637 15487 21695 15493
rect 21637 15453 21649 15487
rect 21683 15484 21695 15487
rect 22462 15484 22468 15496
rect 21683 15456 22468 15484
rect 21683 15453 21695 15456
rect 21637 15447 21695 15453
rect 22462 15444 22468 15456
rect 22520 15444 22526 15496
rect 24305 15487 24363 15493
rect 24305 15453 24317 15487
rect 24351 15453 24363 15487
rect 24578 15484 24584 15496
rect 24539 15456 24584 15484
rect 24305 15447 24363 15453
rect 15841 15419 15899 15425
rect 15841 15385 15853 15419
rect 15887 15416 15899 15419
rect 16945 15419 17003 15425
rect 16945 15416 16957 15419
rect 15887 15388 16957 15416
rect 15887 15385 15899 15388
rect 15841 15379 15899 15385
rect 16945 15385 16957 15388
rect 16991 15416 17003 15419
rect 17218 15416 17224 15428
rect 16991 15388 17224 15416
rect 16991 15385 17003 15388
rect 16945 15379 17003 15385
rect 17218 15376 17224 15388
rect 17276 15376 17282 15428
rect 24320 15416 24348 15447
rect 24578 15444 24584 15456
rect 24636 15484 24642 15496
rect 24762 15484 24768 15496
rect 24636 15456 24768 15484
rect 24636 15444 24642 15456
rect 24762 15444 24768 15456
rect 24820 15444 24826 15496
rect 24854 15416 24860 15428
rect 24320 15388 24860 15416
rect 24854 15376 24860 15388
rect 24912 15376 24918 15428
rect 12989 15351 13047 15357
rect 12989 15348 13001 15351
rect 12952 15320 13001 15348
rect 12952 15308 12958 15320
rect 12989 15317 13001 15320
rect 13035 15317 13047 15351
rect 13446 15348 13452 15360
rect 13407 15320 13452 15348
rect 12989 15311 13047 15317
rect 13446 15308 13452 15320
rect 13504 15348 13510 15360
rect 13679 15351 13737 15357
rect 13679 15348 13691 15351
rect 13504 15320 13691 15348
rect 13504 15308 13510 15320
rect 13679 15317 13691 15320
rect 13725 15317 13737 15351
rect 13679 15311 13737 15317
rect 13817 15351 13875 15357
rect 13817 15317 13829 15351
rect 13863 15348 13875 15351
rect 13998 15348 14004 15360
rect 13863 15320 14004 15348
rect 13863 15317 13875 15320
rect 13817 15311 13875 15317
rect 13998 15308 14004 15320
rect 14056 15308 14062 15360
rect 14642 15308 14648 15360
rect 14700 15348 14706 15360
rect 15013 15351 15071 15357
rect 15013 15348 15025 15351
rect 14700 15320 15025 15348
rect 14700 15308 14706 15320
rect 15013 15317 15025 15320
rect 15059 15317 15071 15351
rect 18046 15348 18052 15360
rect 18007 15320 18052 15348
rect 15013 15311 15071 15317
rect 18046 15308 18052 15320
rect 18104 15308 18110 15360
rect 18322 15308 18328 15360
rect 18380 15348 18386 15360
rect 18417 15351 18475 15357
rect 18417 15348 18429 15351
rect 18380 15320 18429 15348
rect 18380 15308 18386 15320
rect 18417 15317 18429 15320
rect 18463 15317 18475 15351
rect 18417 15311 18475 15317
rect 19426 15308 19432 15360
rect 19484 15348 19490 15360
rect 19705 15351 19763 15357
rect 19705 15348 19717 15351
rect 19484 15320 19717 15348
rect 19484 15308 19490 15320
rect 19705 15317 19717 15320
rect 19751 15317 19763 15351
rect 19705 15311 19763 15317
rect 19794 15308 19800 15360
rect 19852 15348 19858 15360
rect 22278 15348 22284 15360
rect 19852 15320 22284 15348
rect 19852 15308 19858 15320
rect 22278 15308 22284 15320
rect 22336 15308 22342 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 11422 15144 11428 15156
rect 11383 15116 11428 15144
rect 11422 15104 11428 15116
rect 11480 15104 11486 15156
rect 11790 15144 11796 15156
rect 11751 15116 11796 15144
rect 11790 15104 11796 15116
rect 11848 15144 11854 15156
rect 13906 15144 13912 15156
rect 11848 15116 12480 15144
rect 13867 15116 13912 15144
rect 11848 15104 11854 15116
rect 9766 15036 9772 15088
rect 9824 15076 9830 15088
rect 9953 15079 10011 15085
rect 9953 15076 9965 15079
rect 9824 15048 9965 15076
rect 9824 15036 9830 15048
rect 9953 15045 9965 15048
rect 9999 15076 10011 15079
rect 11149 15079 11207 15085
rect 9999 15048 10593 15076
rect 9999 15045 10011 15048
rect 9953 15039 10011 15045
rect 8573 15011 8631 15017
rect 8573 14977 8585 15011
rect 8619 15008 8631 15011
rect 8619 14980 9260 15008
rect 8619 14977 8631 14980
rect 8573 14971 8631 14977
rect 8941 14943 8999 14949
rect 8941 14909 8953 14943
rect 8987 14940 8999 14943
rect 9030 14940 9036 14952
rect 8987 14912 9036 14940
rect 8987 14909 8999 14912
rect 8941 14903 8999 14909
rect 9030 14900 9036 14912
rect 9088 14900 9094 14952
rect 9232 14949 9260 14980
rect 10134 14968 10140 15020
rect 10192 15008 10198 15020
rect 10229 15011 10287 15017
rect 10229 15008 10241 15011
rect 10192 14980 10241 15008
rect 10192 14968 10198 14980
rect 10229 14977 10241 14980
rect 10275 14977 10287 15011
rect 10229 14971 10287 14977
rect 9217 14943 9275 14949
rect 9217 14909 9229 14943
rect 9263 14940 9275 14943
rect 10042 14940 10048 14952
rect 9263 14912 10048 14940
rect 9263 14909 9275 14912
rect 9217 14903 9275 14909
rect 10042 14900 10048 14912
rect 10100 14900 10106 14952
rect 9398 14872 9404 14884
rect 9359 14844 9404 14872
rect 9398 14832 9404 14844
rect 9456 14832 9462 14884
rect 9674 14832 9680 14884
rect 9732 14872 9738 14884
rect 10565 14881 10593 15048
rect 11149 15045 11161 15079
rect 11195 15076 11207 15079
rect 11514 15076 11520 15088
rect 11195 15048 11520 15076
rect 11195 15045 11207 15048
rect 11149 15039 11207 15045
rect 11514 15036 11520 15048
rect 11572 15036 11578 15088
rect 12452 15017 12480 15116
rect 13906 15104 13912 15116
rect 13964 15104 13970 15156
rect 15470 15144 15476 15156
rect 15431 15116 15476 15144
rect 15470 15104 15476 15116
rect 15528 15104 15534 15156
rect 16758 15144 16764 15156
rect 16719 15116 16764 15144
rect 16758 15104 16764 15116
rect 16816 15104 16822 15156
rect 18046 15104 18052 15156
rect 18104 15144 18110 15156
rect 18325 15147 18383 15153
rect 18325 15144 18337 15147
rect 18104 15116 18337 15144
rect 18104 15104 18110 15116
rect 18325 15113 18337 15116
rect 18371 15113 18383 15147
rect 18325 15107 18383 15113
rect 18693 15147 18751 15153
rect 18693 15113 18705 15147
rect 18739 15144 18751 15147
rect 20806 15144 20812 15156
rect 18739 15116 20812 15144
rect 18739 15113 18751 15116
rect 18693 15107 18751 15113
rect 20806 15104 20812 15116
rect 20864 15104 20870 15156
rect 20993 15147 21051 15153
rect 20993 15113 21005 15147
rect 21039 15144 21051 15147
rect 21266 15144 21272 15156
rect 21039 15116 21272 15144
rect 21039 15113 21051 15116
rect 20993 15107 21051 15113
rect 21266 15104 21272 15116
rect 21324 15104 21330 15156
rect 23382 15144 23388 15156
rect 23343 15116 23388 15144
rect 23382 15104 23388 15116
rect 23440 15104 23446 15156
rect 24026 15144 24032 15156
rect 23987 15116 24032 15144
rect 24026 15104 24032 15116
rect 24084 15104 24090 15156
rect 24854 15104 24860 15156
rect 24912 15144 24918 15156
rect 25225 15147 25283 15153
rect 25225 15144 25237 15147
rect 24912 15116 25237 15144
rect 24912 15104 24918 15116
rect 25225 15113 25237 15116
rect 25271 15113 25283 15147
rect 25225 15107 25283 15113
rect 12989 15079 13047 15085
rect 12989 15045 13001 15079
rect 13035 15076 13047 15079
rect 13725 15079 13783 15085
rect 13725 15076 13737 15079
rect 13035 15048 13737 15076
rect 13035 15045 13047 15048
rect 12989 15039 13047 15045
rect 13725 15045 13737 15048
rect 13771 15076 13783 15079
rect 13998 15076 14004 15088
rect 13771 15048 14004 15076
rect 13771 15045 13783 15048
rect 13725 15039 13783 15045
rect 13998 15036 14004 15048
rect 14056 15076 14062 15088
rect 14737 15079 14795 15085
rect 14737 15076 14749 15079
rect 14056 15048 14749 15076
rect 14056 15036 14062 15048
rect 14737 15045 14749 15048
rect 14783 15076 14795 15079
rect 15289 15079 15347 15085
rect 15289 15076 15301 15079
rect 14783 15048 15301 15076
rect 14783 15045 14795 15048
rect 14737 15039 14795 15045
rect 15289 15045 15301 15048
rect 15335 15045 15347 15079
rect 19150 15076 19156 15088
rect 19063 15048 19156 15076
rect 15289 15039 15347 15045
rect 19150 15036 19156 15048
rect 19208 15076 19214 15088
rect 19794 15076 19800 15088
rect 19208 15048 19800 15076
rect 19208 15036 19214 15048
rect 19794 15036 19800 15048
rect 19852 15036 19858 15088
rect 20530 15076 20536 15088
rect 20491 15048 20536 15076
rect 20530 15036 20536 15048
rect 20588 15036 20594 15088
rect 12437 15011 12495 15017
rect 12437 14977 12449 15011
rect 12483 14977 12495 15011
rect 12437 14971 12495 14977
rect 13446 14968 13452 15020
rect 13504 15008 13510 15020
rect 13596 15011 13654 15017
rect 13596 15008 13608 15011
rect 13504 14980 13608 15008
rect 13504 14968 13510 14980
rect 13596 14977 13608 14980
rect 13642 14977 13654 15011
rect 13814 15008 13820 15020
rect 13775 14980 13820 15008
rect 13596 14971 13654 14977
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 15010 14968 15016 15020
rect 15068 15008 15074 15020
rect 15160 15011 15218 15017
rect 15160 15008 15172 15011
rect 15068 14980 15172 15008
rect 15068 14968 15074 14980
rect 15160 14977 15172 14980
rect 15206 14977 15218 15011
rect 15160 14971 15218 14977
rect 15381 15011 15439 15017
rect 15381 14977 15393 15011
rect 15427 15008 15439 15011
rect 15562 15008 15568 15020
rect 15427 14980 15568 15008
rect 15427 14977 15439 14980
rect 15381 14971 15439 14977
rect 15562 14968 15568 14980
rect 15620 14968 15626 15020
rect 15838 14968 15844 15020
rect 15896 15008 15902 15020
rect 17405 15011 17463 15017
rect 17405 15008 17417 15011
rect 15896 14980 17417 15008
rect 15896 14968 15902 14980
rect 17405 14977 17417 14980
rect 17451 15008 17463 15011
rect 18414 15008 18420 15020
rect 17451 14980 18420 15008
rect 17451 14977 17463 14980
rect 17405 14971 17463 14977
rect 18414 14968 18420 14980
rect 18472 14968 18478 15020
rect 19978 15008 19984 15020
rect 19939 14980 19984 15008
rect 19978 14968 19984 14980
rect 20036 14968 20042 15020
rect 22094 15008 22100 15020
rect 22055 14980 22100 15008
rect 22094 14968 22100 14980
rect 22152 14968 22158 15020
rect 22370 15008 22376 15020
rect 22331 14980 22376 15008
rect 22370 14968 22376 14980
rect 22428 14968 22434 15020
rect 24302 15008 24308 15020
rect 24215 14980 24308 15008
rect 24302 14968 24308 14980
rect 24360 15008 24366 15020
rect 24670 15008 24676 15020
rect 24360 14980 24676 15008
rect 24360 14968 24366 14980
rect 24670 14968 24676 14980
rect 24728 14968 24734 15020
rect 24762 14968 24768 15020
rect 24820 15008 24826 15020
rect 24820 14980 24865 15008
rect 24820 14968 24826 14980
rect 12250 14940 12256 14952
rect 12163 14912 12256 14940
rect 12250 14900 12256 14912
rect 12308 14940 12314 14952
rect 13078 14940 13084 14952
rect 12308 14912 13084 14940
rect 12308 14900 12314 14912
rect 13078 14900 13084 14912
rect 13136 14900 13142 14952
rect 15286 14900 15292 14952
rect 15344 14940 15350 14952
rect 16577 14943 16635 14949
rect 16577 14940 16589 14943
rect 15344 14912 16589 14940
rect 15344 14900 15350 14912
rect 16577 14909 16589 14912
rect 16623 14940 16635 14943
rect 17037 14943 17095 14949
rect 17037 14940 17049 14943
rect 16623 14912 17049 14940
rect 16623 14909 16635 14912
rect 16577 14903 16635 14909
rect 17037 14909 17049 14912
rect 17083 14909 17095 14943
rect 17037 14903 17095 14909
rect 18196 14943 18254 14949
rect 18196 14909 18208 14943
rect 18242 14940 18254 14943
rect 18322 14940 18328 14952
rect 18242 14912 18328 14940
rect 18242 14909 18254 14912
rect 18196 14903 18254 14909
rect 18322 14900 18328 14912
rect 18380 14900 18386 14952
rect 9769 14875 9827 14881
rect 9769 14872 9781 14875
rect 9732 14844 9781 14872
rect 9732 14832 9738 14844
rect 9769 14841 9781 14844
rect 9815 14872 9827 14875
rect 10550 14875 10608 14881
rect 9815 14844 10180 14872
rect 9815 14841 9827 14844
rect 9769 14835 9827 14841
rect 9953 14807 10011 14813
rect 9953 14773 9965 14807
rect 9999 14804 10011 14807
rect 10042 14804 10048 14816
rect 9999 14776 10048 14804
rect 9999 14773 10011 14776
rect 9953 14767 10011 14773
rect 10042 14764 10048 14776
rect 10100 14764 10106 14816
rect 10152 14804 10180 14844
rect 10550 14841 10562 14875
rect 10596 14841 10608 14875
rect 10550 14835 10608 14841
rect 12894 14832 12900 14884
rect 12952 14872 12958 14884
rect 13449 14875 13507 14881
rect 13449 14872 13461 14875
rect 12952 14844 13461 14872
rect 12952 14832 12958 14844
rect 13449 14841 13461 14844
rect 13495 14841 13507 14875
rect 13449 14835 13507 14841
rect 14642 14832 14648 14884
rect 14700 14872 14706 14884
rect 15013 14875 15071 14881
rect 15013 14872 15025 14875
rect 14700 14844 15025 14872
rect 14700 14832 14706 14844
rect 15013 14841 15025 14844
rect 15059 14841 15071 14875
rect 15013 14835 15071 14841
rect 15378 14832 15384 14884
rect 15436 14872 15442 14884
rect 16025 14875 16083 14881
rect 16025 14872 16037 14875
rect 15436 14844 16037 14872
rect 15436 14832 15442 14844
rect 16025 14841 16037 14844
rect 16071 14841 16083 14875
rect 18049 14875 18107 14881
rect 18049 14872 18061 14875
rect 16025 14835 16083 14841
rect 17788 14844 18061 14872
rect 17788 14816 17816 14844
rect 18049 14841 18061 14844
rect 18095 14841 18107 14875
rect 18049 14835 18107 14841
rect 20073 14875 20131 14881
rect 20073 14841 20085 14875
rect 20119 14841 20131 14875
rect 20073 14835 20131 14841
rect 22189 14875 22247 14881
rect 22189 14841 22201 14875
rect 22235 14841 22247 14875
rect 22189 14835 22247 14841
rect 24397 14875 24455 14881
rect 24397 14841 24409 14875
rect 24443 14841 24455 14875
rect 24397 14835 24455 14841
rect 10778 14804 10784 14816
rect 10152 14776 10784 14804
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 13357 14807 13415 14813
rect 13357 14773 13369 14807
rect 13403 14804 13415 14807
rect 13814 14804 13820 14816
rect 13403 14776 13820 14804
rect 13403 14773 13415 14776
rect 13357 14767 13415 14773
rect 13814 14764 13820 14776
rect 13872 14764 13878 14816
rect 14550 14804 14556 14816
rect 14511 14776 14556 14804
rect 14550 14764 14556 14776
rect 14608 14804 14614 14816
rect 14737 14807 14795 14813
rect 14737 14804 14749 14807
rect 14608 14776 14749 14804
rect 14608 14764 14614 14776
rect 14737 14773 14749 14776
rect 14783 14804 14795 14807
rect 14829 14807 14887 14813
rect 14829 14804 14841 14807
rect 14783 14776 14841 14804
rect 14783 14773 14795 14776
rect 14737 14767 14795 14773
rect 14829 14773 14841 14776
rect 14875 14773 14887 14807
rect 16482 14804 16488 14816
rect 16443 14776 16488 14804
rect 14829 14767 14887 14773
rect 16482 14764 16488 14776
rect 16540 14764 16546 14816
rect 17770 14804 17776 14816
rect 17731 14776 17776 14804
rect 17770 14764 17776 14776
rect 17828 14764 17834 14816
rect 19518 14764 19524 14816
rect 19576 14804 19582 14816
rect 19705 14807 19763 14813
rect 19705 14804 19717 14807
rect 19576 14776 19717 14804
rect 19576 14764 19582 14776
rect 19705 14773 19717 14776
rect 19751 14804 19763 14807
rect 20088 14804 20116 14835
rect 19751 14776 20116 14804
rect 19751 14773 19763 14776
rect 19705 14767 19763 14773
rect 21174 14764 21180 14816
rect 21232 14804 21238 14816
rect 21269 14807 21327 14813
rect 21269 14804 21281 14807
rect 21232 14776 21281 14804
rect 21232 14764 21238 14776
rect 21269 14773 21281 14776
rect 21315 14773 21327 14807
rect 21910 14804 21916 14816
rect 21871 14776 21916 14804
rect 21269 14767 21327 14773
rect 21910 14764 21916 14776
rect 21968 14804 21974 14816
rect 22204 14804 22232 14835
rect 21968 14776 22232 14804
rect 21968 14764 21974 14776
rect 22278 14764 22284 14816
rect 22336 14804 22342 14816
rect 23017 14807 23075 14813
rect 23017 14804 23029 14807
rect 22336 14776 23029 14804
rect 22336 14764 22342 14776
rect 23017 14773 23029 14776
rect 23063 14773 23075 14807
rect 23017 14767 23075 14773
rect 24026 14764 24032 14816
rect 24084 14804 24090 14816
rect 24412 14804 24440 14835
rect 24084 14776 24440 14804
rect 24084 14764 24090 14776
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 8757 14603 8815 14609
rect 8757 14569 8769 14603
rect 8803 14600 8815 14603
rect 9030 14600 9036 14612
rect 8803 14572 9036 14600
rect 8803 14569 8815 14572
rect 8757 14563 8815 14569
rect 9030 14560 9036 14572
rect 9088 14560 9094 14612
rect 10134 14560 10140 14612
rect 10192 14600 10198 14612
rect 10229 14603 10287 14609
rect 10229 14600 10241 14603
rect 10192 14572 10241 14600
rect 10192 14560 10198 14572
rect 10229 14569 10241 14572
rect 10275 14569 10287 14603
rect 12894 14600 12900 14612
rect 12855 14572 12900 14600
rect 10229 14563 10287 14569
rect 12894 14560 12900 14572
rect 12952 14560 12958 14612
rect 14461 14603 14519 14609
rect 14461 14569 14473 14603
rect 14507 14600 14519 14603
rect 14826 14600 14832 14612
rect 14507 14572 14832 14600
rect 14507 14569 14519 14572
rect 14461 14563 14519 14569
rect 14826 14560 14832 14572
rect 14884 14600 14890 14612
rect 15010 14600 15016 14612
rect 14884 14572 15016 14600
rect 14884 14560 14890 14572
rect 15010 14560 15016 14572
rect 15068 14560 15074 14612
rect 15562 14560 15568 14612
rect 15620 14600 15626 14612
rect 16393 14603 16451 14609
rect 16393 14600 16405 14603
rect 15620 14572 16405 14600
rect 15620 14560 15626 14572
rect 16393 14569 16405 14572
rect 16439 14600 16451 14603
rect 18509 14603 18567 14609
rect 18509 14600 18521 14603
rect 16439 14572 18521 14600
rect 16439 14569 16451 14572
rect 16393 14563 16451 14569
rect 11241 14535 11299 14541
rect 11241 14501 11253 14535
rect 11287 14532 11299 14535
rect 11514 14532 11520 14544
rect 11287 14504 11520 14532
rect 11287 14501 11299 14504
rect 11241 14495 11299 14501
rect 11514 14492 11520 14504
rect 11572 14492 11578 14544
rect 11606 14492 11612 14544
rect 11664 14532 11670 14544
rect 14093 14535 14151 14541
rect 14093 14532 14105 14535
rect 11664 14504 14105 14532
rect 11664 14492 11670 14504
rect 14093 14501 14105 14504
rect 14139 14501 14151 14535
rect 14093 14495 14151 14501
rect 13265 14467 13323 14473
rect 13265 14433 13277 14467
rect 13311 14464 13323 14467
rect 13357 14467 13415 14473
rect 13357 14464 13369 14467
rect 13311 14436 13369 14464
rect 13311 14433 13323 14436
rect 13265 14427 13323 14433
rect 13357 14433 13369 14436
rect 13403 14433 13415 14467
rect 15378 14464 15384 14476
rect 15339 14436 15384 14464
rect 13357 14427 13415 14433
rect 11149 14399 11207 14405
rect 11149 14365 11161 14399
rect 11195 14396 11207 14399
rect 11330 14396 11336 14408
rect 11195 14368 11336 14396
rect 11195 14365 11207 14368
rect 11149 14359 11207 14365
rect 11330 14356 11336 14368
rect 11388 14356 11394 14408
rect 11698 14328 11704 14340
rect 11659 14300 11704 14328
rect 11698 14288 11704 14300
rect 11756 14288 11762 14340
rect 13262 14288 13268 14340
rect 13320 14328 13326 14340
rect 13372 14328 13400 14427
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 17129 14467 17187 14473
rect 17129 14433 17141 14467
rect 17175 14433 17187 14467
rect 17129 14427 17187 14433
rect 13725 14399 13783 14405
rect 13725 14365 13737 14399
rect 13771 14396 13783 14399
rect 13814 14396 13820 14408
rect 13771 14368 13820 14396
rect 13771 14365 13783 14368
rect 13725 14359 13783 14365
rect 13814 14356 13820 14368
rect 13872 14356 13878 14408
rect 15286 14396 15292 14408
rect 15247 14368 15292 14396
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 14642 14328 14648 14340
rect 13320 14300 14648 14328
rect 13320 14288 13326 14300
rect 14642 14288 14648 14300
rect 14700 14288 14706 14340
rect 17037 14331 17095 14337
rect 17037 14297 17049 14331
rect 17083 14328 17095 14331
rect 17144 14328 17172 14427
rect 17512 14405 17540 14572
rect 18509 14569 18521 14572
rect 18555 14569 18567 14603
rect 18874 14600 18880 14612
rect 18835 14572 18880 14600
rect 18509 14563 18567 14569
rect 18874 14560 18880 14572
rect 18932 14560 18938 14612
rect 19518 14600 19524 14612
rect 19479 14572 19524 14600
rect 19518 14560 19524 14572
rect 19576 14560 19582 14612
rect 22462 14600 22468 14612
rect 22423 14572 22468 14600
rect 22462 14560 22468 14572
rect 22520 14560 22526 14612
rect 24302 14600 24308 14612
rect 24263 14572 24308 14600
rect 24302 14560 24308 14572
rect 24360 14560 24366 14612
rect 17865 14535 17923 14541
rect 17865 14501 17877 14535
rect 17911 14532 17923 14535
rect 21174 14532 21180 14544
rect 17911 14504 21180 14532
rect 17911 14501 17923 14504
rect 17865 14495 17923 14501
rect 21174 14492 21180 14504
rect 21232 14492 21238 14544
rect 21453 14535 21511 14541
rect 21453 14501 21465 14535
rect 21499 14532 21511 14535
rect 21818 14532 21824 14544
rect 21499 14504 21824 14532
rect 21499 14501 21511 14504
rect 21453 14495 21511 14501
rect 21818 14492 21824 14504
rect 21876 14492 21882 14544
rect 22005 14535 22063 14541
rect 22005 14501 22017 14535
rect 22051 14532 22063 14535
rect 22370 14532 22376 14544
rect 22051 14504 22376 14532
rect 22051 14501 22063 14504
rect 22005 14495 22063 14501
rect 22370 14492 22376 14504
rect 22428 14492 22434 14544
rect 19518 14464 19524 14476
rect 19479 14436 19524 14464
rect 19518 14424 19524 14436
rect 19576 14424 19582 14476
rect 22922 14464 22928 14476
rect 22883 14436 22928 14464
rect 22922 14424 22928 14436
rect 22980 14424 22986 14476
rect 23566 14424 23572 14476
rect 23624 14464 23630 14476
rect 24581 14467 24639 14473
rect 24581 14464 24593 14467
rect 23624 14436 24593 14464
rect 23624 14424 23630 14436
rect 24581 14433 24593 14436
rect 24627 14464 24639 14467
rect 24670 14464 24676 14476
rect 24627 14436 24676 14464
rect 24627 14433 24639 14436
rect 24581 14427 24639 14433
rect 24670 14424 24676 14436
rect 24728 14424 24734 14476
rect 17497 14399 17555 14405
rect 17497 14365 17509 14399
rect 17543 14365 17555 14399
rect 17497 14359 17555 14365
rect 20346 14356 20352 14408
rect 20404 14396 20410 14408
rect 21361 14399 21419 14405
rect 21361 14396 21373 14399
rect 20404 14368 21373 14396
rect 20404 14356 20410 14368
rect 21361 14365 21373 14368
rect 21407 14365 21419 14399
rect 21361 14359 21419 14365
rect 17862 14328 17868 14340
rect 17083 14300 17868 14328
rect 17083 14297 17095 14300
rect 17037 14291 17095 14297
rect 17862 14288 17868 14300
rect 17920 14288 17926 14340
rect 24762 14328 24768 14340
rect 24723 14300 24768 14328
rect 24762 14288 24768 14300
rect 24820 14288 24826 14340
rect 13446 14220 13452 14272
rect 13504 14269 13510 14272
rect 13504 14263 13553 14269
rect 13504 14229 13507 14263
rect 13541 14229 13553 14263
rect 13504 14223 13553 14229
rect 13633 14263 13691 14269
rect 13633 14229 13645 14263
rect 13679 14260 13691 14263
rect 14550 14260 14556 14272
rect 13679 14232 14556 14260
rect 13679 14229 13691 14232
rect 13633 14223 13691 14229
rect 13504 14220 13510 14223
rect 14550 14220 14556 14232
rect 14608 14220 14614 14272
rect 16482 14220 16488 14272
rect 16540 14260 16546 14272
rect 17267 14263 17325 14269
rect 17267 14260 17279 14263
rect 16540 14232 17279 14260
rect 16540 14220 16546 14232
rect 17267 14229 17279 14232
rect 17313 14229 17325 14263
rect 17402 14260 17408 14272
rect 17363 14232 17408 14260
rect 17267 14223 17325 14229
rect 17402 14220 17408 14232
rect 17460 14220 17466 14272
rect 18046 14220 18052 14272
rect 18104 14260 18110 14272
rect 18141 14263 18199 14269
rect 18141 14260 18153 14263
rect 18104 14232 18153 14260
rect 18104 14220 18110 14232
rect 18141 14229 18153 14232
rect 18187 14229 18199 14263
rect 23290 14260 23296 14272
rect 23251 14232 23296 14260
rect 18141 14223 18199 14229
rect 23290 14220 23296 14232
rect 23348 14220 23354 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 9309 14059 9367 14065
rect 9309 14025 9321 14059
rect 9355 14056 9367 14059
rect 9398 14056 9404 14068
rect 9355 14028 9404 14056
rect 9355 14025 9367 14028
rect 9309 14019 9367 14025
rect 9398 14016 9404 14028
rect 9456 14016 9462 14068
rect 9677 14059 9735 14065
rect 9677 14025 9689 14059
rect 9723 14056 9735 14059
rect 10042 14056 10048 14068
rect 9723 14028 10048 14056
rect 9723 14025 9735 14028
rect 9677 14019 9735 14025
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 11149 14059 11207 14065
rect 11149 14025 11161 14059
rect 11195 14056 11207 14059
rect 11514 14056 11520 14068
rect 11195 14028 11520 14056
rect 11195 14025 11207 14028
rect 11149 14019 11207 14025
rect 11514 14016 11520 14028
rect 11572 14016 11578 14068
rect 13446 14016 13452 14068
rect 13504 14056 13510 14068
rect 13614 14059 13672 14065
rect 13614 14056 13626 14059
rect 13504 14028 13626 14056
rect 13504 14016 13510 14028
rect 13614 14025 13626 14028
rect 13660 14056 13672 14059
rect 14826 14056 14832 14068
rect 13660 14028 14832 14056
rect 13660 14025 13672 14028
rect 13614 14019 13672 14025
rect 14826 14016 14832 14028
rect 14884 14016 14890 14068
rect 15378 14016 15384 14068
rect 15436 14056 15442 14068
rect 15841 14059 15899 14065
rect 15841 14056 15853 14059
rect 15436 14028 15853 14056
rect 15436 14016 15442 14028
rect 15841 14025 15853 14028
rect 15887 14025 15899 14059
rect 15841 14019 15899 14025
rect 16206 14016 16212 14068
rect 16264 14056 16270 14068
rect 16669 14059 16727 14065
rect 16669 14056 16681 14059
rect 16264 14028 16681 14056
rect 16264 14016 16270 14028
rect 16669 14025 16681 14028
rect 16715 14056 16727 14059
rect 17402 14056 17408 14068
rect 16715 14028 17408 14056
rect 16715 14025 16727 14028
rect 16669 14019 16727 14025
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 18046 14056 18052 14068
rect 17959 14028 18052 14056
rect 18046 14016 18052 14028
rect 18104 14056 18110 14068
rect 18325 14059 18383 14065
rect 18325 14056 18337 14059
rect 18104 14028 18337 14056
rect 18104 14016 18110 14028
rect 18325 14025 18337 14028
rect 18371 14025 18383 14059
rect 19518 14056 19524 14068
rect 19479 14028 19524 14056
rect 18325 14019 18383 14025
rect 19518 14016 19524 14028
rect 19576 14016 19582 14068
rect 20346 14016 20352 14068
rect 20404 14056 20410 14068
rect 20533 14059 20591 14065
rect 20533 14056 20545 14059
rect 20404 14028 20545 14056
rect 20404 14016 20410 14028
rect 20533 14025 20545 14028
rect 20579 14025 20591 14059
rect 21910 14056 21916 14068
rect 21871 14028 21916 14056
rect 20533 14019 20591 14025
rect 21910 14016 21916 14028
rect 21968 14016 21974 14068
rect 22922 14056 22928 14068
rect 22883 14028 22928 14056
rect 22922 14016 22928 14028
rect 22980 14016 22986 14068
rect 23290 14016 23296 14068
rect 23348 14056 23354 14068
rect 23385 14059 23443 14065
rect 23385 14056 23397 14059
rect 23348 14028 23397 14056
rect 23348 14016 23354 14028
rect 23385 14025 23397 14028
rect 23431 14025 23443 14059
rect 24670 14056 24676 14068
rect 24631 14028 24676 14056
rect 23385 14019 23443 14025
rect 24670 14016 24676 14028
rect 24728 14016 24734 14068
rect 25406 14056 25412 14068
rect 25367 14028 25412 14056
rect 25406 14016 25412 14028
rect 25464 14016 25470 14068
rect 9416 13920 9444 14016
rect 12989 13991 13047 13997
rect 12989 13957 13001 13991
rect 13035 13988 13047 13991
rect 13357 13991 13415 13997
rect 13357 13988 13369 13991
rect 13035 13960 13369 13988
rect 13035 13957 13047 13960
rect 12989 13951 13047 13957
rect 13357 13957 13369 13960
rect 13403 13988 13415 13991
rect 13403 13960 13676 13988
rect 13403 13957 13415 13960
rect 13357 13951 13415 13957
rect 9769 13923 9827 13929
rect 9769 13920 9781 13923
rect 9416 13892 9781 13920
rect 9769 13889 9781 13892
rect 9815 13889 9827 13923
rect 13648 13920 13676 13960
rect 13722 13948 13728 14000
rect 13780 13988 13786 14000
rect 13780 13960 13825 13988
rect 13780 13948 13786 13960
rect 14642 13948 14648 14000
rect 14700 13988 14706 14000
rect 15197 13991 15255 13997
rect 15197 13988 15209 13991
rect 14700 13960 15209 13988
rect 14700 13948 14706 13960
rect 15197 13957 15209 13960
rect 15243 13957 15255 13991
rect 15562 13988 15568 14000
rect 15523 13960 15568 13988
rect 15197 13951 15255 13957
rect 15562 13948 15568 13960
rect 15620 13948 15626 14000
rect 16482 13948 16488 14000
rect 16540 13997 16546 14000
rect 16540 13991 16589 13997
rect 16540 13957 16543 13991
rect 16577 13957 16589 13991
rect 16540 13951 16589 13957
rect 16540 13948 16546 13951
rect 17126 13948 17132 14000
rect 17184 13988 17190 14000
rect 18064 13988 18092 14016
rect 17184 13960 18092 13988
rect 17184 13948 17190 13960
rect 13814 13920 13820 13932
rect 13648 13892 13820 13920
rect 9769 13883 9827 13889
rect 13814 13880 13820 13892
rect 13872 13880 13878 13932
rect 15580 13920 15608 13948
rect 16758 13920 16764 13932
rect 15580 13892 16764 13920
rect 16758 13880 16764 13892
rect 16816 13880 16822 13932
rect 13262 13812 13268 13864
rect 13320 13852 13326 13864
rect 13449 13855 13507 13861
rect 13449 13852 13461 13855
rect 13320 13824 13461 13852
rect 13320 13812 13326 13824
rect 13449 13821 13461 13824
rect 13495 13821 13507 13855
rect 13449 13815 13507 13821
rect 15381 13855 15439 13861
rect 15381 13821 15393 13855
rect 15427 13852 15439 13855
rect 15838 13852 15844 13864
rect 15427 13824 15844 13852
rect 15427 13821 15439 13824
rect 15381 13815 15439 13821
rect 15838 13812 15844 13824
rect 15896 13812 15902 13864
rect 17129 13855 17187 13861
rect 17129 13821 17141 13855
rect 17175 13852 17187 13855
rect 17954 13852 17960 13864
rect 17175 13824 17960 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 17954 13812 17960 13824
rect 18012 13812 18018 13864
rect 18064 13852 18092 13960
rect 22554 13948 22560 14000
rect 22612 13988 22618 14000
rect 22612 13960 25268 13988
rect 22612 13948 22618 13960
rect 18196 13923 18254 13929
rect 18196 13889 18208 13923
rect 18242 13920 18254 13923
rect 18322 13920 18328 13932
rect 18242 13892 18328 13920
rect 18242 13889 18254 13892
rect 18196 13883 18254 13889
rect 18322 13880 18328 13892
rect 18380 13880 18386 13932
rect 18414 13880 18420 13932
rect 18472 13920 18478 13932
rect 18785 13923 18843 13929
rect 18472 13892 18517 13920
rect 18472 13880 18478 13892
rect 18785 13889 18797 13923
rect 18831 13920 18843 13923
rect 20898 13920 20904 13932
rect 18831 13892 20904 13920
rect 18831 13889 18843 13892
rect 18785 13883 18843 13889
rect 20898 13880 20904 13892
rect 20956 13880 20962 13932
rect 20993 13923 21051 13929
rect 20993 13889 21005 13923
rect 21039 13920 21051 13923
rect 21361 13923 21419 13929
rect 21361 13920 21373 13923
rect 21039 13892 21373 13920
rect 21039 13889 21051 13892
rect 20993 13883 21051 13889
rect 21361 13889 21373 13892
rect 21407 13920 21419 13923
rect 21407 13892 21864 13920
rect 21407 13889 21419 13892
rect 21361 13883 21419 13889
rect 18340 13852 18368 13880
rect 21836 13864 21864 13892
rect 22738 13880 22744 13932
rect 22796 13920 22802 13932
rect 24029 13923 24087 13929
rect 24029 13920 24041 13923
rect 22796 13892 24041 13920
rect 22796 13880 22802 13892
rect 24029 13889 24041 13892
rect 24075 13889 24087 13923
rect 24029 13883 24087 13889
rect 25240 13920 25268 13960
rect 25777 13923 25835 13929
rect 25777 13920 25789 13923
rect 25240 13892 25789 13920
rect 19058 13852 19064 13864
rect 18064 13824 18276 13852
rect 18340 13824 19064 13852
rect 11054 13744 11060 13796
rect 11112 13784 11118 13796
rect 14185 13787 14243 13793
rect 14185 13784 14197 13787
rect 11112 13756 14197 13784
rect 11112 13744 11118 13756
rect 14185 13753 14197 13756
rect 14231 13753 14243 13787
rect 16390 13784 16396 13796
rect 16351 13756 16396 13784
rect 14185 13747 14243 13753
rect 16390 13744 16396 13756
rect 16448 13744 16454 13796
rect 18049 13787 18107 13793
rect 18049 13753 18061 13787
rect 18095 13753 18107 13787
rect 18049 13747 18107 13753
rect 10134 13716 10140 13728
rect 10095 13688 10140 13716
rect 10134 13676 10140 13688
rect 10192 13676 10198 13728
rect 10686 13716 10692 13728
rect 10647 13688 10692 13716
rect 10686 13676 10692 13688
rect 10744 13676 10750 13728
rect 11330 13676 11336 13728
rect 11388 13716 11394 13728
rect 11425 13719 11483 13725
rect 11425 13716 11437 13719
rect 11388 13688 11437 13716
rect 11388 13676 11394 13688
rect 11425 13685 11437 13688
rect 11471 13685 11483 13719
rect 11425 13679 11483 13685
rect 12253 13719 12311 13725
rect 12253 13685 12265 13719
rect 12299 13716 12311 13719
rect 12894 13716 12900 13728
rect 12299 13688 12900 13716
rect 12299 13685 12311 13688
rect 12253 13679 12311 13685
rect 12894 13676 12900 13688
rect 12952 13676 12958 13728
rect 14550 13716 14556 13728
rect 14463 13688 14556 13716
rect 14550 13676 14556 13688
rect 14608 13716 14614 13728
rect 14826 13716 14832 13728
rect 14608 13688 14832 13716
rect 14608 13676 14614 13688
rect 14826 13676 14832 13688
rect 14884 13676 14890 13728
rect 16206 13716 16212 13728
rect 16167 13688 16212 13716
rect 16206 13676 16212 13688
rect 16264 13676 16270 13728
rect 17862 13716 17868 13728
rect 17823 13688 17868 13716
rect 17862 13676 17868 13688
rect 17920 13716 17926 13728
rect 18064 13716 18092 13747
rect 17920 13688 18092 13716
rect 18248 13716 18276 13824
rect 19058 13812 19064 13824
rect 19116 13852 19122 13864
rect 19334 13852 19340 13864
rect 19116 13824 19340 13852
rect 19116 13812 19122 13824
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 19613 13855 19671 13861
rect 19613 13821 19625 13855
rect 19659 13852 19671 13855
rect 20073 13855 20131 13861
rect 20073 13852 20085 13855
rect 19659 13824 20085 13852
rect 19659 13821 19671 13824
rect 19613 13815 19671 13821
rect 20073 13821 20085 13824
rect 20119 13821 20131 13855
rect 21818 13852 21824 13864
rect 21779 13824 21824 13852
rect 20073 13815 20131 13821
rect 19628 13716 19656 13815
rect 21818 13812 21824 13824
rect 21876 13812 21882 13864
rect 25240 13861 25268 13892
rect 25777 13889 25789 13892
rect 25823 13889 25835 13923
rect 25777 13883 25835 13889
rect 25225 13855 25283 13861
rect 25225 13821 25237 13855
rect 25271 13821 25283 13855
rect 25225 13815 25283 13821
rect 23750 13784 23756 13796
rect 23711 13756 23756 13784
rect 23750 13744 23756 13756
rect 23808 13744 23814 13796
rect 23845 13787 23903 13793
rect 23845 13753 23857 13787
rect 23891 13753 23903 13787
rect 23845 13747 23903 13753
rect 18248 13688 19656 13716
rect 19797 13719 19855 13725
rect 17920 13676 17926 13688
rect 19797 13685 19809 13719
rect 19843 13716 19855 13719
rect 19978 13716 19984 13728
rect 19843 13688 19984 13716
rect 19843 13685 19855 13688
rect 19797 13679 19855 13685
rect 19978 13676 19984 13688
rect 20036 13676 20042 13728
rect 23290 13676 23296 13728
rect 23348 13716 23354 13728
rect 23860 13716 23888 13747
rect 23348 13688 23888 13716
rect 23348 13676 23354 13688
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 12621 13515 12679 13521
rect 12621 13481 12633 13515
rect 12667 13481 12679 13515
rect 12894 13512 12900 13524
rect 12855 13484 12900 13512
rect 12621 13475 12679 13481
rect 11057 13447 11115 13453
rect 11057 13413 11069 13447
rect 11103 13444 11115 13447
rect 11146 13444 11152 13456
rect 11103 13416 11152 13444
rect 11103 13413 11115 13416
rect 11057 13407 11115 13413
rect 11146 13404 11152 13416
rect 11204 13404 11210 13456
rect 12636 13444 12664 13475
rect 12894 13472 12900 13484
rect 12952 13472 12958 13524
rect 13078 13472 13084 13524
rect 13136 13512 13142 13524
rect 14093 13515 14151 13521
rect 14093 13512 14105 13515
rect 13136 13484 14105 13512
rect 13136 13472 13142 13484
rect 14093 13481 14105 13484
rect 14139 13481 14151 13515
rect 14093 13475 14151 13481
rect 14734 13472 14740 13524
rect 14792 13512 14798 13524
rect 16298 13512 16304 13524
rect 14792 13484 16304 13512
rect 14792 13472 14798 13484
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 16390 13472 16396 13524
rect 16448 13512 16454 13524
rect 16485 13515 16543 13521
rect 16485 13512 16497 13515
rect 16448 13484 16497 13512
rect 16448 13472 16454 13484
rect 16485 13481 16497 13484
rect 16531 13512 16543 13515
rect 17770 13512 17776 13524
rect 16531 13484 17776 13512
rect 16531 13481 16543 13484
rect 16485 13475 16543 13481
rect 17770 13472 17776 13484
rect 17828 13512 17834 13524
rect 18046 13512 18052 13524
rect 17828 13484 18052 13512
rect 17828 13472 17834 13484
rect 18046 13472 18052 13484
rect 18104 13472 18110 13524
rect 18506 13512 18512 13524
rect 18467 13484 18512 13512
rect 18506 13472 18512 13484
rect 18564 13472 18570 13524
rect 21266 13512 21272 13524
rect 21227 13484 21272 13512
rect 21266 13472 21272 13484
rect 21324 13472 21330 13524
rect 21818 13512 21824 13524
rect 21779 13484 21824 13512
rect 21818 13472 21824 13484
rect 21876 13472 21882 13524
rect 13449 13447 13507 13453
rect 13449 13444 13461 13447
rect 12636 13416 13461 13444
rect 13449 13413 13461 13416
rect 13495 13444 13507 13447
rect 13998 13444 14004 13456
rect 13495 13416 14004 13444
rect 13495 13413 13507 13416
rect 13449 13407 13507 13413
rect 13998 13404 14004 13416
rect 14056 13444 14062 13456
rect 16666 13444 16672 13456
rect 14056 13416 16672 13444
rect 14056 13404 14062 13416
rect 16666 13404 16672 13416
rect 16724 13444 16730 13456
rect 16850 13444 16856 13456
rect 16724 13416 16856 13444
rect 16724 13404 16730 13416
rect 16850 13404 16856 13416
rect 16908 13444 16914 13456
rect 17037 13447 17095 13453
rect 17037 13444 17049 13447
rect 16908 13416 17049 13444
rect 16908 13404 16914 13416
rect 17037 13413 17049 13416
rect 17083 13413 17095 13447
rect 21284 13444 21312 13472
rect 22278 13444 22284 13456
rect 21284 13416 22284 13444
rect 17037 13407 17095 13413
rect 22278 13404 22284 13416
rect 22336 13404 22342 13456
rect 22370 13404 22376 13456
rect 22428 13444 22434 13456
rect 22741 13447 22799 13453
rect 22741 13444 22753 13447
rect 22428 13416 22753 13444
rect 22428 13404 22434 13416
rect 22741 13413 22753 13416
rect 22787 13413 22799 13447
rect 22741 13407 22799 13413
rect 22833 13447 22891 13453
rect 22833 13413 22845 13447
rect 22879 13444 22891 13447
rect 22922 13444 22928 13456
rect 22879 13416 22928 13444
rect 22879 13413 22891 13416
rect 22833 13407 22891 13413
rect 22922 13404 22928 13416
rect 22980 13404 22986 13456
rect 24397 13447 24455 13453
rect 24397 13413 24409 13447
rect 24443 13444 24455 13447
rect 24670 13444 24676 13456
rect 24443 13416 24676 13444
rect 24443 13413 24455 13416
rect 24397 13407 24455 13413
rect 24670 13404 24676 13416
rect 24728 13404 24734 13456
rect 12434 13376 12440 13388
rect 12395 13348 12440 13376
rect 12434 13336 12440 13348
rect 12492 13336 12498 13388
rect 13354 13376 13360 13388
rect 13315 13348 13360 13376
rect 13354 13336 13360 13348
rect 13412 13376 13418 13388
rect 13630 13385 13636 13388
rect 13596 13379 13636 13385
rect 13596 13376 13608 13379
rect 13412 13348 13608 13376
rect 13412 13336 13418 13348
rect 13596 13345 13608 13348
rect 13596 13339 13636 13345
rect 13630 13336 13636 13339
rect 13688 13336 13694 13388
rect 15286 13376 15292 13388
rect 15199 13348 15292 13376
rect 15286 13336 15292 13348
rect 15344 13376 15350 13388
rect 15562 13376 15568 13388
rect 15344 13348 15568 13376
rect 15344 13336 15350 13348
rect 15562 13336 15568 13348
rect 15620 13336 15626 13388
rect 19242 13376 19248 13388
rect 19203 13348 19248 13376
rect 19242 13336 19248 13348
rect 19300 13336 19306 13388
rect 19518 13336 19524 13388
rect 19576 13376 19582 13388
rect 19705 13379 19763 13385
rect 19705 13376 19717 13379
rect 19576 13348 19717 13376
rect 19576 13336 19582 13348
rect 19705 13345 19717 13348
rect 19751 13345 19763 13379
rect 19705 13339 19763 13345
rect 10965 13311 11023 13317
rect 10965 13277 10977 13311
rect 11011 13308 11023 13311
rect 11422 13308 11428 13320
rect 11011 13280 11428 13308
rect 11011 13277 11023 13280
rect 10965 13271 11023 13277
rect 11422 13268 11428 13280
rect 11480 13268 11486 13320
rect 13814 13308 13820 13320
rect 13727 13280 13820 13308
rect 13814 13268 13820 13280
rect 13872 13308 13878 13320
rect 14366 13308 14372 13320
rect 13872 13280 14372 13308
rect 13872 13268 13878 13280
rect 14366 13268 14372 13280
rect 14424 13268 14430 13320
rect 14660 13280 16620 13308
rect 10870 13200 10876 13252
rect 10928 13240 10934 13252
rect 11330 13240 11336 13252
rect 10928 13212 11336 13240
rect 10928 13200 10934 13212
rect 11330 13200 11336 13212
rect 11388 13240 11394 13252
rect 11517 13243 11575 13249
rect 11517 13240 11529 13243
rect 11388 13212 11529 13240
rect 11388 13200 11394 13212
rect 11517 13209 11529 13212
rect 11563 13209 11575 13243
rect 11517 13203 11575 13209
rect 12894 13200 12900 13252
rect 12952 13240 12958 13252
rect 13262 13240 13268 13252
rect 12952 13212 13268 13240
rect 12952 13200 12958 13212
rect 13262 13200 13268 13212
rect 13320 13240 13326 13252
rect 13722 13240 13728 13252
rect 13320 13212 13728 13240
rect 13320 13200 13326 13212
rect 13722 13200 13728 13212
rect 13780 13240 13786 13252
rect 14660 13240 14688 13280
rect 13780 13212 14688 13240
rect 13780 13200 13786 13212
rect 14734 13200 14740 13252
rect 14792 13240 14798 13252
rect 15013 13243 15071 13249
rect 15013 13240 15025 13243
rect 14792 13212 15025 13240
rect 14792 13200 14798 13212
rect 15013 13209 15025 13212
rect 15059 13240 15071 13243
rect 16482 13240 16488 13252
rect 15059 13212 16488 13240
rect 15059 13209 15071 13212
rect 15013 13203 15071 13209
rect 16482 13200 16488 13212
rect 16540 13200 16546 13252
rect 16592 13240 16620 13280
rect 16758 13268 16764 13320
rect 16816 13308 16822 13320
rect 17405 13311 17463 13317
rect 17405 13308 17417 13311
rect 16816 13280 17417 13308
rect 16816 13268 16822 13280
rect 17405 13277 17417 13280
rect 17451 13277 17463 13311
rect 17405 13271 17463 13277
rect 19981 13311 20039 13317
rect 19981 13277 19993 13311
rect 20027 13308 20039 13311
rect 20901 13311 20959 13317
rect 20901 13308 20913 13311
rect 20027 13280 20913 13308
rect 20027 13277 20039 13280
rect 19981 13271 20039 13277
rect 20901 13277 20913 13280
rect 20947 13308 20959 13311
rect 21082 13308 21088 13320
rect 20947 13280 21088 13308
rect 20947 13277 20959 13280
rect 20901 13271 20959 13277
rect 21082 13268 21088 13280
rect 21140 13268 21146 13320
rect 22830 13268 22836 13320
rect 22888 13308 22894 13320
rect 23017 13311 23075 13317
rect 23017 13308 23029 13311
rect 22888 13280 23029 13308
rect 22888 13268 22894 13280
rect 23017 13277 23029 13280
rect 23063 13277 23075 13311
rect 23017 13271 23075 13277
rect 24305 13311 24363 13317
rect 24305 13277 24317 13311
rect 24351 13308 24363 13311
rect 25130 13308 25136 13320
rect 24351 13280 25136 13308
rect 24351 13277 24363 13280
rect 24305 13271 24363 13277
rect 25130 13268 25136 13280
rect 25188 13268 25194 13320
rect 16853 13243 16911 13249
rect 16853 13240 16865 13243
rect 16592 13212 16865 13240
rect 16853 13209 16865 13212
rect 16899 13240 16911 13243
rect 17313 13243 17371 13249
rect 17313 13240 17325 13243
rect 16899 13212 17325 13240
rect 16899 13209 16911 13212
rect 16853 13203 16911 13209
rect 17313 13209 17325 13212
rect 17359 13240 17371 13243
rect 17494 13240 17500 13252
rect 17359 13212 17500 13240
rect 17359 13209 17371 13212
rect 17313 13203 17371 13209
rect 17494 13200 17500 13212
rect 17552 13200 17558 13252
rect 24854 13240 24860 13252
rect 24815 13212 24860 13240
rect 24854 13200 24860 13212
rect 24912 13200 24918 13252
rect 12342 13132 12348 13184
rect 12400 13172 12406 13184
rect 14645 13175 14703 13181
rect 14645 13172 14657 13175
rect 12400 13144 14657 13172
rect 12400 13132 12406 13144
rect 14645 13141 14657 13144
rect 14691 13172 14703 13175
rect 14826 13172 14832 13184
rect 14691 13144 14832 13172
rect 14691 13141 14703 13144
rect 14645 13135 14703 13141
rect 14826 13132 14832 13144
rect 14884 13132 14890 13184
rect 15470 13172 15476 13184
rect 15431 13144 15476 13172
rect 15470 13132 15476 13144
rect 15528 13132 15534 13184
rect 15838 13172 15844 13184
rect 15799 13144 15844 13172
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 17202 13175 17260 13181
rect 17202 13141 17214 13175
rect 17248 13172 17260 13175
rect 17402 13172 17408 13184
rect 17248 13144 17408 13172
rect 17248 13141 17260 13144
rect 17202 13135 17260 13141
rect 17402 13132 17408 13144
rect 17460 13132 17466 13184
rect 17678 13172 17684 13184
rect 17639 13144 17684 13172
rect 17678 13132 17684 13144
rect 17736 13132 17742 13184
rect 18598 13132 18604 13184
rect 18656 13172 18662 13184
rect 18785 13175 18843 13181
rect 18785 13172 18797 13175
rect 18656 13144 18797 13172
rect 18656 13132 18662 13144
rect 18785 13141 18797 13144
rect 18831 13141 18843 13175
rect 23750 13172 23756 13184
rect 23711 13144 23756 13172
rect 18785 13135 18843 13141
rect 23750 13132 23756 13144
rect 23808 13132 23814 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 13262 12968 13268 12980
rect 13223 12940 13268 12968
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 14734 12977 14740 12980
rect 14718 12971 14740 12977
rect 14718 12937 14730 12971
rect 14718 12931 14740 12937
rect 14734 12928 14740 12931
rect 14792 12928 14798 12980
rect 15562 12968 15568 12980
rect 15523 12940 15568 12968
rect 15562 12928 15568 12940
rect 15620 12928 15626 12980
rect 16482 12928 16488 12980
rect 16540 12968 16546 12980
rect 18187 12971 18245 12977
rect 18187 12968 18199 12971
rect 16540 12940 18199 12968
rect 16540 12928 16546 12940
rect 18187 12937 18199 12940
rect 18233 12968 18245 12971
rect 18598 12968 18604 12980
rect 18233 12940 18604 12968
rect 18233 12937 18245 12940
rect 18187 12931 18245 12937
rect 18598 12928 18604 12940
rect 18656 12928 18662 12980
rect 18874 12928 18880 12980
rect 18932 12968 18938 12980
rect 19978 12968 19984 12980
rect 18932 12940 19984 12968
rect 18932 12928 18938 12940
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 22370 12968 22376 12980
rect 22331 12940 22376 12968
rect 22370 12928 22376 12940
rect 22428 12928 22434 12980
rect 23106 12968 23112 12980
rect 23067 12940 23112 12968
rect 23106 12928 23112 12940
rect 23164 12928 23170 12980
rect 25130 12968 25136 12980
rect 25091 12940 25136 12968
rect 25130 12928 25136 12940
rect 25188 12928 25194 12980
rect 12434 12860 12440 12912
rect 12492 12900 12498 12912
rect 14277 12903 14335 12909
rect 14277 12900 14289 12903
rect 12492 12872 14289 12900
rect 12492 12860 12498 12872
rect 14277 12869 14289 12872
rect 14323 12869 14335 12903
rect 14277 12863 14335 12869
rect 14826 12860 14832 12912
rect 14884 12900 14890 12912
rect 15654 12900 15660 12912
rect 14884 12872 15660 12900
rect 14884 12860 14890 12872
rect 15654 12860 15660 12872
rect 15712 12860 15718 12912
rect 17494 12860 17500 12912
rect 17552 12900 17558 12912
rect 18325 12903 18383 12909
rect 18325 12900 18337 12903
rect 17552 12872 18337 12900
rect 17552 12860 17558 12872
rect 18325 12869 18337 12872
rect 18371 12869 18383 12903
rect 18616 12900 18644 12928
rect 19797 12903 19855 12909
rect 19797 12900 19809 12903
rect 18616 12872 19809 12900
rect 18325 12863 18383 12869
rect 19797 12869 19809 12872
rect 19843 12869 19855 12903
rect 19797 12863 19855 12869
rect 21913 12903 21971 12909
rect 21913 12869 21925 12903
rect 21959 12869 21971 12903
rect 21913 12863 21971 12869
rect 10870 12832 10876 12844
rect 10831 12804 10876 12832
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 11885 12835 11943 12841
rect 11885 12801 11897 12835
rect 11931 12832 11943 12835
rect 12250 12832 12256 12844
rect 11931 12804 12256 12832
rect 11931 12801 11943 12804
rect 11885 12795 11943 12801
rect 12250 12792 12256 12804
rect 12308 12832 12314 12844
rect 13357 12835 13415 12841
rect 13357 12832 13369 12835
rect 12308 12804 13369 12832
rect 12308 12792 12314 12804
rect 13357 12801 13369 12804
rect 13403 12801 13415 12835
rect 13357 12795 13415 12801
rect 14918 12792 14924 12844
rect 14976 12832 14982 12844
rect 15746 12832 15752 12844
rect 14976 12804 15752 12832
rect 14976 12792 14982 12804
rect 15746 12792 15752 12804
rect 15804 12792 15810 12844
rect 17126 12832 17132 12844
rect 17087 12804 17132 12832
rect 17126 12792 17132 12804
rect 17184 12792 17190 12844
rect 18417 12835 18475 12841
rect 18417 12832 18429 12835
rect 17788 12804 18429 12832
rect 13136 12767 13194 12773
rect 13136 12733 13148 12767
rect 13182 12733 13194 12767
rect 13136 12727 13194 12733
rect 14093 12767 14151 12773
rect 14093 12733 14105 12767
rect 14139 12764 14151 12767
rect 14366 12764 14372 12776
rect 14139 12736 14372 12764
rect 14139 12733 14151 12736
rect 14093 12727 14151 12733
rect 10042 12696 10048 12708
rect 4126 12668 10048 12696
rect 1578 12588 1584 12640
rect 1636 12628 1642 12640
rect 4126 12628 4154 12668
rect 10042 12656 10048 12668
rect 10100 12696 10106 12708
rect 10229 12699 10287 12705
rect 10229 12696 10241 12699
rect 10100 12668 10241 12696
rect 10100 12656 10106 12668
rect 10229 12665 10241 12668
rect 10275 12665 10287 12699
rect 10229 12659 10287 12665
rect 10321 12699 10379 12705
rect 10321 12665 10333 12699
rect 10367 12696 10379 12699
rect 10686 12696 10692 12708
rect 10367 12668 10692 12696
rect 10367 12665 10379 12668
rect 10321 12659 10379 12665
rect 1636 12600 4154 12628
rect 1636 12588 1642 12600
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 9953 12631 10011 12637
rect 9953 12628 9965 12631
rect 9732 12600 9965 12628
rect 9732 12588 9738 12600
rect 9953 12597 9965 12600
rect 9999 12628 10011 12631
rect 10336 12628 10364 12659
rect 10686 12656 10692 12668
rect 10744 12656 10750 12708
rect 10870 12656 10876 12708
rect 10928 12696 10934 12708
rect 12161 12699 12219 12705
rect 12161 12696 12173 12699
rect 10928 12668 12173 12696
rect 10928 12656 10934 12668
rect 12161 12665 12173 12668
rect 12207 12696 12219 12699
rect 12434 12696 12440 12708
rect 12207 12668 12440 12696
rect 12207 12665 12219 12668
rect 12161 12659 12219 12665
rect 12434 12656 12440 12668
rect 12492 12656 12498 12708
rect 12986 12696 12992 12708
rect 12947 12668 12992 12696
rect 12986 12656 12992 12668
rect 13044 12656 13050 12708
rect 11146 12628 11152 12640
rect 9999 12600 10364 12628
rect 11107 12600 11152 12628
rect 9999 12597 10011 12600
rect 9953 12591 10011 12597
rect 11146 12588 11152 12600
rect 11204 12588 11210 12640
rect 12897 12631 12955 12637
rect 12897 12597 12909 12631
rect 12943 12628 12955 12631
rect 13151 12628 13179 12727
rect 14366 12724 14372 12736
rect 14424 12724 14430 12776
rect 16390 12764 16396 12776
rect 14936 12736 16396 12764
rect 13722 12696 13728 12708
rect 13683 12668 13728 12696
rect 13722 12656 13728 12668
rect 13780 12656 13786 12708
rect 14277 12699 14335 12705
rect 14277 12665 14289 12699
rect 14323 12696 14335 12699
rect 14553 12699 14611 12705
rect 14553 12696 14565 12699
rect 14323 12668 14565 12696
rect 14323 12665 14335 12668
rect 14277 12659 14335 12665
rect 14553 12665 14565 12668
rect 14599 12696 14611 12699
rect 14734 12696 14740 12708
rect 14599 12668 14740 12696
rect 14599 12665 14611 12668
rect 14553 12659 14611 12665
rect 14734 12656 14740 12668
rect 14792 12696 14798 12708
rect 14936 12696 14964 12736
rect 16390 12724 16396 12736
rect 16448 12724 16454 12776
rect 16485 12767 16543 12773
rect 16485 12733 16497 12767
rect 16531 12733 16543 12767
rect 16485 12727 16543 12733
rect 15286 12696 15292 12708
rect 14792 12668 14964 12696
rect 15247 12668 15292 12696
rect 14792 12656 14798 12668
rect 15286 12656 15292 12668
rect 15344 12656 15350 12708
rect 16500 12696 16528 12727
rect 16224 12668 16528 12696
rect 16224 12640 16252 12668
rect 14182 12628 14188 12640
rect 12943 12600 14188 12628
rect 12943 12597 12955 12600
rect 12897 12591 12955 12597
rect 14182 12588 14188 12600
rect 14240 12588 14246 12640
rect 14366 12588 14372 12640
rect 14424 12628 14430 12640
rect 14461 12631 14519 12637
rect 14461 12628 14473 12631
rect 14424 12600 14473 12628
rect 14424 12588 14430 12600
rect 14461 12597 14473 12600
rect 14507 12628 14519 12631
rect 14918 12628 14924 12640
rect 14507 12600 14924 12628
rect 14507 12597 14519 12600
rect 14461 12591 14519 12597
rect 14918 12588 14924 12600
rect 14976 12588 14982 12640
rect 16206 12628 16212 12640
rect 16167 12600 16212 12628
rect 16206 12588 16212 12600
rect 16264 12588 16270 12640
rect 17402 12628 17408 12640
rect 17363 12600 17408 12628
rect 17402 12588 17408 12600
rect 17460 12588 17466 12640
rect 17586 12588 17592 12640
rect 17644 12628 17650 12640
rect 17788 12637 17816 12804
rect 18417 12801 18429 12804
rect 18463 12801 18475 12835
rect 19242 12832 19248 12844
rect 19203 12804 19248 12832
rect 18417 12795 18475 12801
rect 19242 12792 19248 12804
rect 19300 12792 19306 12844
rect 21928 12832 21956 12863
rect 22741 12835 22799 12841
rect 22741 12832 22753 12835
rect 21928 12804 22753 12832
rect 22741 12801 22753 12804
rect 22787 12832 22799 12835
rect 22922 12832 22928 12844
rect 22787 12804 22928 12832
rect 22787 12801 22799 12804
rect 22741 12795 22799 12801
rect 22922 12792 22928 12804
rect 22980 12792 22986 12844
rect 23750 12792 23756 12844
rect 23808 12832 23814 12844
rect 25225 12835 25283 12841
rect 25225 12832 25237 12835
rect 23808 12804 25237 12832
rect 23808 12792 23814 12804
rect 25225 12801 25237 12804
rect 25271 12801 25283 12835
rect 25225 12795 25283 12801
rect 18046 12764 18052 12776
rect 18007 12736 18052 12764
rect 18046 12724 18052 12736
rect 18104 12724 18110 12776
rect 19334 12724 19340 12776
rect 19392 12764 19398 12776
rect 19613 12767 19671 12773
rect 19613 12764 19625 12767
rect 19392 12736 19625 12764
rect 19392 12724 19398 12736
rect 19613 12733 19625 12736
rect 19659 12764 19671 12767
rect 20073 12767 20131 12773
rect 20073 12764 20085 12767
rect 19659 12736 20085 12764
rect 19659 12733 19671 12736
rect 19613 12727 19671 12733
rect 20073 12733 20085 12736
rect 20119 12733 20131 12767
rect 20990 12764 20996 12776
rect 20951 12736 20996 12764
rect 20073 12727 20131 12733
rect 20990 12724 20996 12736
rect 21048 12724 21054 12776
rect 18785 12699 18843 12705
rect 18785 12665 18797 12699
rect 18831 12696 18843 12699
rect 19518 12696 19524 12708
rect 18831 12668 19524 12696
rect 18831 12665 18843 12668
rect 18785 12659 18843 12665
rect 19518 12656 19524 12668
rect 19576 12656 19582 12708
rect 21266 12696 21272 12708
rect 21224 12668 21272 12696
rect 21266 12656 21272 12668
rect 21324 12705 21330 12708
rect 21324 12699 21372 12705
rect 21324 12665 21326 12699
rect 21360 12665 21372 12699
rect 21324 12659 21372 12665
rect 21324 12656 21357 12659
rect 23106 12656 23112 12708
rect 23164 12696 23170 12708
rect 23753 12699 23811 12705
rect 23753 12696 23765 12699
rect 23164 12668 23765 12696
rect 23164 12656 23170 12668
rect 23753 12665 23765 12668
rect 23799 12665 23811 12699
rect 23753 12659 23811 12665
rect 23845 12699 23903 12705
rect 23845 12665 23857 12699
rect 23891 12696 23903 12699
rect 24210 12696 24216 12708
rect 23891 12668 24216 12696
rect 23891 12665 23903 12668
rect 23845 12659 23903 12665
rect 17773 12631 17831 12637
rect 17773 12628 17785 12631
rect 17644 12600 17785 12628
rect 17644 12588 17650 12600
rect 17773 12597 17785 12600
rect 17819 12597 17831 12631
rect 17773 12591 17831 12597
rect 20533 12631 20591 12637
rect 20533 12597 20545 12631
rect 20579 12628 20591 12631
rect 20809 12631 20867 12637
rect 20809 12628 20821 12631
rect 20579 12600 20821 12628
rect 20579 12597 20591 12600
rect 20533 12591 20591 12597
rect 20809 12597 20821 12600
rect 20855 12628 20867 12631
rect 21329 12628 21357 12656
rect 21634 12628 21640 12640
rect 20855 12600 21640 12628
rect 20855 12597 20867 12600
rect 20809 12591 20867 12597
rect 21634 12588 21640 12600
rect 21692 12588 21698 12640
rect 23477 12631 23535 12637
rect 23477 12597 23489 12631
rect 23523 12628 23535 12631
rect 23860 12628 23888 12659
rect 24210 12656 24216 12668
rect 24268 12656 24274 12708
rect 24397 12699 24455 12705
rect 24397 12665 24409 12699
rect 24443 12696 24455 12699
rect 24578 12696 24584 12708
rect 24443 12668 24584 12696
rect 24443 12665 24455 12668
rect 24397 12659 24455 12665
rect 24578 12656 24584 12668
rect 24636 12696 24642 12708
rect 24854 12696 24860 12708
rect 24636 12668 24860 12696
rect 24636 12656 24642 12668
rect 24854 12656 24860 12668
rect 24912 12656 24918 12708
rect 24670 12628 24676 12640
rect 23523 12600 23888 12628
rect 24631 12600 24676 12628
rect 23523 12597 23535 12600
rect 23477 12591 23535 12597
rect 24670 12588 24676 12600
rect 24728 12588 24734 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 10137 12427 10195 12433
rect 10137 12424 10149 12427
rect 10100 12396 10149 12424
rect 10100 12384 10106 12396
rect 10137 12393 10149 12396
rect 10183 12393 10195 12427
rect 12342 12424 12348 12436
rect 12303 12396 12348 12424
rect 10137 12387 10195 12393
rect 12342 12384 12348 12396
rect 12400 12384 12406 12436
rect 12713 12427 12771 12433
rect 12713 12393 12725 12427
rect 12759 12424 12771 12427
rect 12894 12424 12900 12436
rect 12759 12396 12900 12424
rect 12759 12393 12771 12396
rect 12713 12387 12771 12393
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 12986 12384 12992 12436
rect 13044 12424 13050 12436
rect 13081 12427 13139 12433
rect 13081 12424 13093 12427
rect 13044 12396 13093 12424
rect 13044 12384 13050 12396
rect 13081 12393 13093 12396
rect 13127 12424 13139 12427
rect 13357 12427 13415 12433
rect 13357 12424 13369 12427
rect 13127 12396 13369 12424
rect 13127 12393 13139 12396
rect 13081 12387 13139 12393
rect 13357 12393 13369 12396
rect 13403 12424 13415 12427
rect 13446 12424 13452 12436
rect 13403 12396 13452 12424
rect 13403 12393 13415 12396
rect 13357 12387 13415 12393
rect 13446 12384 13452 12396
rect 13504 12384 13510 12436
rect 13630 12424 13636 12436
rect 13591 12396 13636 12424
rect 13630 12384 13636 12396
rect 13688 12384 13694 12436
rect 13722 12384 13728 12436
rect 13780 12424 13786 12436
rect 14826 12424 14832 12436
rect 13780 12396 14832 12424
rect 13780 12384 13786 12396
rect 14826 12384 14832 12396
rect 14884 12384 14890 12436
rect 16393 12427 16451 12433
rect 16393 12393 16405 12427
rect 16439 12424 16451 12427
rect 16482 12424 16488 12436
rect 16439 12396 16488 12424
rect 16439 12393 16451 12396
rect 16393 12387 16451 12393
rect 16482 12384 16488 12396
rect 16540 12384 16546 12436
rect 16758 12424 16764 12436
rect 16719 12396 16764 12424
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 16850 12384 16856 12436
rect 16908 12424 16914 12436
rect 17037 12427 17095 12433
rect 17037 12424 17049 12427
rect 16908 12396 17049 12424
rect 16908 12384 16914 12396
rect 17037 12393 17049 12396
rect 17083 12393 17095 12427
rect 18598 12424 18604 12436
rect 18559 12396 18604 12424
rect 17037 12387 17095 12393
rect 18598 12384 18604 12396
rect 18656 12384 18662 12436
rect 21082 12424 21088 12436
rect 21043 12396 21088 12424
rect 21082 12384 21088 12396
rect 21140 12384 21146 12436
rect 11146 12356 11152 12368
rect 11107 12328 11152 12356
rect 11146 12316 11152 12328
rect 11204 12316 11210 12368
rect 13998 12356 14004 12368
rect 13959 12328 14004 12356
rect 13998 12316 14004 12328
rect 14056 12316 14062 12368
rect 14734 12356 14740 12368
rect 14695 12328 14740 12356
rect 14734 12316 14740 12328
rect 14792 12316 14798 12368
rect 17221 12359 17279 12365
rect 17221 12356 17233 12359
rect 15396 12328 17233 12356
rect 15396 12300 15424 12328
rect 17221 12325 17233 12328
rect 17267 12356 17279 12359
rect 17770 12356 17776 12368
rect 17267 12328 17776 12356
rect 17267 12325 17279 12328
rect 17221 12319 17279 12325
rect 17770 12316 17776 12328
rect 17828 12316 17834 12368
rect 19981 12359 20039 12365
rect 19981 12325 19993 12359
rect 20027 12356 20039 12359
rect 20990 12356 20996 12368
rect 20027 12328 20996 12356
rect 20027 12325 20039 12328
rect 19981 12319 20039 12325
rect 20990 12316 20996 12328
rect 21048 12356 21054 12368
rect 21453 12359 21511 12365
rect 21453 12356 21465 12359
rect 21048 12328 21465 12356
rect 21048 12316 21054 12328
rect 21453 12325 21465 12328
rect 21499 12325 21511 12359
rect 21453 12319 21511 12325
rect 21634 12316 21640 12368
rect 21692 12356 21698 12368
rect 22050 12359 22108 12365
rect 22050 12356 22062 12359
rect 21692 12328 22062 12356
rect 21692 12316 21698 12328
rect 22050 12325 22062 12328
rect 22096 12325 22108 12359
rect 22050 12319 22108 12325
rect 24397 12359 24455 12365
rect 24397 12325 24409 12359
rect 24443 12356 24455 12359
rect 24670 12356 24676 12368
rect 24443 12328 24676 12356
rect 24443 12325 24455 12328
rect 24397 12319 24455 12325
rect 24670 12316 24676 12328
rect 24728 12316 24734 12368
rect 9674 12248 9680 12300
rect 9732 12288 9738 12300
rect 10505 12291 10563 12297
rect 10505 12288 10517 12291
rect 9732 12260 10517 12288
rect 9732 12248 9738 12260
rect 10505 12257 10517 12260
rect 10551 12257 10563 12291
rect 10505 12251 10563 12257
rect 12161 12291 12219 12297
rect 12161 12257 12173 12291
rect 12207 12288 12219 12291
rect 12342 12288 12348 12300
rect 12207 12260 12348 12288
rect 12207 12257 12219 12260
rect 12161 12251 12219 12257
rect 12342 12248 12348 12260
rect 12400 12248 12406 12300
rect 12986 12248 12992 12300
rect 13044 12288 13050 12300
rect 13173 12291 13231 12297
rect 13173 12288 13185 12291
rect 13044 12260 13185 12288
rect 13044 12248 13050 12260
rect 13173 12257 13185 12260
rect 13219 12257 13231 12291
rect 14182 12288 14188 12300
rect 14143 12260 14188 12288
rect 13173 12251 13231 12257
rect 14182 12248 14188 12260
rect 14240 12248 14246 12300
rect 15289 12291 15347 12297
rect 15289 12257 15301 12291
rect 15335 12288 15347 12291
rect 15378 12288 15384 12300
rect 15335 12260 15384 12288
rect 15335 12257 15347 12260
rect 15289 12251 15347 12257
rect 15378 12248 15384 12260
rect 15436 12248 15442 12300
rect 16482 12288 16488 12300
rect 15488 12260 16488 12288
rect 13630 12112 13636 12164
rect 13688 12152 13694 12164
rect 15488 12161 15516 12260
rect 16482 12248 16488 12260
rect 16540 12248 16546 12300
rect 19242 12288 19248 12300
rect 19203 12260 19248 12288
rect 19242 12248 19248 12260
rect 19300 12248 19306 12300
rect 19518 12248 19524 12300
rect 19576 12288 19582 12300
rect 19705 12291 19763 12297
rect 19705 12288 19717 12291
rect 19576 12260 19717 12288
rect 19576 12248 19582 12260
rect 19705 12257 19717 12260
rect 19751 12257 19763 12291
rect 19705 12251 19763 12257
rect 22649 12291 22707 12297
rect 22649 12257 22661 12291
rect 22695 12288 22707 12291
rect 24210 12288 24216 12300
rect 22695 12260 24216 12288
rect 22695 12257 22707 12260
rect 22649 12251 22707 12257
rect 24210 12248 24216 12260
rect 24268 12248 24274 12300
rect 25222 12288 25228 12300
rect 25183 12260 25228 12288
rect 25222 12248 25228 12260
rect 25280 12248 25286 12300
rect 15657 12223 15715 12229
rect 15657 12189 15669 12223
rect 15703 12220 15715 12223
rect 15746 12220 15752 12232
rect 15703 12192 15752 12220
rect 15703 12189 15715 12192
rect 15657 12183 15715 12189
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 17586 12220 17592 12232
rect 17547 12192 17592 12220
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 19153 12223 19211 12229
rect 19153 12189 19165 12223
rect 19199 12220 19211 12223
rect 19536 12220 19564 12248
rect 19199 12192 19564 12220
rect 21729 12223 21787 12229
rect 19199 12189 19211 12192
rect 19153 12183 19211 12189
rect 21729 12189 21741 12223
rect 21775 12220 21787 12223
rect 22094 12220 22100 12232
rect 21775 12192 22100 12220
rect 21775 12189 21787 12192
rect 21729 12183 21787 12189
rect 22094 12180 22100 12192
rect 22152 12180 22158 12232
rect 14369 12155 14427 12161
rect 14369 12152 14381 12155
rect 13688 12124 14381 12152
rect 13688 12112 13694 12124
rect 14369 12121 14381 12124
rect 14415 12121 14427 12155
rect 14369 12115 14427 12121
rect 15454 12155 15516 12161
rect 15454 12121 15466 12155
rect 15500 12124 15516 12155
rect 15500 12121 15512 12124
rect 15454 12115 15512 12121
rect 16482 12112 16488 12164
rect 16540 12152 16546 12164
rect 17494 12152 17500 12164
rect 16540 12124 17080 12152
rect 17455 12124 17500 12152
rect 16540 12112 16546 12124
rect 11514 12084 11520 12096
rect 11475 12056 11520 12084
rect 11514 12044 11520 12056
rect 11572 12044 11578 12096
rect 14826 12044 14832 12096
rect 14884 12084 14890 12096
rect 15013 12087 15071 12093
rect 15013 12084 15025 12087
rect 14884 12056 15025 12084
rect 14884 12044 14890 12056
rect 15013 12053 15025 12056
rect 15059 12053 15071 12087
rect 15013 12047 15071 12053
rect 15565 12087 15623 12093
rect 15565 12053 15577 12087
rect 15611 12084 15623 12087
rect 15654 12084 15660 12096
rect 15611 12056 15660 12084
rect 15611 12053 15623 12056
rect 15565 12047 15623 12053
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 15933 12087 15991 12093
rect 15933 12053 15945 12087
rect 15979 12084 15991 12087
rect 16850 12084 16856 12096
rect 15979 12056 16856 12084
rect 15979 12053 15991 12056
rect 15933 12047 15991 12053
rect 16850 12044 16856 12056
rect 16908 12044 16914 12096
rect 17052 12084 17080 12124
rect 17494 12112 17500 12124
rect 17552 12112 17558 12164
rect 17865 12155 17923 12161
rect 17865 12121 17877 12155
rect 17911 12152 17923 12155
rect 20530 12152 20536 12164
rect 17911 12124 20536 12152
rect 17911 12121 17923 12124
rect 17865 12115 17923 12121
rect 20530 12112 20536 12124
rect 20588 12112 20594 12164
rect 25406 12152 25412 12164
rect 25367 12124 25412 12152
rect 25406 12112 25412 12124
rect 25464 12112 25470 12164
rect 17359 12087 17417 12093
rect 17359 12084 17371 12087
rect 17052 12056 17371 12084
rect 17359 12053 17371 12056
rect 17405 12053 17417 12087
rect 17512 12084 17540 12112
rect 18233 12087 18291 12093
rect 18233 12084 18245 12087
rect 17512 12056 18245 12084
rect 17359 12047 17417 12053
rect 18233 12053 18245 12056
rect 18279 12084 18291 12087
rect 18874 12084 18880 12096
rect 18279 12056 18880 12084
rect 18279 12053 18291 12056
rect 18233 12047 18291 12053
rect 18874 12044 18880 12056
rect 18932 12044 18938 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 9674 11880 9680 11892
rect 9635 11852 9680 11880
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 13909 11883 13967 11889
rect 13909 11849 13921 11883
rect 13955 11880 13967 11883
rect 14182 11880 14188 11892
rect 13955 11852 14188 11880
rect 13955 11849 13967 11852
rect 13909 11843 13967 11849
rect 14182 11840 14188 11852
rect 14240 11840 14246 11892
rect 15654 11880 15660 11892
rect 15615 11852 15660 11880
rect 15654 11840 15660 11852
rect 15712 11840 15718 11892
rect 17770 11880 17776 11892
rect 17731 11852 17776 11880
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 18874 11880 18880 11892
rect 18835 11852 18880 11880
rect 18874 11840 18880 11852
rect 18932 11840 18938 11892
rect 23658 11840 23664 11892
rect 23716 11880 23722 11892
rect 23799 11883 23857 11889
rect 23799 11880 23811 11883
rect 23716 11852 23811 11880
rect 23716 11840 23722 11852
rect 23799 11849 23811 11852
rect 23845 11849 23857 11883
rect 24210 11880 24216 11892
rect 24171 11852 24216 11880
rect 23799 11843 23857 11849
rect 24210 11840 24216 11852
rect 24268 11840 24274 11892
rect 25222 11840 25228 11892
rect 25280 11880 25286 11892
rect 25501 11883 25559 11889
rect 25501 11880 25513 11883
rect 25280 11852 25513 11880
rect 25280 11840 25286 11852
rect 25501 11849 25513 11852
rect 25547 11849 25559 11883
rect 25501 11843 25559 11849
rect 15381 11815 15439 11821
rect 15381 11781 15393 11815
rect 15427 11812 15439 11815
rect 15746 11812 15752 11824
rect 15427 11784 15752 11812
rect 15427 11781 15439 11784
rect 15381 11775 15439 11781
rect 15746 11772 15752 11784
rect 15804 11812 15810 11824
rect 18233 11815 18291 11821
rect 18233 11812 18245 11815
rect 15804 11784 18245 11812
rect 15804 11772 15810 11784
rect 18233 11781 18245 11784
rect 18279 11781 18291 11815
rect 18233 11775 18291 11781
rect 21358 11772 21364 11824
rect 21416 11812 21422 11824
rect 24811 11815 24869 11821
rect 24811 11812 24823 11815
rect 21416 11784 24823 11812
rect 21416 11772 21422 11784
rect 24811 11781 24823 11784
rect 24857 11781 24869 11815
rect 24811 11775 24869 11781
rect 8938 11704 8944 11756
rect 8996 11744 9002 11756
rect 10321 11747 10379 11753
rect 10321 11744 10333 11747
rect 8996 11716 10333 11744
rect 8996 11704 9002 11716
rect 10321 11713 10333 11716
rect 10367 11744 10379 11747
rect 14458 11744 14464 11756
rect 10367 11716 11100 11744
rect 10367 11713 10379 11716
rect 10321 11707 10379 11713
rect 10505 11679 10563 11685
rect 10505 11676 10517 11679
rect 10152 11648 10517 11676
rect 10152 11552 10180 11648
rect 10505 11645 10517 11648
rect 10551 11645 10563 11679
rect 10870 11676 10876 11688
rect 10831 11648 10876 11676
rect 10505 11639 10563 11645
rect 10870 11636 10876 11648
rect 10928 11636 10934 11688
rect 11072 11685 11100 11716
rect 14292 11716 14464 11744
rect 14292 11685 14320 11716
rect 14458 11704 14464 11716
rect 14516 11744 14522 11756
rect 15470 11744 15476 11756
rect 14516 11716 15476 11744
rect 14516 11704 14522 11716
rect 15470 11704 15476 11716
rect 15528 11704 15534 11756
rect 15838 11704 15844 11756
rect 15896 11744 15902 11756
rect 16393 11747 16451 11753
rect 16393 11744 16405 11747
rect 15896 11716 16405 11744
rect 15896 11704 15902 11716
rect 16393 11713 16405 11716
rect 16439 11713 16451 11747
rect 16393 11707 16451 11713
rect 11057 11679 11115 11685
rect 11057 11645 11069 11679
rect 11103 11676 11115 11679
rect 12621 11679 12679 11685
rect 12621 11676 12633 11679
rect 11103 11648 12633 11676
rect 11103 11645 11115 11648
rect 11057 11639 11115 11645
rect 12621 11645 12633 11648
rect 12667 11676 12679 11679
rect 13265 11679 13323 11685
rect 13265 11676 13277 11679
rect 12667 11648 13277 11676
rect 12667 11645 12679 11648
rect 12621 11639 12679 11645
rect 13265 11645 13277 11648
rect 13311 11645 13323 11679
rect 13265 11639 13323 11645
rect 14277 11679 14335 11685
rect 14277 11645 14289 11679
rect 14323 11645 14335 11679
rect 14277 11639 14335 11645
rect 14553 11679 14611 11685
rect 14553 11645 14565 11679
rect 14599 11676 14611 11679
rect 14826 11676 14832 11688
rect 14599 11648 14832 11676
rect 14599 11645 14611 11648
rect 14553 11639 14611 11645
rect 14826 11636 14832 11648
rect 14884 11636 14890 11688
rect 16485 11679 16543 11685
rect 16485 11676 16497 11679
rect 16408 11648 16497 11676
rect 12434 11608 12440 11620
rect 12395 11580 12440 11608
rect 12434 11568 12440 11580
rect 12492 11568 12498 11620
rect 12986 11608 12992 11620
rect 12947 11580 12992 11608
rect 12986 11568 12992 11580
rect 13044 11568 13050 11620
rect 14734 11608 14740 11620
rect 14695 11580 14740 11608
rect 14734 11568 14740 11580
rect 14792 11568 14798 11620
rect 16408 11552 16436 11648
rect 16485 11645 16497 11648
rect 16531 11676 16543 11679
rect 17405 11679 17463 11685
rect 17405 11676 17417 11679
rect 16531 11648 17417 11676
rect 16531 11645 16543 11648
rect 16485 11639 16543 11645
rect 17405 11645 17417 11648
rect 17451 11676 17463 11679
rect 17586 11676 17592 11688
rect 17451 11648 17592 11676
rect 17451 11645 17463 11648
rect 17405 11639 17463 11645
rect 17586 11636 17592 11648
rect 17644 11676 17650 11688
rect 18049 11679 18107 11685
rect 18049 11676 18061 11679
rect 17644 11648 18061 11676
rect 17644 11636 17650 11648
rect 18049 11645 18061 11648
rect 18095 11676 18107 11679
rect 18509 11679 18567 11685
rect 18509 11676 18521 11679
rect 18095 11648 18521 11676
rect 18095 11645 18107 11648
rect 18049 11639 18107 11645
rect 18509 11645 18521 11648
rect 18555 11645 18567 11679
rect 20073 11679 20131 11685
rect 20073 11676 20085 11679
rect 18509 11639 18567 11645
rect 19904 11648 20085 11676
rect 10045 11543 10103 11549
rect 10045 11509 10057 11543
rect 10091 11540 10103 11543
rect 10134 11540 10140 11552
rect 10091 11512 10140 11540
rect 10091 11509 10103 11512
rect 10045 11503 10103 11509
rect 10134 11500 10140 11512
rect 10192 11500 10198 11552
rect 12253 11543 12311 11549
rect 12253 11509 12265 11543
rect 12299 11540 12311 11543
rect 12342 11540 12348 11552
rect 12299 11512 12348 11540
rect 12299 11509 12311 11512
rect 12253 11503 12311 11509
rect 12342 11500 12348 11512
rect 12400 11500 12406 11552
rect 16301 11543 16359 11549
rect 16301 11509 16313 11543
rect 16347 11540 16359 11543
rect 16390 11540 16396 11552
rect 16347 11512 16396 11540
rect 16347 11509 16359 11512
rect 16301 11503 16359 11509
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 18690 11500 18696 11552
rect 18748 11540 18754 11552
rect 19242 11540 19248 11552
rect 18748 11512 19248 11540
rect 18748 11500 18754 11512
rect 19242 11500 19248 11512
rect 19300 11540 19306 11552
rect 19904 11549 19932 11648
rect 20073 11645 20085 11648
rect 20119 11645 20131 11679
rect 20530 11676 20536 11688
rect 20491 11648 20536 11676
rect 20073 11639 20131 11645
rect 20530 11636 20536 11648
rect 20588 11636 20594 11688
rect 22646 11636 22652 11688
rect 22704 11676 22710 11688
rect 23728 11679 23786 11685
rect 23728 11676 23740 11679
rect 22704 11648 23740 11676
rect 22704 11636 22710 11648
rect 23728 11645 23740 11648
rect 23774 11676 23786 11679
rect 24489 11679 24547 11685
rect 24489 11676 24501 11679
rect 23774 11648 24501 11676
rect 23774 11645 23786 11648
rect 23728 11639 23786 11645
rect 24489 11645 24501 11648
rect 24535 11645 24547 11679
rect 24489 11639 24547 11645
rect 24740 11679 24798 11685
rect 24740 11645 24752 11679
rect 24786 11676 24798 11679
rect 24786 11648 25268 11676
rect 24786 11645 24798 11648
rect 24740 11639 24798 11645
rect 20809 11611 20867 11617
rect 20809 11577 20821 11611
rect 20855 11608 20867 11611
rect 22738 11608 22744 11620
rect 20855 11580 22744 11608
rect 20855 11577 20867 11580
rect 20809 11571 20867 11577
rect 22738 11568 22744 11580
rect 22796 11568 22802 11620
rect 25240 11552 25268 11648
rect 19889 11543 19947 11549
rect 19889 11540 19901 11543
rect 19300 11512 19901 11540
rect 19300 11500 19306 11512
rect 19889 11509 19901 11512
rect 19935 11509 19947 11543
rect 19889 11503 19947 11509
rect 21634 11500 21640 11552
rect 21692 11540 21698 11552
rect 21729 11543 21787 11549
rect 21729 11540 21741 11543
rect 21692 11512 21741 11540
rect 21692 11500 21698 11512
rect 21729 11509 21741 11512
rect 21775 11509 21787 11543
rect 22094 11540 22100 11552
rect 22055 11512 22100 11540
rect 21729 11503 21787 11509
rect 22094 11500 22100 11512
rect 22152 11500 22158 11552
rect 22557 11543 22615 11549
rect 22557 11509 22569 11543
rect 22603 11540 22615 11543
rect 23934 11540 23940 11552
rect 22603 11512 23940 11540
rect 22603 11509 22615 11512
rect 22557 11503 22615 11509
rect 23934 11500 23940 11512
rect 23992 11500 23998 11552
rect 25222 11540 25228 11552
rect 25183 11512 25228 11540
rect 25222 11500 25228 11512
rect 25280 11500 25286 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 13173 11339 13231 11345
rect 13173 11336 13185 11339
rect 13044 11308 13185 11336
rect 13044 11296 13050 11308
rect 13173 11305 13185 11308
rect 13219 11305 13231 11339
rect 13538 11336 13544 11348
rect 13499 11308 13544 11336
rect 13173 11299 13231 11305
rect 13188 11268 13216 11299
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 14458 11336 14464 11348
rect 14419 11308 14464 11336
rect 14458 11296 14464 11308
rect 14516 11296 14522 11348
rect 16482 11296 16488 11348
rect 16540 11336 16546 11348
rect 16945 11339 17003 11345
rect 16945 11336 16957 11339
rect 16540 11308 16957 11336
rect 16540 11296 16546 11308
rect 16945 11305 16957 11308
rect 16991 11305 17003 11339
rect 16945 11299 17003 11305
rect 17034 11296 17040 11348
rect 17092 11336 17098 11348
rect 18831 11339 18889 11345
rect 18831 11336 18843 11339
rect 17092 11308 18843 11336
rect 17092 11296 17098 11308
rect 18831 11305 18843 11308
rect 18877 11305 18889 11339
rect 18831 11299 18889 11305
rect 19337 11339 19395 11345
rect 19337 11305 19349 11339
rect 19383 11336 19395 11339
rect 19518 11336 19524 11348
rect 19383 11308 19524 11336
rect 19383 11305 19395 11308
rect 19337 11299 19395 11305
rect 19518 11296 19524 11308
rect 19576 11296 19582 11348
rect 20349 11339 20407 11345
rect 20349 11305 20361 11339
rect 20395 11336 20407 11339
rect 20530 11336 20536 11348
rect 20395 11308 20536 11336
rect 20395 11305 20407 11308
rect 20349 11299 20407 11305
rect 20530 11296 20536 11308
rect 20588 11296 20594 11348
rect 23661 11339 23719 11345
rect 23661 11305 23673 11339
rect 23707 11336 23719 11339
rect 24210 11336 24216 11348
rect 23707 11308 24216 11336
rect 23707 11305 23719 11308
rect 23661 11299 23719 11305
rect 24210 11296 24216 11308
rect 24268 11336 24274 11348
rect 24268 11308 24716 11336
rect 24268 11296 24274 11308
rect 15013 11271 15071 11277
rect 15013 11268 15025 11271
rect 13188 11240 15025 11268
rect 15013 11237 15025 11240
rect 15059 11268 15071 11271
rect 15378 11268 15384 11280
rect 15059 11240 15384 11268
rect 15059 11237 15071 11240
rect 15013 11231 15071 11237
rect 15378 11228 15384 11240
rect 15436 11228 15442 11280
rect 19150 11228 19156 11280
rect 19208 11268 19214 11280
rect 20548 11268 20576 11296
rect 21637 11271 21695 11277
rect 19208 11240 20484 11268
rect 20548 11240 21404 11268
rect 19208 11228 19214 11240
rect 10134 11160 10140 11212
rect 10192 11200 10198 11212
rect 10321 11203 10379 11209
rect 10321 11200 10333 11203
rect 10192 11172 10333 11200
rect 10192 11160 10198 11172
rect 10321 11169 10333 11172
rect 10367 11169 10379 11203
rect 10321 11163 10379 11169
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11200 11023 11203
rect 12434 11200 12440 11212
rect 11011 11172 12440 11200
rect 11011 11169 11023 11172
rect 10965 11163 11023 11169
rect 12434 11160 12440 11172
rect 12492 11160 12498 11212
rect 13725 11203 13783 11209
rect 13725 11169 13737 11203
rect 13771 11169 13783 11203
rect 13725 11163 13783 11169
rect 14001 11203 14059 11209
rect 14001 11169 14013 11203
rect 14047 11200 14059 11203
rect 14182 11200 14188 11212
rect 14047 11172 14188 11200
rect 14047 11169 14059 11172
rect 14001 11163 14059 11169
rect 13740 11132 13768 11163
rect 14182 11160 14188 11172
rect 14240 11200 14246 11212
rect 14826 11200 14832 11212
rect 14240 11172 14832 11200
rect 14240 11160 14246 11172
rect 14826 11160 14832 11172
rect 14884 11160 14890 11212
rect 15470 11200 15476 11212
rect 15431 11172 15476 11200
rect 15470 11160 15476 11172
rect 15528 11160 15534 11212
rect 17126 11200 17132 11212
rect 17087 11172 17132 11200
rect 17126 11160 17132 11172
rect 17184 11160 17190 11212
rect 17681 11203 17739 11209
rect 17681 11169 17693 11203
rect 17727 11169 17739 11203
rect 18728 11203 18786 11209
rect 18728 11200 18740 11203
rect 17681 11163 17739 11169
rect 18524 11172 18740 11200
rect 14090 11132 14096 11144
rect 13740 11104 14096 11132
rect 14090 11092 14096 11104
rect 14148 11092 14154 11144
rect 16485 11135 16543 11141
rect 16485 11101 16497 11135
rect 16531 11132 16543 11135
rect 17402 11132 17408 11144
rect 16531 11104 17408 11132
rect 16531 11101 16543 11104
rect 16485 11095 16543 11101
rect 17402 11092 17408 11104
rect 17460 11132 17466 11144
rect 17696 11132 17724 11163
rect 17460 11104 17724 11132
rect 17460 11092 17466 11104
rect 15654 11024 15660 11076
rect 15712 11064 15718 11076
rect 18524 11073 18552 11172
rect 18728 11169 18740 11172
rect 18774 11169 18786 11203
rect 18728 11163 18786 11169
rect 19864 11203 19922 11209
rect 19864 11169 19876 11203
rect 19910 11200 19922 11203
rect 20456 11200 20484 11240
rect 20901 11203 20959 11209
rect 20901 11200 20913 11203
rect 19910 11172 20024 11200
rect 20456 11172 20913 11200
rect 19910 11169 19922 11172
rect 19864 11163 19922 11169
rect 19996 11076 20024 11172
rect 20901 11169 20913 11172
rect 20947 11200 20959 11203
rect 21266 11200 21272 11212
rect 20947 11172 21272 11200
rect 20947 11169 20959 11172
rect 20901 11163 20959 11169
rect 21266 11160 21272 11172
rect 21324 11160 21330 11212
rect 21376 11209 21404 11240
rect 21637 11237 21649 11271
rect 21683 11268 21695 11271
rect 22094 11268 22100 11280
rect 21683 11240 22100 11268
rect 21683 11237 21695 11240
rect 21637 11231 21695 11237
rect 22094 11228 22100 11240
rect 22152 11228 22158 11280
rect 22922 11228 22928 11280
rect 22980 11268 22986 11280
rect 24688 11277 24716 11308
rect 23062 11271 23120 11277
rect 23062 11268 23074 11271
rect 22980 11240 23074 11268
rect 22980 11228 22986 11240
rect 23062 11237 23074 11240
rect 23108 11237 23120 11271
rect 23062 11231 23120 11237
rect 24673 11271 24731 11277
rect 24673 11237 24685 11271
rect 24719 11237 24731 11271
rect 24673 11231 24731 11237
rect 21361 11203 21419 11209
rect 21361 11169 21373 11203
rect 21407 11200 21419 11203
rect 21542 11200 21548 11212
rect 21407 11172 21548 11200
rect 21407 11169 21419 11172
rect 21361 11163 21419 11169
rect 21542 11160 21548 11172
rect 21600 11160 21606 11212
rect 22738 11200 22744 11212
rect 22699 11172 22744 11200
rect 22738 11160 22744 11172
rect 22796 11160 22802 11212
rect 20073 11135 20131 11141
rect 20073 11101 20085 11135
rect 20119 11132 20131 11135
rect 21726 11132 21732 11144
rect 20119 11104 21732 11132
rect 20119 11101 20131 11104
rect 20073 11095 20131 11101
rect 21726 11092 21732 11104
rect 21784 11092 21790 11144
rect 24581 11135 24639 11141
rect 24581 11101 24593 11135
rect 24627 11132 24639 11135
rect 24670 11132 24676 11144
rect 24627 11104 24676 11132
rect 24627 11101 24639 11104
rect 24581 11095 24639 11101
rect 24670 11092 24676 11104
rect 24728 11092 24734 11144
rect 18509 11067 18567 11073
rect 18509 11064 18521 11067
rect 15712 11036 18521 11064
rect 15712 11024 15718 11036
rect 18509 11033 18521 11036
rect 18555 11033 18567 11067
rect 18509 11027 18567 11033
rect 19978 11024 19984 11076
rect 20036 11064 20042 11076
rect 25130 11064 25136 11076
rect 20036 11036 22140 11064
rect 25091 11036 25136 11064
rect 20036 11024 20042 11036
rect 15562 10996 15568 11008
rect 15523 10968 15568 10996
rect 15562 10956 15568 10968
rect 15620 10956 15626 11008
rect 17221 10999 17279 11005
rect 17221 10965 17233 10999
rect 17267 10996 17279 10999
rect 19058 10996 19064 11008
rect 17267 10968 19064 10996
rect 17267 10965 17279 10968
rect 17221 10959 17279 10965
rect 19058 10956 19064 10968
rect 19116 10956 19122 11008
rect 22002 10996 22008 11008
rect 21963 10968 22008 10996
rect 22002 10956 22008 10968
rect 22060 10956 22066 11008
rect 22112 10996 22140 11036
rect 25130 11024 25136 11036
rect 25188 11024 25194 11076
rect 25148 10996 25176 11024
rect 22112 10968 25176 10996
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 12713 10795 12771 10801
rect 12713 10761 12725 10795
rect 12759 10761 12771 10795
rect 14182 10792 14188 10804
rect 14143 10764 14188 10792
rect 12713 10755 12771 10761
rect 12728 10724 12756 10755
rect 14182 10752 14188 10764
rect 14240 10752 14246 10804
rect 15470 10752 15476 10804
rect 15528 10792 15534 10804
rect 15565 10795 15623 10801
rect 15565 10792 15577 10795
rect 15528 10764 15577 10792
rect 15528 10752 15534 10764
rect 15565 10761 15577 10764
rect 15611 10761 15623 10795
rect 15565 10755 15623 10761
rect 16853 10795 16911 10801
rect 16853 10761 16865 10795
rect 16899 10792 16911 10795
rect 16942 10792 16948 10804
rect 16899 10764 16948 10792
rect 16899 10761 16911 10764
rect 16853 10755 16911 10761
rect 16942 10752 16948 10764
rect 17000 10752 17006 10804
rect 19797 10795 19855 10801
rect 19797 10761 19809 10795
rect 19843 10792 19855 10795
rect 19978 10792 19984 10804
rect 19843 10764 19984 10792
rect 19843 10761 19855 10764
rect 19797 10755 19855 10761
rect 19978 10752 19984 10764
rect 20036 10752 20042 10804
rect 21266 10792 21272 10804
rect 21227 10764 21272 10792
rect 21266 10752 21272 10764
rect 21324 10752 21330 10804
rect 21542 10752 21548 10804
rect 21600 10792 21606 10804
rect 21637 10795 21695 10801
rect 21637 10792 21649 10795
rect 21600 10764 21649 10792
rect 21600 10752 21606 10764
rect 21637 10761 21649 10764
rect 21683 10761 21695 10795
rect 21637 10755 21695 10761
rect 22738 10752 22744 10804
rect 22796 10792 22802 10804
rect 23293 10795 23351 10801
rect 23293 10792 23305 10795
rect 22796 10764 23305 10792
rect 22796 10752 22802 10764
rect 23293 10761 23305 10764
rect 23339 10761 23351 10795
rect 23934 10792 23940 10804
rect 23895 10764 23940 10792
rect 23293 10755 23351 10761
rect 23934 10752 23940 10764
rect 23992 10752 23998 10804
rect 24670 10752 24676 10804
rect 24728 10792 24734 10804
rect 25501 10795 25559 10801
rect 25501 10792 25513 10795
rect 24728 10764 25513 10792
rect 24728 10752 24734 10764
rect 25501 10761 25513 10764
rect 25547 10761 25559 10795
rect 25501 10755 25559 10761
rect 14461 10727 14519 10733
rect 14461 10724 14473 10727
rect 12728 10696 14473 10724
rect 12728 10520 12756 10696
rect 14461 10693 14473 10696
rect 14507 10693 14519 10727
rect 14461 10687 14519 10693
rect 12897 10659 12955 10665
rect 12897 10625 12909 10659
rect 12943 10656 12955 10659
rect 12986 10656 12992 10668
rect 12943 10628 12992 10656
rect 12943 10625 12955 10628
rect 12897 10619 12955 10625
rect 12986 10616 12992 10628
rect 13044 10656 13050 10668
rect 13538 10656 13544 10668
rect 13044 10628 13544 10656
rect 13044 10616 13050 10628
rect 13538 10616 13544 10628
rect 13596 10616 13602 10668
rect 13218 10523 13276 10529
rect 13218 10520 13230 10523
rect 12728 10492 13230 10520
rect 13218 10489 13230 10492
rect 13264 10489 13276 10523
rect 14476 10520 14504 10687
rect 16206 10684 16212 10736
rect 16264 10724 16270 10736
rect 16669 10727 16727 10733
rect 16669 10724 16681 10727
rect 16264 10696 16681 10724
rect 16264 10684 16270 10696
rect 16669 10693 16681 10696
rect 16715 10693 16727 10727
rect 22922 10724 22928 10736
rect 16669 10687 16727 10693
rect 22065 10696 22928 10724
rect 14645 10659 14703 10665
rect 14645 10625 14657 10659
rect 14691 10656 14703 10659
rect 14734 10656 14740 10668
rect 14691 10628 14740 10656
rect 14691 10625 14703 10628
rect 14645 10619 14703 10625
rect 14734 10616 14740 10628
rect 14792 10616 14798 10668
rect 16390 10616 16396 10668
rect 16448 10656 16454 10668
rect 16761 10659 16819 10665
rect 16761 10656 16773 10659
rect 16448 10628 16773 10656
rect 16448 10616 16454 10628
rect 16761 10625 16773 10628
rect 16807 10625 16819 10659
rect 19150 10656 19156 10668
rect 16761 10619 16819 10625
rect 18708 10628 19156 10656
rect 16540 10591 16598 10597
rect 16540 10557 16552 10591
rect 16586 10588 16598 10591
rect 17402 10588 17408 10600
rect 16586 10560 17408 10588
rect 16586 10557 16598 10560
rect 16540 10551 16598 10557
rect 17402 10548 17408 10560
rect 17460 10548 17466 10600
rect 18708 10597 18736 10628
rect 19150 10616 19156 10628
rect 19208 10616 19214 10668
rect 21634 10616 21640 10668
rect 21692 10656 21698 10668
rect 22065 10656 22093 10696
rect 22922 10684 22928 10696
rect 22980 10684 22986 10736
rect 22646 10656 22652 10668
rect 21692 10628 22093 10656
rect 22607 10628 22652 10656
rect 21692 10616 21698 10628
rect 22646 10616 22652 10628
rect 22704 10616 22710 10668
rect 23952 10656 23980 10752
rect 25130 10724 25136 10736
rect 25091 10696 25136 10724
rect 25130 10684 25136 10696
rect 25188 10684 25194 10736
rect 24581 10659 24639 10665
rect 24581 10656 24593 10659
rect 23952 10628 24593 10656
rect 24581 10625 24593 10628
rect 24627 10625 24639 10659
rect 24581 10619 24639 10625
rect 18325 10591 18383 10597
rect 18325 10557 18337 10591
rect 18371 10588 18383 10591
rect 18693 10591 18751 10597
rect 18693 10588 18705 10591
rect 18371 10560 18705 10588
rect 18371 10557 18383 10560
rect 18325 10551 18383 10557
rect 18693 10557 18705 10560
rect 18739 10557 18751 10591
rect 18874 10588 18880 10600
rect 18835 10560 18880 10588
rect 18693 10551 18751 10557
rect 18874 10548 18880 10560
rect 18932 10548 18938 10600
rect 14966 10523 15024 10529
rect 14966 10520 14978 10523
rect 14476 10492 14978 10520
rect 13218 10483 13276 10489
rect 14966 10489 14978 10492
rect 15012 10520 15024 10523
rect 15838 10520 15844 10532
rect 15012 10492 15844 10520
rect 15012 10489 15024 10492
rect 14966 10483 15024 10489
rect 15838 10480 15844 10492
rect 15896 10480 15902 10532
rect 15933 10523 15991 10529
rect 15933 10489 15945 10523
rect 15979 10520 15991 10523
rect 16393 10523 16451 10529
rect 16393 10520 16405 10523
rect 15979 10492 16405 10520
rect 15979 10489 15991 10492
rect 15933 10483 15991 10489
rect 16393 10489 16405 10492
rect 16439 10520 16451 10523
rect 17126 10520 17132 10532
rect 16439 10492 17132 10520
rect 16439 10489 16451 10492
rect 16393 10483 16451 10489
rect 17126 10480 17132 10492
rect 17184 10520 17190 10532
rect 19150 10520 19156 10532
rect 17184 10492 17816 10520
rect 19111 10492 19156 10520
rect 17184 10480 17190 10492
rect 17788 10464 17816 10492
rect 19150 10480 19156 10492
rect 19208 10480 19214 10532
rect 20346 10520 20352 10532
rect 20307 10492 20352 10520
rect 20346 10480 20352 10492
rect 20404 10480 20410 10532
rect 20441 10523 20499 10529
rect 20441 10489 20453 10523
rect 20487 10489 20499 10523
rect 20441 10483 20499 10489
rect 20993 10523 21051 10529
rect 20993 10489 21005 10523
rect 21039 10520 21051 10523
rect 22002 10520 22008 10532
rect 21039 10492 22008 10520
rect 21039 10489 21051 10492
rect 20993 10483 21051 10489
rect 9582 10412 9588 10464
rect 9640 10452 9646 10464
rect 10134 10452 10140 10464
rect 9640 10424 10140 10452
rect 9640 10412 9646 10424
rect 10134 10412 10140 10424
rect 10192 10452 10198 10464
rect 10229 10455 10287 10461
rect 10229 10452 10241 10455
rect 10192 10424 10241 10452
rect 10192 10412 10198 10424
rect 10229 10421 10241 10424
rect 10275 10421 10287 10455
rect 10229 10415 10287 10421
rect 13814 10412 13820 10464
rect 13872 10452 13878 10464
rect 16206 10452 16212 10464
rect 13872 10424 13917 10452
rect 16167 10424 16212 10452
rect 13872 10412 13878 10424
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 17402 10452 17408 10464
rect 17363 10424 17408 10452
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 17770 10452 17776 10464
rect 17731 10424 17776 10452
rect 17770 10412 17776 10424
rect 17828 10412 17834 10464
rect 20070 10452 20076 10464
rect 20031 10424 20076 10452
rect 20070 10412 20076 10424
rect 20128 10452 20134 10464
rect 20456 10452 20484 10483
rect 22002 10480 22008 10492
rect 22060 10480 22066 10532
rect 22097 10523 22155 10529
rect 22097 10489 22109 10523
rect 22143 10489 22155 10523
rect 22097 10483 22155 10489
rect 24673 10523 24731 10529
rect 24673 10489 24685 10523
rect 24719 10489 24731 10523
rect 24673 10483 24731 10489
rect 20128 10424 20484 10452
rect 20128 10412 20134 10424
rect 21910 10412 21916 10464
rect 21968 10452 21974 10464
rect 22112 10452 22140 10483
rect 24394 10452 24400 10464
rect 21968 10424 22140 10452
rect 24355 10424 24400 10452
rect 21968 10412 21974 10424
rect 24394 10412 24400 10424
rect 24452 10452 24458 10464
rect 24688 10452 24716 10483
rect 24452 10424 24716 10452
rect 24452 10412 24458 10424
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 12986 10248 12992 10260
rect 12947 10220 12992 10248
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 14734 10248 14740 10260
rect 14695 10220 14740 10248
rect 14734 10208 14740 10220
rect 14792 10208 14798 10260
rect 15105 10251 15163 10257
rect 15105 10217 15117 10251
rect 15151 10248 15163 10251
rect 15378 10248 15384 10260
rect 15151 10220 15384 10248
rect 15151 10217 15163 10220
rect 15105 10211 15163 10217
rect 15378 10208 15384 10220
rect 15436 10208 15442 10260
rect 17678 10208 17684 10260
rect 17736 10248 17742 10260
rect 18322 10248 18328 10260
rect 17736 10220 18328 10248
rect 17736 10208 17742 10220
rect 18322 10208 18328 10220
rect 18380 10248 18386 10260
rect 18417 10251 18475 10257
rect 18417 10248 18429 10251
rect 18380 10220 18429 10248
rect 18380 10208 18386 10220
rect 18417 10217 18429 10220
rect 18463 10248 18475 10251
rect 18874 10248 18880 10260
rect 18463 10220 18880 10248
rect 18463 10217 18475 10220
rect 18417 10211 18475 10217
rect 18874 10208 18880 10220
rect 18932 10208 18938 10260
rect 19150 10208 19156 10260
rect 19208 10248 19214 10260
rect 19705 10251 19763 10257
rect 19705 10248 19717 10251
rect 19208 10220 19717 10248
rect 19208 10208 19214 10220
rect 19705 10217 19717 10220
rect 19751 10217 19763 10251
rect 20346 10248 20352 10260
rect 20307 10220 20352 10248
rect 19705 10211 19763 10217
rect 20346 10208 20352 10220
rect 20404 10208 20410 10260
rect 24394 10248 24400 10260
rect 24355 10220 24400 10248
rect 24394 10208 24400 10220
rect 24452 10208 24458 10260
rect 12894 10140 12900 10192
rect 12952 10180 12958 10192
rect 13265 10183 13323 10189
rect 13265 10180 13277 10183
rect 12952 10152 13277 10180
rect 12952 10140 12958 10152
rect 13265 10149 13277 10152
rect 13311 10180 13323 10183
rect 13814 10180 13820 10192
rect 13311 10152 13820 10180
rect 13311 10149 13323 10152
rect 13265 10143 13323 10149
rect 13814 10140 13820 10152
rect 13872 10140 13878 10192
rect 15473 10183 15531 10189
rect 15473 10149 15485 10183
rect 15519 10180 15531 10183
rect 15562 10180 15568 10192
rect 15519 10152 15568 10180
rect 15519 10149 15531 10152
rect 15473 10143 15531 10149
rect 15562 10140 15568 10152
rect 15620 10140 15626 10192
rect 17770 10180 17776 10192
rect 17731 10152 17776 10180
rect 17770 10140 17776 10152
rect 17828 10140 17834 10192
rect 17218 10112 17224 10124
rect 17179 10084 17224 10112
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 18690 10112 18696 10124
rect 18651 10084 18696 10112
rect 18690 10072 18696 10084
rect 18748 10072 18754 10124
rect 18892 10112 18920 10208
rect 22554 10180 22560 10192
rect 22515 10152 22560 10180
rect 22554 10140 22560 10152
rect 22612 10140 22618 10192
rect 22646 10140 22652 10192
rect 22704 10180 22710 10192
rect 23109 10183 23167 10189
rect 23109 10180 23121 10183
rect 22704 10152 23121 10180
rect 22704 10140 22710 10152
rect 23109 10149 23121 10152
rect 23155 10149 23167 10183
rect 23109 10143 23167 10149
rect 19153 10115 19211 10121
rect 19153 10112 19165 10115
rect 18892 10084 19165 10112
rect 19153 10081 19165 10084
rect 19199 10081 19211 10115
rect 24210 10112 24216 10124
rect 24171 10084 24216 10112
rect 19153 10075 19211 10081
rect 24210 10072 24216 10084
rect 24268 10112 24274 10124
rect 24949 10115 25007 10121
rect 24949 10112 24961 10115
rect 24268 10084 24961 10112
rect 24268 10072 24274 10084
rect 24949 10081 24961 10084
rect 24995 10081 25007 10115
rect 24949 10075 25007 10081
rect 12158 10004 12164 10056
rect 12216 10044 12222 10056
rect 13173 10047 13231 10053
rect 13173 10044 13185 10047
rect 12216 10016 13185 10044
rect 12216 10004 12222 10016
rect 13173 10013 13185 10016
rect 13219 10013 13231 10047
rect 15378 10044 15384 10056
rect 15339 10016 15384 10044
rect 13173 10007 13231 10013
rect 15378 10004 15384 10016
rect 15436 10004 15442 10056
rect 15654 10044 15660 10056
rect 15615 10016 15660 10044
rect 15654 10004 15660 10016
rect 15712 10004 15718 10056
rect 19429 10047 19487 10053
rect 19429 10013 19441 10047
rect 19475 10044 19487 10047
rect 20346 10044 20352 10056
rect 19475 10016 20352 10044
rect 19475 10013 19487 10016
rect 19429 10007 19487 10013
rect 20346 10004 20352 10016
rect 20404 10004 20410 10056
rect 21361 10047 21419 10053
rect 21361 10013 21373 10047
rect 21407 10044 21419 10047
rect 22465 10047 22523 10053
rect 22465 10044 22477 10047
rect 21407 10016 22477 10044
rect 21407 10013 21419 10016
rect 21361 10007 21419 10013
rect 22465 10013 22477 10016
rect 22511 10044 22523 10047
rect 22738 10044 22744 10056
rect 22511 10016 22744 10044
rect 22511 10013 22523 10016
rect 22465 10007 22523 10013
rect 22738 10004 22744 10016
rect 22796 10004 22802 10056
rect 13722 9976 13728 9988
rect 13683 9948 13728 9976
rect 13722 9936 13728 9948
rect 13780 9936 13786 9988
rect 14182 9908 14188 9920
rect 14143 9880 14188 9908
rect 14182 9868 14188 9880
rect 14240 9868 14246 9920
rect 16390 9908 16396 9920
rect 16351 9880 16396 9908
rect 16390 9868 16396 9880
rect 16448 9868 16454 9920
rect 21910 9908 21916 9920
rect 21871 9880 21916 9908
rect 21910 9868 21916 9880
rect 21968 9868 21974 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 6822 9664 6828 9716
rect 6880 9704 6886 9716
rect 12158 9704 12164 9716
rect 6880 9676 12164 9704
rect 6880 9664 6886 9676
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 12894 9704 12900 9716
rect 12855 9676 12900 9704
rect 12894 9664 12900 9676
rect 12952 9664 12958 9716
rect 14829 9707 14887 9713
rect 14829 9673 14841 9707
rect 14875 9704 14887 9707
rect 15378 9704 15384 9716
rect 14875 9676 15384 9704
rect 14875 9673 14887 9676
rect 14829 9667 14887 9673
rect 15378 9664 15384 9676
rect 15436 9664 15442 9716
rect 15562 9664 15568 9716
rect 15620 9704 15626 9716
rect 15933 9707 15991 9713
rect 15933 9704 15945 9707
rect 15620 9676 15945 9704
rect 15620 9664 15626 9676
rect 15933 9673 15945 9676
rect 15979 9673 15991 9707
rect 18322 9704 18328 9716
rect 18283 9676 18328 9704
rect 15933 9667 15991 9673
rect 18322 9664 18328 9676
rect 18380 9664 18386 9716
rect 20346 9704 20352 9716
rect 20307 9676 20352 9704
rect 20346 9664 20352 9676
rect 20404 9704 20410 9716
rect 22738 9704 22744 9716
rect 20404 9676 20944 9704
rect 22699 9676 22744 9704
rect 20404 9664 20410 9676
rect 12342 9596 12348 9648
rect 12400 9636 12406 9648
rect 16206 9636 16212 9648
rect 12400 9608 16212 9636
rect 12400 9596 12406 9608
rect 16206 9596 16212 9608
rect 16264 9596 16270 9648
rect 13265 9571 13323 9577
rect 13265 9537 13277 9571
rect 13311 9568 13323 9571
rect 13538 9568 13544 9580
rect 13311 9540 13544 9568
rect 13311 9537 13323 9540
rect 13265 9531 13323 9537
rect 13538 9528 13544 9540
rect 13596 9528 13602 9580
rect 15654 9568 15660 9580
rect 15615 9540 15660 9568
rect 15654 9528 15660 9540
rect 15712 9528 15718 9580
rect 19150 9568 19156 9580
rect 19111 9540 19156 9568
rect 19150 9528 19156 9540
rect 19208 9528 19214 9580
rect 20916 9577 20944 9676
rect 22738 9664 22744 9676
rect 22796 9664 22802 9716
rect 24029 9707 24087 9713
rect 24029 9673 24041 9707
rect 24075 9704 24087 9707
rect 24210 9704 24216 9716
rect 24075 9676 24216 9704
rect 24075 9673 24087 9676
rect 24029 9667 24087 9673
rect 24210 9664 24216 9676
rect 24268 9664 24274 9716
rect 24765 9707 24823 9713
rect 24765 9673 24777 9707
rect 24811 9704 24823 9707
rect 24946 9704 24952 9716
rect 24811 9676 24952 9704
rect 24811 9673 24823 9676
rect 24765 9667 24823 9673
rect 24946 9664 24952 9676
rect 25004 9664 25010 9716
rect 21726 9596 21732 9648
rect 21784 9636 21790 9648
rect 21784 9608 23474 9636
rect 21784 9596 21790 9608
rect 20901 9571 20959 9577
rect 20901 9537 20913 9571
rect 20947 9537 20959 9571
rect 20901 9531 20959 9537
rect 21821 9503 21879 9509
rect 21821 9469 21833 9503
rect 21867 9500 21879 9503
rect 21910 9500 21916 9512
rect 21867 9472 21916 9500
rect 21867 9469 21879 9472
rect 21821 9463 21879 9469
rect 21910 9460 21916 9472
rect 21968 9500 21974 9512
rect 23014 9500 23020 9512
rect 21968 9472 23020 9500
rect 21968 9460 21974 9472
rect 23014 9460 23020 9472
rect 23072 9460 23078 9512
rect 23446 9500 23474 9608
rect 24581 9503 24639 9509
rect 24581 9500 24593 9503
rect 23446 9472 24593 9500
rect 24581 9469 24593 9472
rect 24627 9500 24639 9503
rect 25133 9503 25191 9509
rect 25133 9500 25145 9503
rect 24627 9472 25145 9500
rect 24627 9469 24639 9472
rect 24581 9463 24639 9469
rect 25133 9469 25145 9472
rect 25179 9469 25191 9503
rect 25133 9463 25191 9469
rect 13449 9435 13507 9441
rect 13449 9401 13461 9435
rect 13495 9401 13507 9435
rect 13449 9395 13507 9401
rect 13464 9364 13492 9395
rect 13538 9392 13544 9444
rect 13596 9432 13602 9444
rect 13596 9404 13641 9432
rect 13596 9392 13602 9404
rect 13722 9392 13728 9444
rect 13780 9432 13786 9444
rect 14093 9435 14151 9441
rect 14093 9432 14105 9435
rect 13780 9404 14105 9432
rect 13780 9392 13786 9404
rect 14093 9401 14105 9404
rect 14139 9432 14151 9435
rect 15010 9432 15016 9444
rect 14139 9404 15016 9432
rect 14139 9401 14151 9404
rect 14093 9395 14151 9401
rect 15010 9392 15016 9404
rect 15068 9392 15074 9444
rect 15102 9392 15108 9444
rect 15160 9432 15166 9444
rect 15470 9432 15476 9444
rect 15160 9404 15476 9432
rect 15160 9392 15166 9404
rect 15470 9392 15476 9404
rect 15528 9392 15534 9444
rect 18601 9435 18659 9441
rect 18601 9432 18613 9435
rect 16085 9404 18613 9432
rect 14458 9364 14464 9376
rect 13464 9336 14464 9364
rect 14458 9324 14464 9336
rect 14516 9324 14522 9376
rect 14550 9324 14556 9376
rect 14608 9364 14614 9376
rect 16085 9364 16113 9404
rect 18601 9401 18613 9404
rect 18647 9432 18659 9435
rect 18690 9432 18696 9444
rect 18647 9404 18696 9432
rect 18647 9401 18659 9404
rect 18601 9395 18659 9401
rect 18690 9392 18696 9404
rect 18748 9392 18754 9444
rect 19474 9435 19532 9441
rect 19474 9432 19486 9435
rect 18984 9404 19486 9432
rect 14608 9336 16113 9364
rect 17129 9367 17187 9373
rect 14608 9324 14614 9336
rect 17129 9333 17141 9367
rect 17175 9364 17187 9367
rect 17218 9364 17224 9376
rect 17175 9336 17224 9364
rect 17175 9333 17187 9336
rect 17129 9327 17187 9333
rect 17218 9324 17224 9336
rect 17276 9324 17282 9376
rect 17862 9324 17868 9376
rect 17920 9364 17926 9376
rect 18984 9373 19012 9404
rect 19474 9401 19486 9404
rect 19520 9432 19532 9435
rect 20717 9435 20775 9441
rect 20717 9432 20729 9435
rect 19520 9404 20729 9432
rect 19520 9401 19532 9404
rect 19474 9395 19532 9401
rect 20717 9401 20729 9404
rect 20763 9432 20775 9435
rect 21222 9435 21280 9441
rect 21222 9432 21234 9435
rect 20763 9404 21234 9432
rect 20763 9401 20775 9404
rect 20717 9395 20775 9401
rect 21222 9401 21234 9404
rect 21268 9432 21280 9435
rect 21542 9432 21548 9444
rect 21268 9404 21548 9432
rect 21268 9401 21280 9404
rect 21222 9395 21280 9401
rect 21542 9392 21548 9404
rect 21600 9392 21606 9444
rect 18969 9367 19027 9373
rect 18969 9364 18981 9367
rect 17920 9336 18981 9364
rect 17920 9324 17926 9336
rect 18969 9333 18981 9336
rect 19015 9333 19027 9367
rect 18969 9327 19027 9333
rect 19334 9324 19340 9376
rect 19392 9364 19398 9376
rect 20070 9364 20076 9376
rect 19392 9336 20076 9364
rect 19392 9324 19398 9336
rect 20070 9324 20076 9336
rect 20128 9324 20134 9376
rect 22465 9367 22523 9373
rect 22465 9333 22477 9367
rect 22511 9364 22523 9367
rect 22554 9364 22560 9376
rect 22511 9336 22560 9364
rect 22511 9333 22523 9336
rect 22465 9327 22523 9333
rect 22554 9324 22560 9336
rect 22612 9364 22618 9376
rect 22738 9364 22744 9376
rect 22612 9336 22744 9364
rect 22612 9324 22618 9336
rect 22738 9324 22744 9336
rect 22796 9324 22802 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 13449 9163 13507 9169
rect 13449 9129 13461 9163
rect 13495 9160 13507 9163
rect 13538 9160 13544 9172
rect 13495 9132 13544 9160
rect 13495 9129 13507 9132
rect 13449 9123 13507 9129
rect 13538 9120 13544 9132
rect 13596 9120 13602 9172
rect 14921 9163 14979 9169
rect 14921 9129 14933 9163
rect 14967 9160 14979 9163
rect 15102 9160 15108 9172
rect 14967 9132 15108 9160
rect 14967 9129 14979 9132
rect 14921 9123 14979 9129
rect 15102 9120 15108 9132
rect 15160 9120 15166 9172
rect 15289 9163 15347 9169
rect 15289 9129 15301 9163
rect 15335 9160 15347 9163
rect 15378 9160 15384 9172
rect 15335 9132 15384 9160
rect 15335 9129 15347 9132
rect 15289 9123 15347 9129
rect 15378 9120 15384 9132
rect 15436 9120 15442 9172
rect 17310 9120 17316 9172
rect 17368 9160 17374 9172
rect 17497 9163 17555 9169
rect 17497 9160 17509 9163
rect 17368 9132 17509 9160
rect 17368 9120 17374 9132
rect 17497 9129 17509 9132
rect 17543 9129 17555 9163
rect 24118 9160 24124 9172
rect 24079 9132 24124 9160
rect 17497 9123 17555 9129
rect 24118 9120 24124 9132
rect 24176 9120 24182 9172
rect 24762 9160 24768 9172
rect 24723 9132 24768 9160
rect 24762 9120 24768 9132
rect 24820 9120 24826 9172
rect 15010 9052 15016 9104
rect 15068 9092 15074 9104
rect 15749 9095 15807 9101
rect 15749 9092 15761 9095
rect 15068 9064 15761 9092
rect 15068 9052 15074 9064
rect 15749 9061 15761 9064
rect 15795 9061 15807 9095
rect 15749 9055 15807 9061
rect 19981 9095 20039 9101
rect 19981 9061 19993 9095
rect 20027 9092 20039 9095
rect 21266 9092 21272 9104
rect 20027 9064 21272 9092
rect 20027 9061 20039 9064
rect 19981 9055 20039 9061
rect 21266 9052 21272 9064
rect 21324 9092 21330 9104
rect 21361 9095 21419 9101
rect 21361 9092 21373 9095
rect 21324 9064 21373 9092
rect 21324 9052 21330 9064
rect 21361 9061 21373 9064
rect 21407 9061 21419 9095
rect 21361 9055 21419 9061
rect 21913 9095 21971 9101
rect 21913 9061 21925 9095
rect 21959 9092 21971 9095
rect 22002 9092 22008 9104
rect 21959 9064 22008 9092
rect 21959 9061 21971 9064
rect 21913 9055 21971 9061
rect 22002 9052 22008 9064
rect 22060 9052 22066 9104
rect 22738 9092 22744 9104
rect 22699 9064 22744 9092
rect 22738 9052 22744 9064
rect 22796 9052 22802 9104
rect 12894 8984 12900 9036
rect 12952 9024 12958 9036
rect 13265 9027 13323 9033
rect 13265 9024 13277 9027
rect 12952 8996 13277 9024
rect 12952 8984 12958 8996
rect 13265 8993 13277 8996
rect 13311 8993 13323 9027
rect 17218 9024 17224 9036
rect 17179 8996 17224 9024
rect 13265 8987 13323 8993
rect 17218 8984 17224 8996
rect 17276 8984 17282 9036
rect 17402 9024 17408 9036
rect 17363 8996 17408 9024
rect 17402 8984 17408 8996
rect 17460 8984 17466 9036
rect 19334 9024 19340 9036
rect 19295 8996 19340 9024
rect 19334 8984 19340 8996
rect 19392 8984 19398 9036
rect 23014 9024 23020 9036
rect 22975 8996 23020 9024
rect 23014 8984 23020 8996
rect 23072 8984 23078 9036
rect 24581 9027 24639 9033
rect 24581 8993 24593 9027
rect 24627 9024 24639 9027
rect 25038 9024 25044 9036
rect 24627 8996 25044 9024
rect 24627 8993 24639 8996
rect 24581 8987 24639 8993
rect 25038 8984 25044 8996
rect 25096 8984 25102 9036
rect 21269 8959 21327 8965
rect 21269 8925 21281 8959
rect 21315 8956 21327 8959
rect 21358 8956 21364 8968
rect 21315 8928 21364 8956
rect 21315 8925 21327 8928
rect 21269 8919 21327 8925
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 18138 8820 18144 8832
rect 18099 8792 18144 8820
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 12894 8576 12900 8628
rect 12952 8616 12958 8628
rect 13173 8619 13231 8625
rect 13173 8616 13185 8619
rect 12952 8588 13185 8616
rect 12952 8576 12958 8588
rect 13173 8585 13185 8588
rect 13219 8585 13231 8619
rect 13173 8579 13231 8585
rect 14093 8619 14151 8625
rect 14093 8585 14105 8619
rect 14139 8616 14151 8619
rect 14182 8616 14188 8628
rect 14139 8588 14188 8616
rect 14139 8585 14151 8588
rect 14093 8579 14151 8585
rect 14182 8576 14188 8588
rect 14240 8576 14246 8628
rect 14550 8576 14556 8628
rect 14608 8616 14614 8628
rect 15013 8619 15071 8625
rect 15013 8616 15025 8619
rect 14608 8588 15025 8616
rect 14608 8576 14614 8588
rect 15013 8585 15025 8588
rect 15059 8585 15071 8619
rect 19334 8616 19340 8628
rect 19295 8588 19340 8616
rect 15013 8579 15071 8585
rect 5166 8372 5172 8424
rect 5224 8412 5230 8424
rect 10778 8412 10784 8424
rect 5224 8384 10784 8412
rect 5224 8372 5230 8384
rect 10778 8372 10784 8384
rect 10836 8412 10842 8424
rect 13909 8415 13967 8421
rect 13909 8412 13921 8415
rect 10836 8384 13921 8412
rect 10836 8372 10842 8384
rect 13909 8381 13921 8384
rect 13955 8412 13967 8415
rect 14369 8415 14427 8421
rect 14369 8412 14381 8415
rect 13955 8384 14381 8412
rect 13955 8381 13967 8384
rect 13909 8375 13967 8381
rect 14369 8381 14381 8384
rect 14415 8381 14427 8415
rect 15028 8412 15056 8579
rect 19334 8576 19340 8588
rect 19392 8576 19398 8628
rect 21266 8616 21272 8628
rect 21227 8588 21272 8616
rect 21266 8576 21272 8588
rect 21324 8576 21330 8628
rect 21358 8576 21364 8628
rect 21416 8616 21422 8628
rect 21637 8619 21695 8625
rect 21637 8616 21649 8619
rect 21416 8588 21649 8616
rect 21416 8576 21422 8588
rect 21637 8585 21649 8588
rect 21683 8585 21695 8619
rect 21637 8579 21695 8585
rect 22695 8619 22753 8625
rect 22695 8585 22707 8619
rect 22741 8616 22753 8619
rect 23474 8616 23480 8628
rect 22741 8588 23480 8616
rect 22741 8585 22753 8588
rect 22695 8579 22753 8585
rect 23474 8576 23480 8588
rect 23532 8576 23538 8628
rect 26145 8619 26203 8625
rect 26145 8585 26157 8619
rect 26191 8616 26203 8619
rect 27614 8616 27620 8628
rect 26191 8588 27620 8616
rect 26191 8585 26203 8588
rect 26145 8579 26203 8585
rect 17218 8508 17224 8560
rect 17276 8548 17282 8560
rect 17681 8551 17739 8557
rect 17681 8548 17693 8551
rect 17276 8520 17693 8548
rect 17276 8508 17282 8520
rect 17681 8517 17693 8520
rect 17727 8548 17739 8551
rect 22462 8548 22468 8560
rect 17727 8520 22468 8548
rect 17727 8517 17739 8520
rect 17681 8511 17739 8517
rect 22462 8508 22468 8520
rect 22520 8508 22526 8560
rect 23014 8548 23020 8560
rect 22975 8520 23020 8548
rect 23014 8508 23020 8520
rect 23072 8508 23078 8560
rect 23106 8508 23112 8560
rect 23164 8548 23170 8560
rect 23845 8551 23903 8557
rect 23845 8548 23857 8551
rect 23164 8520 23857 8548
rect 23164 8508 23170 8520
rect 23845 8517 23857 8520
rect 23891 8548 23903 8551
rect 24210 8548 24216 8560
rect 23891 8520 24216 8548
rect 23891 8517 23903 8520
rect 23845 8511 23903 8517
rect 24210 8508 24216 8520
rect 24268 8508 24274 8560
rect 17313 8483 17371 8489
rect 17313 8449 17325 8483
rect 17359 8480 17371 8483
rect 17402 8480 17408 8492
rect 17359 8452 17408 8480
rect 17359 8449 17371 8452
rect 17313 8443 17371 8449
rect 17402 8440 17408 8452
rect 17460 8480 17466 8492
rect 18966 8480 18972 8492
rect 17460 8452 18972 8480
rect 17460 8440 17466 8452
rect 18966 8440 18972 8452
rect 19024 8440 19030 8492
rect 24118 8480 24124 8492
rect 24079 8452 24124 8480
rect 24118 8440 24124 8452
rect 24176 8440 24182 8492
rect 24302 8440 24308 8492
rect 24360 8480 24366 8492
rect 24397 8483 24455 8489
rect 24397 8480 24409 8483
rect 24360 8452 24409 8480
rect 24360 8440 24366 8452
rect 24397 8449 24409 8452
rect 24443 8449 24455 8483
rect 24397 8443 24455 8449
rect 15197 8415 15255 8421
rect 15197 8412 15209 8415
rect 15028 8384 15209 8412
rect 14369 8375 14427 8381
rect 15197 8381 15209 8384
rect 15243 8381 15255 8415
rect 15197 8375 15255 8381
rect 15286 8372 15292 8424
rect 15344 8412 15350 8424
rect 15657 8415 15715 8421
rect 15657 8412 15669 8415
rect 15344 8384 15669 8412
rect 15344 8372 15350 8384
rect 15657 8381 15669 8384
rect 15703 8381 15715 8415
rect 18138 8412 18144 8424
rect 18099 8384 18144 8412
rect 15657 8375 15715 8381
rect 18138 8372 18144 8384
rect 18196 8372 18202 8424
rect 18690 8372 18696 8424
rect 18748 8412 18754 8424
rect 20073 8415 20131 8421
rect 20073 8412 20085 8415
rect 18748 8384 20085 8412
rect 18748 8372 18754 8384
rect 20073 8381 20085 8384
rect 20119 8412 20131 8415
rect 20257 8415 20315 8421
rect 20257 8412 20269 8415
rect 20119 8384 20269 8412
rect 20119 8381 20131 8384
rect 20073 8375 20131 8381
rect 20257 8381 20269 8384
rect 20303 8381 20315 8415
rect 20714 8412 20720 8424
rect 20675 8384 20720 8412
rect 20257 8375 20315 8381
rect 20714 8372 20720 8384
rect 20772 8372 20778 8424
rect 22624 8415 22682 8421
rect 22624 8381 22636 8415
rect 22670 8381 22682 8415
rect 22624 8375 22682 8381
rect 25660 8415 25718 8421
rect 25660 8381 25672 8415
rect 25706 8412 25718 8415
rect 26160 8412 26188 8579
rect 27614 8576 27620 8588
rect 27672 8576 27678 8628
rect 25706 8384 26188 8412
rect 25706 8381 25718 8384
rect 25660 8375 25718 8381
rect 15930 8344 15936 8356
rect 15891 8316 15936 8344
rect 15930 8304 15936 8316
rect 15988 8304 15994 8356
rect 18782 8344 18788 8356
rect 18743 8316 18788 8344
rect 18782 8304 18788 8316
rect 18840 8304 18846 8356
rect 20993 8347 21051 8353
rect 20993 8313 21005 8347
rect 21039 8344 21051 8347
rect 21726 8344 21732 8356
rect 21039 8316 21732 8344
rect 21039 8313 21051 8316
rect 20993 8307 21051 8313
rect 21726 8304 21732 8316
rect 21784 8304 21790 8356
rect 22639 8344 22667 8375
rect 23385 8347 23443 8353
rect 23385 8344 23397 8347
rect 22639 8316 23397 8344
rect 23385 8313 23397 8316
rect 23431 8313 23443 8347
rect 23385 8307 23443 8313
rect 23400 8276 23428 8307
rect 24210 8304 24216 8356
rect 24268 8344 24274 8356
rect 24268 8316 24313 8344
rect 24268 8304 24274 8316
rect 24394 8276 24400 8288
rect 23400 8248 24400 8276
rect 24394 8236 24400 8248
rect 24452 8236 24458 8288
rect 25038 8276 25044 8288
rect 24999 8248 25044 8276
rect 25038 8236 25044 8248
rect 25096 8236 25102 8288
rect 25130 8236 25136 8288
rect 25188 8276 25194 8288
rect 25731 8279 25789 8285
rect 25731 8276 25743 8279
rect 25188 8248 25743 8276
rect 25188 8236 25194 8248
rect 25731 8245 25743 8248
rect 25777 8245 25789 8279
rect 25731 8239 25789 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 15286 8032 15292 8084
rect 15344 8072 15350 8084
rect 15473 8075 15531 8081
rect 15473 8072 15485 8075
rect 15344 8044 15485 8072
rect 15344 8032 15350 8044
rect 15473 8041 15485 8044
rect 15519 8041 15531 8075
rect 15473 8035 15531 8041
rect 16206 8032 16212 8084
rect 16264 8072 16270 8084
rect 16945 8075 17003 8081
rect 16945 8072 16957 8075
rect 16264 8044 16957 8072
rect 16264 8032 16270 8044
rect 16945 8041 16957 8044
rect 16991 8041 17003 8075
rect 17862 8072 17868 8084
rect 17823 8044 17868 8072
rect 16945 8035 17003 8041
rect 17862 8032 17868 8044
rect 17920 8032 17926 8084
rect 18138 8032 18144 8084
rect 18196 8072 18202 8084
rect 18417 8075 18475 8081
rect 18417 8072 18429 8075
rect 18196 8044 18429 8072
rect 18196 8032 18202 8044
rect 18417 8041 18429 8044
rect 18463 8041 18475 8075
rect 18417 8035 18475 8041
rect 15838 7964 15844 8016
rect 15896 8004 15902 8016
rect 16070 8007 16128 8013
rect 16070 8004 16082 8007
rect 15896 7976 16082 8004
rect 15896 7964 15902 7976
rect 16070 7973 16082 7976
rect 16116 7973 16128 8007
rect 16070 7967 16128 7973
rect 21542 7964 21548 8016
rect 21600 8004 21606 8016
rect 22050 8007 22108 8013
rect 22050 8004 22062 8007
rect 21600 7976 22062 8004
rect 21600 7964 21606 7976
rect 22050 7973 22062 7976
rect 22096 7973 22108 8007
rect 22050 7967 22108 7973
rect 23934 7964 23940 8016
rect 23992 8004 23998 8016
rect 24213 8007 24271 8013
rect 24213 8004 24225 8007
rect 23992 7976 24225 8004
rect 23992 7964 23998 7976
rect 24213 7973 24225 7976
rect 24259 7973 24271 8007
rect 24213 7967 24271 7973
rect 15930 7896 15936 7948
rect 15988 7936 15994 7948
rect 17402 7936 17408 7948
rect 15988 7908 17408 7936
rect 15988 7896 15994 7908
rect 17402 7896 17408 7908
rect 17460 7936 17466 7948
rect 17497 7939 17555 7945
rect 17497 7936 17509 7939
rect 17460 7908 17509 7936
rect 17460 7896 17466 7908
rect 17497 7905 17509 7908
rect 17543 7905 17555 7939
rect 19242 7936 19248 7948
rect 19203 7908 19248 7936
rect 17497 7899 17555 7905
rect 19242 7896 19248 7908
rect 19300 7896 19306 7948
rect 19705 7939 19763 7945
rect 19705 7905 19717 7939
rect 19751 7936 19763 7939
rect 20257 7939 20315 7945
rect 20257 7936 20269 7939
rect 19751 7908 20269 7936
rect 19751 7905 19763 7908
rect 19705 7899 19763 7905
rect 20257 7905 20269 7908
rect 20303 7936 20315 7939
rect 20714 7936 20720 7948
rect 20303 7908 20720 7936
rect 20303 7905 20315 7908
rect 20257 7899 20315 7905
rect 15746 7868 15752 7880
rect 15707 7840 15752 7868
rect 15746 7828 15752 7840
rect 15804 7828 15810 7880
rect 16850 7828 16856 7880
rect 16908 7868 16914 7880
rect 19518 7868 19524 7880
rect 16908 7840 19524 7868
rect 16908 7828 16914 7840
rect 19518 7828 19524 7840
rect 19576 7868 19582 7880
rect 19720 7868 19748 7899
rect 20714 7896 20720 7908
rect 20772 7896 20778 7948
rect 19576 7840 19748 7868
rect 19981 7871 20039 7877
rect 19576 7828 19582 7840
rect 19981 7837 19993 7871
rect 20027 7868 20039 7871
rect 21174 7868 21180 7880
rect 20027 7840 21180 7868
rect 20027 7837 20039 7840
rect 19981 7831 20039 7837
rect 21174 7828 21180 7840
rect 21232 7828 21238 7880
rect 21726 7868 21732 7880
rect 21687 7840 21732 7868
rect 21726 7828 21732 7840
rect 21784 7828 21790 7880
rect 24118 7868 24124 7880
rect 24079 7840 24124 7868
rect 24118 7828 24124 7840
rect 24176 7828 24182 7880
rect 24394 7868 24400 7880
rect 24355 7840 24400 7868
rect 24394 7828 24400 7840
rect 24452 7868 24458 7880
rect 24452 7840 24716 7868
rect 24452 7828 24458 7840
rect 24688 7812 24716 7840
rect 24670 7760 24676 7812
rect 24728 7760 24734 7812
rect 16666 7732 16672 7744
rect 16627 7704 16672 7732
rect 16666 7692 16672 7704
rect 16724 7692 16730 7744
rect 18230 7692 18236 7744
rect 18288 7732 18294 7744
rect 18693 7735 18751 7741
rect 18693 7732 18705 7735
rect 18288 7704 18705 7732
rect 18288 7692 18294 7704
rect 18693 7701 18705 7704
rect 18739 7701 18751 7735
rect 22646 7732 22652 7744
rect 22607 7704 22652 7732
rect 18693 7695 18751 7701
rect 22646 7692 22652 7704
rect 22704 7692 22710 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 15838 7528 15844 7540
rect 15799 7500 15844 7528
rect 15838 7488 15844 7500
rect 15896 7528 15902 7540
rect 17497 7531 17555 7537
rect 17497 7528 17509 7531
rect 15896 7500 17509 7528
rect 15896 7488 15902 7500
rect 17497 7497 17509 7500
rect 17543 7528 17555 7531
rect 17862 7528 17868 7540
rect 17543 7500 17868 7528
rect 17543 7497 17555 7500
rect 17497 7491 17555 7497
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 18782 7488 18788 7540
rect 18840 7528 18846 7540
rect 19429 7531 19487 7537
rect 19429 7528 19441 7531
rect 18840 7500 19441 7528
rect 18840 7488 18846 7500
rect 19429 7497 19441 7500
rect 19475 7528 19487 7531
rect 19794 7528 19800 7540
rect 19475 7500 19800 7528
rect 19475 7497 19487 7500
rect 19429 7491 19487 7497
rect 19794 7488 19800 7500
rect 19852 7488 19858 7540
rect 21174 7528 21180 7540
rect 21135 7500 21180 7528
rect 21174 7488 21180 7500
rect 21232 7528 21238 7540
rect 22649 7531 22707 7537
rect 21232 7500 21772 7528
rect 21232 7488 21238 7500
rect 14182 7420 14188 7472
rect 14240 7460 14246 7472
rect 14737 7463 14795 7469
rect 14737 7460 14749 7463
rect 14240 7432 14749 7460
rect 14240 7420 14246 7432
rect 14737 7429 14749 7432
rect 14783 7460 14795 7463
rect 19153 7463 19211 7469
rect 19153 7460 19165 7463
rect 14783 7432 19165 7460
rect 14783 7429 14795 7432
rect 14737 7423 14795 7429
rect 15120 7333 15148 7432
rect 19153 7429 19165 7432
rect 19199 7460 19211 7463
rect 19242 7460 19248 7472
rect 19199 7432 19248 7460
rect 19199 7429 19211 7432
rect 19153 7423 19211 7429
rect 19242 7420 19248 7432
rect 19300 7420 19306 7472
rect 21542 7460 21548 7472
rect 21503 7432 21548 7460
rect 21542 7420 21548 7432
rect 21600 7420 21606 7472
rect 15565 7395 15623 7401
rect 15565 7361 15577 7395
rect 15611 7392 15623 7395
rect 15746 7392 15752 7404
rect 15611 7364 15752 7392
rect 15611 7361 15623 7364
rect 15565 7355 15623 7361
rect 15746 7352 15752 7364
rect 15804 7352 15810 7404
rect 16206 7352 16212 7404
rect 16264 7392 16270 7404
rect 16485 7395 16543 7401
rect 16485 7392 16497 7395
rect 16264 7364 16497 7392
rect 16264 7352 16270 7364
rect 16485 7361 16497 7364
rect 16531 7361 16543 7395
rect 16485 7355 16543 7361
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7392 17187 7395
rect 18141 7395 18199 7401
rect 18141 7392 18153 7395
rect 17175 7364 18153 7392
rect 17175 7361 17187 7364
rect 17129 7355 17187 7361
rect 18141 7361 18153 7364
rect 18187 7392 18199 7395
rect 18230 7392 18236 7404
rect 18187 7364 18236 7392
rect 18187 7361 18199 7364
rect 18141 7355 18199 7361
rect 18230 7352 18236 7364
rect 18288 7352 18294 7404
rect 21744 7401 21772 7500
rect 22649 7497 22661 7531
rect 22695 7528 22707 7531
rect 23106 7528 23112 7540
rect 22695 7500 23112 7528
rect 22695 7497 22707 7500
rect 22649 7491 22707 7497
rect 23106 7488 23112 7500
rect 23164 7488 23170 7540
rect 23474 7488 23480 7540
rect 23532 7528 23538 7540
rect 24118 7528 24124 7540
rect 23532 7500 24124 7528
rect 23532 7488 23538 7500
rect 24118 7488 24124 7500
rect 24176 7488 24182 7540
rect 25406 7488 25412 7540
rect 25464 7528 25470 7540
rect 25731 7531 25789 7537
rect 25731 7528 25743 7531
rect 25464 7500 25743 7528
rect 25464 7488 25470 7500
rect 25731 7497 25743 7500
rect 25777 7497 25789 7531
rect 25731 7491 25789 7497
rect 26145 7531 26203 7537
rect 26145 7497 26157 7531
rect 26191 7528 26203 7531
rect 27614 7528 27620 7540
rect 26191 7500 27620 7528
rect 26191 7497 26203 7500
rect 26145 7491 26203 7497
rect 23934 7460 23940 7472
rect 23895 7432 23940 7460
rect 23934 7420 23940 7432
rect 23992 7420 23998 7472
rect 24670 7460 24676 7472
rect 24631 7432 24676 7460
rect 24670 7420 24676 7432
rect 24728 7420 24734 7472
rect 19981 7395 20039 7401
rect 19981 7392 19993 7395
rect 18800 7364 19993 7392
rect 15105 7327 15163 7333
rect 15105 7293 15117 7327
rect 15151 7293 15163 7327
rect 15286 7324 15292 7336
rect 15247 7296 15292 7324
rect 15105 7287 15163 7293
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 18800 7268 18828 7364
rect 19981 7361 19993 7364
rect 20027 7361 20039 7395
rect 19981 7355 20039 7361
rect 21729 7395 21787 7401
rect 21729 7361 21741 7395
rect 21775 7361 21787 7395
rect 21729 7355 21787 7361
rect 24121 7395 24179 7401
rect 24121 7361 24133 7395
rect 24167 7392 24179 7395
rect 24210 7392 24216 7404
rect 24167 7364 24216 7392
rect 24167 7361 24179 7364
rect 24121 7355 24179 7361
rect 24210 7352 24216 7364
rect 24268 7392 24274 7404
rect 25409 7395 25467 7401
rect 25409 7392 25421 7395
rect 24268 7364 25421 7392
rect 24268 7352 24274 7364
rect 25409 7361 25421 7364
rect 25455 7361 25467 7395
rect 25409 7355 25467 7361
rect 25660 7327 25718 7333
rect 25660 7293 25672 7327
rect 25706 7324 25718 7327
rect 26160 7324 26188 7491
rect 27614 7488 27620 7500
rect 27672 7488 27678 7540
rect 25706 7296 26188 7324
rect 25706 7293 25718 7296
rect 25660 7287 25718 7293
rect 16577 7259 16635 7265
rect 16577 7225 16589 7259
rect 16623 7256 16635 7259
rect 16666 7256 16672 7268
rect 16623 7228 16672 7256
rect 16623 7225 16635 7228
rect 16577 7219 16635 7225
rect 16301 7191 16359 7197
rect 16301 7157 16313 7191
rect 16347 7188 16359 7191
rect 16592 7188 16620 7219
rect 16666 7216 16672 7228
rect 16724 7216 16730 7268
rect 18230 7216 18236 7268
rect 18288 7256 18294 7268
rect 18782 7256 18788 7268
rect 18288 7228 18333 7256
rect 18743 7228 18788 7256
rect 18288 7216 18294 7228
rect 18782 7216 18788 7228
rect 18840 7216 18846 7268
rect 19705 7259 19763 7265
rect 19705 7225 19717 7259
rect 19751 7225 19763 7259
rect 19705 7219 19763 7225
rect 16347 7160 16620 7188
rect 19720 7188 19748 7219
rect 19794 7216 19800 7268
rect 19852 7256 19858 7268
rect 19852 7228 19897 7256
rect 19852 7216 19858 7228
rect 21542 7216 21548 7268
rect 21600 7256 21606 7268
rect 22050 7259 22108 7265
rect 22050 7256 22062 7259
rect 21600 7228 22062 7256
rect 21600 7216 21606 7228
rect 22050 7225 22062 7228
rect 22096 7225 22108 7259
rect 22050 7219 22108 7225
rect 22738 7216 22744 7268
rect 22796 7256 22802 7268
rect 24213 7259 24271 7265
rect 22796 7228 24072 7256
rect 22796 7216 22802 7228
rect 20070 7188 20076 7200
rect 19720 7160 20076 7188
rect 16347 7157 16359 7160
rect 16301 7151 16359 7157
rect 20070 7148 20076 7160
rect 20128 7148 20134 7200
rect 23290 7148 23296 7200
rect 23348 7188 23354 7200
rect 23934 7188 23940 7200
rect 23348 7160 23940 7188
rect 23348 7148 23354 7160
rect 23934 7148 23940 7160
rect 23992 7148 23998 7200
rect 24044 7188 24072 7228
rect 24213 7225 24225 7259
rect 24259 7225 24271 7259
rect 24213 7219 24271 7225
rect 24228 7188 24256 7219
rect 25041 7191 25099 7197
rect 25041 7188 25053 7191
rect 24044 7160 25053 7188
rect 25041 7157 25053 7160
rect 25087 7157 25099 7191
rect 25041 7151 25099 7157
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 14921 6987 14979 6993
rect 14921 6953 14933 6987
rect 14967 6984 14979 6987
rect 15286 6984 15292 6996
rect 14967 6956 15292 6984
rect 14967 6953 14979 6956
rect 14921 6947 14979 6953
rect 15286 6944 15292 6956
rect 15344 6944 15350 6996
rect 15746 6984 15752 6996
rect 15707 6956 15752 6984
rect 15746 6944 15752 6956
rect 15804 6944 15810 6996
rect 17402 6984 17408 6996
rect 17363 6956 17408 6984
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 18230 6944 18236 6996
rect 18288 6984 18294 6996
rect 18601 6987 18659 6993
rect 18601 6984 18613 6987
rect 18288 6956 18613 6984
rect 18288 6944 18294 6956
rect 18601 6953 18613 6956
rect 18647 6953 18659 6987
rect 18601 6947 18659 6953
rect 19383 6987 19441 6993
rect 19383 6953 19395 6987
rect 19429 6984 19441 6987
rect 25038 6984 25044 6996
rect 19429 6956 25044 6984
rect 19429 6953 19441 6956
rect 19383 6947 19441 6953
rect 25038 6944 25044 6956
rect 25096 6944 25102 6996
rect 16761 6919 16819 6925
rect 16761 6885 16773 6919
rect 16807 6916 16819 6919
rect 17678 6916 17684 6928
rect 16807 6888 17684 6916
rect 16807 6885 16819 6888
rect 16761 6879 16819 6885
rect 17678 6876 17684 6888
rect 17736 6916 17742 6928
rect 17773 6919 17831 6925
rect 17773 6916 17785 6919
rect 17736 6888 17785 6916
rect 17736 6876 17742 6888
rect 17773 6885 17785 6888
rect 17819 6885 17831 6919
rect 18322 6916 18328 6928
rect 18283 6888 18328 6916
rect 17773 6879 17831 6885
rect 18322 6876 18328 6888
rect 18380 6876 18386 6928
rect 19518 6876 19524 6928
rect 19576 6916 19582 6928
rect 19705 6919 19763 6925
rect 19705 6916 19717 6919
rect 19576 6888 19717 6916
rect 19576 6876 19582 6888
rect 19705 6885 19717 6888
rect 19751 6885 19763 6919
rect 19705 6879 19763 6885
rect 21726 6876 21732 6928
rect 21784 6916 21790 6928
rect 22097 6919 22155 6925
rect 22097 6916 22109 6919
rect 21784 6888 22109 6916
rect 21784 6876 21790 6888
rect 22097 6885 22109 6888
rect 22143 6885 22155 6919
rect 23290 6916 23296 6928
rect 23251 6888 23296 6916
rect 22097 6879 22155 6885
rect 23290 6876 23296 6888
rect 23348 6876 23354 6928
rect 24305 6919 24363 6925
rect 24305 6885 24317 6919
rect 24351 6916 24363 6919
rect 24670 6916 24676 6928
rect 24351 6888 24676 6916
rect 24351 6885 24363 6888
rect 24305 6879 24363 6885
rect 24670 6876 24676 6888
rect 24728 6876 24734 6928
rect 16666 6848 16672 6860
rect 16627 6820 16672 6848
rect 16666 6808 16672 6820
rect 16724 6808 16730 6860
rect 18782 6808 18788 6860
rect 18840 6848 18846 6860
rect 19242 6848 19248 6860
rect 19300 6857 19306 6860
rect 19300 6851 19338 6857
rect 18840 6820 19248 6848
rect 18840 6808 18846 6820
rect 19242 6808 19248 6820
rect 19326 6817 19338 6851
rect 22646 6848 22652 6860
rect 22607 6820 22652 6848
rect 19300 6811 19338 6817
rect 19300 6808 19306 6811
rect 22646 6808 22652 6820
rect 22704 6808 22710 6860
rect 17310 6740 17316 6792
rect 17368 6780 17374 6792
rect 17681 6783 17739 6789
rect 17681 6780 17693 6783
rect 17368 6752 17693 6780
rect 17368 6740 17374 6752
rect 17681 6749 17693 6752
rect 17727 6749 17739 6783
rect 17681 6743 17739 6749
rect 21542 6740 21548 6792
rect 21600 6780 21606 6792
rect 21729 6783 21787 6789
rect 21729 6780 21741 6783
rect 21600 6752 21741 6780
rect 21600 6740 21606 6752
rect 21729 6749 21741 6752
rect 21775 6780 21787 6783
rect 24210 6780 24216 6792
rect 21775 6752 23474 6780
rect 24171 6752 24216 6780
rect 21775 6749 21787 6752
rect 21729 6743 21787 6749
rect 23446 6712 23474 6752
rect 24210 6740 24216 6752
rect 24268 6740 24274 6792
rect 24302 6740 24308 6792
rect 24360 6780 24366 6792
rect 24489 6783 24547 6789
rect 24489 6780 24501 6783
rect 24360 6752 24501 6780
rect 24360 6740 24366 6752
rect 24489 6749 24501 6752
rect 24535 6749 24547 6783
rect 24489 6743 24547 6749
rect 25958 6712 25964 6724
rect 23446 6684 25964 6712
rect 25958 6672 25964 6684
rect 26016 6672 26022 6724
rect 20070 6644 20076 6656
rect 20031 6616 20076 6644
rect 20070 6604 20076 6616
rect 20128 6604 20134 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 16117 6443 16175 6449
rect 16117 6409 16129 6443
rect 16163 6440 16175 6443
rect 16666 6440 16672 6452
rect 16163 6412 16672 6440
rect 16163 6409 16175 6412
rect 16117 6403 16175 6409
rect 16666 6400 16672 6412
rect 16724 6400 16730 6452
rect 17678 6440 17684 6452
rect 17639 6412 17684 6440
rect 17678 6400 17684 6412
rect 17736 6400 17742 6452
rect 19242 6440 19248 6452
rect 19203 6412 19248 6440
rect 19242 6400 19248 6412
rect 19300 6400 19306 6452
rect 22646 6440 22652 6452
rect 22607 6412 22652 6440
rect 22646 6400 22652 6412
rect 22704 6400 22710 6452
rect 23106 6400 23112 6452
rect 23164 6440 23170 6452
rect 23385 6443 23443 6449
rect 23385 6440 23397 6443
rect 23164 6412 23397 6440
rect 23164 6400 23170 6412
rect 23385 6409 23397 6412
rect 23431 6440 23443 6443
rect 23431 6412 23796 6440
rect 23431 6409 23443 6412
rect 23385 6403 23443 6409
rect 18141 6307 18199 6313
rect 18141 6273 18153 6307
rect 18187 6304 18199 6307
rect 20070 6304 20076 6316
rect 18187 6276 20076 6304
rect 18187 6273 18199 6276
rect 18141 6267 18199 6273
rect 20070 6264 20076 6276
rect 20128 6264 20134 6316
rect 23768 6245 23796 6412
rect 25222 6400 25228 6452
rect 25280 6440 25286 6452
rect 25363 6443 25421 6449
rect 25363 6440 25375 6443
rect 25280 6412 25375 6440
rect 25280 6400 25286 6412
rect 25363 6409 25375 6412
rect 25409 6409 25421 6443
rect 25363 6403 25421 6409
rect 25777 6443 25835 6449
rect 25777 6409 25789 6443
rect 25823 6440 25835 6443
rect 27614 6440 27620 6452
rect 25823 6412 27620 6440
rect 25823 6409 25835 6412
rect 25777 6403 25835 6409
rect 24397 6307 24455 6313
rect 24397 6273 24409 6307
rect 24443 6304 24455 6307
rect 24670 6304 24676 6316
rect 24443 6276 24676 6304
rect 24443 6273 24455 6276
rect 24397 6267 24455 6273
rect 24670 6264 24676 6276
rect 24728 6264 24734 6316
rect 23753 6239 23811 6245
rect 23753 6205 23765 6239
rect 23799 6205 23811 6239
rect 23753 6199 23811 6205
rect 25292 6239 25350 6245
rect 25292 6205 25304 6239
rect 25338 6236 25350 6239
rect 25792 6236 25820 6403
rect 27614 6400 27620 6412
rect 27672 6400 27678 6452
rect 25338 6208 25820 6236
rect 25338 6205 25350 6208
rect 25292 6199 25350 6205
rect 17310 6100 17316 6112
rect 17271 6072 17316 6100
rect 17310 6060 17316 6072
rect 17368 6060 17374 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 17310 5856 17316 5908
rect 17368 5896 17374 5908
rect 18187 5899 18245 5905
rect 18187 5896 18199 5899
rect 17368 5868 18199 5896
rect 17368 5856 17374 5868
rect 18187 5865 18199 5868
rect 18233 5865 18245 5899
rect 18187 5859 18245 5865
rect 23474 5856 23480 5908
rect 23532 5896 23538 5908
rect 23532 5868 23577 5896
rect 23532 5856 23538 5868
rect 18116 5763 18174 5769
rect 18116 5729 18128 5763
rect 18162 5760 18174 5763
rect 18322 5760 18328 5772
rect 18162 5732 18328 5760
rect 18162 5729 18174 5732
rect 18116 5723 18174 5729
rect 18322 5720 18328 5732
rect 18380 5720 18386 5772
rect 24670 5769 24676 5772
rect 24648 5763 24676 5769
rect 24648 5760 24660 5763
rect 24583 5732 24660 5760
rect 24648 5729 24660 5732
rect 24728 5760 24734 5772
rect 27614 5760 27620 5772
rect 24728 5732 27620 5760
rect 24648 5723 24676 5729
rect 24670 5720 24676 5723
rect 24728 5720 24734 5732
rect 27614 5720 27620 5732
rect 27672 5720 27678 5772
rect 24578 5584 24584 5636
rect 24636 5624 24642 5636
rect 24719 5627 24777 5633
rect 24719 5624 24731 5627
rect 24636 5596 24731 5624
rect 24636 5584 24642 5596
rect 24719 5593 24731 5596
rect 24765 5593 24777 5627
rect 24719 5587 24777 5593
rect 24210 5556 24216 5568
rect 24171 5528 24216 5556
rect 24210 5516 24216 5528
rect 24268 5516 24274 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 24670 5352 24676 5364
rect 24631 5324 24676 5352
rect 24670 5312 24676 5324
rect 24728 5312 24734 5364
rect 18322 5012 18328 5024
rect 18283 4984 18328 5012
rect 18322 4972 18328 4984
rect 18380 4972 18386 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 24394 4700 24400 4752
rect 24452 4740 24458 4752
rect 24719 4743 24777 4749
rect 24719 4740 24731 4743
rect 24452 4712 24731 4740
rect 24452 4700 24458 4712
rect 24719 4709 24731 4712
rect 24765 4709 24777 4743
rect 24719 4703 24777 4709
rect 24578 4672 24584 4684
rect 24539 4644 24584 4672
rect 24578 4632 24584 4644
rect 24636 4632 24642 4684
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 24670 4264 24676 4276
rect 24583 4236 24676 4264
rect 24670 4224 24676 4236
rect 24728 4264 24734 4276
rect 27614 4264 27620 4276
rect 24728 4236 27620 4264
rect 24728 4224 24734 4236
rect 27614 4224 27620 4236
rect 27672 4224 27678 4276
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 24486 3612 24492 3664
rect 24544 3652 24550 3664
rect 24719 3655 24777 3661
rect 24719 3652 24731 3655
rect 24544 3624 24731 3652
rect 24544 3612 24550 3624
rect 24719 3621 24731 3624
rect 24765 3621 24777 3655
rect 24719 3615 24777 3621
rect 24578 3584 24584 3596
rect 24539 3556 24584 3584
rect 24578 3544 24584 3556
rect 24636 3544 24642 3596
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 24670 3176 24676 3188
rect 24583 3148 24676 3176
rect 24670 3136 24676 3148
rect 24728 3176 24734 3188
rect 27614 3176 27620 3188
rect 24728 3148 27620 3176
rect 24728 3136 24734 3148
rect 27614 3136 27620 3148
rect 27672 3136 27678 3188
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 11514 2592 11520 2644
rect 11572 2632 11578 2644
rect 11609 2635 11667 2641
rect 11609 2632 11621 2635
rect 11572 2604 11621 2632
rect 11572 2592 11578 2604
rect 11609 2601 11621 2604
rect 11655 2601 11667 2635
rect 11609 2595 11667 2601
rect 24210 2592 24216 2644
rect 24268 2632 24274 2644
rect 24719 2635 24777 2641
rect 24719 2632 24731 2635
rect 24268 2604 24731 2632
rect 24268 2592 24274 2604
rect 24719 2601 24731 2604
rect 24765 2601 24777 2635
rect 24719 2595 24777 2601
rect 11400 2499 11458 2505
rect 11400 2465 11412 2499
rect 11446 2465 11458 2499
rect 11400 2459 11458 2465
rect 24648 2499 24706 2505
rect 24648 2465 24660 2499
rect 24694 2496 24706 2499
rect 25130 2496 25136 2508
rect 24694 2468 25136 2496
rect 24694 2465 24706 2468
rect 24648 2459 24706 2465
rect 11415 2428 11443 2459
rect 25130 2456 25136 2468
rect 25188 2456 25194 2508
rect 11882 2428 11888 2440
rect 11415 2400 11888 2428
rect 11882 2388 11888 2400
rect 11940 2388 11946 2440
rect 25130 2292 25136 2304
rect 25091 2264 25136 2292
rect 25130 2252 25136 2264
rect 25188 2252 25194 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 1762 76 1768 128
rect 1820 116 1826 128
rect 9582 116 9588 128
rect 1820 88 9588 116
rect 1820 76 1826 88
rect 9582 76 9588 88
rect 9640 76 9646 128
rect 15746 76 15752 128
rect 15804 116 15810 128
rect 16390 116 16396 128
rect 15804 88 16396 116
rect 15804 76 15810 88
rect 16390 76 16396 88
rect 16448 76 16454 128
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 13912 25440 13964 25492
rect 20076 25440 20128 25492
rect 25504 25304 25556 25356
rect 23848 25100 23900 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 9956 24939 10008 24948
rect 9956 24905 9965 24939
rect 9965 24905 9999 24939
rect 9999 24905 10008 24939
rect 9956 24896 10008 24905
rect 12900 24939 12952 24948
rect 12900 24905 12909 24939
rect 12909 24905 12943 24939
rect 12943 24905 12952 24939
rect 12900 24896 12952 24905
rect 14832 24896 14884 24948
rect 17316 24939 17368 24948
rect 17316 24905 17325 24939
rect 17325 24905 17359 24939
rect 17359 24905 17368 24939
rect 17316 24896 17368 24905
rect 25136 24939 25188 24948
rect 25136 24905 25145 24939
rect 25145 24905 25179 24939
rect 25179 24905 25188 24939
rect 25136 24896 25188 24905
rect 16212 24828 16264 24880
rect 9956 24692 10008 24744
rect 12900 24692 12952 24744
rect 14832 24692 14884 24744
rect 15568 24692 15620 24744
rect 17316 24692 17368 24744
rect 25136 24692 25188 24744
rect 17960 24624 18012 24676
rect 18144 24667 18196 24676
rect 18144 24633 18153 24667
rect 18153 24633 18187 24667
rect 18187 24633 18196 24667
rect 18144 24624 18196 24633
rect 11704 24556 11756 24608
rect 13636 24556 13688 24608
rect 14740 24556 14792 24608
rect 15752 24556 15804 24608
rect 17868 24599 17920 24608
rect 17868 24565 17877 24599
rect 17877 24565 17911 24599
rect 17911 24565 17920 24599
rect 20352 24624 20404 24676
rect 25504 24667 25556 24676
rect 25504 24633 25513 24667
rect 25513 24633 25547 24667
rect 25547 24633 25556 24667
rect 25504 24624 25556 24633
rect 17868 24556 17920 24565
rect 22008 24556 22060 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 6644 24216 6696 24268
rect 10416 24216 10468 24268
rect 11796 24284 11848 24336
rect 18144 24395 18196 24404
rect 18144 24361 18153 24395
rect 18153 24361 18187 24395
rect 18187 24361 18196 24395
rect 18144 24352 18196 24361
rect 19064 24352 19116 24404
rect 22192 24352 22244 24404
rect 25320 24352 25372 24404
rect 18880 24327 18932 24336
rect 18880 24293 18889 24327
rect 18889 24293 18923 24327
rect 18923 24293 18932 24327
rect 18880 24284 18932 24293
rect 11336 24216 11388 24268
rect 12808 24259 12860 24268
rect 12808 24225 12817 24259
rect 12817 24225 12851 24259
rect 12851 24225 12860 24259
rect 12808 24216 12860 24225
rect 13544 24216 13596 24268
rect 14188 24216 14240 24268
rect 15844 24259 15896 24268
rect 15844 24225 15853 24259
rect 15853 24225 15887 24259
rect 15887 24225 15896 24259
rect 15844 24216 15896 24225
rect 15936 24216 15988 24268
rect 17408 24216 17460 24268
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 23664 24259 23716 24268
rect 23664 24225 23673 24259
rect 23673 24225 23707 24259
rect 23707 24225 23716 24259
rect 23664 24216 23716 24225
rect 24860 24259 24912 24268
rect 24860 24225 24878 24259
rect 24878 24225 24912 24259
rect 24860 24216 24912 24225
rect 27344 24216 27396 24268
rect 11704 24148 11756 24200
rect 15292 24191 15344 24200
rect 13452 24080 13504 24132
rect 15292 24157 15301 24191
rect 15301 24157 15335 24191
rect 15335 24157 15344 24191
rect 15292 24148 15344 24157
rect 18788 24191 18840 24200
rect 18788 24157 18797 24191
rect 18797 24157 18831 24191
rect 18831 24157 18840 24191
rect 18788 24148 18840 24157
rect 18972 24148 19024 24200
rect 18328 24080 18380 24132
rect 6828 24012 6880 24064
rect 13728 24055 13780 24064
rect 13728 24021 13737 24055
rect 13737 24021 13771 24055
rect 13771 24021 13780 24055
rect 13728 24012 13780 24021
rect 18512 24012 18564 24064
rect 19800 24055 19852 24064
rect 19800 24021 19809 24055
rect 19809 24021 19843 24055
rect 19843 24021 19852 24055
rect 19800 24012 19852 24021
rect 24124 24012 24176 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 3700 23851 3752 23860
rect 3700 23817 3709 23851
rect 3709 23817 3743 23851
rect 3743 23817 3752 23851
rect 3700 23808 3752 23817
rect 5540 23808 5592 23860
rect 6644 23808 6696 23860
rect 7840 23851 7892 23860
rect 7840 23817 7849 23851
rect 7849 23817 7883 23851
rect 7883 23817 7892 23851
rect 7840 23808 7892 23817
rect 8944 23851 8996 23860
rect 8944 23817 8953 23851
rect 8953 23817 8987 23851
rect 8987 23817 8996 23851
rect 8944 23808 8996 23817
rect 10416 23851 10468 23860
rect 10416 23817 10425 23851
rect 10425 23817 10459 23851
rect 10459 23817 10468 23851
rect 10416 23808 10468 23817
rect 13544 23851 13596 23860
rect 13544 23817 13553 23851
rect 13553 23817 13587 23851
rect 13587 23817 13596 23851
rect 13544 23808 13596 23817
rect 13912 23851 13964 23860
rect 13912 23817 13921 23851
rect 13921 23817 13955 23851
rect 13955 23817 13964 23851
rect 13912 23808 13964 23817
rect 14188 23808 14240 23860
rect 15476 23808 15528 23860
rect 15844 23851 15896 23860
rect 15844 23817 15853 23851
rect 15853 23817 15887 23851
rect 15887 23817 15896 23851
rect 15844 23808 15896 23817
rect 17408 23851 17460 23860
rect 17408 23817 17417 23851
rect 17417 23817 17451 23851
rect 17451 23817 17460 23851
rect 17408 23808 17460 23817
rect 17868 23851 17920 23860
rect 17868 23817 17877 23851
rect 17877 23817 17911 23851
rect 17911 23817 17920 23851
rect 17868 23808 17920 23817
rect 18880 23808 18932 23860
rect 19156 23851 19208 23860
rect 19156 23817 19165 23851
rect 19165 23817 19199 23851
rect 19199 23817 19208 23851
rect 19156 23808 19208 23817
rect 20904 23851 20956 23860
rect 20904 23817 20913 23851
rect 20913 23817 20947 23851
rect 20947 23817 20956 23851
rect 20904 23808 20956 23817
rect 23204 23808 23256 23860
rect 24860 23851 24912 23860
rect 24860 23817 24869 23851
rect 24869 23817 24903 23851
rect 24903 23817 24912 23851
rect 24860 23808 24912 23817
rect 26332 23808 26384 23860
rect 480 23604 532 23656
rect 3700 23604 3752 23656
rect 5540 23604 5592 23656
rect 7840 23604 7892 23656
rect 8944 23604 8996 23656
rect 10784 23740 10836 23792
rect 17040 23783 17092 23792
rect 14740 23672 14792 23724
rect 15568 23715 15620 23724
rect 15568 23681 15577 23715
rect 15577 23681 15611 23715
rect 15611 23681 15620 23715
rect 15568 23672 15620 23681
rect 17040 23749 17049 23783
rect 17049 23749 17083 23783
rect 17083 23749 17092 23783
rect 17040 23740 17092 23749
rect 20352 23783 20404 23792
rect 20352 23749 20361 23783
rect 20361 23749 20395 23783
rect 20395 23749 20404 23783
rect 20352 23740 20404 23749
rect 18052 23672 18104 23724
rect 19800 23715 19852 23724
rect 19800 23681 19809 23715
rect 19809 23681 19843 23715
rect 19843 23681 19852 23715
rect 19800 23672 19852 23681
rect 21364 23672 21416 23724
rect 11060 23647 11112 23656
rect 11060 23613 11069 23647
rect 11069 23613 11103 23647
rect 11103 23613 11112 23647
rect 11060 23604 11112 23613
rect 12624 23647 12676 23656
rect 12624 23613 12633 23647
rect 12633 23613 12667 23647
rect 12667 23613 12676 23647
rect 12624 23604 12676 23613
rect 13728 23647 13780 23656
rect 13728 23613 13737 23647
rect 13737 23613 13771 23647
rect 13771 23613 13780 23647
rect 13728 23604 13780 23613
rect 17040 23604 17092 23656
rect 17868 23604 17920 23656
rect 18144 23604 18196 23656
rect 21272 23647 21324 23656
rect 21272 23613 21281 23647
rect 21281 23613 21315 23647
rect 21315 23613 21324 23647
rect 21272 23604 21324 23613
rect 22192 23604 22244 23656
rect 25228 23647 25280 23656
rect 25228 23613 25237 23647
rect 25237 23613 25271 23647
rect 25271 23613 25280 23647
rect 25228 23604 25280 23613
rect 1676 23468 1728 23520
rect 5356 23468 5408 23520
rect 7380 23468 7432 23520
rect 7656 23468 7708 23520
rect 8760 23468 8812 23520
rect 9496 23468 9548 23520
rect 10784 23511 10836 23520
rect 10784 23477 10793 23511
rect 10793 23477 10827 23511
rect 10827 23477 10836 23511
rect 10784 23468 10836 23477
rect 11336 23468 11388 23520
rect 15292 23536 15344 23588
rect 23664 23536 23716 23588
rect 23940 23511 23992 23520
rect 23940 23477 23949 23511
rect 23949 23477 23983 23511
rect 23983 23477 23992 23511
rect 23940 23468 23992 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 12624 23264 12676 23316
rect 14740 23264 14792 23316
rect 18788 23264 18840 23316
rect 10600 23196 10652 23248
rect 10784 23196 10836 23248
rect 13176 23196 13228 23248
rect 15476 23239 15528 23248
rect 15476 23205 15485 23239
rect 15485 23205 15519 23239
rect 15519 23205 15528 23239
rect 15476 23196 15528 23205
rect 19156 23196 19208 23248
rect 20812 23264 20864 23316
rect 21272 23264 21324 23316
rect 21364 23264 21416 23316
rect 22008 23196 22060 23248
rect 22192 23196 22244 23248
rect 23756 23196 23808 23248
rect 23940 23196 23992 23248
rect 2504 23128 2556 23180
rect 8300 23171 8352 23180
rect 8300 23137 8344 23171
rect 8344 23137 8352 23171
rect 12256 23171 12308 23180
rect 8300 23128 8352 23137
rect 12256 23137 12265 23171
rect 12265 23137 12299 23171
rect 12299 23137 12308 23171
rect 12256 23128 12308 23137
rect 18236 23171 18288 23180
rect 10140 23060 10192 23112
rect 13360 23103 13412 23112
rect 5356 22992 5408 23044
rect 13360 23069 13369 23103
rect 13369 23069 13403 23103
rect 13403 23069 13412 23103
rect 13360 23060 13412 23069
rect 14280 23060 14332 23112
rect 15384 23103 15436 23112
rect 15384 23069 15393 23103
rect 15393 23069 15427 23103
rect 15427 23069 15436 23103
rect 15384 23060 15436 23069
rect 15568 23060 15620 23112
rect 11336 23035 11388 23044
rect 11336 23001 11345 23035
rect 11345 23001 11379 23035
rect 11379 23001 11388 23035
rect 11336 22992 11388 23001
rect 18236 23137 18245 23171
rect 18245 23137 18279 23171
rect 18279 23137 18288 23171
rect 18236 23128 18288 23137
rect 19708 23171 19760 23180
rect 19708 23137 19717 23171
rect 19717 23137 19751 23171
rect 19751 23137 19760 23171
rect 19708 23128 19760 23137
rect 20812 23128 20864 23180
rect 26148 23128 26200 23180
rect 18512 23060 18564 23112
rect 22468 23060 22520 23112
rect 24032 23060 24084 23112
rect 20904 22992 20956 23044
rect 23940 22992 23992 23044
rect 9220 22924 9272 22976
rect 11060 22924 11112 22976
rect 14372 22967 14424 22976
rect 14372 22933 14381 22967
rect 14381 22933 14415 22967
rect 14415 22933 14424 22967
rect 14372 22924 14424 22933
rect 16488 22967 16540 22976
rect 16488 22933 16497 22967
rect 16497 22933 16531 22967
rect 16531 22933 16540 22967
rect 16488 22924 16540 22933
rect 17132 22924 17184 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 8300 22763 8352 22772
rect 8300 22729 8309 22763
rect 8309 22729 8343 22763
rect 8343 22729 8352 22763
rect 8300 22720 8352 22729
rect 10140 22763 10192 22772
rect 10140 22729 10149 22763
rect 10149 22729 10183 22763
rect 10183 22729 10192 22763
rect 10140 22720 10192 22729
rect 10600 22763 10652 22772
rect 10600 22729 10609 22763
rect 10609 22729 10643 22763
rect 10643 22729 10652 22763
rect 10600 22720 10652 22729
rect 12808 22720 12860 22772
rect 13360 22720 13412 22772
rect 15384 22720 15436 22772
rect 15844 22720 15896 22772
rect 11336 22695 11388 22704
rect 11336 22661 11345 22695
rect 11345 22661 11379 22695
rect 11379 22661 11388 22695
rect 11336 22652 11388 22661
rect 9220 22627 9272 22636
rect 9220 22593 9229 22627
rect 9229 22593 9263 22627
rect 9263 22593 9272 22627
rect 9220 22584 9272 22593
rect 11704 22584 11756 22636
rect 12256 22584 12308 22636
rect 14372 22652 14424 22704
rect 14740 22652 14792 22704
rect 14280 22627 14332 22636
rect 14280 22593 14289 22627
rect 14289 22593 14323 22627
rect 14323 22593 14332 22627
rect 14280 22584 14332 22593
rect 17960 22720 18012 22772
rect 19708 22720 19760 22772
rect 25780 22763 25832 22772
rect 25780 22729 25789 22763
rect 25789 22729 25823 22763
rect 25823 22729 25832 22763
rect 25780 22720 25832 22729
rect 26148 22763 26200 22772
rect 26148 22729 26157 22763
rect 26157 22729 26191 22763
rect 26191 22729 26200 22763
rect 26148 22720 26200 22729
rect 23572 22652 23624 22704
rect 23848 22584 23900 22636
rect 10784 22491 10836 22500
rect 9036 22423 9088 22432
rect 9036 22389 9045 22423
rect 9045 22389 9079 22423
rect 9079 22389 9088 22423
rect 10784 22457 10793 22491
rect 10793 22457 10827 22491
rect 10827 22457 10836 22491
rect 10784 22448 10836 22457
rect 11060 22448 11112 22500
rect 19432 22516 19484 22568
rect 25780 22516 25832 22568
rect 9036 22380 9088 22389
rect 12256 22423 12308 22432
rect 12256 22389 12265 22423
rect 12265 22389 12299 22423
rect 12299 22389 12308 22423
rect 12256 22380 12308 22389
rect 13176 22380 13228 22432
rect 13820 22423 13872 22432
rect 13820 22389 13829 22423
rect 13829 22389 13863 22423
rect 13863 22389 13872 22423
rect 15384 22448 15436 22500
rect 16488 22491 16540 22500
rect 16488 22457 16497 22491
rect 16497 22457 16531 22491
rect 16531 22457 16540 22491
rect 16488 22448 16540 22457
rect 17132 22491 17184 22500
rect 13820 22380 13872 22389
rect 14372 22380 14424 22432
rect 15476 22380 15528 22432
rect 16304 22423 16356 22432
rect 16304 22389 16313 22423
rect 16313 22389 16347 22423
rect 16347 22389 16356 22423
rect 17132 22457 17141 22491
rect 17141 22457 17175 22491
rect 17175 22457 17184 22491
rect 17132 22448 17184 22457
rect 18236 22491 18288 22500
rect 18236 22457 18245 22491
rect 18245 22457 18279 22491
rect 18279 22457 18288 22491
rect 18788 22491 18840 22500
rect 18236 22448 18288 22457
rect 18788 22457 18797 22491
rect 18797 22457 18831 22491
rect 18831 22457 18840 22491
rect 18788 22448 18840 22457
rect 19248 22448 19300 22500
rect 20812 22448 20864 22500
rect 16304 22380 16356 22389
rect 20076 22423 20128 22432
rect 20076 22389 20085 22423
rect 20085 22389 20119 22423
rect 20119 22389 20128 22423
rect 20076 22380 20128 22389
rect 21456 22423 21508 22432
rect 21456 22389 21465 22423
rect 21465 22389 21499 22423
rect 21499 22389 21508 22423
rect 21456 22380 21508 22389
rect 22744 22380 22796 22432
rect 23388 22423 23440 22432
rect 23388 22389 23397 22423
rect 23397 22389 23431 22423
rect 23431 22389 23440 22423
rect 23388 22380 23440 22389
rect 24032 22380 24084 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 9220 22219 9272 22228
rect 9220 22185 9229 22219
rect 9229 22185 9263 22219
rect 9263 22185 9272 22219
rect 9220 22176 9272 22185
rect 13820 22219 13872 22228
rect 13820 22185 13829 22219
rect 13829 22185 13863 22219
rect 13863 22185 13872 22219
rect 17500 22219 17552 22228
rect 13820 22176 13872 22185
rect 17500 22185 17509 22219
rect 17509 22185 17543 22219
rect 17543 22185 17552 22219
rect 17500 22176 17552 22185
rect 18236 22176 18288 22228
rect 22468 22219 22520 22228
rect 22468 22185 22477 22219
rect 22477 22185 22511 22219
rect 22511 22185 22520 22219
rect 22468 22176 22520 22185
rect 23756 22219 23808 22228
rect 23756 22185 23765 22219
rect 23765 22185 23799 22219
rect 23799 22185 23808 22219
rect 23756 22176 23808 22185
rect 24032 22219 24084 22228
rect 24032 22185 24041 22219
rect 24041 22185 24075 22219
rect 24075 22185 24084 22219
rect 24032 22176 24084 22185
rect 9680 22108 9732 22160
rect 16304 22151 16356 22160
rect 16304 22117 16313 22151
rect 16313 22117 16347 22151
rect 16347 22117 16356 22151
rect 16304 22108 16356 22117
rect 19432 22151 19484 22160
rect 19432 22117 19441 22151
rect 19441 22117 19475 22151
rect 19475 22117 19484 22151
rect 19432 22108 19484 22117
rect 23388 22151 23440 22160
rect 23388 22117 23397 22151
rect 23397 22117 23431 22151
rect 23431 22117 23440 22151
rect 23388 22108 23440 22117
rect 13176 22040 13228 22092
rect 15936 22083 15988 22092
rect 15936 22049 15945 22083
rect 15945 22049 15979 22083
rect 15979 22049 15988 22083
rect 15936 22040 15988 22049
rect 22744 22083 22796 22092
rect 22744 22049 22753 22083
rect 22753 22049 22787 22083
rect 22787 22049 22796 22083
rect 22744 22040 22796 22049
rect 24768 22040 24820 22092
rect 9956 21972 10008 22024
rect 17684 21972 17736 22024
rect 18880 21972 18932 22024
rect 20536 21972 20588 22024
rect 10784 21947 10836 21956
rect 10784 21913 10793 21947
rect 10793 21913 10827 21947
rect 10827 21913 10836 21947
rect 10784 21904 10836 21913
rect 20352 21947 20404 21956
rect 20352 21913 20361 21947
rect 20361 21913 20395 21947
rect 20395 21913 20404 21947
rect 20352 21904 20404 21913
rect 11060 21836 11112 21888
rect 21824 21879 21876 21888
rect 21824 21845 21833 21879
rect 21833 21845 21867 21879
rect 21867 21845 21876 21879
rect 21824 21836 21876 21845
rect 22192 21879 22244 21888
rect 22192 21845 22201 21879
rect 22201 21845 22235 21879
rect 22235 21845 22244 21879
rect 22192 21836 22244 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 4804 21675 4856 21684
rect 4804 21641 4813 21675
rect 4813 21641 4847 21675
rect 4847 21641 4856 21675
rect 4804 21632 4856 21641
rect 9680 21675 9732 21684
rect 9680 21641 9689 21675
rect 9689 21641 9723 21675
rect 9723 21641 9732 21675
rect 9680 21632 9732 21641
rect 11060 21675 11112 21684
rect 11060 21641 11069 21675
rect 11069 21641 11103 21675
rect 11103 21641 11112 21675
rect 11060 21632 11112 21641
rect 14372 21675 14424 21684
rect 14372 21641 14381 21675
rect 14381 21641 14415 21675
rect 14415 21641 14424 21675
rect 14372 21632 14424 21641
rect 15936 21675 15988 21684
rect 15936 21641 15945 21675
rect 15945 21641 15979 21675
rect 15979 21641 15988 21675
rect 15936 21632 15988 21641
rect 19432 21632 19484 21684
rect 20076 21632 20128 21684
rect 22192 21632 22244 21684
rect 22744 21632 22796 21684
rect 24768 21675 24820 21684
rect 24768 21641 24777 21675
rect 24777 21641 24811 21675
rect 24811 21641 24820 21675
rect 24768 21632 24820 21641
rect 13544 21564 13596 21616
rect 18880 21607 18932 21616
rect 18880 21573 18889 21607
rect 18889 21573 18923 21607
rect 18923 21573 18932 21607
rect 18880 21564 18932 21573
rect 25780 21607 25832 21616
rect 25780 21573 25789 21607
rect 25789 21573 25823 21607
rect 25823 21573 25832 21607
rect 25780 21564 25832 21573
rect 10232 21496 10284 21548
rect 15384 21539 15436 21548
rect 15384 21505 15393 21539
rect 15393 21505 15427 21539
rect 15427 21505 15436 21539
rect 15384 21496 15436 21505
rect 17132 21539 17184 21548
rect 17132 21505 17141 21539
rect 17141 21505 17175 21539
rect 17175 21505 17184 21539
rect 17132 21496 17184 21505
rect 20352 21496 20404 21548
rect 20536 21539 20588 21548
rect 20536 21505 20545 21539
rect 20545 21505 20579 21539
rect 20579 21505 20588 21539
rect 20536 21496 20588 21505
rect 4804 21428 4856 21480
rect 9036 21428 9088 21480
rect 9220 21471 9272 21480
rect 9220 21437 9229 21471
rect 9229 21437 9263 21471
rect 9263 21437 9272 21471
rect 9220 21428 9272 21437
rect 10692 21428 10744 21480
rect 13912 21428 13964 21480
rect 21824 21428 21876 21480
rect 22284 21428 22336 21480
rect 23480 21471 23532 21480
rect 23480 21437 23489 21471
rect 23489 21437 23523 21471
rect 23523 21437 23532 21471
rect 23480 21428 23532 21437
rect 10232 21360 10284 21412
rect 13360 21403 13412 21412
rect 13360 21369 13369 21403
rect 13369 21369 13403 21403
rect 13403 21369 13412 21403
rect 13360 21360 13412 21369
rect 14004 21360 14056 21412
rect 16488 21403 16540 21412
rect 16488 21369 16497 21403
rect 16497 21369 16531 21403
rect 16531 21369 16540 21403
rect 16488 21360 16540 21369
rect 17500 21403 17552 21412
rect 9128 21292 9180 21344
rect 13176 21292 13228 21344
rect 15936 21292 15988 21344
rect 17500 21369 17509 21403
rect 17509 21369 17543 21403
rect 17543 21369 17552 21403
rect 17500 21360 17552 21369
rect 19340 21360 19392 21412
rect 20168 21403 20220 21412
rect 20168 21369 20177 21403
rect 20177 21369 20211 21403
rect 20211 21369 20220 21403
rect 20168 21360 20220 21369
rect 24400 21403 24452 21412
rect 17684 21292 17736 21344
rect 21640 21335 21692 21344
rect 21640 21301 21649 21335
rect 21649 21301 21683 21335
rect 21683 21301 21692 21335
rect 24400 21369 24409 21403
rect 24409 21369 24443 21403
rect 24443 21369 24452 21403
rect 24400 21360 24452 21369
rect 21640 21292 21692 21301
rect 25044 21292 25096 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 9220 21088 9272 21140
rect 13176 21088 13228 21140
rect 13912 21131 13964 21140
rect 13912 21097 13921 21131
rect 13921 21097 13955 21131
rect 13955 21097 13964 21131
rect 13912 21088 13964 21097
rect 15660 21131 15712 21140
rect 15660 21097 15669 21131
rect 15669 21097 15703 21131
rect 15703 21097 15712 21131
rect 15660 21088 15712 21097
rect 15936 21088 15988 21140
rect 16488 21131 16540 21140
rect 16488 21097 16497 21131
rect 16497 21097 16531 21131
rect 16531 21097 16540 21131
rect 16488 21088 16540 21097
rect 10140 21020 10192 21072
rect 13360 21020 13412 21072
rect 17224 21063 17276 21072
rect 17224 21029 17233 21063
rect 17233 21029 17267 21063
rect 17267 21029 17276 21063
rect 17224 21020 17276 21029
rect 19432 21088 19484 21140
rect 22744 21088 22796 21140
rect 19340 21020 19392 21072
rect 21640 21020 21692 21072
rect 23480 21063 23532 21072
rect 23480 21029 23489 21063
rect 23489 21029 23523 21063
rect 23523 21029 23532 21063
rect 23480 21020 23532 21029
rect 24400 21020 24452 21072
rect 24952 21020 25004 21072
rect 9680 20927 9732 20936
rect 9680 20893 9689 20927
rect 9689 20893 9723 20927
rect 9723 20893 9732 20927
rect 9680 20884 9732 20893
rect 12716 20927 12768 20936
rect 12716 20893 12725 20927
rect 12725 20893 12759 20927
rect 12759 20893 12768 20927
rect 12716 20884 12768 20893
rect 15384 20884 15436 20936
rect 17132 20927 17184 20936
rect 17132 20893 17141 20927
rect 17141 20893 17175 20927
rect 17175 20893 17184 20927
rect 17132 20884 17184 20893
rect 18696 20884 18748 20936
rect 21916 20884 21968 20936
rect 23388 20927 23440 20936
rect 23388 20893 23397 20927
rect 23397 20893 23431 20927
rect 23431 20893 23440 20927
rect 23388 20884 23440 20893
rect 25044 20884 25096 20936
rect 24860 20816 24912 20868
rect 9956 20748 10008 20800
rect 19984 20791 20036 20800
rect 19984 20757 19993 20791
rect 19993 20757 20027 20791
rect 20027 20757 20036 20791
rect 19984 20748 20036 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 10140 20544 10192 20596
rect 16304 20544 16356 20596
rect 17224 20587 17276 20596
rect 17224 20553 17233 20587
rect 17233 20553 17267 20587
rect 17267 20553 17276 20587
rect 17224 20544 17276 20553
rect 22744 20544 22796 20596
rect 23480 20544 23532 20596
rect 24952 20587 25004 20596
rect 24952 20553 24961 20587
rect 24961 20553 24995 20587
rect 24995 20553 25004 20587
rect 24952 20544 25004 20553
rect 1492 20340 1544 20392
rect 7380 20340 7432 20392
rect 9680 20408 9732 20460
rect 9864 20383 9916 20392
rect 9864 20349 9873 20383
rect 9873 20349 9907 20383
rect 9907 20349 9916 20383
rect 9864 20340 9916 20349
rect 10140 20340 10192 20392
rect 10692 20340 10744 20392
rect 14004 20476 14056 20528
rect 13912 20408 13964 20460
rect 13084 20340 13136 20392
rect 13820 20383 13872 20392
rect 13820 20349 13829 20383
rect 13829 20349 13863 20383
rect 13863 20349 13872 20383
rect 14280 20383 14332 20392
rect 13820 20340 13872 20349
rect 14280 20349 14289 20383
rect 14289 20349 14323 20383
rect 14323 20349 14332 20383
rect 14280 20340 14332 20349
rect 15660 20476 15712 20528
rect 16488 20408 16540 20460
rect 17132 20476 17184 20528
rect 19340 20519 19392 20528
rect 19340 20485 19349 20519
rect 19349 20485 19383 20519
rect 19383 20485 19392 20519
rect 19340 20476 19392 20485
rect 21640 20476 21692 20528
rect 25780 20519 25832 20528
rect 25780 20485 25789 20519
rect 25789 20485 25823 20519
rect 25823 20485 25832 20519
rect 25780 20476 25832 20485
rect 19984 20408 20036 20460
rect 17592 20340 17644 20392
rect 16028 20272 16080 20324
rect 20536 20315 20588 20324
rect 16120 20247 16172 20256
rect 16120 20213 16129 20247
rect 16129 20213 16163 20247
rect 16163 20213 16172 20247
rect 18696 20247 18748 20256
rect 16120 20204 16172 20213
rect 18696 20213 18705 20247
rect 18705 20213 18739 20247
rect 18739 20213 18748 20247
rect 18696 20204 18748 20213
rect 19524 20204 19576 20256
rect 20536 20281 20545 20315
rect 20545 20281 20579 20315
rect 20579 20281 20588 20315
rect 23388 20340 23440 20392
rect 20536 20272 20588 20281
rect 23940 20272 23992 20324
rect 21640 20247 21692 20256
rect 21640 20213 21649 20247
rect 21649 20213 21683 20247
rect 21683 20213 21692 20247
rect 21640 20204 21692 20213
rect 21916 20247 21968 20256
rect 21916 20213 21925 20247
rect 21925 20213 21959 20247
rect 21959 20213 21968 20247
rect 21916 20204 21968 20213
rect 23112 20204 23164 20256
rect 23756 20204 23808 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 9680 20000 9732 20052
rect 12716 20000 12768 20052
rect 14280 20000 14332 20052
rect 17592 20043 17644 20052
rect 17592 20009 17601 20043
rect 17601 20009 17635 20043
rect 17635 20009 17644 20043
rect 17592 20000 17644 20009
rect 18144 20043 18196 20052
rect 18144 20009 18153 20043
rect 18153 20009 18187 20043
rect 18187 20009 18196 20043
rect 18144 20000 18196 20009
rect 19524 20043 19576 20052
rect 19524 20009 19533 20043
rect 19533 20009 19567 20043
rect 19567 20009 19576 20043
rect 19524 20000 19576 20009
rect 22744 20043 22796 20052
rect 22744 20009 22753 20043
rect 22753 20009 22787 20043
rect 22787 20009 22796 20043
rect 22744 20000 22796 20009
rect 23296 20043 23348 20052
rect 23296 20009 23305 20043
rect 23305 20009 23339 20043
rect 23339 20009 23348 20043
rect 23296 20000 23348 20009
rect 25044 20000 25096 20052
rect 9772 19907 9824 19916
rect 9772 19873 9781 19907
rect 9781 19873 9815 19907
rect 9815 19873 9824 19907
rect 9772 19864 9824 19873
rect 10140 19907 10192 19916
rect 10140 19873 10149 19907
rect 10149 19873 10183 19907
rect 10183 19873 10192 19907
rect 10140 19864 10192 19873
rect 12716 19864 12768 19916
rect 21640 19932 21692 19984
rect 22376 19932 22428 19984
rect 23940 19975 23992 19984
rect 23940 19941 23949 19975
rect 23949 19941 23983 19975
rect 23983 19941 23992 19975
rect 23940 19932 23992 19941
rect 24032 19932 24084 19984
rect 13820 19864 13872 19916
rect 15292 19907 15344 19916
rect 15292 19873 15301 19907
rect 15301 19873 15335 19907
rect 15335 19873 15344 19907
rect 15292 19864 15344 19873
rect 15476 19864 15528 19916
rect 19340 19907 19392 19916
rect 19340 19873 19349 19907
rect 19349 19873 19383 19907
rect 19383 19873 19392 19907
rect 19340 19864 19392 19873
rect 11336 19796 11388 19848
rect 14556 19796 14608 19848
rect 15384 19796 15436 19848
rect 16764 19796 16816 19848
rect 21548 19796 21600 19848
rect 23848 19839 23900 19848
rect 23848 19805 23857 19839
rect 23857 19805 23891 19839
rect 23891 19805 23900 19839
rect 23848 19796 23900 19805
rect 24216 19839 24268 19848
rect 24216 19805 24225 19839
rect 24225 19805 24259 19839
rect 24259 19805 24268 19839
rect 24216 19796 24268 19805
rect 16028 19660 16080 19712
rect 20812 19660 20864 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 9036 19456 9088 19508
rect 9772 19499 9824 19508
rect 9772 19465 9781 19499
rect 9781 19465 9815 19499
rect 9815 19465 9824 19499
rect 9772 19456 9824 19465
rect 12348 19456 12400 19508
rect 12716 19499 12768 19508
rect 12716 19465 12725 19499
rect 12725 19465 12759 19499
rect 12759 19465 12768 19499
rect 12716 19456 12768 19465
rect 15292 19499 15344 19508
rect 15292 19465 15301 19499
rect 15301 19465 15335 19499
rect 15335 19465 15344 19499
rect 15292 19456 15344 19465
rect 16120 19499 16172 19508
rect 16120 19465 16129 19499
rect 16129 19465 16163 19499
rect 16163 19465 16172 19499
rect 16120 19456 16172 19465
rect 19340 19499 19392 19508
rect 19340 19465 19349 19499
rect 19349 19465 19383 19499
rect 19383 19465 19392 19499
rect 19340 19456 19392 19465
rect 19984 19456 20036 19508
rect 23020 19456 23072 19508
rect 23940 19456 23992 19508
rect 7380 19320 7432 19372
rect 13084 19320 13136 19372
rect 14556 19363 14608 19372
rect 10876 19295 10928 19304
rect 10876 19261 10885 19295
rect 10885 19261 10919 19295
rect 10919 19261 10928 19295
rect 10876 19252 10928 19261
rect 14556 19329 14565 19363
rect 14565 19329 14599 19363
rect 14599 19329 14608 19363
rect 14556 19320 14608 19329
rect 20444 19388 20496 19440
rect 24032 19388 24084 19440
rect 26056 19431 26108 19440
rect 26056 19397 26065 19431
rect 26065 19397 26099 19431
rect 26099 19397 26108 19431
rect 26056 19388 26108 19397
rect 20536 19363 20588 19372
rect 20536 19329 20545 19363
rect 20545 19329 20579 19363
rect 20579 19329 20588 19363
rect 20536 19320 20588 19329
rect 20996 19320 21048 19372
rect 22008 19320 22060 19372
rect 24216 19320 24268 19372
rect 13912 19252 13964 19304
rect 16304 19295 16356 19304
rect 8852 19116 8904 19168
rect 10140 19159 10192 19168
rect 10140 19125 10149 19159
rect 10149 19125 10183 19159
rect 10183 19125 10192 19159
rect 10140 19116 10192 19125
rect 11060 19116 11112 19168
rect 11244 19159 11296 19168
rect 11244 19125 11253 19159
rect 11253 19125 11287 19159
rect 11287 19125 11296 19159
rect 11244 19116 11296 19125
rect 13176 19116 13228 19168
rect 13820 19116 13872 19168
rect 16304 19261 16313 19295
rect 16313 19261 16347 19295
rect 16347 19261 16356 19295
rect 16304 19252 16356 19261
rect 17960 19252 18012 19304
rect 21272 19295 21324 19304
rect 21272 19261 21281 19295
rect 21281 19261 21315 19295
rect 21315 19261 21324 19295
rect 21272 19252 21324 19261
rect 19984 19227 20036 19236
rect 19984 19193 19993 19227
rect 19993 19193 20027 19227
rect 20027 19193 20036 19227
rect 19984 19184 20036 19193
rect 20812 19184 20864 19236
rect 22100 19227 22152 19236
rect 22100 19193 22109 19227
rect 22109 19193 22143 19227
rect 22143 19193 22152 19227
rect 22100 19184 22152 19193
rect 24032 19227 24084 19236
rect 24032 19193 24041 19227
rect 24041 19193 24075 19227
rect 24075 19193 24084 19227
rect 24032 19184 24084 19193
rect 15476 19116 15528 19168
rect 16764 19116 16816 19168
rect 17592 19116 17644 19168
rect 18144 19116 18196 19168
rect 22376 19159 22428 19168
rect 22376 19125 22385 19159
rect 22385 19125 22419 19159
rect 22419 19125 22428 19159
rect 22376 19116 22428 19125
rect 22468 19116 22520 19168
rect 23756 19116 23808 19168
rect 23940 19116 23992 19168
rect 25136 19116 25188 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 11244 18844 11296 18896
rect 12256 18912 12308 18964
rect 13912 18955 13964 18964
rect 12900 18887 12952 18896
rect 12900 18853 12909 18887
rect 12909 18853 12943 18887
rect 12943 18853 12952 18887
rect 12900 18844 12952 18853
rect 13912 18921 13921 18955
rect 13921 18921 13955 18955
rect 13955 18921 13964 18955
rect 13912 18912 13964 18921
rect 16304 18955 16356 18964
rect 16304 18921 16313 18955
rect 16313 18921 16347 18955
rect 16347 18921 16356 18955
rect 16304 18912 16356 18921
rect 20444 18912 20496 18964
rect 22376 18912 22428 18964
rect 23020 18955 23072 18964
rect 23020 18921 23029 18955
rect 23029 18921 23063 18955
rect 23063 18921 23072 18955
rect 23020 18912 23072 18921
rect 23388 18912 23440 18964
rect 23940 18955 23992 18964
rect 23940 18921 23949 18955
rect 23949 18921 23983 18955
rect 23983 18921 23992 18955
rect 23940 18912 23992 18921
rect 27620 18912 27672 18964
rect 15752 18844 15804 18896
rect 18972 18887 19024 18896
rect 18972 18853 18981 18887
rect 18981 18853 19015 18887
rect 19015 18853 19024 18887
rect 18972 18844 19024 18853
rect 23848 18844 23900 18896
rect 20996 18819 21048 18828
rect 20996 18785 21005 18819
rect 21005 18785 21039 18819
rect 21039 18785 21048 18819
rect 20996 18776 21048 18785
rect 22100 18819 22152 18828
rect 22100 18785 22109 18819
rect 22109 18785 22143 18819
rect 22143 18785 22152 18819
rect 22100 18776 22152 18785
rect 23112 18776 23164 18828
rect 24676 18776 24728 18828
rect 11336 18708 11388 18760
rect 16120 18708 16172 18760
rect 17776 18751 17828 18760
rect 17776 18717 17785 18751
rect 17785 18717 17819 18751
rect 17819 18717 17828 18751
rect 17776 18708 17828 18717
rect 18880 18751 18932 18760
rect 18880 18717 18889 18751
rect 18889 18717 18923 18751
rect 18923 18717 18932 18751
rect 18880 18708 18932 18717
rect 23480 18708 23532 18760
rect 25228 18708 25280 18760
rect 15936 18683 15988 18692
rect 15936 18649 15945 18683
rect 15945 18649 15979 18683
rect 15979 18649 15988 18683
rect 15936 18640 15988 18649
rect 19248 18640 19300 18692
rect 19432 18683 19484 18692
rect 19432 18649 19441 18683
rect 19441 18649 19475 18683
rect 19475 18649 19484 18683
rect 19432 18640 19484 18649
rect 10140 18572 10192 18624
rect 12532 18615 12584 18624
rect 12532 18581 12541 18615
rect 12541 18581 12575 18615
rect 12575 18581 12584 18615
rect 12532 18572 12584 18581
rect 17960 18572 18012 18624
rect 21548 18572 21600 18624
rect 25228 18572 25280 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 11244 18368 11296 18420
rect 16120 18411 16172 18420
rect 16120 18377 16129 18411
rect 16129 18377 16163 18411
rect 16163 18377 16172 18411
rect 16120 18368 16172 18377
rect 7472 18300 7524 18352
rect 8852 18275 8904 18284
rect 8852 18241 8861 18275
rect 8861 18241 8895 18275
rect 8895 18241 8904 18275
rect 8852 18232 8904 18241
rect 11336 18300 11388 18352
rect 15936 18232 15988 18284
rect 18880 18368 18932 18420
rect 22100 18368 22152 18420
rect 24676 18411 24728 18420
rect 24676 18377 24685 18411
rect 24685 18377 24719 18411
rect 24719 18377 24728 18411
rect 24676 18368 24728 18377
rect 27620 18300 27672 18352
rect 10140 18164 10192 18216
rect 10876 18164 10928 18216
rect 12900 18164 12952 18216
rect 18972 18207 19024 18216
rect 18972 18173 18981 18207
rect 18981 18173 19015 18207
rect 19015 18173 19024 18207
rect 18972 18164 19024 18173
rect 20352 18164 20404 18216
rect 21916 18232 21968 18284
rect 22284 18232 22336 18284
rect 21088 18207 21140 18216
rect 21088 18173 21097 18207
rect 21097 18173 21131 18207
rect 21131 18173 21140 18207
rect 21088 18164 21140 18173
rect 8944 18139 8996 18148
rect 8944 18105 8953 18139
rect 8953 18105 8987 18139
rect 8987 18105 8996 18139
rect 8944 18096 8996 18105
rect 9496 18139 9548 18148
rect 9496 18105 9505 18139
rect 9505 18105 9539 18139
rect 9539 18105 9548 18139
rect 9496 18096 9548 18105
rect 9772 18028 9824 18080
rect 14832 18139 14884 18148
rect 14832 18105 14841 18139
rect 14841 18105 14875 18139
rect 14875 18105 14884 18139
rect 14832 18096 14884 18105
rect 19156 18139 19208 18148
rect 13636 18028 13688 18080
rect 19156 18105 19165 18139
rect 19165 18105 19199 18139
rect 19199 18105 19208 18139
rect 19156 18096 19208 18105
rect 19524 18096 19576 18148
rect 24032 18164 24084 18216
rect 25228 18207 25280 18216
rect 25228 18173 25237 18207
rect 25237 18173 25271 18207
rect 25271 18173 25280 18207
rect 25228 18164 25280 18173
rect 25044 18096 25096 18148
rect 15384 18028 15436 18080
rect 15752 18071 15804 18080
rect 15752 18037 15761 18071
rect 15761 18037 15795 18071
rect 15795 18037 15804 18071
rect 15752 18028 15804 18037
rect 16948 18071 17000 18080
rect 16948 18037 16957 18071
rect 16957 18037 16991 18071
rect 16991 18037 17000 18071
rect 16948 18028 17000 18037
rect 22284 18028 22336 18080
rect 23388 18028 23440 18080
rect 24032 18028 24084 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 8852 17867 8904 17876
rect 8852 17833 8861 17867
rect 8861 17833 8895 17867
rect 8895 17833 8904 17867
rect 8852 17824 8904 17833
rect 8944 17824 8996 17876
rect 14832 17867 14884 17876
rect 9772 17756 9824 17808
rect 14832 17833 14841 17867
rect 14841 17833 14875 17867
rect 14875 17833 14884 17867
rect 14832 17824 14884 17833
rect 15752 17867 15804 17876
rect 15752 17833 15761 17867
rect 15761 17833 15795 17867
rect 15795 17833 15804 17867
rect 15752 17824 15804 17833
rect 17960 17867 18012 17876
rect 17960 17833 17969 17867
rect 17969 17833 18003 17867
rect 18003 17833 18012 17867
rect 17960 17824 18012 17833
rect 22008 17867 22060 17876
rect 22008 17833 22017 17867
rect 22017 17833 22051 17867
rect 22051 17833 22060 17867
rect 22008 17824 22060 17833
rect 14004 17756 14056 17808
rect 11520 17731 11572 17740
rect 11520 17697 11529 17731
rect 11529 17697 11563 17731
rect 11563 17697 11572 17731
rect 11520 17688 11572 17697
rect 15384 17731 15436 17740
rect 15384 17697 15393 17731
rect 15393 17697 15427 17731
rect 15427 17697 15436 17731
rect 15384 17688 15436 17697
rect 16856 17731 16908 17740
rect 16856 17697 16865 17731
rect 16865 17697 16899 17731
rect 16899 17697 16908 17731
rect 16856 17688 16908 17697
rect 16948 17688 17000 17740
rect 17776 17756 17828 17808
rect 18788 17756 18840 17808
rect 19156 17756 19208 17808
rect 20812 17756 20864 17808
rect 17868 17688 17920 17740
rect 22284 17756 22336 17808
rect 24768 17756 24820 17808
rect 9680 17663 9732 17672
rect 9680 17629 9689 17663
rect 9689 17629 9723 17663
rect 9723 17629 9732 17663
rect 9680 17620 9732 17629
rect 10416 17620 10468 17672
rect 19432 17663 19484 17672
rect 19432 17629 19441 17663
rect 19441 17629 19475 17663
rect 19475 17629 19484 17663
rect 19432 17620 19484 17629
rect 21088 17552 21140 17604
rect 21364 17552 21416 17604
rect 23388 17688 23440 17740
rect 22100 17663 22152 17672
rect 22100 17629 22109 17663
rect 22109 17629 22143 17663
rect 22143 17629 22152 17663
rect 22100 17620 22152 17629
rect 23572 17620 23624 17672
rect 23756 17620 23808 17672
rect 24032 17552 24084 17604
rect 24676 17620 24728 17672
rect 12624 17484 12676 17536
rect 13268 17527 13320 17536
rect 13268 17493 13277 17527
rect 13277 17493 13311 17527
rect 13311 17493 13320 17527
rect 13268 17484 13320 17493
rect 18236 17527 18288 17536
rect 18236 17493 18245 17527
rect 18245 17493 18279 17527
rect 18279 17493 18288 17527
rect 18236 17484 18288 17493
rect 21824 17484 21876 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 11520 17323 11572 17332
rect 11520 17289 11529 17323
rect 11529 17289 11563 17323
rect 11563 17289 11572 17323
rect 11520 17280 11572 17289
rect 13636 17323 13688 17332
rect 13636 17289 13645 17323
rect 13645 17289 13679 17323
rect 13679 17289 13688 17323
rect 13636 17280 13688 17289
rect 17684 17280 17736 17332
rect 18972 17323 19024 17332
rect 18972 17289 18981 17323
rect 18981 17289 19015 17323
rect 19015 17289 19024 17323
rect 18972 17280 19024 17289
rect 19156 17280 19208 17332
rect 20352 17323 20404 17332
rect 20352 17289 20361 17323
rect 20361 17289 20395 17323
rect 20395 17289 20404 17323
rect 20352 17280 20404 17289
rect 9496 17212 9548 17264
rect 12532 17212 12584 17264
rect 18788 17212 18840 17264
rect 9680 17144 9732 17196
rect 10968 17144 11020 17196
rect 14832 17187 14884 17196
rect 14832 17153 14841 17187
rect 14841 17153 14875 17187
rect 14875 17153 14884 17187
rect 14832 17144 14884 17153
rect 16948 17187 17000 17196
rect 9036 17076 9088 17128
rect 9220 17119 9272 17128
rect 9220 17085 9229 17119
rect 9229 17085 9263 17119
rect 9263 17085 9272 17119
rect 9220 17076 9272 17085
rect 12624 17076 12676 17128
rect 13636 17076 13688 17128
rect 14188 17076 14240 17128
rect 10416 17051 10468 17060
rect 10416 17017 10425 17051
rect 10425 17017 10459 17051
rect 10459 17017 10468 17051
rect 10416 17008 10468 17017
rect 14280 17008 14332 17060
rect 9772 16983 9824 16992
rect 9772 16949 9781 16983
rect 9781 16949 9815 16983
rect 9815 16949 9824 16983
rect 9772 16940 9824 16949
rect 12716 16940 12768 16992
rect 14004 16940 14056 16992
rect 14372 16983 14424 16992
rect 14372 16949 14381 16983
rect 14381 16949 14415 16983
rect 14415 16949 14424 16983
rect 16948 17153 16957 17187
rect 16957 17153 16991 17187
rect 16991 17153 17000 17187
rect 16948 17144 17000 17153
rect 18328 17144 18380 17196
rect 20352 17144 20404 17196
rect 17132 17076 17184 17128
rect 18236 17076 18288 17128
rect 25228 17280 25280 17332
rect 25412 17323 25464 17332
rect 25412 17289 25421 17323
rect 25421 17289 25455 17323
rect 25455 17289 25464 17323
rect 25412 17280 25464 17289
rect 21548 17187 21600 17196
rect 21548 17153 21557 17187
rect 21557 17153 21591 17187
rect 21591 17153 21600 17187
rect 21548 17144 21600 17153
rect 24676 17212 24728 17264
rect 24768 17255 24820 17264
rect 24768 17221 24777 17255
rect 24777 17221 24811 17255
rect 24811 17221 24820 17255
rect 24768 17212 24820 17221
rect 24032 17187 24084 17196
rect 24032 17153 24041 17187
rect 24041 17153 24075 17187
rect 24075 17153 24084 17187
rect 24032 17144 24084 17153
rect 17224 17008 17276 17060
rect 18144 17008 18196 17060
rect 19156 17008 19208 17060
rect 22744 17076 22796 17128
rect 25044 17076 25096 17128
rect 15844 16983 15896 16992
rect 14372 16940 14424 16949
rect 15844 16949 15853 16983
rect 15853 16949 15887 16983
rect 15887 16949 15896 16983
rect 15844 16940 15896 16949
rect 16488 16940 16540 16992
rect 16856 16940 16908 16992
rect 19984 16940 20036 16992
rect 21180 16940 21232 16992
rect 22284 16940 22336 16992
rect 23572 16940 23624 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 9680 16736 9732 16788
rect 10140 16779 10192 16788
rect 10140 16745 10149 16779
rect 10149 16745 10183 16779
rect 10183 16745 10192 16779
rect 10140 16736 10192 16745
rect 13268 16779 13320 16788
rect 13268 16745 13277 16779
rect 13277 16745 13311 16779
rect 13311 16745 13320 16779
rect 13268 16736 13320 16745
rect 15384 16736 15436 16788
rect 16764 16779 16816 16788
rect 16764 16745 16773 16779
rect 16773 16745 16807 16779
rect 16807 16745 16816 16779
rect 16764 16736 16816 16745
rect 18696 16779 18748 16788
rect 18696 16745 18705 16779
rect 18705 16745 18739 16779
rect 18739 16745 18748 16779
rect 18696 16736 18748 16745
rect 20076 16779 20128 16788
rect 20076 16745 20085 16779
rect 20085 16745 20119 16779
rect 20119 16745 20128 16779
rect 20076 16736 20128 16745
rect 20628 16736 20680 16788
rect 22744 16736 22796 16788
rect 23572 16779 23624 16788
rect 23572 16745 23581 16779
rect 23581 16745 23615 16779
rect 23615 16745 23624 16779
rect 23572 16736 23624 16745
rect 23756 16736 23808 16788
rect 9220 16668 9272 16720
rect 9864 16643 9916 16652
rect 9864 16609 9873 16643
rect 9873 16609 9907 16643
rect 9907 16609 9916 16643
rect 9864 16600 9916 16609
rect 13912 16668 13964 16720
rect 11520 16643 11572 16652
rect 11520 16609 11529 16643
rect 11529 16609 11563 16643
rect 11563 16609 11572 16643
rect 11520 16600 11572 16609
rect 13084 16643 13136 16652
rect 13084 16609 13093 16643
rect 13093 16609 13127 16643
rect 13127 16609 13136 16643
rect 13084 16600 13136 16609
rect 13452 16643 13504 16652
rect 13452 16609 13461 16643
rect 13461 16609 13495 16643
rect 13495 16609 13504 16643
rect 13452 16600 13504 16609
rect 15292 16643 15344 16652
rect 15292 16609 15301 16643
rect 15301 16609 15335 16643
rect 15335 16609 15344 16643
rect 15292 16600 15344 16609
rect 16488 16643 16540 16652
rect 16488 16609 16497 16643
rect 16497 16609 16531 16643
rect 16531 16609 16540 16643
rect 16488 16600 16540 16609
rect 16948 16643 17000 16652
rect 16948 16609 16957 16643
rect 16957 16609 16991 16643
rect 16991 16609 17000 16643
rect 16948 16600 17000 16609
rect 17224 16600 17276 16652
rect 18696 16643 18748 16652
rect 18696 16609 18705 16643
rect 18705 16609 18739 16643
rect 18739 16609 18748 16643
rect 18696 16600 18748 16609
rect 21272 16668 21324 16720
rect 22100 16711 22152 16720
rect 22100 16677 22109 16711
rect 22109 16677 22143 16711
rect 22143 16677 22152 16711
rect 22100 16668 22152 16677
rect 21364 16643 21416 16652
rect 11428 16575 11480 16584
rect 11428 16541 11437 16575
rect 11437 16541 11471 16575
rect 11471 16541 11480 16575
rect 11428 16532 11480 16541
rect 13544 16532 13596 16584
rect 21364 16609 21373 16643
rect 21373 16609 21407 16643
rect 21407 16609 21416 16643
rect 21364 16600 21416 16609
rect 23388 16600 23440 16652
rect 24768 16600 24820 16652
rect 9772 16464 9824 16516
rect 12716 16507 12768 16516
rect 12716 16473 12725 16507
rect 12725 16473 12759 16507
rect 12759 16473 12768 16507
rect 12716 16464 12768 16473
rect 10968 16439 11020 16448
rect 10968 16405 10977 16439
rect 10977 16405 11011 16439
rect 11011 16405 11020 16439
rect 10968 16396 11020 16405
rect 14188 16439 14240 16448
rect 14188 16405 14197 16439
rect 14197 16405 14231 16439
rect 14231 16405 14240 16439
rect 14188 16396 14240 16405
rect 14280 16396 14332 16448
rect 16764 16396 16816 16448
rect 17960 16396 18012 16448
rect 24676 16532 24728 16584
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 9220 16192 9272 16244
rect 9864 16192 9916 16244
rect 11520 16235 11572 16244
rect 11520 16201 11529 16235
rect 11529 16201 11563 16235
rect 11563 16201 11572 16235
rect 11520 16192 11572 16201
rect 12348 16192 12400 16244
rect 13544 16235 13596 16244
rect 13544 16201 13553 16235
rect 13553 16201 13587 16235
rect 13587 16201 13596 16235
rect 13544 16192 13596 16201
rect 14372 16235 14424 16244
rect 14372 16201 14381 16235
rect 14381 16201 14415 16235
rect 14415 16201 14424 16235
rect 14372 16192 14424 16201
rect 17132 16235 17184 16244
rect 17132 16201 17141 16235
rect 17141 16201 17175 16235
rect 17175 16201 17184 16235
rect 17132 16192 17184 16201
rect 16948 16099 17000 16108
rect 16948 16065 16957 16099
rect 16957 16065 16991 16099
rect 16991 16065 17000 16099
rect 16948 16056 17000 16065
rect 9864 16031 9916 16040
rect 9864 15997 9873 16031
rect 9873 15997 9907 16031
rect 9907 15997 9916 16031
rect 9864 15988 9916 15997
rect 10692 15988 10744 16040
rect 12348 15988 12400 16040
rect 12992 16031 13044 16040
rect 12992 15997 13001 16031
rect 13001 15997 13035 16031
rect 13035 15997 13044 16031
rect 12992 15988 13044 15997
rect 13452 15988 13504 16040
rect 14188 16031 14240 16040
rect 14188 15997 14197 16031
rect 14197 15997 14231 16031
rect 14231 15997 14240 16031
rect 14188 15988 14240 15997
rect 14648 15920 14700 15972
rect 15844 15963 15896 15972
rect 15844 15929 15853 15963
rect 15853 15929 15887 15963
rect 15887 15929 15896 15963
rect 16764 15988 16816 16040
rect 17868 16031 17920 16040
rect 17868 15997 17877 16031
rect 17877 15997 17911 16031
rect 17911 15997 17920 16031
rect 17868 15988 17920 15997
rect 21272 16192 21324 16244
rect 21824 16192 21876 16244
rect 23388 16235 23440 16244
rect 18696 16124 18748 16176
rect 20260 16124 20312 16176
rect 20076 16099 20128 16108
rect 20076 16065 20085 16099
rect 20085 16065 20119 16099
rect 20119 16065 20128 16099
rect 20076 16056 20128 16065
rect 20536 16099 20588 16108
rect 20536 16065 20545 16099
rect 20545 16065 20579 16099
rect 20579 16065 20588 16099
rect 20536 16056 20588 16065
rect 15844 15920 15896 15929
rect 17960 15920 18012 15972
rect 19432 15988 19484 16040
rect 23388 16201 23397 16235
rect 23397 16201 23431 16235
rect 23431 16201 23440 16235
rect 23388 16192 23440 16201
rect 27620 16124 27672 16176
rect 23940 16031 23992 16040
rect 18880 15920 18932 15972
rect 10140 15895 10192 15904
rect 10140 15861 10149 15895
rect 10149 15861 10183 15895
rect 10183 15861 10192 15895
rect 10140 15852 10192 15861
rect 12624 15895 12676 15904
rect 12624 15861 12633 15895
rect 12633 15861 12667 15895
rect 12667 15861 12676 15895
rect 12624 15852 12676 15861
rect 15292 15895 15344 15904
rect 15292 15861 15301 15895
rect 15301 15861 15335 15895
rect 15335 15861 15344 15895
rect 15292 15852 15344 15861
rect 20904 15920 20956 15972
rect 21364 15963 21416 15972
rect 21364 15929 21373 15963
rect 21373 15929 21407 15963
rect 21407 15929 21416 15963
rect 21364 15920 21416 15929
rect 23572 15920 23624 15972
rect 23940 15997 23949 16031
rect 23949 15997 23983 16031
rect 23983 15997 23992 16031
rect 23940 15988 23992 15997
rect 24584 15920 24636 15972
rect 22560 15852 22612 15904
rect 24032 15852 24084 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 9036 15648 9088 15700
rect 12992 15648 13044 15700
rect 16948 15648 17000 15700
rect 19156 15691 19208 15700
rect 19156 15657 19165 15691
rect 19165 15657 19199 15691
rect 19199 15657 19208 15691
rect 19156 15648 19208 15657
rect 19984 15691 20036 15700
rect 19984 15657 19993 15691
rect 19993 15657 20027 15691
rect 20027 15657 20036 15691
rect 19984 15648 20036 15657
rect 22100 15691 22152 15700
rect 22100 15657 22109 15691
rect 22109 15657 22143 15691
rect 22143 15657 22152 15691
rect 22100 15648 22152 15657
rect 22468 15648 22520 15700
rect 23388 15691 23440 15700
rect 23388 15657 23397 15691
rect 23397 15657 23431 15691
rect 23431 15657 23440 15691
rect 23940 15691 23992 15700
rect 23388 15648 23440 15657
rect 23940 15657 23949 15691
rect 23949 15657 23983 15691
rect 23983 15657 23992 15691
rect 23940 15648 23992 15657
rect 11428 15580 11480 15632
rect 16488 15623 16540 15632
rect 9680 15555 9732 15564
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 11796 15444 11848 15496
rect 11704 15419 11756 15428
rect 11704 15385 11713 15419
rect 11713 15385 11747 15419
rect 11747 15385 11756 15419
rect 11704 15376 11756 15385
rect 10048 15308 10100 15360
rect 10692 15308 10744 15360
rect 11612 15308 11664 15360
rect 12900 15308 12952 15360
rect 16488 15589 16497 15623
rect 16497 15589 16531 15623
rect 16531 15589 16540 15623
rect 16488 15580 16540 15589
rect 15384 15512 15436 15564
rect 16948 15512 17000 15564
rect 21272 15580 21324 15632
rect 22284 15580 22336 15632
rect 21180 15512 21232 15564
rect 13084 15444 13136 15496
rect 15568 15444 15620 15496
rect 18880 15444 18932 15496
rect 22468 15487 22520 15496
rect 22468 15453 22477 15487
rect 22477 15453 22511 15487
rect 22511 15453 22520 15487
rect 22468 15444 22520 15453
rect 24584 15487 24636 15496
rect 17224 15376 17276 15428
rect 24584 15453 24593 15487
rect 24593 15453 24627 15487
rect 24627 15453 24636 15487
rect 24584 15444 24636 15453
rect 24768 15444 24820 15496
rect 24860 15376 24912 15428
rect 13452 15351 13504 15360
rect 13452 15317 13461 15351
rect 13461 15317 13495 15351
rect 13495 15317 13504 15351
rect 13452 15308 13504 15317
rect 14004 15308 14056 15360
rect 14648 15308 14700 15360
rect 18052 15351 18104 15360
rect 18052 15317 18061 15351
rect 18061 15317 18095 15351
rect 18095 15317 18104 15351
rect 18052 15308 18104 15317
rect 18328 15308 18380 15360
rect 19432 15308 19484 15360
rect 19800 15308 19852 15360
rect 22284 15308 22336 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 11428 15147 11480 15156
rect 11428 15113 11437 15147
rect 11437 15113 11471 15147
rect 11471 15113 11480 15147
rect 11428 15104 11480 15113
rect 11796 15147 11848 15156
rect 11796 15113 11805 15147
rect 11805 15113 11839 15147
rect 11839 15113 11848 15147
rect 13912 15147 13964 15156
rect 11796 15104 11848 15113
rect 9772 15036 9824 15088
rect 9036 14900 9088 14952
rect 10140 14968 10192 15020
rect 10048 14900 10100 14952
rect 9404 14875 9456 14884
rect 9404 14841 9413 14875
rect 9413 14841 9447 14875
rect 9447 14841 9456 14875
rect 9404 14832 9456 14841
rect 9680 14832 9732 14884
rect 11520 15036 11572 15088
rect 13912 15113 13921 15147
rect 13921 15113 13955 15147
rect 13955 15113 13964 15147
rect 13912 15104 13964 15113
rect 15476 15147 15528 15156
rect 15476 15113 15485 15147
rect 15485 15113 15519 15147
rect 15519 15113 15528 15147
rect 15476 15104 15528 15113
rect 16764 15147 16816 15156
rect 16764 15113 16773 15147
rect 16773 15113 16807 15147
rect 16807 15113 16816 15147
rect 16764 15104 16816 15113
rect 18052 15104 18104 15156
rect 20812 15104 20864 15156
rect 21272 15104 21324 15156
rect 23388 15147 23440 15156
rect 23388 15113 23397 15147
rect 23397 15113 23431 15147
rect 23431 15113 23440 15147
rect 23388 15104 23440 15113
rect 24032 15147 24084 15156
rect 24032 15113 24041 15147
rect 24041 15113 24075 15147
rect 24075 15113 24084 15147
rect 24032 15104 24084 15113
rect 24860 15104 24912 15156
rect 14004 15036 14056 15088
rect 19156 15079 19208 15088
rect 19156 15045 19165 15079
rect 19165 15045 19199 15079
rect 19199 15045 19208 15079
rect 19156 15036 19208 15045
rect 19800 15036 19852 15088
rect 20536 15079 20588 15088
rect 20536 15045 20545 15079
rect 20545 15045 20579 15079
rect 20579 15045 20588 15079
rect 20536 15036 20588 15045
rect 13452 14968 13504 15020
rect 13820 15011 13872 15020
rect 13820 14977 13829 15011
rect 13829 14977 13863 15011
rect 13863 14977 13872 15011
rect 13820 14968 13872 14977
rect 15016 14968 15068 15020
rect 15568 14968 15620 15020
rect 15844 14968 15896 15020
rect 18420 15011 18472 15020
rect 18420 14977 18429 15011
rect 18429 14977 18463 15011
rect 18463 14977 18472 15011
rect 18420 14968 18472 14977
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 22100 15011 22152 15020
rect 22100 14977 22109 15011
rect 22109 14977 22143 15011
rect 22143 14977 22152 15011
rect 22100 14968 22152 14977
rect 22376 15011 22428 15020
rect 22376 14977 22385 15011
rect 22385 14977 22419 15011
rect 22419 14977 22428 15011
rect 22376 14968 22428 14977
rect 24308 15011 24360 15020
rect 24308 14977 24317 15011
rect 24317 14977 24351 15011
rect 24351 14977 24360 15011
rect 24308 14968 24360 14977
rect 24676 14968 24728 15020
rect 24768 15011 24820 15020
rect 24768 14977 24777 15011
rect 24777 14977 24811 15011
rect 24811 14977 24820 15011
rect 24768 14968 24820 14977
rect 12256 14943 12308 14952
rect 12256 14909 12265 14943
rect 12265 14909 12299 14943
rect 12299 14909 12308 14943
rect 12256 14900 12308 14909
rect 13084 14900 13136 14952
rect 15292 14900 15344 14952
rect 18328 14900 18380 14952
rect 10048 14807 10100 14816
rect 10048 14773 10057 14807
rect 10057 14773 10091 14807
rect 10091 14773 10100 14807
rect 10048 14764 10100 14773
rect 12900 14832 12952 14884
rect 14648 14832 14700 14884
rect 15384 14832 15436 14884
rect 10784 14764 10836 14816
rect 13820 14764 13872 14816
rect 14556 14807 14608 14816
rect 14556 14773 14565 14807
rect 14565 14773 14599 14807
rect 14599 14773 14608 14807
rect 14556 14764 14608 14773
rect 16488 14807 16540 14816
rect 16488 14773 16497 14807
rect 16497 14773 16531 14807
rect 16531 14773 16540 14807
rect 16488 14764 16540 14773
rect 17776 14807 17828 14816
rect 17776 14773 17785 14807
rect 17785 14773 17819 14807
rect 17819 14773 17828 14807
rect 17776 14764 17828 14773
rect 19524 14764 19576 14816
rect 21180 14764 21232 14816
rect 21916 14807 21968 14816
rect 21916 14773 21925 14807
rect 21925 14773 21959 14807
rect 21959 14773 21968 14807
rect 21916 14764 21968 14773
rect 22284 14764 22336 14816
rect 24032 14764 24084 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 9036 14560 9088 14612
rect 10140 14560 10192 14612
rect 12900 14603 12952 14612
rect 12900 14569 12909 14603
rect 12909 14569 12943 14603
rect 12943 14569 12952 14603
rect 12900 14560 12952 14569
rect 14832 14560 14884 14612
rect 15016 14603 15068 14612
rect 15016 14569 15025 14603
rect 15025 14569 15059 14603
rect 15059 14569 15068 14603
rect 15016 14560 15068 14569
rect 15568 14560 15620 14612
rect 11520 14492 11572 14544
rect 11612 14492 11664 14544
rect 15384 14467 15436 14476
rect 11336 14356 11388 14408
rect 11704 14331 11756 14340
rect 11704 14297 11713 14331
rect 11713 14297 11747 14331
rect 11747 14297 11756 14331
rect 11704 14288 11756 14297
rect 13268 14288 13320 14340
rect 15384 14433 15393 14467
rect 15393 14433 15427 14467
rect 15427 14433 15436 14467
rect 15384 14424 15436 14433
rect 13820 14356 13872 14408
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 14648 14288 14700 14340
rect 18880 14603 18932 14612
rect 18880 14569 18889 14603
rect 18889 14569 18923 14603
rect 18923 14569 18932 14603
rect 18880 14560 18932 14569
rect 19524 14603 19576 14612
rect 19524 14569 19533 14603
rect 19533 14569 19567 14603
rect 19567 14569 19576 14603
rect 19524 14560 19576 14569
rect 22468 14603 22520 14612
rect 22468 14569 22477 14603
rect 22477 14569 22511 14603
rect 22511 14569 22520 14603
rect 22468 14560 22520 14569
rect 24308 14603 24360 14612
rect 24308 14569 24317 14603
rect 24317 14569 24351 14603
rect 24351 14569 24360 14603
rect 24308 14560 24360 14569
rect 21180 14492 21232 14544
rect 21824 14492 21876 14544
rect 22376 14492 22428 14544
rect 19524 14467 19576 14476
rect 19524 14433 19533 14467
rect 19533 14433 19567 14467
rect 19567 14433 19576 14467
rect 19524 14424 19576 14433
rect 22928 14467 22980 14476
rect 22928 14433 22937 14467
rect 22937 14433 22971 14467
rect 22971 14433 22980 14467
rect 22928 14424 22980 14433
rect 23572 14424 23624 14476
rect 24676 14424 24728 14476
rect 20352 14356 20404 14408
rect 17868 14288 17920 14340
rect 24768 14331 24820 14340
rect 24768 14297 24777 14331
rect 24777 14297 24811 14331
rect 24811 14297 24820 14331
rect 24768 14288 24820 14297
rect 13452 14220 13504 14272
rect 14556 14220 14608 14272
rect 16488 14220 16540 14272
rect 17408 14263 17460 14272
rect 17408 14229 17417 14263
rect 17417 14229 17451 14263
rect 17451 14229 17460 14263
rect 17408 14220 17460 14229
rect 18052 14220 18104 14272
rect 23296 14263 23348 14272
rect 23296 14229 23305 14263
rect 23305 14229 23339 14263
rect 23339 14229 23348 14263
rect 23296 14220 23348 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 9404 14016 9456 14068
rect 10048 14016 10100 14068
rect 11520 14016 11572 14068
rect 13452 14016 13504 14068
rect 14832 14059 14884 14068
rect 14832 14025 14841 14059
rect 14841 14025 14875 14059
rect 14875 14025 14884 14059
rect 14832 14016 14884 14025
rect 15384 14016 15436 14068
rect 16212 14016 16264 14068
rect 17408 14059 17460 14068
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 18052 14016 18104 14068
rect 19524 14059 19576 14068
rect 19524 14025 19533 14059
rect 19533 14025 19567 14059
rect 19567 14025 19576 14059
rect 19524 14016 19576 14025
rect 20352 14016 20404 14068
rect 21916 14059 21968 14068
rect 21916 14025 21925 14059
rect 21925 14025 21959 14059
rect 21959 14025 21968 14059
rect 21916 14016 21968 14025
rect 22928 14059 22980 14068
rect 22928 14025 22937 14059
rect 22937 14025 22971 14059
rect 22971 14025 22980 14059
rect 22928 14016 22980 14025
rect 23296 14016 23348 14068
rect 24676 14059 24728 14068
rect 24676 14025 24685 14059
rect 24685 14025 24719 14059
rect 24719 14025 24728 14059
rect 24676 14016 24728 14025
rect 25412 14059 25464 14068
rect 25412 14025 25421 14059
rect 25421 14025 25455 14059
rect 25455 14025 25464 14059
rect 25412 14016 25464 14025
rect 13728 13991 13780 14000
rect 13728 13957 13737 13991
rect 13737 13957 13771 13991
rect 13771 13957 13780 13991
rect 13728 13948 13780 13957
rect 14648 13948 14700 14000
rect 15568 13991 15620 14000
rect 15568 13957 15577 13991
rect 15577 13957 15611 13991
rect 15611 13957 15620 13991
rect 15568 13948 15620 13957
rect 16488 13948 16540 14000
rect 17132 13948 17184 14000
rect 13820 13923 13872 13932
rect 13820 13889 13829 13923
rect 13829 13889 13863 13923
rect 13863 13889 13872 13923
rect 13820 13880 13872 13889
rect 16764 13923 16816 13932
rect 16764 13889 16773 13923
rect 16773 13889 16807 13923
rect 16807 13889 16816 13923
rect 16764 13880 16816 13889
rect 13268 13812 13320 13864
rect 15844 13812 15896 13864
rect 17960 13812 18012 13864
rect 22560 13948 22612 14000
rect 18328 13880 18380 13932
rect 18420 13923 18472 13932
rect 18420 13889 18429 13923
rect 18429 13889 18463 13923
rect 18463 13889 18472 13923
rect 18420 13880 18472 13889
rect 20904 13880 20956 13932
rect 22744 13880 22796 13932
rect 19064 13855 19116 13864
rect 11060 13744 11112 13796
rect 16396 13787 16448 13796
rect 16396 13753 16405 13787
rect 16405 13753 16439 13787
rect 16439 13753 16448 13787
rect 16396 13744 16448 13753
rect 10140 13719 10192 13728
rect 10140 13685 10149 13719
rect 10149 13685 10183 13719
rect 10183 13685 10192 13719
rect 10140 13676 10192 13685
rect 10692 13719 10744 13728
rect 10692 13685 10701 13719
rect 10701 13685 10735 13719
rect 10735 13685 10744 13719
rect 10692 13676 10744 13685
rect 11336 13676 11388 13728
rect 12900 13676 12952 13728
rect 14556 13719 14608 13728
rect 14556 13685 14565 13719
rect 14565 13685 14599 13719
rect 14599 13685 14608 13719
rect 14556 13676 14608 13685
rect 14832 13676 14884 13728
rect 16212 13719 16264 13728
rect 16212 13685 16221 13719
rect 16221 13685 16255 13719
rect 16255 13685 16264 13719
rect 16212 13676 16264 13685
rect 17868 13719 17920 13728
rect 17868 13685 17877 13719
rect 17877 13685 17911 13719
rect 17911 13685 17920 13719
rect 19064 13821 19073 13855
rect 19073 13821 19107 13855
rect 19107 13821 19116 13855
rect 19064 13812 19116 13821
rect 19340 13812 19392 13864
rect 21824 13855 21876 13864
rect 21824 13821 21833 13855
rect 21833 13821 21867 13855
rect 21867 13821 21876 13855
rect 21824 13812 21876 13821
rect 23756 13787 23808 13796
rect 23756 13753 23765 13787
rect 23765 13753 23799 13787
rect 23799 13753 23808 13787
rect 23756 13744 23808 13753
rect 17868 13676 17920 13685
rect 19984 13676 20036 13728
rect 23296 13676 23348 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 12900 13515 12952 13524
rect 11152 13404 11204 13456
rect 12900 13481 12909 13515
rect 12909 13481 12943 13515
rect 12943 13481 12952 13515
rect 12900 13472 12952 13481
rect 13084 13472 13136 13524
rect 14740 13472 14792 13524
rect 16304 13472 16356 13524
rect 16396 13472 16448 13524
rect 17776 13472 17828 13524
rect 18052 13515 18104 13524
rect 18052 13481 18061 13515
rect 18061 13481 18095 13515
rect 18095 13481 18104 13515
rect 18052 13472 18104 13481
rect 18512 13515 18564 13524
rect 18512 13481 18521 13515
rect 18521 13481 18555 13515
rect 18555 13481 18564 13515
rect 18512 13472 18564 13481
rect 21272 13515 21324 13524
rect 21272 13481 21281 13515
rect 21281 13481 21315 13515
rect 21315 13481 21324 13515
rect 21272 13472 21324 13481
rect 21824 13515 21876 13524
rect 21824 13481 21833 13515
rect 21833 13481 21867 13515
rect 21867 13481 21876 13515
rect 21824 13472 21876 13481
rect 14004 13404 14056 13456
rect 16672 13404 16724 13456
rect 16856 13404 16908 13456
rect 22284 13404 22336 13456
rect 22376 13404 22428 13456
rect 22928 13404 22980 13456
rect 24676 13404 24728 13456
rect 12440 13379 12492 13388
rect 12440 13345 12449 13379
rect 12449 13345 12483 13379
rect 12483 13345 12492 13379
rect 12440 13336 12492 13345
rect 13360 13379 13412 13388
rect 13360 13345 13369 13379
rect 13369 13345 13403 13379
rect 13403 13345 13412 13379
rect 13636 13379 13688 13388
rect 13360 13336 13412 13345
rect 13636 13345 13642 13379
rect 13642 13345 13688 13379
rect 13636 13336 13688 13345
rect 15292 13379 15344 13388
rect 15292 13345 15301 13379
rect 15301 13345 15335 13379
rect 15335 13345 15344 13379
rect 15292 13336 15344 13345
rect 15568 13336 15620 13388
rect 19248 13379 19300 13388
rect 19248 13345 19257 13379
rect 19257 13345 19291 13379
rect 19291 13345 19300 13379
rect 19248 13336 19300 13345
rect 19524 13336 19576 13388
rect 11428 13268 11480 13320
rect 13820 13311 13872 13320
rect 13820 13277 13829 13311
rect 13829 13277 13863 13311
rect 13863 13277 13872 13311
rect 13820 13268 13872 13277
rect 14372 13268 14424 13320
rect 10876 13200 10928 13252
rect 11336 13200 11388 13252
rect 12900 13200 12952 13252
rect 13268 13200 13320 13252
rect 13728 13243 13780 13252
rect 13728 13209 13737 13243
rect 13737 13209 13771 13243
rect 13771 13209 13780 13243
rect 13728 13200 13780 13209
rect 14740 13200 14792 13252
rect 16488 13200 16540 13252
rect 16764 13268 16816 13320
rect 21088 13268 21140 13320
rect 22836 13268 22888 13320
rect 25136 13268 25188 13320
rect 17500 13200 17552 13252
rect 24860 13243 24912 13252
rect 24860 13209 24869 13243
rect 24869 13209 24903 13243
rect 24903 13209 24912 13243
rect 24860 13200 24912 13209
rect 12348 13132 12400 13184
rect 14832 13132 14884 13184
rect 15476 13175 15528 13184
rect 15476 13141 15485 13175
rect 15485 13141 15519 13175
rect 15519 13141 15528 13175
rect 15476 13132 15528 13141
rect 15844 13175 15896 13184
rect 15844 13141 15853 13175
rect 15853 13141 15887 13175
rect 15887 13141 15896 13175
rect 15844 13132 15896 13141
rect 17408 13132 17460 13184
rect 17684 13175 17736 13184
rect 17684 13141 17693 13175
rect 17693 13141 17727 13175
rect 17727 13141 17736 13175
rect 17684 13132 17736 13141
rect 18604 13132 18656 13184
rect 23756 13175 23808 13184
rect 23756 13141 23765 13175
rect 23765 13141 23799 13175
rect 23799 13141 23808 13175
rect 23756 13132 23808 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 13268 12971 13320 12980
rect 13268 12937 13277 12971
rect 13277 12937 13311 12971
rect 13311 12937 13320 12971
rect 13268 12928 13320 12937
rect 14740 12971 14792 12980
rect 14740 12937 14764 12971
rect 14764 12937 14792 12971
rect 14740 12928 14792 12937
rect 15568 12971 15620 12980
rect 15568 12937 15577 12971
rect 15577 12937 15611 12971
rect 15611 12937 15620 12971
rect 15568 12928 15620 12937
rect 16488 12928 16540 12980
rect 18604 12928 18656 12980
rect 18880 12928 18932 12980
rect 19984 12928 20036 12980
rect 22376 12971 22428 12980
rect 22376 12937 22385 12971
rect 22385 12937 22419 12971
rect 22419 12937 22428 12971
rect 22376 12928 22428 12937
rect 23112 12971 23164 12980
rect 23112 12937 23121 12971
rect 23121 12937 23155 12971
rect 23155 12937 23164 12971
rect 23112 12928 23164 12937
rect 25136 12971 25188 12980
rect 25136 12937 25145 12971
rect 25145 12937 25179 12971
rect 25179 12937 25188 12971
rect 25136 12928 25188 12937
rect 12440 12860 12492 12912
rect 14832 12903 14884 12912
rect 14832 12869 14841 12903
rect 14841 12869 14875 12903
rect 14875 12869 14884 12903
rect 14832 12860 14884 12869
rect 15660 12860 15712 12912
rect 17500 12860 17552 12912
rect 10876 12835 10928 12844
rect 10876 12801 10885 12835
rect 10885 12801 10919 12835
rect 10919 12801 10928 12835
rect 10876 12792 10928 12801
rect 12256 12792 12308 12844
rect 14924 12835 14976 12844
rect 14924 12801 14933 12835
rect 14933 12801 14967 12835
rect 14967 12801 14976 12835
rect 14924 12792 14976 12801
rect 15752 12792 15804 12844
rect 17132 12835 17184 12844
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 1584 12588 1636 12640
rect 10048 12656 10100 12708
rect 9680 12588 9732 12640
rect 10692 12656 10744 12708
rect 10876 12656 10928 12708
rect 12440 12656 12492 12708
rect 12992 12699 13044 12708
rect 12992 12665 13001 12699
rect 13001 12665 13035 12699
rect 13035 12665 13044 12699
rect 12992 12656 13044 12665
rect 11152 12631 11204 12640
rect 11152 12597 11161 12631
rect 11161 12597 11195 12631
rect 11195 12597 11204 12631
rect 11152 12588 11204 12597
rect 14372 12724 14424 12776
rect 13728 12699 13780 12708
rect 13728 12665 13737 12699
rect 13737 12665 13771 12699
rect 13771 12665 13780 12699
rect 13728 12656 13780 12665
rect 14740 12656 14792 12708
rect 16396 12724 16448 12776
rect 15292 12699 15344 12708
rect 15292 12665 15301 12699
rect 15301 12665 15335 12699
rect 15335 12665 15344 12699
rect 15292 12656 15344 12665
rect 14188 12588 14240 12640
rect 14372 12588 14424 12640
rect 14924 12588 14976 12640
rect 16212 12631 16264 12640
rect 16212 12597 16221 12631
rect 16221 12597 16255 12631
rect 16255 12597 16264 12631
rect 16212 12588 16264 12597
rect 17408 12631 17460 12640
rect 17408 12597 17417 12631
rect 17417 12597 17451 12631
rect 17451 12597 17460 12631
rect 17408 12588 17460 12597
rect 17592 12588 17644 12640
rect 19248 12835 19300 12844
rect 19248 12801 19257 12835
rect 19257 12801 19291 12835
rect 19291 12801 19300 12835
rect 19248 12792 19300 12801
rect 22928 12792 22980 12844
rect 23756 12792 23808 12844
rect 18052 12767 18104 12776
rect 18052 12733 18061 12767
rect 18061 12733 18095 12767
rect 18095 12733 18104 12767
rect 18052 12724 18104 12733
rect 19340 12724 19392 12776
rect 20996 12767 21048 12776
rect 20996 12733 21005 12767
rect 21005 12733 21039 12767
rect 21039 12733 21048 12767
rect 20996 12724 21048 12733
rect 19524 12656 19576 12708
rect 21272 12656 21324 12708
rect 23112 12656 23164 12708
rect 21640 12588 21692 12640
rect 24216 12656 24268 12708
rect 24584 12656 24636 12708
rect 24860 12656 24912 12708
rect 24676 12631 24728 12640
rect 24676 12597 24685 12631
rect 24685 12597 24719 12631
rect 24719 12597 24728 12631
rect 24676 12588 24728 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 10048 12384 10100 12436
rect 12348 12427 12400 12436
rect 12348 12393 12357 12427
rect 12357 12393 12391 12427
rect 12391 12393 12400 12427
rect 12348 12384 12400 12393
rect 12900 12384 12952 12436
rect 12992 12384 13044 12436
rect 13452 12384 13504 12436
rect 13636 12427 13688 12436
rect 13636 12393 13645 12427
rect 13645 12393 13679 12427
rect 13679 12393 13688 12427
rect 13636 12384 13688 12393
rect 13728 12384 13780 12436
rect 14832 12384 14884 12436
rect 16488 12384 16540 12436
rect 16764 12427 16816 12436
rect 16764 12393 16773 12427
rect 16773 12393 16807 12427
rect 16807 12393 16816 12427
rect 16764 12384 16816 12393
rect 16856 12384 16908 12436
rect 18604 12427 18656 12436
rect 18604 12393 18613 12427
rect 18613 12393 18647 12427
rect 18647 12393 18656 12427
rect 18604 12384 18656 12393
rect 21088 12427 21140 12436
rect 21088 12393 21097 12427
rect 21097 12393 21131 12427
rect 21131 12393 21140 12427
rect 21088 12384 21140 12393
rect 11152 12359 11204 12368
rect 11152 12325 11161 12359
rect 11161 12325 11195 12359
rect 11195 12325 11204 12359
rect 11152 12316 11204 12325
rect 14004 12359 14056 12368
rect 14004 12325 14013 12359
rect 14013 12325 14047 12359
rect 14047 12325 14056 12359
rect 14004 12316 14056 12325
rect 14740 12359 14792 12368
rect 14740 12325 14749 12359
rect 14749 12325 14783 12359
rect 14783 12325 14792 12359
rect 14740 12316 14792 12325
rect 17776 12316 17828 12368
rect 20996 12316 21048 12368
rect 21640 12316 21692 12368
rect 24676 12316 24728 12368
rect 9680 12248 9732 12300
rect 12348 12248 12400 12300
rect 12992 12248 13044 12300
rect 14188 12291 14240 12300
rect 14188 12257 14197 12291
rect 14197 12257 14231 12291
rect 14231 12257 14240 12291
rect 14188 12248 14240 12257
rect 15384 12248 15436 12300
rect 13636 12112 13688 12164
rect 16488 12248 16540 12300
rect 19248 12291 19300 12300
rect 19248 12257 19257 12291
rect 19257 12257 19291 12291
rect 19291 12257 19300 12291
rect 19248 12248 19300 12257
rect 19524 12248 19576 12300
rect 24216 12291 24268 12300
rect 24216 12257 24225 12291
rect 24225 12257 24259 12291
rect 24259 12257 24268 12291
rect 24216 12248 24268 12257
rect 25228 12291 25280 12300
rect 25228 12257 25237 12291
rect 25237 12257 25271 12291
rect 25271 12257 25280 12291
rect 25228 12248 25280 12257
rect 15752 12180 15804 12232
rect 17592 12223 17644 12232
rect 17592 12189 17601 12223
rect 17601 12189 17635 12223
rect 17635 12189 17644 12223
rect 17592 12180 17644 12189
rect 22100 12180 22152 12232
rect 16488 12112 16540 12164
rect 17500 12155 17552 12164
rect 11520 12087 11572 12096
rect 11520 12053 11529 12087
rect 11529 12053 11563 12087
rect 11563 12053 11572 12087
rect 11520 12044 11572 12053
rect 14832 12044 14884 12096
rect 15660 12044 15712 12096
rect 16856 12044 16908 12096
rect 17500 12121 17509 12155
rect 17509 12121 17543 12155
rect 17543 12121 17552 12155
rect 17500 12112 17552 12121
rect 20536 12112 20588 12164
rect 25412 12155 25464 12164
rect 25412 12121 25421 12155
rect 25421 12121 25455 12155
rect 25455 12121 25464 12155
rect 25412 12112 25464 12121
rect 18880 12044 18932 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 9680 11883 9732 11892
rect 9680 11849 9689 11883
rect 9689 11849 9723 11883
rect 9723 11849 9732 11883
rect 9680 11840 9732 11849
rect 14188 11840 14240 11892
rect 15660 11883 15712 11892
rect 15660 11849 15669 11883
rect 15669 11849 15703 11883
rect 15703 11849 15712 11883
rect 15660 11840 15712 11849
rect 17776 11883 17828 11892
rect 17776 11849 17785 11883
rect 17785 11849 17819 11883
rect 17819 11849 17828 11883
rect 17776 11840 17828 11849
rect 18880 11883 18932 11892
rect 18880 11849 18889 11883
rect 18889 11849 18923 11883
rect 18923 11849 18932 11883
rect 18880 11840 18932 11849
rect 23664 11840 23716 11892
rect 24216 11883 24268 11892
rect 24216 11849 24225 11883
rect 24225 11849 24259 11883
rect 24259 11849 24268 11883
rect 24216 11840 24268 11849
rect 25228 11840 25280 11892
rect 15752 11772 15804 11824
rect 21364 11772 21416 11824
rect 8944 11704 8996 11756
rect 10876 11679 10928 11688
rect 10876 11645 10885 11679
rect 10885 11645 10919 11679
rect 10919 11645 10928 11679
rect 10876 11636 10928 11645
rect 14464 11704 14516 11756
rect 15476 11704 15528 11756
rect 15844 11704 15896 11756
rect 14832 11636 14884 11688
rect 12440 11611 12492 11620
rect 12440 11577 12449 11611
rect 12449 11577 12483 11611
rect 12483 11577 12492 11611
rect 12440 11568 12492 11577
rect 12992 11611 13044 11620
rect 12992 11577 13001 11611
rect 13001 11577 13035 11611
rect 13035 11577 13044 11611
rect 12992 11568 13044 11577
rect 14740 11611 14792 11620
rect 14740 11577 14749 11611
rect 14749 11577 14783 11611
rect 14783 11577 14792 11611
rect 14740 11568 14792 11577
rect 17592 11636 17644 11688
rect 10140 11500 10192 11552
rect 12348 11500 12400 11552
rect 16396 11500 16448 11552
rect 18696 11500 18748 11552
rect 19248 11543 19300 11552
rect 19248 11509 19257 11543
rect 19257 11509 19291 11543
rect 19291 11509 19300 11543
rect 20536 11679 20588 11688
rect 20536 11645 20545 11679
rect 20545 11645 20579 11679
rect 20579 11645 20588 11679
rect 20536 11636 20588 11645
rect 22652 11636 22704 11688
rect 22744 11568 22796 11620
rect 19248 11500 19300 11509
rect 21640 11500 21692 11552
rect 22100 11543 22152 11552
rect 22100 11509 22109 11543
rect 22109 11509 22143 11543
rect 22143 11509 22152 11543
rect 22100 11500 22152 11509
rect 23940 11500 23992 11552
rect 25228 11543 25280 11552
rect 25228 11509 25237 11543
rect 25237 11509 25271 11543
rect 25271 11509 25280 11543
rect 25228 11500 25280 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 12992 11296 13044 11348
rect 13544 11339 13596 11348
rect 13544 11305 13553 11339
rect 13553 11305 13587 11339
rect 13587 11305 13596 11339
rect 13544 11296 13596 11305
rect 14464 11339 14516 11348
rect 14464 11305 14473 11339
rect 14473 11305 14507 11339
rect 14507 11305 14516 11339
rect 14464 11296 14516 11305
rect 16488 11296 16540 11348
rect 17040 11296 17092 11348
rect 19524 11296 19576 11348
rect 20536 11296 20588 11348
rect 24216 11296 24268 11348
rect 15384 11228 15436 11280
rect 19156 11228 19208 11280
rect 10140 11160 10192 11212
rect 12440 11203 12492 11212
rect 12440 11169 12449 11203
rect 12449 11169 12483 11203
rect 12483 11169 12492 11203
rect 12440 11160 12492 11169
rect 14188 11160 14240 11212
rect 14832 11160 14884 11212
rect 15476 11203 15528 11212
rect 15476 11169 15485 11203
rect 15485 11169 15519 11203
rect 15519 11169 15528 11203
rect 15476 11160 15528 11169
rect 17132 11203 17184 11212
rect 17132 11169 17141 11203
rect 17141 11169 17175 11203
rect 17175 11169 17184 11203
rect 17132 11160 17184 11169
rect 14096 11092 14148 11144
rect 17408 11092 17460 11144
rect 15660 11024 15712 11076
rect 21272 11160 21324 11212
rect 22100 11228 22152 11280
rect 22928 11228 22980 11280
rect 21548 11160 21600 11212
rect 22744 11203 22796 11212
rect 22744 11169 22753 11203
rect 22753 11169 22787 11203
rect 22787 11169 22796 11203
rect 22744 11160 22796 11169
rect 21732 11092 21784 11144
rect 24676 11092 24728 11144
rect 19984 11024 20036 11076
rect 25136 11067 25188 11076
rect 15568 10999 15620 11008
rect 15568 10965 15577 10999
rect 15577 10965 15611 10999
rect 15611 10965 15620 10999
rect 15568 10956 15620 10965
rect 19064 10956 19116 11008
rect 22008 10999 22060 11008
rect 22008 10965 22017 10999
rect 22017 10965 22051 10999
rect 22051 10965 22060 10999
rect 22008 10956 22060 10965
rect 25136 11033 25145 11067
rect 25145 11033 25179 11067
rect 25179 11033 25188 11067
rect 25136 11024 25188 11033
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 14188 10795 14240 10804
rect 14188 10761 14197 10795
rect 14197 10761 14231 10795
rect 14231 10761 14240 10795
rect 14188 10752 14240 10761
rect 15476 10752 15528 10804
rect 16948 10752 17000 10804
rect 19984 10752 20036 10804
rect 21272 10795 21324 10804
rect 21272 10761 21281 10795
rect 21281 10761 21315 10795
rect 21315 10761 21324 10795
rect 21272 10752 21324 10761
rect 21548 10752 21600 10804
rect 22744 10752 22796 10804
rect 23940 10795 23992 10804
rect 23940 10761 23949 10795
rect 23949 10761 23983 10795
rect 23983 10761 23992 10795
rect 23940 10752 23992 10761
rect 24676 10752 24728 10804
rect 12992 10616 13044 10668
rect 13544 10616 13596 10668
rect 16212 10684 16264 10736
rect 22928 10727 22980 10736
rect 14740 10616 14792 10668
rect 16396 10616 16448 10668
rect 17408 10548 17460 10600
rect 19156 10616 19208 10668
rect 21640 10616 21692 10668
rect 22928 10693 22937 10727
rect 22937 10693 22971 10727
rect 22971 10693 22980 10727
rect 22928 10684 22980 10693
rect 22652 10659 22704 10668
rect 22652 10625 22661 10659
rect 22661 10625 22695 10659
rect 22695 10625 22704 10659
rect 22652 10616 22704 10625
rect 25136 10727 25188 10736
rect 25136 10693 25145 10727
rect 25145 10693 25179 10727
rect 25179 10693 25188 10727
rect 25136 10684 25188 10693
rect 18880 10591 18932 10600
rect 18880 10557 18889 10591
rect 18889 10557 18923 10591
rect 18923 10557 18932 10591
rect 18880 10548 18932 10557
rect 15844 10480 15896 10532
rect 17132 10480 17184 10532
rect 19156 10523 19208 10532
rect 19156 10489 19165 10523
rect 19165 10489 19199 10523
rect 19199 10489 19208 10523
rect 19156 10480 19208 10489
rect 20352 10523 20404 10532
rect 20352 10489 20361 10523
rect 20361 10489 20395 10523
rect 20395 10489 20404 10523
rect 20352 10480 20404 10489
rect 22008 10523 22060 10532
rect 9588 10412 9640 10464
rect 10140 10412 10192 10464
rect 13820 10455 13872 10464
rect 13820 10421 13829 10455
rect 13829 10421 13863 10455
rect 13863 10421 13872 10455
rect 16212 10455 16264 10464
rect 13820 10412 13872 10421
rect 16212 10421 16221 10455
rect 16221 10421 16255 10455
rect 16255 10421 16264 10455
rect 16212 10412 16264 10421
rect 17408 10455 17460 10464
rect 17408 10421 17417 10455
rect 17417 10421 17451 10455
rect 17451 10421 17460 10455
rect 17408 10412 17460 10421
rect 17776 10455 17828 10464
rect 17776 10421 17785 10455
rect 17785 10421 17819 10455
rect 17819 10421 17828 10455
rect 17776 10412 17828 10421
rect 20076 10455 20128 10464
rect 20076 10421 20085 10455
rect 20085 10421 20119 10455
rect 20119 10421 20128 10455
rect 22008 10489 22017 10523
rect 22017 10489 22051 10523
rect 22051 10489 22060 10523
rect 22008 10480 22060 10489
rect 20076 10412 20128 10421
rect 21916 10412 21968 10464
rect 24400 10455 24452 10464
rect 24400 10421 24409 10455
rect 24409 10421 24443 10455
rect 24443 10421 24452 10455
rect 24400 10412 24452 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 12992 10251 13044 10260
rect 12992 10217 13001 10251
rect 13001 10217 13035 10251
rect 13035 10217 13044 10251
rect 12992 10208 13044 10217
rect 14740 10251 14792 10260
rect 14740 10217 14749 10251
rect 14749 10217 14783 10251
rect 14783 10217 14792 10251
rect 14740 10208 14792 10217
rect 15384 10208 15436 10260
rect 17684 10208 17736 10260
rect 18328 10208 18380 10260
rect 18880 10208 18932 10260
rect 19156 10208 19208 10260
rect 20352 10251 20404 10260
rect 20352 10217 20361 10251
rect 20361 10217 20395 10251
rect 20395 10217 20404 10251
rect 20352 10208 20404 10217
rect 24400 10251 24452 10260
rect 24400 10217 24409 10251
rect 24409 10217 24443 10251
rect 24443 10217 24452 10251
rect 24400 10208 24452 10217
rect 12900 10140 12952 10192
rect 13820 10140 13872 10192
rect 15568 10140 15620 10192
rect 17776 10183 17828 10192
rect 17776 10149 17785 10183
rect 17785 10149 17819 10183
rect 17819 10149 17828 10183
rect 17776 10140 17828 10149
rect 17224 10115 17276 10124
rect 17224 10081 17233 10115
rect 17233 10081 17267 10115
rect 17267 10081 17276 10115
rect 17224 10072 17276 10081
rect 18696 10115 18748 10124
rect 18696 10081 18705 10115
rect 18705 10081 18739 10115
rect 18739 10081 18748 10115
rect 18696 10072 18748 10081
rect 22560 10183 22612 10192
rect 22560 10149 22569 10183
rect 22569 10149 22603 10183
rect 22603 10149 22612 10183
rect 22560 10140 22612 10149
rect 22652 10140 22704 10192
rect 24216 10115 24268 10124
rect 24216 10081 24225 10115
rect 24225 10081 24259 10115
rect 24259 10081 24268 10115
rect 24216 10072 24268 10081
rect 12164 10004 12216 10056
rect 15384 10047 15436 10056
rect 15384 10013 15393 10047
rect 15393 10013 15427 10047
rect 15427 10013 15436 10047
rect 15384 10004 15436 10013
rect 15660 10047 15712 10056
rect 15660 10013 15669 10047
rect 15669 10013 15703 10047
rect 15703 10013 15712 10047
rect 15660 10004 15712 10013
rect 20352 10004 20404 10056
rect 22744 10004 22796 10056
rect 13728 9979 13780 9988
rect 13728 9945 13737 9979
rect 13737 9945 13771 9979
rect 13771 9945 13780 9979
rect 13728 9936 13780 9945
rect 14188 9911 14240 9920
rect 14188 9877 14197 9911
rect 14197 9877 14231 9911
rect 14231 9877 14240 9911
rect 14188 9868 14240 9877
rect 16396 9911 16448 9920
rect 16396 9877 16405 9911
rect 16405 9877 16439 9911
rect 16439 9877 16448 9911
rect 16396 9868 16448 9877
rect 21916 9911 21968 9920
rect 21916 9877 21925 9911
rect 21925 9877 21959 9911
rect 21959 9877 21968 9911
rect 21916 9868 21968 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 6828 9664 6880 9716
rect 12164 9707 12216 9716
rect 12164 9673 12173 9707
rect 12173 9673 12207 9707
rect 12207 9673 12216 9707
rect 12164 9664 12216 9673
rect 12900 9707 12952 9716
rect 12900 9673 12909 9707
rect 12909 9673 12943 9707
rect 12943 9673 12952 9707
rect 12900 9664 12952 9673
rect 15384 9664 15436 9716
rect 15568 9664 15620 9716
rect 18328 9707 18380 9716
rect 18328 9673 18337 9707
rect 18337 9673 18371 9707
rect 18371 9673 18380 9707
rect 18328 9664 18380 9673
rect 20352 9707 20404 9716
rect 20352 9673 20361 9707
rect 20361 9673 20395 9707
rect 20395 9673 20404 9707
rect 22744 9707 22796 9716
rect 20352 9664 20404 9673
rect 12348 9596 12400 9648
rect 16212 9596 16264 9648
rect 13544 9528 13596 9580
rect 15660 9571 15712 9580
rect 15660 9537 15669 9571
rect 15669 9537 15703 9571
rect 15703 9537 15712 9571
rect 15660 9528 15712 9537
rect 19156 9571 19208 9580
rect 19156 9537 19165 9571
rect 19165 9537 19199 9571
rect 19199 9537 19208 9571
rect 19156 9528 19208 9537
rect 22744 9673 22753 9707
rect 22753 9673 22787 9707
rect 22787 9673 22796 9707
rect 22744 9664 22796 9673
rect 24216 9664 24268 9716
rect 24952 9664 25004 9716
rect 21732 9596 21784 9648
rect 21916 9460 21968 9512
rect 23020 9460 23072 9512
rect 13544 9435 13596 9444
rect 13544 9401 13553 9435
rect 13553 9401 13587 9435
rect 13587 9401 13596 9435
rect 13544 9392 13596 9401
rect 13728 9392 13780 9444
rect 15016 9435 15068 9444
rect 15016 9401 15025 9435
rect 15025 9401 15059 9435
rect 15059 9401 15068 9435
rect 15016 9392 15068 9401
rect 15108 9435 15160 9444
rect 15108 9401 15117 9435
rect 15117 9401 15151 9435
rect 15151 9401 15160 9435
rect 15108 9392 15160 9401
rect 15476 9392 15528 9444
rect 14464 9367 14516 9376
rect 14464 9333 14473 9367
rect 14473 9333 14507 9367
rect 14507 9333 14516 9367
rect 14464 9324 14516 9333
rect 14556 9324 14608 9376
rect 18696 9392 18748 9444
rect 17224 9324 17276 9376
rect 17868 9324 17920 9376
rect 21548 9392 21600 9444
rect 19340 9324 19392 9376
rect 20076 9367 20128 9376
rect 20076 9333 20085 9367
rect 20085 9333 20119 9367
rect 20119 9333 20128 9367
rect 20076 9324 20128 9333
rect 22560 9324 22612 9376
rect 22744 9324 22796 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 13544 9120 13596 9172
rect 15108 9120 15160 9172
rect 15384 9120 15436 9172
rect 17316 9120 17368 9172
rect 24124 9163 24176 9172
rect 24124 9129 24133 9163
rect 24133 9129 24167 9163
rect 24167 9129 24176 9163
rect 24124 9120 24176 9129
rect 24768 9163 24820 9172
rect 24768 9129 24777 9163
rect 24777 9129 24811 9163
rect 24811 9129 24820 9163
rect 24768 9120 24820 9129
rect 15016 9052 15068 9104
rect 21272 9052 21324 9104
rect 22008 9052 22060 9104
rect 22744 9095 22796 9104
rect 22744 9061 22753 9095
rect 22753 9061 22787 9095
rect 22787 9061 22796 9095
rect 22744 9052 22796 9061
rect 12900 8984 12952 9036
rect 17224 9027 17276 9036
rect 17224 8993 17233 9027
rect 17233 8993 17267 9027
rect 17267 8993 17276 9027
rect 17224 8984 17276 8993
rect 17408 9027 17460 9036
rect 17408 8993 17417 9027
rect 17417 8993 17451 9027
rect 17451 8993 17460 9027
rect 17408 8984 17460 8993
rect 19340 9027 19392 9036
rect 19340 8993 19349 9027
rect 19349 8993 19383 9027
rect 19383 8993 19392 9027
rect 19340 8984 19392 8993
rect 23020 9027 23072 9036
rect 23020 8993 23029 9027
rect 23029 8993 23063 9027
rect 23063 8993 23072 9027
rect 23020 8984 23072 8993
rect 25044 8984 25096 9036
rect 21364 8916 21416 8968
rect 18144 8823 18196 8832
rect 18144 8789 18153 8823
rect 18153 8789 18187 8823
rect 18187 8789 18196 8823
rect 18144 8780 18196 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 12900 8576 12952 8628
rect 14188 8576 14240 8628
rect 14556 8576 14608 8628
rect 19340 8619 19392 8628
rect 5172 8372 5224 8424
rect 10784 8372 10836 8424
rect 19340 8585 19349 8619
rect 19349 8585 19383 8619
rect 19383 8585 19392 8619
rect 19340 8576 19392 8585
rect 21272 8619 21324 8628
rect 21272 8585 21281 8619
rect 21281 8585 21315 8619
rect 21315 8585 21324 8619
rect 21272 8576 21324 8585
rect 21364 8576 21416 8628
rect 23480 8576 23532 8628
rect 17224 8508 17276 8560
rect 22468 8508 22520 8560
rect 23020 8551 23072 8560
rect 23020 8517 23029 8551
rect 23029 8517 23063 8551
rect 23063 8517 23072 8551
rect 23020 8508 23072 8517
rect 23112 8508 23164 8560
rect 24216 8508 24268 8560
rect 17408 8440 17460 8492
rect 18972 8440 19024 8492
rect 24124 8483 24176 8492
rect 24124 8449 24133 8483
rect 24133 8449 24167 8483
rect 24167 8449 24176 8483
rect 24124 8440 24176 8449
rect 24308 8440 24360 8492
rect 15292 8372 15344 8424
rect 18144 8415 18196 8424
rect 18144 8381 18153 8415
rect 18153 8381 18187 8415
rect 18187 8381 18196 8415
rect 18144 8372 18196 8381
rect 18696 8372 18748 8424
rect 20720 8415 20772 8424
rect 20720 8381 20729 8415
rect 20729 8381 20763 8415
rect 20763 8381 20772 8415
rect 20720 8372 20772 8381
rect 27620 8576 27672 8628
rect 15936 8347 15988 8356
rect 15936 8313 15945 8347
rect 15945 8313 15979 8347
rect 15979 8313 15988 8347
rect 15936 8304 15988 8313
rect 18788 8347 18840 8356
rect 18788 8313 18797 8347
rect 18797 8313 18831 8347
rect 18831 8313 18840 8347
rect 18788 8304 18840 8313
rect 21732 8304 21784 8356
rect 24216 8347 24268 8356
rect 24216 8313 24225 8347
rect 24225 8313 24259 8347
rect 24259 8313 24268 8347
rect 24216 8304 24268 8313
rect 24400 8236 24452 8288
rect 25044 8279 25096 8288
rect 25044 8245 25053 8279
rect 25053 8245 25087 8279
rect 25087 8245 25096 8279
rect 25044 8236 25096 8245
rect 25136 8236 25188 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 15292 8032 15344 8084
rect 16212 8032 16264 8084
rect 17868 8075 17920 8084
rect 17868 8041 17877 8075
rect 17877 8041 17911 8075
rect 17911 8041 17920 8075
rect 17868 8032 17920 8041
rect 18144 8032 18196 8084
rect 15844 7964 15896 8016
rect 21548 7964 21600 8016
rect 23940 7964 23992 8016
rect 15936 7896 15988 7948
rect 17408 7896 17460 7948
rect 19248 7939 19300 7948
rect 19248 7905 19257 7939
rect 19257 7905 19291 7939
rect 19291 7905 19300 7939
rect 19248 7896 19300 7905
rect 15752 7871 15804 7880
rect 15752 7837 15761 7871
rect 15761 7837 15795 7871
rect 15795 7837 15804 7871
rect 15752 7828 15804 7837
rect 16856 7828 16908 7880
rect 19524 7828 19576 7880
rect 20720 7896 20772 7948
rect 21180 7828 21232 7880
rect 21732 7871 21784 7880
rect 21732 7837 21741 7871
rect 21741 7837 21775 7871
rect 21775 7837 21784 7871
rect 21732 7828 21784 7837
rect 24124 7871 24176 7880
rect 24124 7837 24133 7871
rect 24133 7837 24167 7871
rect 24167 7837 24176 7871
rect 24124 7828 24176 7837
rect 24400 7871 24452 7880
rect 24400 7837 24409 7871
rect 24409 7837 24443 7871
rect 24443 7837 24452 7871
rect 24400 7828 24452 7837
rect 24676 7760 24728 7812
rect 16672 7735 16724 7744
rect 16672 7701 16681 7735
rect 16681 7701 16715 7735
rect 16715 7701 16724 7735
rect 16672 7692 16724 7701
rect 18236 7692 18288 7744
rect 22652 7735 22704 7744
rect 22652 7701 22661 7735
rect 22661 7701 22695 7735
rect 22695 7701 22704 7735
rect 22652 7692 22704 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 15844 7531 15896 7540
rect 15844 7497 15853 7531
rect 15853 7497 15887 7531
rect 15887 7497 15896 7531
rect 15844 7488 15896 7497
rect 17868 7488 17920 7540
rect 18788 7488 18840 7540
rect 19800 7488 19852 7540
rect 21180 7531 21232 7540
rect 21180 7497 21189 7531
rect 21189 7497 21223 7531
rect 21223 7497 21232 7531
rect 21180 7488 21232 7497
rect 14188 7420 14240 7472
rect 19248 7420 19300 7472
rect 21548 7463 21600 7472
rect 21548 7429 21557 7463
rect 21557 7429 21591 7463
rect 21591 7429 21600 7463
rect 21548 7420 21600 7429
rect 15752 7352 15804 7404
rect 16212 7352 16264 7404
rect 18236 7352 18288 7404
rect 23112 7488 23164 7540
rect 23480 7531 23532 7540
rect 23480 7497 23489 7531
rect 23489 7497 23523 7531
rect 23523 7497 23532 7531
rect 23480 7488 23532 7497
rect 24124 7488 24176 7540
rect 25412 7488 25464 7540
rect 23940 7463 23992 7472
rect 23940 7429 23949 7463
rect 23949 7429 23983 7463
rect 23983 7429 23992 7463
rect 23940 7420 23992 7429
rect 24676 7463 24728 7472
rect 24676 7429 24685 7463
rect 24685 7429 24719 7463
rect 24719 7429 24728 7463
rect 24676 7420 24728 7429
rect 15292 7327 15344 7336
rect 15292 7293 15301 7327
rect 15301 7293 15335 7327
rect 15335 7293 15344 7327
rect 15292 7284 15344 7293
rect 24216 7352 24268 7404
rect 27620 7488 27672 7540
rect 16672 7216 16724 7268
rect 18236 7259 18288 7268
rect 18236 7225 18245 7259
rect 18245 7225 18279 7259
rect 18279 7225 18288 7259
rect 18788 7259 18840 7268
rect 18236 7216 18288 7225
rect 18788 7225 18797 7259
rect 18797 7225 18831 7259
rect 18831 7225 18840 7259
rect 18788 7216 18840 7225
rect 19800 7259 19852 7268
rect 19800 7225 19809 7259
rect 19809 7225 19843 7259
rect 19843 7225 19852 7259
rect 19800 7216 19852 7225
rect 21548 7216 21600 7268
rect 22744 7216 22796 7268
rect 20076 7148 20128 7200
rect 23296 7148 23348 7200
rect 23940 7148 23992 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 15292 6944 15344 6996
rect 15752 6987 15804 6996
rect 15752 6953 15761 6987
rect 15761 6953 15795 6987
rect 15795 6953 15804 6987
rect 15752 6944 15804 6953
rect 17408 6987 17460 6996
rect 17408 6953 17417 6987
rect 17417 6953 17451 6987
rect 17451 6953 17460 6987
rect 17408 6944 17460 6953
rect 18236 6944 18288 6996
rect 25044 6944 25096 6996
rect 17684 6876 17736 6928
rect 18328 6919 18380 6928
rect 18328 6885 18337 6919
rect 18337 6885 18371 6919
rect 18371 6885 18380 6919
rect 18328 6876 18380 6885
rect 19524 6876 19576 6928
rect 21732 6876 21784 6928
rect 23296 6919 23348 6928
rect 23296 6885 23305 6919
rect 23305 6885 23339 6919
rect 23339 6885 23348 6919
rect 23296 6876 23348 6885
rect 24676 6876 24728 6928
rect 16672 6851 16724 6860
rect 16672 6817 16681 6851
rect 16681 6817 16715 6851
rect 16715 6817 16724 6851
rect 16672 6808 16724 6817
rect 18788 6808 18840 6860
rect 19248 6851 19300 6860
rect 19248 6817 19292 6851
rect 19292 6817 19300 6851
rect 22652 6851 22704 6860
rect 19248 6808 19300 6817
rect 22652 6817 22661 6851
rect 22661 6817 22695 6851
rect 22695 6817 22704 6851
rect 22652 6808 22704 6817
rect 17316 6740 17368 6792
rect 21548 6740 21600 6792
rect 24216 6783 24268 6792
rect 24216 6749 24225 6783
rect 24225 6749 24259 6783
rect 24259 6749 24268 6783
rect 24216 6740 24268 6749
rect 24308 6740 24360 6792
rect 25964 6672 26016 6724
rect 20076 6647 20128 6656
rect 20076 6613 20085 6647
rect 20085 6613 20119 6647
rect 20119 6613 20128 6647
rect 20076 6604 20128 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 16672 6400 16724 6452
rect 17684 6443 17736 6452
rect 17684 6409 17693 6443
rect 17693 6409 17727 6443
rect 17727 6409 17736 6443
rect 17684 6400 17736 6409
rect 19248 6443 19300 6452
rect 19248 6409 19257 6443
rect 19257 6409 19291 6443
rect 19291 6409 19300 6443
rect 19248 6400 19300 6409
rect 22652 6443 22704 6452
rect 22652 6409 22661 6443
rect 22661 6409 22695 6443
rect 22695 6409 22704 6443
rect 22652 6400 22704 6409
rect 23112 6400 23164 6452
rect 20076 6264 20128 6316
rect 25228 6400 25280 6452
rect 24676 6307 24728 6316
rect 24676 6273 24685 6307
rect 24685 6273 24719 6307
rect 24719 6273 24728 6307
rect 24676 6264 24728 6273
rect 27620 6400 27672 6452
rect 17316 6103 17368 6112
rect 17316 6069 17325 6103
rect 17325 6069 17359 6103
rect 17359 6069 17368 6103
rect 17316 6060 17368 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 17316 5856 17368 5908
rect 23480 5899 23532 5908
rect 23480 5865 23489 5899
rect 23489 5865 23523 5899
rect 23523 5865 23532 5899
rect 23480 5856 23532 5865
rect 18328 5720 18380 5772
rect 24676 5763 24728 5772
rect 24676 5729 24694 5763
rect 24694 5729 24728 5763
rect 24676 5720 24728 5729
rect 27620 5720 27672 5772
rect 24584 5584 24636 5636
rect 24216 5559 24268 5568
rect 24216 5525 24225 5559
rect 24225 5525 24259 5559
rect 24259 5525 24268 5559
rect 24216 5516 24268 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 24676 5355 24728 5364
rect 24676 5321 24685 5355
rect 24685 5321 24719 5355
rect 24719 5321 24728 5355
rect 24676 5312 24728 5321
rect 18328 5015 18380 5024
rect 18328 4981 18337 5015
rect 18337 4981 18371 5015
rect 18371 4981 18380 5015
rect 18328 4972 18380 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 24400 4700 24452 4752
rect 24584 4675 24636 4684
rect 24584 4641 24593 4675
rect 24593 4641 24627 4675
rect 24627 4641 24636 4675
rect 24584 4632 24636 4641
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 24676 4267 24728 4276
rect 24676 4233 24685 4267
rect 24685 4233 24719 4267
rect 24719 4233 24728 4267
rect 24676 4224 24728 4233
rect 27620 4224 27672 4276
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 24492 3612 24544 3664
rect 24584 3587 24636 3596
rect 24584 3553 24593 3587
rect 24593 3553 24627 3587
rect 24627 3553 24636 3587
rect 24584 3544 24636 3553
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 24676 3179 24728 3188
rect 24676 3145 24685 3179
rect 24685 3145 24719 3179
rect 24719 3145 24728 3179
rect 24676 3136 24728 3145
rect 27620 3136 27672 3188
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 11520 2592 11572 2644
rect 24216 2592 24268 2644
rect 25136 2456 25188 2508
rect 11888 2431 11940 2440
rect 11888 2397 11897 2431
rect 11897 2397 11931 2431
rect 11931 2397 11940 2431
rect 11888 2388 11940 2397
rect 25136 2295 25188 2304
rect 25136 2261 25145 2295
rect 25145 2261 25179 2295
rect 25179 2261 25188 2295
rect 25136 2252 25188 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 1768 76 1820 128
rect 9588 76 9640 128
rect 15752 76 15804 128
rect 16396 76 16448 128
<< metal2 >>
rect 478 27520 534 28000
rect 1490 27520 1546 28000
rect 2502 27520 2558 28000
rect 3514 27554 3570 28000
rect 4618 27554 4674 28000
rect 5630 27554 5686 28000
rect 3514 27526 3740 27554
rect 3514 27520 3570 27526
rect 492 23662 520 27520
rect 480 23656 532 23662
rect 480 23598 532 23604
rect 1504 20398 1532 27520
rect 1676 23520 1728 23526
rect 1676 23462 1728 23468
rect 1492 20392 1544 20398
rect 1492 20334 1544 20340
rect 1688 13814 1716 23462
rect 2516 23186 2544 27520
rect 3712 23866 3740 27526
rect 4618 27526 4844 27554
rect 4618 27520 4674 27526
rect 3700 23860 3752 23866
rect 3700 23802 3752 23808
rect 3712 23662 3740 23802
rect 3700 23656 3752 23662
rect 3700 23598 3752 23604
rect 2504 23180 2556 23186
rect 2504 23122 2556 23128
rect 4816 21690 4844 27526
rect 5552 27526 5686 27554
rect 5552 23866 5580 27526
rect 5630 27520 5686 27526
rect 6642 27520 6698 28000
rect 7654 27554 7710 28000
rect 8758 27554 8814 28000
rect 9770 27554 9826 28000
rect 7654 27526 7880 27554
rect 7654 27520 7710 27526
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6656 24274 6684 27520
rect 6644 24268 6696 24274
rect 6644 24210 6696 24216
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 6656 23866 6684 24210
rect 6828 24064 6880 24070
rect 6828 24006 6880 24012
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 6644 23860 6696 23866
rect 6644 23802 6696 23808
rect 5552 23662 5580 23802
rect 5540 23656 5592 23662
rect 5540 23598 5592 23604
rect 5356 23520 5408 23526
rect 5356 23462 5408 23468
rect 5368 23050 5396 23462
rect 5356 23044 5408 23050
rect 5356 22986 5408 22992
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 4816 21486 4844 21626
rect 4804 21480 4856 21486
rect 4804 21422 4856 21428
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 1596 13786 1716 13814
rect 1596 12646 1624 13786
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6840 9722 6868 24006
rect 7852 23866 7880 27526
rect 8758 27526 8984 27554
rect 8758 27520 8814 27526
rect 8956 23866 8984 27526
rect 9770 27526 9996 27554
rect 9770 27520 9826 27526
rect 9968 24954 9996 27526
rect 10782 27520 10838 28000
rect 11794 27520 11850 28000
rect 12898 27520 12954 28000
rect 13910 27554 13966 28000
rect 14922 27554 14978 28000
rect 13910 27526 14228 27554
rect 13910 27520 13966 27526
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 9956 24948 10008 24954
rect 9956 24890 10008 24896
rect 9968 24750 9996 24890
rect 9956 24744 10008 24750
rect 9956 24686 10008 24692
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10416 24268 10468 24274
rect 10416 24210 10468 24216
rect 10428 23866 10456 24210
rect 7840 23860 7892 23866
rect 7840 23802 7892 23808
rect 8944 23860 8996 23866
rect 8944 23802 8996 23808
rect 10416 23860 10468 23866
rect 10416 23802 10468 23808
rect 7852 23662 7880 23802
rect 8956 23662 8984 23802
rect 10796 23798 10824 27520
rect 11704 24608 11756 24614
rect 11704 24550 11756 24556
rect 11336 24268 11388 24274
rect 11336 24210 11388 24216
rect 10784 23792 10836 23798
rect 10784 23734 10836 23740
rect 7840 23656 7892 23662
rect 7840 23598 7892 23604
rect 8944 23656 8996 23662
rect 8944 23598 8996 23604
rect 11060 23656 11112 23662
rect 11060 23598 11112 23604
rect 7380 23520 7432 23526
rect 7656 23520 7708 23526
rect 7432 23480 7512 23508
rect 7380 23462 7432 23468
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 7392 19378 7420 20334
rect 7380 19372 7432 19378
rect 7380 19314 7432 19320
rect 7484 18358 7512 23480
rect 7656 23462 7708 23468
rect 8760 23520 8812 23526
rect 8760 23462 8812 23468
rect 9496 23520 9548 23526
rect 9496 23462 9548 23468
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 7472 18352 7524 18358
rect 7472 18294 7524 18300
rect 7668 13814 7696 23462
rect 8300 23180 8352 23186
rect 8300 23122 8352 23128
rect 8312 22778 8340 23122
rect 8300 22772 8352 22778
rect 8300 22714 8352 22720
rect 7576 13786 7696 13814
rect 8772 13814 8800 23462
rect 9220 22976 9272 22982
rect 9220 22918 9272 22924
rect 9232 22642 9260 22918
rect 9220 22636 9272 22642
rect 9220 22578 9272 22584
rect 9036 22432 9088 22438
rect 9036 22374 9088 22380
rect 9048 21486 9076 22374
rect 9232 22234 9260 22578
rect 9220 22228 9272 22234
rect 9220 22170 9272 22176
rect 9036 21480 9088 21486
rect 9036 21422 9088 21428
rect 9220 21480 9272 21486
rect 9508 21457 9536 23462
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10796 23254 10824 23462
rect 10600 23248 10652 23254
rect 10600 23190 10652 23196
rect 10784 23248 10836 23254
rect 10784 23190 10836 23196
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 10152 22778 10180 23054
rect 10612 22778 10640 23190
rect 11072 22982 11100 23598
rect 11348 23526 11376 24210
rect 11716 24206 11744 24550
rect 11808 24342 11836 27520
rect 12912 24954 12940 27520
rect 13912 25492 13964 25498
rect 13912 25434 13964 25440
rect 12900 24948 12952 24954
rect 12900 24890 12952 24896
rect 12912 24750 12940 24890
rect 12900 24744 12952 24750
rect 12900 24686 12952 24692
rect 13636 24608 13688 24614
rect 13636 24550 13688 24556
rect 11796 24336 11848 24342
rect 11796 24278 11848 24284
rect 12808 24268 12860 24274
rect 12808 24210 12860 24216
rect 13544 24268 13596 24274
rect 13544 24210 13596 24216
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 12624 23656 12676 23662
rect 12624 23598 12676 23604
rect 11336 23520 11388 23526
rect 11336 23462 11388 23468
rect 11348 23050 11376 23462
rect 12636 23322 12664 23598
rect 12624 23316 12676 23322
rect 12624 23258 12676 23264
rect 12256 23180 12308 23186
rect 12256 23122 12308 23128
rect 11336 23044 11388 23050
rect 11336 22986 11388 22992
rect 11060 22976 11112 22982
rect 11060 22918 11112 22924
rect 10140 22772 10192 22778
rect 10140 22714 10192 22720
rect 10600 22772 10652 22778
rect 10600 22714 10652 22720
rect 11072 22506 11100 22918
rect 11348 22710 11376 22986
rect 11336 22704 11388 22710
rect 11336 22646 11388 22652
rect 12268 22642 12296 23122
rect 12820 22778 12848 24210
rect 13452 24132 13504 24138
rect 13452 24074 13504 24080
rect 13464 23474 13492 24074
rect 13556 23866 13584 24210
rect 13544 23860 13596 23866
rect 13544 23802 13596 23808
rect 13464 23446 13584 23474
rect 13176 23248 13228 23254
rect 13176 23190 13228 23196
rect 12808 22772 12860 22778
rect 12808 22714 12860 22720
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 12256 22636 12308 22642
rect 12256 22578 12308 22584
rect 10784 22500 10836 22506
rect 10784 22442 10836 22448
rect 11060 22500 11112 22506
rect 11060 22442 11112 22448
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 9680 22160 9732 22166
rect 9680 22102 9732 22108
rect 9692 21690 9720 22102
rect 9956 22024 10008 22030
rect 9956 21966 10008 21972
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9220 21422 9272 21428
rect 9494 21448 9550 21457
rect 9128 21344 9180 21350
rect 9128 21286 9180 21292
rect 9140 20505 9168 21286
rect 9232 21146 9260 21422
rect 9494 21383 9550 21392
rect 9220 21140 9272 21146
rect 9220 21082 9272 21088
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 9126 20496 9182 20505
rect 9692 20466 9720 20878
rect 9968 20806 9996 21966
rect 10796 21962 10824 22442
rect 10784 21956 10836 21962
rect 10784 21898 10836 21904
rect 11072 21894 11100 22442
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 11072 21690 11100 21830
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 10232 21548 10284 21554
rect 10232 21490 10284 21496
rect 10244 21418 10272 21490
rect 10692 21480 10744 21486
rect 10692 21422 10744 21428
rect 10232 21412 10284 21418
rect 10152 21372 10232 21400
rect 10152 21078 10180 21372
rect 10232 21354 10284 21360
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10140 21072 10192 21078
rect 10140 21014 10192 21020
rect 9956 20800 10008 20806
rect 9956 20742 10008 20748
rect 9126 20431 9182 20440
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9692 20058 9720 20402
rect 9864 20392 9916 20398
rect 9864 20334 9916 20340
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 9784 19514 9812 19858
rect 9036 19508 9088 19514
rect 9036 19450 9088 19456
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8864 18290 8892 19110
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 8864 17882 8892 18226
rect 8944 18148 8996 18154
rect 8944 18090 8996 18096
rect 8956 17882 8984 18090
rect 8852 17876 8904 17882
rect 8852 17818 8904 17824
rect 8944 17876 8996 17882
rect 8944 17818 8996 17824
rect 9048 17134 9076 19450
rect 9496 18148 9548 18154
rect 9496 18090 9548 18096
rect 9508 17270 9536 18090
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9784 17814 9812 18022
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9496 17264 9548 17270
rect 9496 17206 9548 17212
rect 9692 17202 9720 17614
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 9220 17128 9272 17134
rect 9220 17070 9272 17076
rect 9048 15706 9076 17070
rect 9232 16726 9260 17070
rect 9692 16794 9720 17138
rect 9784 16998 9812 17750
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9220 16720 9272 16726
rect 9220 16662 9272 16668
rect 9232 16250 9260 16662
rect 9784 16522 9812 16934
rect 9876 16658 9904 20334
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9048 14958 9076 15642
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9036 14952 9088 14958
rect 9036 14894 9088 14900
rect 9048 14618 9076 14894
rect 9692 14890 9720 15506
rect 9784 15094 9812 16458
rect 9876 16250 9904 16594
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9876 16046 9904 16186
rect 9864 16040 9916 16046
rect 9864 15982 9916 15988
rect 9772 15088 9824 15094
rect 9772 15030 9824 15036
rect 9404 14884 9456 14890
rect 9404 14826 9456 14832
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 9416 14074 9444 14826
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 8772 13786 8892 13814
rect 7576 10713 7604 13786
rect 8864 13433 8892 13786
rect 8850 13424 8906 13433
rect 8850 13359 8906 13368
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 12306 9720 12582
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9692 11898 9720 12242
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 7562 10704 7618 10713
rect 7562 10639 7618 10648
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5172 8424 5224 8430
rect 5172 8366 5224 8372
rect 1766 128 1822 480
rect 1766 76 1768 128
rect 1820 76 1822 128
rect 1766 0 1822 76
rect 5184 82 5212 8366
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5262 82 5318 480
rect 5184 54 5318 82
rect 5262 0 5318 54
rect 8758 82 8814 480
rect 8956 82 8984 11698
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9600 134 9628 10406
rect 9968 5273 9996 20742
rect 10152 20602 10180 21014
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 10704 20398 10732 21422
rect 10140 20392 10192 20398
rect 10140 20334 10192 20340
rect 10692 20392 10744 20398
rect 10692 20334 10744 20340
rect 10152 19922 10180 20334
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10140 19916 10192 19922
rect 10140 19858 10192 19864
rect 10152 19174 10180 19858
rect 11336 19848 11388 19854
rect 11336 19790 11388 19796
rect 10876 19304 10928 19310
rect 10876 19246 10928 19252
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 10152 18222 10180 18566
rect 10888 18222 10916 19246
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 10876 18216 10928 18222
rect 10876 18158 10928 18164
rect 10152 16794 10180 18158
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 10428 17066 10456 17614
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 10416 17060 10468 17066
rect 10416 17002 10468 17008
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 10980 16454 11008 17138
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 10060 14958 10088 15302
rect 10152 15026 10180 15846
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10704 15366 10732 15982
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 10048 14952 10100 14958
rect 10048 14894 10100 14900
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10060 14074 10088 14758
rect 10152 14618 10180 14962
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 10796 14385 10824 14758
rect 10782 14376 10838 14385
rect 10782 14311 10838 14320
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10060 13814 10088 14010
rect 10060 13786 10180 13814
rect 10152 13734 10180 13786
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10704 12714 10732 13670
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 10692 12708 10744 12714
rect 10692 12650 10744 12656
rect 10060 12442 10088 12650
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10152 11218 10180 11494
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10152 10470 10180 11154
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10796 8430 10824 14311
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10888 12850 10916 13194
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 10888 11694 10916 12650
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 9954 5264 10010 5273
rect 9954 5199 10010 5208
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10980 4154 11008 16390
rect 11072 13802 11100 19110
rect 11256 18902 11284 19110
rect 11244 18896 11296 18902
rect 11244 18838 11296 18844
rect 11256 18426 11284 18838
rect 11348 18766 11376 19790
rect 11336 18760 11388 18766
rect 11336 18702 11388 18708
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 11348 18358 11376 18702
rect 11336 18352 11388 18358
rect 11336 18294 11388 18300
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11532 17338 11560 17682
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 11428 16584 11480 16590
rect 11428 16526 11480 16532
rect 11440 15638 11468 16526
rect 11532 16250 11560 16594
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11428 15632 11480 15638
rect 11428 15574 11480 15580
rect 11440 15162 11468 15574
rect 11428 15156 11480 15162
rect 11428 15098 11480 15104
rect 11532 15094 11560 16186
rect 11716 15434 11744 22578
rect 13188 22438 13216 23190
rect 13360 23112 13412 23118
rect 13360 23054 13412 23060
rect 13372 22778 13400 23054
rect 13360 22772 13412 22778
rect 13360 22714 13412 22720
rect 12256 22432 12308 22438
rect 12256 22374 12308 22380
rect 13176 22432 13228 22438
rect 13176 22374 13228 22380
rect 12268 18970 12296 22374
rect 13188 22098 13216 22374
rect 13176 22092 13228 22098
rect 13176 22034 13228 22040
rect 13188 21350 13216 22034
rect 13556 21622 13584 23446
rect 13648 22545 13676 24550
rect 13728 24064 13780 24070
rect 13728 24006 13780 24012
rect 13740 23662 13768 24006
rect 13924 23866 13952 25434
rect 14200 24274 14228 27526
rect 14844 27526 14978 27554
rect 14844 24954 14872 27526
rect 14922 27520 14978 27526
rect 15934 27520 15990 28000
rect 17038 27554 17094 28000
rect 17038 27526 17356 27554
rect 17038 27520 17094 27526
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14832 24948 14884 24954
rect 14832 24890 14884 24896
rect 14844 24750 14872 24890
rect 14832 24744 14884 24750
rect 14832 24686 14884 24692
rect 15568 24744 15620 24750
rect 15568 24686 15620 24692
rect 14740 24608 14792 24614
rect 14740 24550 14792 24556
rect 14188 24268 14240 24274
rect 14188 24210 14240 24216
rect 14200 23866 14228 24210
rect 13912 23860 13964 23866
rect 13912 23802 13964 23808
rect 14188 23860 14240 23866
rect 14188 23802 14240 23808
rect 14752 23730 14780 24550
rect 15292 24200 15344 24206
rect 15292 24142 15344 24148
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14740 23724 14792 23730
rect 14740 23666 14792 23672
rect 13728 23656 13780 23662
rect 13728 23598 13780 23604
rect 14752 23322 14780 23666
rect 15304 23594 15332 24142
rect 15476 23860 15528 23866
rect 15476 23802 15528 23808
rect 15292 23588 15344 23594
rect 15292 23530 15344 23536
rect 14740 23316 14792 23322
rect 14740 23258 14792 23264
rect 15488 23254 15516 23802
rect 15580 23730 15608 24686
rect 15752 24608 15804 24614
rect 15752 24550 15804 24556
rect 15568 23724 15620 23730
rect 15568 23666 15620 23672
rect 15476 23248 15528 23254
rect 15476 23190 15528 23196
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 15384 23112 15436 23118
rect 15384 23054 15436 23060
rect 14292 22642 14320 23054
rect 14372 22976 14424 22982
rect 14372 22918 14424 22924
rect 14384 22710 14412 22918
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15396 22778 15424 23054
rect 15384 22772 15436 22778
rect 15384 22714 15436 22720
rect 14372 22704 14424 22710
rect 14372 22646 14424 22652
rect 14740 22704 14792 22710
rect 14740 22646 14792 22652
rect 14280 22636 14332 22642
rect 14280 22578 14332 22584
rect 13634 22536 13690 22545
rect 13634 22471 13690 22480
rect 13820 22432 13872 22438
rect 13820 22374 13872 22380
rect 14372 22432 14424 22438
rect 14372 22374 14424 22380
rect 13832 22234 13860 22374
rect 13820 22228 13872 22234
rect 13820 22170 13872 22176
rect 14384 21690 14412 22374
rect 14372 21684 14424 21690
rect 14372 21626 14424 21632
rect 13544 21616 13596 21622
rect 13544 21558 13596 21564
rect 13912 21480 13964 21486
rect 13912 21422 13964 21428
rect 13360 21412 13412 21418
rect 13360 21354 13412 21360
rect 13176 21344 13228 21350
rect 13176 21286 13228 21292
rect 13188 21146 13216 21286
rect 13176 21140 13228 21146
rect 13176 21082 13228 21088
rect 13372 21078 13400 21354
rect 13924 21146 13952 21422
rect 14004 21412 14056 21418
rect 14004 21354 14056 21360
rect 13912 21140 13964 21146
rect 13912 21082 13964 21088
rect 13360 21072 13412 21078
rect 13360 21014 13412 21020
rect 12716 20936 12768 20942
rect 12716 20878 12768 20884
rect 12728 20058 12756 20878
rect 13924 20466 13952 21082
rect 14016 20534 14044 21354
rect 14004 20528 14056 20534
rect 14004 20470 14056 20476
rect 13912 20460 13964 20466
rect 13912 20402 13964 20408
rect 13084 20392 13136 20398
rect 13084 20334 13136 20340
rect 13820 20392 13872 20398
rect 13820 20334 13872 20340
rect 12716 20052 12768 20058
rect 12716 19994 12768 20000
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 12728 19514 12756 19858
rect 12348 19508 12400 19514
rect 12348 19450 12400 19456
rect 12716 19508 12768 19514
rect 12716 19450 12768 19456
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 12360 16250 12388 19450
rect 13096 19378 13124 20334
rect 13832 19922 13860 20334
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 12900 18896 12952 18902
rect 12900 18838 12952 18844
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12544 17270 12572 18566
rect 12912 18222 12940 18838
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12532 17264 12584 17270
rect 12532 17206 12584 17212
rect 12636 17134 12664 17478
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12360 16046 12388 16186
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12636 15910 12664 17070
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12728 16522 12756 16934
rect 13096 16658 13124 19314
rect 13832 19174 13860 19858
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 13004 15706 13032 15982
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 11704 15428 11756 15434
rect 11704 15370 11756 15376
rect 11612 15360 11664 15366
rect 11612 15302 11664 15308
rect 11520 15088 11572 15094
rect 11520 15030 11572 15036
rect 11532 14550 11560 15030
rect 11624 14550 11652 15302
rect 11520 14544 11572 14550
rect 11520 14486 11572 14492
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11060 13796 11112 13802
rect 11060 13738 11112 13744
rect 11348 13734 11376 14350
rect 11532 14074 11560 14486
rect 11716 14346 11744 15370
rect 11808 15162 11836 15438
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 11704 14340 11756 14346
rect 11704 14282 11756 14288
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11152 13456 11204 13462
rect 11152 13398 11204 13404
rect 11164 12646 11192 13398
rect 11348 13258 11376 13670
rect 11428 13320 11480 13326
rect 11480 13280 11560 13308
rect 11428 13262 11480 13268
rect 11336 13252 11388 13258
rect 11336 13194 11388 13200
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11164 12374 11192 12582
rect 11152 12368 11204 12374
rect 11152 12310 11204 12316
rect 11532 12102 11560 13280
rect 12268 12850 12296 14894
rect 12912 14890 12940 15302
rect 13096 14958 13124 15438
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 12900 14884 12952 14890
rect 12900 14826 12952 14832
rect 12912 14618 12940 14826
rect 12900 14612 12952 14618
rect 12900 14554 12952 14560
rect 13188 13814 13216 19110
rect 13924 18970 13952 19246
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13636 18080 13688 18086
rect 13636 18022 13688 18028
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13280 16794 13308 17478
rect 13648 17338 13676 18022
rect 14016 17814 14044 20470
rect 14280 20392 14332 20398
rect 14280 20334 14332 20340
rect 14292 20058 14320 20334
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14568 19378 14596 19790
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14004 17808 14056 17814
rect 14004 17750 14056 17756
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 13648 17134 13676 17274
rect 13636 17128 13688 17134
rect 13636 17070 13688 17076
rect 14016 16998 14044 17750
rect 14188 17128 14240 17134
rect 14188 17070 14240 17076
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 13464 16046 13492 16594
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13556 16250 13584 16526
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13464 15026 13492 15302
rect 13924 15162 13952 16662
rect 14200 16454 14228 17070
rect 14280 17060 14332 17066
rect 14280 17002 14332 17008
rect 14292 16454 14320 17002
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14188 16448 14240 16454
rect 14188 16390 14240 16396
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14200 16046 14228 16390
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 14004 15360 14056 15366
rect 14004 15302 14056 15308
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 14016 15094 14044 15302
rect 14004 15088 14056 15094
rect 14004 15030 14056 15036
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13268 14340 13320 14346
rect 13268 14282 13320 14288
rect 13280 13870 13308 14282
rect 13464 14278 13492 14962
rect 13832 14822 13860 14962
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13832 14414 13860 14758
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13464 14074 13492 14214
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13464 13920 13492 14010
rect 13728 14000 13780 14006
rect 13728 13942 13780 13948
rect 13372 13892 13492 13920
rect 13268 13864 13320 13870
rect 13096 13786 13216 13814
rect 13266 13832 13268 13841
rect 13320 13832 13322 13841
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12912 13530 12940 13670
rect 13096 13530 13124 13786
rect 13266 13767 13322 13776
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 12360 12442 12388 13126
rect 12452 12918 12480 13330
rect 12912 13258 12940 13466
rect 13372 13394 13400 13892
rect 13450 13832 13506 13841
rect 13450 13767 13506 13776
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12452 12714 12480 12854
rect 12440 12708 12492 12714
rect 12440 12650 12492 12656
rect 12912 12442 12940 13194
rect 13280 12986 13308 13194
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 12992 12708 13044 12714
rect 12992 12650 13044 12656
rect 13004 12442 13032 12650
rect 13464 12442 13492 13767
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13648 12442 13676 13330
rect 13740 13258 13768 13942
rect 13832 13938 13860 14350
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13832 13326 13860 13874
rect 14004 13456 14056 13462
rect 14004 13398 14056 13404
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13728 13252 13780 13258
rect 13728 13194 13780 13200
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13740 12442 13768 12650
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 11520 12096 11572 12102
rect 11520 12038 11572 12044
rect 10888 4126 11008 4154
rect 10888 4049 10916 4126
rect 10874 4040 10930 4049
rect 10874 3975 10930 3984
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 11532 2650 11560 12038
rect 12360 11558 12388 12242
rect 13004 11626 13032 12242
rect 13648 12170 13676 12378
rect 14016 12374 14044 13398
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 14200 12306 14228 12582
rect 14188 12300 14240 12306
rect 14188 12242 14240 12248
rect 14200 12209 14228 12242
rect 14186 12200 14242 12209
rect 13636 12164 13688 12170
rect 14186 12135 14242 12144
rect 13636 12106 13688 12112
rect 14200 11898 14228 12135
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 12440 11620 12492 11626
rect 12440 11562 12492 11568
rect 12992 11620 13044 11626
rect 12992 11562 13044 11568
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 12176 9722 12204 9998
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12360 9654 12388 11494
rect 12452 11218 12480 11562
rect 13004 11354 13032 11562
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 13556 10674 13584 11290
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13004 10266 13032 10610
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 13832 10198 13860 10406
rect 12900 10192 12952 10198
rect 12900 10134 12952 10140
rect 13820 10192 13872 10198
rect 13820 10134 13872 10140
rect 12912 9722 12940 10134
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 12900 9716 12952 9722
rect 12900 9658 12952 9664
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 11886 2544 11942 2553
rect 11886 2479 11942 2488
rect 11900 2446 11928 2479
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 8758 54 8984 82
rect 9588 128 9640 134
rect 9588 70 9640 76
rect 12254 82 12310 480
rect 12360 82 12388 9590
rect 12912 9042 12940 9658
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13556 9450 13584 9522
rect 13740 9450 13768 9930
rect 14108 9908 14136 11086
rect 14200 10810 14228 11154
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14188 9920 14240 9926
rect 14108 9880 14188 9908
rect 14188 9862 14240 9868
rect 13544 9444 13596 9450
rect 13544 9386 13596 9392
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13556 9178 13584 9386
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12912 8634 12940 8978
rect 14200 8634 14228 9862
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 14188 8628 14240 8634
rect 14188 8570 14240 8576
rect 14200 7478 14228 8570
rect 14292 7993 14320 16390
rect 14384 16250 14412 16934
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14648 15972 14700 15978
rect 14648 15914 14700 15920
rect 14660 15366 14688 15914
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14660 14890 14688 15302
rect 14648 14884 14700 14890
rect 14648 14826 14700 14832
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14568 14278 14596 14758
rect 14660 14346 14688 14826
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 14568 13734 14596 14214
rect 14660 14006 14688 14282
rect 14648 14000 14700 14006
rect 14648 13942 14700 13948
rect 14556 13728 14608 13734
rect 14556 13670 14608 13676
rect 14752 13530 14780 22646
rect 15384 22500 15436 22506
rect 15384 22442 15436 22448
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15396 21554 15424 22442
rect 15488 22438 15516 23190
rect 15580 23118 15608 23666
rect 15764 23474 15792 24550
rect 15948 24274 15976 27520
rect 17328 24954 17356 27526
rect 18050 27520 18106 28000
rect 19062 27520 19118 28000
rect 20074 27520 20130 28000
rect 20824 27526 21128 27554
rect 17316 24948 17368 24954
rect 17316 24890 17368 24896
rect 16212 24880 16264 24886
rect 16212 24822 16264 24828
rect 15844 24268 15896 24274
rect 15844 24210 15896 24216
rect 15936 24268 15988 24274
rect 15936 24210 15988 24216
rect 15856 23866 15884 24210
rect 15844 23860 15896 23866
rect 15844 23802 15896 23808
rect 15764 23446 15884 23474
rect 15568 23112 15620 23118
rect 15568 23054 15620 23060
rect 15856 22778 15884 23446
rect 15844 22772 15896 22778
rect 15844 22714 15896 22720
rect 15476 22432 15528 22438
rect 15476 22374 15528 22380
rect 15936 22092 15988 22098
rect 15936 22034 15988 22040
rect 15948 21690 15976 22034
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 15948 21350 15976 21626
rect 15936 21344 15988 21350
rect 15936 21286 15988 21292
rect 15948 21146 15976 21286
rect 15660 21140 15712 21146
rect 15660 21082 15712 21088
rect 15936 21140 15988 21146
rect 15936 21082 15988 21088
rect 15384 20936 15436 20942
rect 15384 20878 15436 20884
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 19514 15332 19858
rect 15396 19854 15424 20878
rect 15672 20534 15700 21082
rect 15660 20528 15712 20534
rect 15660 20470 15712 20476
rect 16028 20324 16080 20330
rect 16028 20266 16080 20272
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15488 19174 15516 19858
rect 16040 19718 16068 20266
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 15476 19168 15528 19174
rect 15476 19110 15528 19116
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14832 18148 14884 18154
rect 14832 18090 14884 18096
rect 14844 17882 14872 18090
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14844 17202 14872 17818
rect 15396 17746 15424 18022
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14832 17196 14884 17202
rect 14832 17138 14884 17144
rect 15396 16794 15424 17682
rect 15384 16788 15436 16794
rect 15384 16730 15436 16736
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 15910 15332 16594
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 15028 14618 15056 14962
rect 15304 14958 15332 15846
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 15016 14612 15068 14618
rect 15016 14554 15068 14560
rect 14844 14074 14872 14554
rect 15304 14414 15332 14894
rect 15396 14890 15424 15506
rect 15488 15162 15516 19110
rect 15752 18896 15804 18902
rect 15752 18838 15804 18844
rect 15764 18086 15792 18838
rect 15936 18692 15988 18698
rect 15936 18634 15988 18640
rect 15948 18290 15976 18634
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 15764 17882 15792 18022
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 15856 15978 15884 16934
rect 15844 15972 15896 15978
rect 15844 15914 15896 15920
rect 15568 15496 15620 15502
rect 15568 15438 15620 15444
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15580 15026 15608 15438
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 15384 14884 15436 14890
rect 15384 14826 15436 14832
rect 15396 14482 15424 14826
rect 15580 14618 15608 14962
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15292 14408 15344 14414
rect 15396 14385 15424 14418
rect 15292 14350 15344 14356
rect 15382 14376 15438 14385
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14384 12782 14412 13262
rect 14740 13252 14792 13258
rect 14740 13194 14792 13200
rect 14752 12986 14780 13194
rect 14844 13190 14872 13670
rect 15304 13394 15332 14350
rect 15382 14311 15438 14320
rect 15396 14074 15424 14311
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15580 14006 15608 14554
rect 15568 14000 15620 14006
rect 15568 13942 15620 13948
rect 15856 13870 15884 14962
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 14844 12918 14872 13126
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14832 12912 14884 12918
rect 14832 12854 14884 12860
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 14384 12646 14412 12718
rect 14740 12708 14792 12714
rect 14740 12650 14792 12656
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14752 12374 14780 12650
rect 14936 12646 14964 12786
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14832 12436 14884 12442
rect 14832 12378 14884 12384
rect 14740 12368 14792 12374
rect 14740 12310 14792 12316
rect 14844 12102 14872 12378
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14476 11354 14504 11698
rect 14844 11694 14872 12038
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14740 11620 14792 11626
rect 14740 11562 14792 11568
rect 14464 11348 14516 11354
rect 14516 11308 14596 11336
rect 14464 11290 14516 11296
rect 14568 9382 14596 11308
rect 14752 10674 14780 11562
rect 14844 11218 14872 11630
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14752 10266 14780 10610
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 15108 9444 15160 9450
rect 15108 9386 15160 9392
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14278 7984 14334 7993
rect 14278 7919 14334 7928
rect 14476 7857 14504 9318
rect 14568 8634 14596 9318
rect 15028 9110 15056 9386
rect 15120 9178 15148 9386
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 15016 9104 15068 9110
rect 15016 9046 15068 9052
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 15304 8430 15332 12650
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15396 11286 15424 12242
rect 15488 11762 15516 13126
rect 15580 12986 15608 13330
rect 15856 13190 15884 13806
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15672 12102 15700 12854
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15764 12238 15792 12786
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15672 11898 15700 12038
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15764 11830 15792 12174
rect 15752 11824 15804 11830
rect 15752 11766 15804 11772
rect 15856 11762 15884 13126
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 15384 11280 15436 11286
rect 15384 11222 15436 11228
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15488 10810 15516 11154
rect 15660 11076 15712 11082
rect 15660 11018 15712 11024
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15384 10260 15436 10266
rect 15488 10248 15516 10746
rect 15436 10220 15516 10248
rect 15384 10202 15436 10208
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15396 9722 15424 9998
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15396 9178 15424 9658
rect 15488 9450 15516 10220
rect 15580 10198 15608 10950
rect 15568 10192 15620 10198
rect 15568 10134 15620 10140
rect 15580 9722 15608 10134
rect 15672 10062 15700 11018
rect 15844 10532 15896 10538
rect 15844 10474 15896 10480
rect 15660 10056 15712 10062
rect 15660 9998 15712 10004
rect 15568 9716 15620 9722
rect 15568 9658 15620 9664
rect 15672 9586 15700 9998
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15304 8090 15332 8366
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 14462 7848 14518 7857
rect 14462 7783 14518 7792
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14188 7472 14240 7478
rect 14188 7414 14240 7420
rect 15304 7342 15332 8026
rect 15856 8022 15884 10474
rect 15936 8356 15988 8362
rect 15936 8298 15988 8304
rect 15844 8016 15896 8022
rect 15844 7958 15896 7964
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15764 7410 15792 7822
rect 15856 7546 15884 7958
rect 15948 7954 15976 8298
rect 15936 7948 15988 7954
rect 15936 7890 15988 7896
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15304 7002 15332 7278
rect 15764 7002 15792 7346
rect 15292 6996 15344 7002
rect 15292 6938 15344 6944
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 16040 6905 16068 19654
rect 16132 19514 16160 20198
rect 16120 19508 16172 19514
rect 16120 19450 16172 19456
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16132 18426 16160 18702
rect 16120 18420 16172 18426
rect 16120 18362 16172 18368
rect 16224 18306 16252 24822
rect 17328 24750 17356 24890
rect 17316 24744 17368 24750
rect 17316 24686 17368 24692
rect 17960 24676 18012 24682
rect 17960 24618 18012 24624
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 17408 24268 17460 24274
rect 17408 24210 17460 24216
rect 17038 23896 17094 23905
rect 17420 23866 17448 24210
rect 17880 23866 17908 24550
rect 17038 23831 17094 23840
rect 17408 23860 17460 23866
rect 17052 23798 17080 23831
rect 17408 23802 17460 23808
rect 17868 23860 17920 23866
rect 17868 23802 17920 23808
rect 17040 23792 17092 23798
rect 17040 23734 17092 23740
rect 17880 23662 17908 23802
rect 17040 23656 17092 23662
rect 17040 23598 17092 23604
rect 17868 23656 17920 23662
rect 17868 23598 17920 23604
rect 16488 22976 16540 22982
rect 16488 22918 16540 22924
rect 16500 22506 16528 22918
rect 16488 22500 16540 22506
rect 16488 22442 16540 22448
rect 16304 22432 16356 22438
rect 16304 22374 16356 22380
rect 16316 22166 16344 22374
rect 16304 22160 16356 22166
rect 16304 22102 16356 22108
rect 16488 21412 16540 21418
rect 16488 21354 16540 21360
rect 16500 21146 16528 21354
rect 16488 21140 16540 21146
rect 16488 21082 16540 21088
rect 16304 20596 16356 20602
rect 16304 20538 16356 20544
rect 16316 19310 16344 20538
rect 16500 20466 16528 21082
rect 16488 20460 16540 20466
rect 16488 20402 16540 20408
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 16316 18970 16344 19246
rect 16776 19174 16804 19790
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16304 18964 16356 18970
rect 16304 18906 16356 18912
rect 16132 18278 16252 18306
rect 16132 8072 16160 18278
rect 16488 16992 16540 16998
rect 16488 16934 16540 16940
rect 16500 16658 16528 16934
rect 16776 16794 16804 19110
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16960 17746 16988 18022
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 16868 16998 16896 17682
rect 16960 17202 16988 17682
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16960 16658 16988 17138
rect 16488 16652 16540 16658
rect 16488 16594 16540 16600
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 16500 15638 16528 16594
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16776 16046 16804 16390
rect 16960 16114 16988 16594
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16764 16040 16816 16046
rect 16764 15982 16816 15988
rect 16488 15632 16540 15638
rect 16540 15592 16712 15620
rect 16488 15574 16540 15580
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16500 14278 16528 14758
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16224 13734 16252 14010
rect 16500 14006 16528 14214
rect 16488 14000 16540 14006
rect 16488 13942 16540 13948
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16224 12646 16252 13670
rect 16408 13530 16436 13738
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16224 10742 16252 12582
rect 16212 10736 16264 10742
rect 16212 10678 16264 10684
rect 16224 10470 16252 10678
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16224 9654 16252 10406
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 16212 8084 16264 8090
rect 16132 8044 16212 8072
rect 16212 8026 16264 8032
rect 16224 7410 16252 8026
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 16026 6896 16082 6905
rect 16026 6831 16082 6840
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 16316 6225 16344 13466
rect 16408 12782 16436 13466
rect 16500 13258 16528 13942
rect 16684 13462 16712 15592
rect 16776 15162 16804 15982
rect 16960 15706 16988 16050
rect 16948 15700 17000 15706
rect 16948 15642 17000 15648
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16672 13456 16724 13462
rect 16672 13398 16724 13404
rect 16776 13326 16804 13874
rect 16856 13456 16908 13462
rect 16856 13398 16908 13404
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16488 13252 16540 13258
rect 16488 13194 16540 13200
rect 16500 12986 16528 13194
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16396 12776 16448 12782
rect 16396 12718 16448 12724
rect 16500 12442 16528 12922
rect 16776 12442 16804 13262
rect 16868 12442 16896 13398
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 16500 12306 16528 12378
rect 16488 12300 16540 12306
rect 16488 12242 16540 12248
rect 16500 12170 16528 12242
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16408 10674 16436 11494
rect 16500 11354 16528 12106
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 16408 9926 16436 10610
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16302 6216 16358 6225
rect 16302 6151 16358 6160
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 12254 54 12388 82
rect 15750 128 15806 480
rect 16408 134 16436 9862
rect 16868 7886 16896 12038
rect 16960 10810 16988 15506
rect 17052 11354 17080 23598
rect 17132 22976 17184 22982
rect 17132 22918 17184 22924
rect 17144 22506 17172 22918
rect 17972 22778 18000 24618
rect 18064 23730 18092 27520
rect 18144 24676 18196 24682
rect 18144 24618 18196 24624
rect 18156 24410 18184 24618
rect 19076 24410 19104 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 20088 25498 20116 27520
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 20352 24676 20404 24682
rect 20352 24618 20404 24624
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 18144 24404 18196 24410
rect 18144 24346 18196 24352
rect 19064 24404 19116 24410
rect 19064 24346 19116 24352
rect 18880 24336 18932 24342
rect 18880 24278 18932 24284
rect 18788 24200 18840 24206
rect 18788 24142 18840 24148
rect 18328 24132 18380 24138
rect 18328 24074 18380 24080
rect 18052 23724 18104 23730
rect 18052 23666 18104 23672
rect 18144 23656 18196 23662
rect 18144 23598 18196 23604
rect 17960 22772 18012 22778
rect 17960 22714 18012 22720
rect 17132 22500 17184 22506
rect 17132 22442 17184 22448
rect 17144 21554 17172 22442
rect 17500 22228 17552 22234
rect 17500 22170 17552 22176
rect 17132 21548 17184 21554
rect 17132 21490 17184 21496
rect 17512 21418 17540 22170
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 17500 21412 17552 21418
rect 17500 21354 17552 21360
rect 17696 21350 17724 21966
rect 17684 21344 17736 21350
rect 17684 21286 17736 21292
rect 17224 21072 17276 21078
rect 17224 21014 17276 21020
rect 17132 20936 17184 20942
rect 17132 20878 17184 20884
rect 17144 20534 17172 20878
rect 17236 20602 17264 21014
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 17132 20528 17184 20534
rect 17130 20496 17132 20505
rect 17184 20496 17186 20505
rect 17130 20431 17186 20440
rect 17144 20405 17172 20431
rect 17592 20392 17644 20398
rect 17592 20334 17644 20340
rect 17604 20058 17632 20334
rect 17592 20052 17644 20058
rect 17592 19994 17644 20000
rect 17604 19174 17632 19994
rect 17592 19168 17644 19174
rect 17592 19110 17644 19116
rect 17696 17338 17724 21286
rect 18156 20058 18184 23598
rect 18236 23180 18288 23186
rect 18236 23122 18288 23128
rect 18248 22506 18276 23122
rect 18236 22500 18288 22506
rect 18236 22442 18288 22448
rect 18248 22234 18276 22442
rect 18236 22228 18288 22234
rect 18236 22170 18288 22176
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17788 17814 17816 18702
rect 17972 18630 18000 19246
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17972 17882 18000 18566
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 17776 17808 17828 17814
rect 17776 17750 17828 17756
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 17684 17332 17736 17338
rect 17684 17274 17736 17280
rect 17132 17128 17184 17134
rect 17132 17070 17184 17076
rect 17144 16250 17172 17070
rect 17224 17060 17276 17066
rect 17224 17002 17276 17008
rect 17236 16658 17264 17002
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17132 16244 17184 16250
rect 17132 16186 17184 16192
rect 17236 15434 17264 16594
rect 17880 16046 17908 17682
rect 18156 17066 18184 19110
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18248 17134 18276 17478
rect 18340 17202 18368 24074
rect 18512 24064 18564 24070
rect 18512 24006 18564 24012
rect 18524 23118 18552 24006
rect 18800 23322 18828 24142
rect 18892 23866 18920 24278
rect 18972 24200 19024 24206
rect 18972 24142 19024 24148
rect 18880 23860 18932 23866
rect 18880 23802 18932 23808
rect 18984 23474 19012 24142
rect 19800 24064 19852 24070
rect 19800 24006 19852 24012
rect 19156 23860 19208 23866
rect 19156 23802 19208 23808
rect 18892 23446 19012 23474
rect 18788 23316 18840 23322
rect 18788 23258 18840 23264
rect 18512 23112 18564 23118
rect 18512 23054 18564 23060
rect 18788 22500 18840 22506
rect 18892 22488 18920 23446
rect 19168 23254 19196 23802
rect 19812 23730 19840 24006
rect 20364 23798 20392 24618
rect 20352 23792 20404 23798
rect 20352 23734 20404 23740
rect 19800 23724 19852 23730
rect 19800 23666 19852 23672
rect 20364 23474 20392 23734
rect 20364 23446 20484 23474
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19156 23248 19208 23254
rect 19156 23190 19208 23196
rect 19708 23180 19760 23186
rect 19708 23122 19760 23128
rect 19720 22778 19748 23122
rect 19708 22772 19760 22778
rect 19708 22714 19760 22720
rect 19432 22568 19484 22574
rect 19432 22510 19484 22516
rect 18840 22460 18920 22488
rect 19248 22500 19300 22506
rect 18788 22442 18840 22448
rect 19248 22442 19300 22448
rect 18696 20936 18748 20942
rect 18696 20878 18748 20884
rect 18708 20262 18736 20878
rect 18696 20256 18748 20262
rect 18696 20198 18748 20204
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 18144 17060 18196 17066
rect 18144 17002 18196 17008
rect 18708 16794 18736 20198
rect 18800 18748 18828 22442
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 18892 21622 18920 21966
rect 18880 21616 18932 21622
rect 18880 21558 18932 21564
rect 18972 18896 19024 18902
rect 18972 18838 19024 18844
rect 18880 18760 18932 18766
rect 18800 18720 18880 18748
rect 18880 18702 18932 18708
rect 18892 18426 18920 18702
rect 18880 18420 18932 18426
rect 18880 18362 18932 18368
rect 18984 18222 19012 18838
rect 19260 18698 19288 22442
rect 19444 22166 19472 22510
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19432 22160 19484 22166
rect 19432 22102 19484 22108
rect 19444 21690 19472 22102
rect 20088 21690 20116 22374
rect 20352 21956 20404 21962
rect 20352 21898 20404 21904
rect 19432 21684 19484 21690
rect 19432 21626 19484 21632
rect 20076 21684 20128 21690
rect 20076 21626 20128 21632
rect 19340 21412 19392 21418
rect 19340 21354 19392 21360
rect 19352 21078 19380 21354
rect 19444 21146 19472 21626
rect 20088 21400 20116 21626
rect 20364 21554 20392 21898
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20168 21412 20220 21418
rect 20088 21372 20168 21400
rect 20168 21354 20220 21360
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19432 21140 19484 21146
rect 19432 21082 19484 21088
rect 19340 21072 19392 21078
rect 19340 21014 19392 21020
rect 19352 20534 19380 21014
rect 19984 20800 20036 20806
rect 19984 20742 20036 20748
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 19996 20466 20024 20742
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19536 20058 19564 20198
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19524 20052 19576 20058
rect 19524 19994 19576 20000
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19352 19514 19380 19858
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19996 19242 20024 19450
rect 20456 19446 20484 23446
rect 20824 23322 20852 27526
rect 21100 27418 21128 27526
rect 21178 27520 21234 28000
rect 22190 27520 22246 28000
rect 23202 27520 23258 28000
rect 24214 27554 24270 28000
rect 24044 27526 24270 27554
rect 21192 27418 21220 27520
rect 21100 27390 21220 27418
rect 22008 24608 22060 24614
rect 22008 24550 22060 24556
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20916 23866 20944 24210
rect 20904 23860 20956 23866
rect 20904 23802 20956 23808
rect 20812 23316 20864 23322
rect 20812 23258 20864 23264
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20824 22506 20852 23122
rect 20916 23050 20944 23802
rect 21364 23724 21416 23730
rect 21364 23666 21416 23672
rect 21272 23656 21324 23662
rect 21272 23598 21324 23604
rect 21284 23322 21312 23598
rect 21376 23322 21404 23666
rect 21272 23316 21324 23322
rect 21272 23258 21324 23264
rect 21364 23316 21416 23322
rect 21364 23258 21416 23264
rect 22020 23254 22048 24550
rect 22204 24410 22232 27520
rect 22192 24404 22244 24410
rect 22192 24346 22244 24352
rect 23216 23866 23244 27520
rect 23848 25152 23900 25158
rect 23848 25094 23900 25100
rect 23664 24268 23716 24274
rect 23664 24210 23716 24216
rect 23204 23860 23256 23866
rect 23204 23802 23256 23808
rect 22192 23656 22244 23662
rect 22192 23598 22244 23604
rect 22204 23254 22232 23598
rect 23676 23594 23704 24210
rect 23664 23588 23716 23594
rect 23664 23530 23716 23536
rect 22008 23248 22060 23254
rect 22008 23190 22060 23196
rect 22192 23248 22244 23254
rect 22192 23190 22244 23196
rect 20904 23044 20956 23050
rect 20904 22986 20956 22992
rect 21454 22536 21510 22545
rect 20812 22500 20864 22506
rect 21454 22471 21510 22480
rect 20812 22442 20864 22448
rect 21468 22438 21496 22471
rect 21456 22432 21508 22438
rect 21456 22374 21508 22380
rect 20536 22024 20588 22030
rect 20536 21966 20588 21972
rect 20548 21554 20576 21966
rect 22204 21894 22232 23190
rect 22468 23112 22520 23118
rect 22468 23054 22520 23060
rect 22480 22234 22508 23054
rect 23572 22704 23624 22710
rect 23572 22646 23624 22652
rect 22744 22432 22796 22438
rect 22744 22374 22796 22380
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 22468 22228 22520 22234
rect 22468 22170 22520 22176
rect 22756 22098 22784 22374
rect 23400 22166 23428 22374
rect 23388 22160 23440 22166
rect 23388 22102 23440 22108
rect 22744 22092 22796 22098
rect 22744 22034 22796 22040
rect 21824 21888 21876 21894
rect 21824 21830 21876 21836
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 20536 21548 20588 21554
rect 20588 21508 20668 21536
rect 20536 21490 20588 21496
rect 20536 20324 20588 20330
rect 20536 20266 20588 20272
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 19984 19236 20036 19242
rect 19984 19178 20036 19184
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 20456 18970 20484 19382
rect 20548 19378 20576 20266
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20444 18964 20496 18970
rect 20444 18906 20496 18912
rect 19248 18692 19300 18698
rect 19248 18634 19300 18640
rect 19432 18692 19484 18698
rect 19432 18634 19484 18640
rect 18972 18216 19024 18222
rect 18972 18158 19024 18164
rect 18788 17808 18840 17814
rect 18788 17750 18840 17756
rect 18800 17270 18828 17750
rect 18984 17338 19012 18158
rect 19156 18148 19208 18154
rect 19156 18090 19208 18096
rect 19444 18136 19472 18634
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 19524 18148 19576 18154
rect 19444 18108 19524 18136
rect 19168 17814 19196 18090
rect 19156 17808 19208 17814
rect 19156 17750 19208 17756
rect 19168 17338 19196 17750
rect 19444 17678 19472 18108
rect 19524 18090 19576 18096
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 20364 17338 20392 18158
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 19156 17332 19208 17338
rect 20352 17332 20404 17338
rect 19156 17274 19208 17280
rect 20272 17292 20352 17320
rect 18788 17264 18840 17270
rect 18788 17206 18840 17212
rect 19156 17060 19208 17066
rect 19156 17002 19208 17008
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18696 16652 18748 16658
rect 18696 16594 18748 16600
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17972 15978 18000 16390
rect 18708 16182 18736 16594
rect 18696 16176 18748 16182
rect 18696 16118 18748 16124
rect 17960 15972 18012 15978
rect 17960 15914 18012 15920
rect 18880 15972 18932 15978
rect 18880 15914 18932 15920
rect 17224 15428 17276 15434
rect 17224 15370 17276 15376
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17420 14074 17448 14214
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17132 14000 17184 14006
rect 17132 13942 17184 13948
rect 17144 12850 17172 13942
rect 17788 13530 17816 14758
rect 17868 14340 17920 14346
rect 17868 14282 17920 14288
rect 17880 13734 17908 14282
rect 17972 13870 18000 15914
rect 18892 15502 18920 15914
rect 19168 15706 19196 17002
rect 19984 16992 20036 16998
rect 19984 16934 20036 16940
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19432 16040 19484 16046
rect 19432 15982 19484 15988
rect 19156 15700 19208 15706
rect 19156 15642 19208 15648
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 18328 15360 18380 15366
rect 18328 15302 18380 15308
rect 18064 15162 18092 15302
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 18064 14278 18092 15098
rect 18340 14958 18368 15302
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 18064 14074 18092 14214
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 18340 13938 18368 14894
rect 18432 13938 18460 14962
rect 18892 14618 18920 15438
rect 19168 15094 19196 15642
rect 19444 15366 19472 15982
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19996 15706 20024 16934
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 20088 16114 20116 16730
rect 20272 16182 20300 17292
rect 20352 17274 20404 17280
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 20260 16176 20312 16182
rect 20260 16118 20312 16124
rect 20076 16108 20128 16114
rect 20076 16050 20128 16056
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19156 15088 19208 15094
rect 19156 15030 19208 15036
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 19444 14464 19472 15302
rect 19812 15094 19840 15302
rect 19800 15088 19852 15094
rect 19800 15030 19852 15036
rect 19996 15026 20024 15642
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19536 14618 19564 14758
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19524 14476 19576 14482
rect 19444 14436 19524 14464
rect 19524 14418 19576 14424
rect 19536 14074 19564 14418
rect 20364 14414 20392 17138
rect 20640 16794 20668 21508
rect 21836 21486 21864 21830
rect 22204 21690 22232 21830
rect 22756 21690 22784 22034
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 22744 21684 22796 21690
rect 22744 21626 22796 21632
rect 21824 21480 21876 21486
rect 21824 21422 21876 21428
rect 22284 21480 22336 21486
rect 22284 21422 22336 21428
rect 21640 21344 21692 21350
rect 21640 21286 21692 21292
rect 21652 21078 21680 21286
rect 21640 21072 21692 21078
rect 21640 21014 21692 21020
rect 21652 20534 21680 21014
rect 21916 20936 21968 20942
rect 21916 20878 21968 20884
rect 21640 20528 21692 20534
rect 21640 20470 21692 20476
rect 21652 20262 21680 20470
rect 21928 20262 21956 20878
rect 21640 20256 21692 20262
rect 21640 20198 21692 20204
rect 21916 20256 21968 20262
rect 21916 20198 21968 20204
rect 21652 19990 21680 20198
rect 21640 19984 21692 19990
rect 21640 19926 21692 19932
rect 21548 19848 21600 19854
rect 21548 19790 21600 19796
rect 20812 19712 20864 19718
rect 20812 19654 20864 19660
rect 20824 19242 20852 19654
rect 20996 19372 21048 19378
rect 20996 19314 21048 19320
rect 20812 19236 20864 19242
rect 20812 19178 20864 19184
rect 20824 17814 20852 19178
rect 21008 18834 21036 19314
rect 21272 19304 21324 19310
rect 21272 19246 21324 19252
rect 20996 18828 21048 18834
rect 20996 18770 21048 18776
rect 21088 18216 21140 18222
rect 21088 18158 21140 18164
rect 20812 17808 20864 17814
rect 20812 17750 20864 17756
rect 20628 16788 20680 16794
rect 20628 16730 20680 16736
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20548 15094 20576 16050
rect 20824 15162 20852 17750
rect 21100 17610 21128 18158
rect 21088 17604 21140 17610
rect 21088 17546 21140 17552
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 20904 15972 20956 15978
rect 20904 15914 20956 15920
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 20536 15088 20588 15094
rect 20536 15030 20588 15036
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20364 14074 20392 14350
rect 19524 14068 19576 14074
rect 19524 14010 19576 14016
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20916 13938 20944 15914
rect 21192 15570 21220 16934
rect 21284 16726 21312 19246
rect 21560 18630 21588 19790
rect 21548 18624 21600 18630
rect 21548 18566 21600 18572
rect 21364 17604 21416 17610
rect 21364 17546 21416 17552
rect 21272 16720 21324 16726
rect 21272 16662 21324 16668
rect 21284 16250 21312 16662
rect 21376 16658 21404 17546
rect 21560 17202 21588 18566
rect 21928 18290 21956 20198
rect 22008 19372 22060 19378
rect 22008 19314 22060 19320
rect 21916 18284 21968 18290
rect 21916 18226 21968 18232
rect 22020 17882 22048 19314
rect 22100 19236 22152 19242
rect 22100 19178 22152 19184
rect 22112 18834 22140 19178
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 22112 18426 22140 18770
rect 22100 18420 22152 18426
rect 22100 18362 22152 18368
rect 22296 18290 22324 21422
rect 22756 21146 22784 21626
rect 23480 21480 23532 21486
rect 23386 21448 23442 21457
rect 23480 21422 23532 21428
rect 23386 21383 23442 21392
rect 22744 21140 22796 21146
rect 22744 21082 22796 21088
rect 23400 20942 23428 21383
rect 23492 21078 23520 21422
rect 23480 21072 23532 21078
rect 23480 21014 23532 21020
rect 23388 20936 23440 20942
rect 23308 20896 23388 20924
rect 22744 20596 22796 20602
rect 22744 20538 22796 20544
rect 22756 20058 22784 20538
rect 23112 20256 23164 20262
rect 23112 20198 23164 20204
rect 22744 20052 22796 20058
rect 22744 19994 22796 20000
rect 22376 19984 22428 19990
rect 22376 19926 22428 19932
rect 22388 19174 22416 19926
rect 23020 19508 23072 19514
rect 23020 19450 23072 19456
rect 22376 19168 22428 19174
rect 22376 19110 22428 19116
rect 22468 19168 22520 19174
rect 22468 19110 22520 19116
rect 22388 18970 22416 19110
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22284 18284 22336 18290
rect 22284 18226 22336 18232
rect 22284 18080 22336 18086
rect 22388 18068 22416 18906
rect 22336 18040 22416 18068
rect 22284 18022 22336 18028
rect 22008 17876 22060 17882
rect 22008 17818 22060 17824
rect 22296 17814 22324 18022
rect 22284 17808 22336 17814
rect 22284 17750 22336 17756
rect 22100 17672 22152 17678
rect 22100 17614 22152 17620
rect 21824 17536 21876 17542
rect 21824 17478 21876 17484
rect 21548 17196 21600 17202
rect 21548 17138 21600 17144
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 21284 15638 21312 16186
rect 21376 15978 21404 16594
rect 21836 16250 21864 17478
rect 22112 16726 22140 17614
rect 22296 16998 22324 17750
rect 22284 16992 22336 16998
rect 22284 16934 22336 16940
rect 22100 16720 22152 16726
rect 22100 16662 22152 16668
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 21364 15972 21416 15978
rect 21364 15914 21416 15920
rect 22100 15700 22152 15706
rect 22100 15642 22152 15648
rect 21272 15632 21324 15638
rect 21272 15574 21324 15580
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21192 14822 21220 15506
rect 21284 15162 21312 15574
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 22112 15026 22140 15642
rect 22296 15638 22324 16934
rect 22480 15706 22508 19110
rect 23032 18970 23060 19450
rect 23020 18964 23072 18970
rect 23020 18906 23072 18912
rect 23124 18834 23152 20198
rect 23308 20058 23336 20896
rect 23388 20878 23440 20884
rect 23492 20602 23520 21014
rect 23480 20596 23532 20602
rect 23480 20538 23532 20544
rect 23388 20392 23440 20398
rect 23388 20334 23440 20340
rect 23296 20052 23348 20058
rect 23296 19994 23348 20000
rect 23400 18970 23428 20334
rect 23388 18964 23440 18970
rect 23388 18906 23440 18912
rect 23112 18828 23164 18834
rect 23112 18770 23164 18776
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 23400 17746 23428 18022
rect 23388 17740 23440 17746
rect 23388 17682 23440 17688
rect 22744 17128 22796 17134
rect 22744 17070 22796 17076
rect 22756 16794 22784 17070
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 22284 15632 22336 15638
rect 22284 15574 22336 15580
rect 22296 15366 22324 15574
rect 22468 15496 22520 15502
rect 22468 15438 22520 15444
rect 22284 15360 22336 15366
rect 22284 15302 22336 15308
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 22296 14822 22324 15302
rect 22376 15020 22428 15026
rect 22376 14962 22428 14968
rect 21180 14816 21232 14822
rect 21180 14758 21232 14764
rect 21916 14816 21968 14822
rect 21916 14758 21968 14764
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 21192 14550 21220 14758
rect 21180 14544 21232 14550
rect 21180 14486 21232 14492
rect 21824 14544 21876 14550
rect 21824 14486 21876 14492
rect 18328 13932 18380 13938
rect 18328 13874 18380 13880
rect 18420 13932 18472 13938
rect 20904 13932 20956 13938
rect 18472 13892 18552 13920
rect 18420 13874 18472 13880
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 17500 13252 17552 13258
rect 17500 13194 17552 13200
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 17420 12646 17448 13126
rect 17512 12918 17540 13194
rect 17684 13184 17736 13190
rect 17684 13126 17736 13132
rect 17500 12912 17552 12918
rect 17500 12854 17552 12860
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17420 12209 17448 12582
rect 17406 12200 17462 12209
rect 17512 12170 17540 12854
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17604 12238 17632 12582
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17406 12135 17462 12144
rect 17500 12164 17552 12170
rect 17420 11880 17448 12135
rect 17500 12106 17552 12112
rect 17328 11852 17448 11880
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 17144 10538 17172 11154
rect 17132 10532 17184 10538
rect 17132 10474 17184 10480
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17236 9382 17264 10066
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17236 9042 17264 9318
rect 17328 9178 17356 11852
rect 17604 11694 17632 12174
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17420 10606 17448 11086
rect 17408 10600 17460 10606
rect 17408 10542 17460 10548
rect 17420 10470 17448 10542
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17420 9042 17448 10406
rect 17696 10266 17724 13126
rect 17776 12368 17828 12374
rect 17880 12356 17908 13670
rect 18524 13530 18552 13892
rect 20904 13874 20956 13880
rect 21836 13870 21864 14486
rect 21928 14074 21956 14758
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 19064 13864 19116 13870
rect 19064 13806 19116 13812
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 21824 13864 21876 13870
rect 21824 13806 21876 13812
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18064 12782 18092 13466
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18616 12986 18644 13126
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 18616 12442 18644 12922
rect 18604 12436 18656 12442
rect 18604 12378 18656 12384
rect 17828 12328 17908 12356
rect 17776 12310 17828 12316
rect 17788 11898 17816 12310
rect 18892 12102 18920 12922
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18892 11898 18920 12038
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 18880 11892 18932 11898
rect 18880 11834 18932 11840
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17788 10198 17816 10406
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 17776 10192 17828 10198
rect 17776 10134 17828 10140
rect 18340 9722 18368 10202
rect 18708 10130 18736 11494
rect 19076 11014 19104 13806
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19260 12850 19288 13330
rect 19248 12844 19300 12850
rect 19168 12804 19248 12832
rect 19168 11286 19196 12804
rect 19248 12786 19300 12792
rect 19352 12782 19380 13806
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19524 13388 19576 13394
rect 19524 13330 19576 13336
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 19536 12714 19564 13330
rect 19996 12986 20024 13670
rect 21836 13530 21864 13806
rect 21272 13524 21324 13530
rect 21272 13466 21324 13472
rect 21824 13524 21876 13530
rect 21824 13466 21876 13472
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 20996 12776 21048 12782
rect 20996 12718 21048 12724
rect 19524 12708 19576 12714
rect 19524 12650 19576 12656
rect 19536 12306 19564 12650
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 21008 12374 21036 12718
rect 21100 12442 21128 13262
rect 21284 12714 21312 13466
rect 22296 13462 22324 14758
rect 22388 14550 22416 14962
rect 22480 14618 22508 15438
rect 22468 14612 22520 14618
rect 22468 14554 22520 14560
rect 22376 14544 22428 14550
rect 22376 14486 22428 14492
rect 22388 13462 22416 14486
rect 22572 14006 22600 15846
rect 22560 14000 22612 14006
rect 22560 13942 22612 13948
rect 22756 13938 22784 16730
rect 23388 16652 23440 16658
rect 23388 16594 23440 16600
rect 23400 16250 23428 16594
rect 23388 16244 23440 16250
rect 23388 16186 23440 16192
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 23400 15162 23428 15642
rect 23388 15156 23440 15162
rect 23388 15098 23440 15104
rect 22928 14476 22980 14482
rect 22928 14418 22980 14424
rect 22940 14074 22968 14418
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 23308 14074 23336 14214
rect 22928 14068 22980 14074
rect 22928 14010 22980 14016
rect 23296 14068 23348 14074
rect 23296 14010 23348 14016
rect 22744 13932 22796 13938
rect 22744 13874 22796 13880
rect 22756 13814 22784 13874
rect 22756 13786 22876 13814
rect 22284 13456 22336 13462
rect 22284 13398 22336 13404
rect 22376 13456 22428 13462
rect 22376 13398 22428 13404
rect 22388 12986 22416 13398
rect 22848 13326 22876 13786
rect 22940 13462 22968 14010
rect 23308 13734 23336 14010
rect 23296 13728 23348 13734
rect 23296 13670 23348 13676
rect 22928 13456 22980 13462
rect 22928 13398 22980 13404
rect 23110 13424 23166 13433
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22376 12980 22428 12986
rect 22376 12922 22428 12928
rect 22940 12850 22968 13398
rect 23110 13359 23166 13368
rect 23124 12986 23152 13359
rect 23112 12980 23164 12986
rect 23112 12922 23164 12928
rect 22928 12844 22980 12850
rect 22928 12786 22980 12792
rect 23124 12714 23152 12922
rect 21272 12708 21324 12714
rect 21272 12650 21324 12656
rect 23112 12708 23164 12714
rect 23112 12650 23164 12656
rect 21640 12640 21692 12646
rect 21640 12582 21692 12588
rect 21088 12436 21140 12442
rect 21088 12378 21140 12384
rect 21652 12374 21680 12582
rect 20996 12368 21048 12374
rect 20996 12310 21048 12316
rect 21640 12368 21692 12374
rect 21640 12310 21692 12316
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19524 12300 19576 12306
rect 19524 12242 19576 12248
rect 19260 11558 19288 12242
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 19536 11354 19564 12242
rect 20536 12164 20588 12170
rect 20536 12106 20588 12112
rect 20548 11694 20576 12106
rect 21364 11824 21416 11830
rect 21364 11766 21416 11772
rect 20536 11688 20588 11694
rect 20536 11630 20588 11636
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 20548 11354 20576 11630
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 19156 11280 19208 11286
rect 19156 11222 19208 11228
rect 19064 11008 19116 11014
rect 19064 10950 19116 10956
rect 19168 10674 19196 11222
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 19984 11076 20036 11082
rect 19984 11018 20036 11024
rect 19996 10810 20024 11018
rect 21284 10810 21312 11154
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 20350 10704 20406 10713
rect 19156 10668 19208 10674
rect 19208 10628 19288 10656
rect 20350 10639 20406 10648
rect 19156 10610 19208 10616
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 18892 10266 18920 10542
rect 19156 10532 19208 10538
rect 19156 10474 19208 10480
rect 19168 10266 19196 10474
rect 18880 10260 18932 10266
rect 18880 10202 18932 10208
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 18328 9716 18380 9722
rect 18328 9658 18380 9664
rect 18708 9450 18736 10066
rect 19168 9586 19196 10202
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 18696 9444 18748 9450
rect 18696 9386 18748 9392
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17224 9036 17276 9042
rect 17224 8978 17276 8984
rect 17408 9036 17460 9042
rect 17408 8978 17460 8984
rect 17236 8566 17264 8978
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 17420 8498 17448 8978
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17880 8090 17908 9318
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18156 8430 18184 8774
rect 18708 8430 18736 9386
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 18144 8424 18196 8430
rect 18144 8366 18196 8372
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18156 8090 18184 8366
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16684 7274 16712 7686
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16684 6866 16712 7210
rect 17420 7002 17448 7890
rect 17880 7546 17908 8026
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 18156 7256 18184 8026
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18248 7410 18276 7686
rect 18800 7546 18828 8298
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18236 7404 18288 7410
rect 18288 7364 18368 7392
rect 18236 7346 18288 7352
rect 18236 7268 18288 7274
rect 18156 7228 18236 7256
rect 18236 7210 18288 7216
rect 18248 7002 18276 7210
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 18236 6996 18288 7002
rect 18236 6938 18288 6944
rect 18340 6934 18368 7364
rect 18788 7268 18840 7274
rect 18788 7210 18840 7216
rect 17684 6928 17736 6934
rect 17684 6870 17736 6876
rect 18328 6928 18380 6934
rect 18328 6870 18380 6876
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16684 6458 16712 6802
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 17328 6118 17356 6734
rect 17696 6458 17724 6870
rect 18800 6866 18828 7210
rect 18788 6860 18840 6866
rect 18788 6802 18840 6808
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 17328 5914 17356 6054
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 18340 5030 18368 5714
rect 18328 5024 18380 5030
rect 18328 4966 18380 4972
rect 18340 2417 18368 4966
rect 18326 2408 18382 2417
rect 18326 2343 18382 2352
rect 15750 76 15752 128
rect 15804 76 15806 128
rect 8758 0 8814 54
rect 12254 0 12310 54
rect 15750 0 15806 76
rect 16396 128 16448 134
rect 16396 70 16448 76
rect 18984 82 19012 8434
rect 19260 7954 19288 10628
rect 20364 10538 20392 10639
rect 20352 10532 20404 10538
rect 20352 10474 20404 10480
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 20088 9382 20116 10406
rect 20364 10266 20392 10474
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 20364 9722 20392 9998
rect 20352 9716 20404 9722
rect 20352 9658 20404 9664
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 19352 9042 19380 9318
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 21272 9104 21324 9110
rect 21272 9046 21324 9052
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19352 8634 19380 8978
rect 21284 8634 21312 9046
rect 21376 8974 21404 11766
rect 21652 11558 21680 12310
rect 22100 12232 22152 12238
rect 22100 12174 22152 12180
rect 22112 11558 22140 12174
rect 22652 11688 22704 11694
rect 22652 11630 22704 11636
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 22100 11552 22152 11558
rect 22100 11494 22152 11500
rect 21548 11212 21600 11218
rect 21548 11154 21600 11160
rect 21560 10810 21588 11154
rect 21548 10804 21600 10810
rect 21548 10746 21600 10752
rect 21652 10674 21680 11494
rect 22112 11286 22140 11494
rect 22100 11280 22152 11286
rect 22100 11222 22152 11228
rect 21732 11144 21784 11150
rect 21732 11086 21784 11092
rect 21640 10668 21692 10674
rect 21640 10610 21692 10616
rect 21548 9444 21600 9450
rect 21652 9432 21680 10610
rect 21744 9654 21772 11086
rect 22008 11008 22060 11014
rect 22008 10950 22060 10956
rect 22020 10538 22048 10950
rect 22664 10674 22692 11630
rect 22744 11620 22796 11626
rect 22744 11562 22796 11568
rect 22756 11218 22784 11562
rect 22928 11280 22980 11286
rect 22928 11222 22980 11228
rect 22744 11212 22796 11218
rect 22744 11154 22796 11160
rect 22756 10810 22784 11154
rect 22744 10804 22796 10810
rect 22744 10746 22796 10752
rect 22940 10742 22968 11222
rect 22928 10736 22980 10742
rect 22928 10678 22980 10684
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 22008 10532 22060 10538
rect 22008 10474 22060 10480
rect 21916 10464 21968 10470
rect 21916 10406 21968 10412
rect 21928 9926 21956 10406
rect 21916 9920 21968 9926
rect 21916 9862 21968 9868
rect 21732 9648 21784 9654
rect 21732 9590 21784 9596
rect 21928 9518 21956 9862
rect 21916 9512 21968 9518
rect 21916 9454 21968 9460
rect 21600 9404 21680 9432
rect 21548 9386 21600 9392
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 21376 8634 21404 8910
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 20732 7954 20760 8366
rect 21560 8022 21588 9386
rect 22020 9110 22048 10474
rect 22664 10198 22692 10610
rect 22560 10192 22612 10198
rect 22560 10134 22612 10140
rect 22652 10192 22704 10198
rect 22652 10134 22704 10140
rect 22572 9382 22600 10134
rect 22744 10056 22796 10062
rect 22744 9998 22796 10004
rect 22756 9722 22784 9998
rect 22744 9716 22796 9722
rect 22744 9658 22796 9664
rect 23020 9512 23072 9518
rect 23020 9454 23072 9460
rect 22560 9376 22612 9382
rect 22560 9318 22612 9324
rect 22744 9376 22796 9382
rect 22744 9318 22796 9324
rect 22756 9110 22784 9318
rect 22008 9104 22060 9110
rect 22008 9046 22060 9052
rect 22744 9104 22796 9110
rect 22744 9046 22796 9052
rect 23032 9042 23060 9454
rect 23020 9036 23072 9042
rect 23020 8978 23072 8984
rect 23032 8566 23060 8978
rect 23492 8634 23520 18702
rect 23584 17678 23612 22646
rect 23572 17672 23624 17678
rect 23572 17614 23624 17620
rect 23572 16992 23624 16998
rect 23572 16934 23624 16940
rect 23584 16794 23612 16934
rect 23572 16788 23624 16794
rect 23572 16730 23624 16736
rect 23572 15972 23624 15978
rect 23572 15914 23624 15920
rect 23584 14482 23612 15914
rect 23572 14476 23624 14482
rect 23572 14418 23624 14424
rect 23676 11898 23704 23530
rect 23756 23248 23808 23254
rect 23756 23190 23808 23196
rect 23768 22234 23796 23190
rect 23860 22642 23888 25094
rect 24044 23905 24072 27526
rect 24214 27520 24270 27526
rect 25318 27520 25374 28000
rect 26330 27520 26386 28000
rect 27342 27520 27398 28000
rect 25134 25800 25190 25809
rect 25134 25735 25190 25744
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 25148 24954 25176 25735
rect 25136 24948 25188 24954
rect 25136 24890 25188 24896
rect 25148 24750 25176 24890
rect 25136 24744 25188 24750
rect 25136 24686 25188 24692
rect 25332 24410 25360 27520
rect 26146 26888 26202 26897
rect 26146 26823 26202 26832
rect 25504 25356 25556 25362
rect 25504 25298 25556 25304
rect 25516 24682 25544 25298
rect 25778 25120 25834 25129
rect 25778 25055 25834 25064
rect 25504 24676 25556 24682
rect 25504 24618 25556 24624
rect 25516 24585 25544 24618
rect 25502 24576 25558 24585
rect 25502 24511 25558 24520
rect 25320 24404 25372 24410
rect 25320 24346 25372 24352
rect 24860 24268 24912 24274
rect 24860 24210 24912 24216
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 24030 23896 24086 23905
rect 24030 23831 24086 23840
rect 23940 23520 23992 23526
rect 23940 23462 23992 23468
rect 23952 23254 23980 23462
rect 23940 23248 23992 23254
rect 23940 23190 23992 23196
rect 24032 23112 24084 23118
rect 24032 23054 24084 23060
rect 23940 23044 23992 23050
rect 23940 22986 23992 22992
rect 23848 22636 23900 22642
rect 23848 22578 23900 22584
rect 23952 22522 23980 22986
rect 23860 22494 23980 22522
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23768 19174 23796 20198
rect 23860 19854 23888 22494
rect 24044 22438 24072 23054
rect 24032 22432 24084 22438
rect 24032 22374 24084 22380
rect 24044 22234 24072 22374
rect 24032 22228 24084 22234
rect 24032 22170 24084 22176
rect 23940 20324 23992 20330
rect 23940 20266 23992 20272
rect 23952 19990 23980 20266
rect 23940 19984 23992 19990
rect 23940 19926 23992 19932
rect 24032 19984 24084 19990
rect 24032 19926 24084 19932
rect 23848 19848 23900 19854
rect 23848 19790 23900 19796
rect 23756 19168 23808 19174
rect 23756 19110 23808 19116
rect 23860 18902 23888 19790
rect 23952 19514 23980 19926
rect 23940 19508 23992 19514
rect 23940 19450 23992 19456
rect 24044 19446 24072 19926
rect 24032 19440 24084 19446
rect 24032 19382 24084 19388
rect 24044 19242 24072 19382
rect 24032 19236 24084 19242
rect 24032 19178 24084 19184
rect 23940 19168 23992 19174
rect 23940 19110 23992 19116
rect 23952 18970 23980 19110
rect 23940 18964 23992 18970
rect 23940 18906 23992 18912
rect 23848 18896 23900 18902
rect 23848 18838 23900 18844
rect 24032 18216 24084 18222
rect 24032 18158 24084 18164
rect 24044 18086 24072 18158
rect 24032 18080 24084 18086
rect 24032 18022 24084 18028
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 23768 16794 23796 17614
rect 24032 17604 24084 17610
rect 24032 17546 24084 17552
rect 24044 17202 24072 17546
rect 24032 17196 24084 17202
rect 24032 17138 24084 17144
rect 23756 16788 23808 16794
rect 23756 16730 23808 16736
rect 23940 16040 23992 16046
rect 23940 15982 23992 15988
rect 23952 15706 23980 15982
rect 24032 15904 24084 15910
rect 24032 15846 24084 15852
rect 23940 15700 23992 15706
rect 23940 15642 23992 15648
rect 24044 15162 24072 15846
rect 24032 15156 24084 15162
rect 24032 15098 24084 15104
rect 24044 14822 24072 15098
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 23756 13796 23808 13802
rect 23756 13738 23808 13744
rect 23768 13190 23796 13738
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23768 12850 23796 13126
rect 23756 12844 23808 12850
rect 23756 12786 23808 12792
rect 23664 11892 23716 11898
rect 23664 11834 23716 11840
rect 23940 11552 23992 11558
rect 23940 11494 23992 11500
rect 23952 10810 23980 11494
rect 23940 10804 23992 10810
rect 23940 10746 23992 10752
rect 24136 9178 24164 24006
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24872 23866 24900 24210
rect 24860 23860 24912 23866
rect 24860 23802 24912 23808
rect 25228 23656 25280 23662
rect 25228 23598 25280 23604
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24766 22672 24822 22681
rect 24766 22607 24822 22616
rect 24780 22098 24808 22607
rect 24768 22092 24820 22098
rect 24768 22034 24820 22040
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24780 21690 24808 22034
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24400 21412 24452 21418
rect 24400 21354 24452 21360
rect 24412 21078 24440 21354
rect 25044 21344 25096 21350
rect 25044 21286 25096 21292
rect 24400 21072 24452 21078
rect 24400 21014 24452 21020
rect 24952 21072 25004 21078
rect 24952 21014 25004 21020
rect 24860 20868 24912 20874
rect 24860 20810 24912 20816
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24216 19848 24268 19854
rect 24216 19790 24268 19796
rect 24228 19378 24256 19790
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24216 19372 24268 19378
rect 24216 19314 24268 19320
rect 24676 18828 24728 18834
rect 24676 18770 24728 18776
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24688 18426 24716 18770
rect 24676 18420 24728 18426
rect 24676 18362 24728 18368
rect 24768 17808 24820 17814
rect 24768 17750 24820 17756
rect 24676 17672 24728 17678
rect 24676 17614 24728 17620
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24688 17270 24716 17614
rect 24780 17270 24808 17750
rect 24676 17264 24728 17270
rect 24676 17206 24728 17212
rect 24768 17264 24820 17270
rect 24768 17206 24820 17212
rect 24780 16658 24808 17206
rect 24768 16652 24820 16658
rect 24768 16594 24820 16600
rect 24676 16584 24728 16590
rect 24676 16526 24728 16532
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24584 15972 24636 15978
rect 24584 15914 24636 15920
rect 24596 15502 24624 15914
rect 24584 15496 24636 15502
rect 24584 15438 24636 15444
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24688 15026 24716 16526
rect 24768 15496 24820 15502
rect 24768 15438 24820 15444
rect 24780 15026 24808 15438
rect 24872 15434 24900 20810
rect 24964 20602 24992 21014
rect 25056 20942 25084 21286
rect 25044 20936 25096 20942
rect 25044 20878 25096 20884
rect 24952 20596 25004 20602
rect 24952 20538 25004 20544
rect 25056 20058 25084 20878
rect 25044 20052 25096 20058
rect 25044 19994 25096 20000
rect 25136 19168 25188 19174
rect 25136 19110 25188 19116
rect 25044 18148 25096 18154
rect 25044 18090 25096 18096
rect 25056 17134 25084 18090
rect 25044 17128 25096 17134
rect 25044 17070 25096 17076
rect 24860 15428 24912 15434
rect 24860 15370 24912 15376
rect 24872 15162 24900 15370
rect 24860 15156 24912 15162
rect 24860 15098 24912 15104
rect 24308 15020 24360 15026
rect 24308 14962 24360 14968
rect 24676 15020 24728 15026
rect 24676 14962 24728 14968
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 24320 14618 24348 14962
rect 24766 14648 24822 14657
rect 24308 14612 24360 14618
rect 24766 14583 24822 14592
rect 24308 14554 24360 14560
rect 24676 14476 24728 14482
rect 24676 14418 24728 14424
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24688 14074 24716 14418
rect 24780 14346 24808 14583
rect 24768 14340 24820 14346
rect 24768 14282 24820 14288
rect 24676 14068 24728 14074
rect 24676 14010 24728 14016
rect 24676 13456 24728 13462
rect 24676 13398 24728 13404
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24216 12708 24268 12714
rect 24216 12650 24268 12656
rect 24584 12708 24636 12714
rect 24584 12650 24636 12656
rect 24228 12306 24256 12650
rect 24216 12300 24268 12306
rect 24216 12242 24268 12248
rect 24228 11898 24256 12242
rect 24596 12186 24624 12650
rect 24688 12646 24716 13398
rect 25148 13326 25176 19110
rect 25240 18766 25268 23598
rect 25792 22778 25820 25055
rect 26160 23186 26188 26823
rect 26344 23866 26372 27520
rect 27356 24274 27384 27520
rect 27344 24268 27396 24274
rect 27344 24210 27396 24216
rect 26332 23860 26384 23866
rect 26332 23802 26384 23808
rect 26148 23180 26200 23186
rect 26148 23122 26200 23128
rect 26160 22778 26188 23122
rect 25780 22772 25832 22778
rect 25780 22714 25832 22720
rect 26148 22772 26200 22778
rect 26148 22714 26200 22720
rect 25792 22574 25820 22714
rect 25780 22568 25832 22574
rect 25780 22510 25832 22516
rect 25778 21720 25834 21729
rect 25778 21655 25834 21664
rect 25792 21622 25820 21655
rect 25780 21616 25832 21622
rect 25780 21558 25832 21564
rect 25778 20632 25834 20641
rect 25778 20567 25834 20576
rect 25792 20534 25820 20567
rect 25780 20528 25832 20534
rect 25780 20470 25832 20476
rect 26054 19544 26110 19553
rect 26054 19479 26110 19488
rect 26068 19446 26096 19479
rect 26056 19440 26108 19446
rect 26056 19382 26108 19388
rect 27618 19136 27674 19145
rect 27618 19071 27674 19080
rect 27632 18970 27660 19071
rect 27620 18964 27672 18970
rect 27620 18906 27672 18912
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 25228 18624 25280 18630
rect 25228 18566 25280 18572
rect 25240 18222 25268 18566
rect 27620 18352 27672 18358
rect 27620 18294 27672 18300
rect 25228 18216 25280 18222
rect 25228 18158 25280 18164
rect 25410 17504 25466 17513
rect 25410 17439 25466 17448
rect 25424 17338 25452 17439
rect 25228 17332 25280 17338
rect 25228 17274 25280 17280
rect 25412 17332 25464 17338
rect 25412 17274 25464 17280
rect 25136 13320 25188 13326
rect 25136 13262 25188 13268
rect 24860 13252 24912 13258
rect 24860 13194 24912 13200
rect 24872 12714 24900 13194
rect 25148 12986 25176 13262
rect 25136 12980 25188 12986
rect 25136 12922 25188 12928
rect 24860 12708 24912 12714
rect 24860 12650 24912 12656
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24688 12374 24716 12582
rect 24676 12368 24728 12374
rect 24676 12310 24728 12316
rect 25240 12306 25268 17274
rect 27632 17105 27660 18294
rect 27618 17096 27674 17105
rect 27618 17031 27674 17040
rect 27620 16176 27672 16182
rect 27620 16118 27672 16124
rect 27632 16017 27660 16118
rect 27618 16008 27674 16017
rect 27618 15943 27674 15952
rect 25410 14240 25466 14249
rect 25410 14175 25466 14184
rect 25424 14074 25452 14175
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 25410 12472 25466 12481
rect 25410 12407 25466 12416
rect 25228 12300 25280 12306
rect 25228 12242 25280 12248
rect 24596 12158 24716 12186
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24216 11892 24268 11898
rect 24216 11834 24268 11840
rect 24216 11348 24268 11354
rect 24216 11290 24268 11296
rect 24228 10130 24256 11290
rect 24688 11150 24716 12158
rect 25240 11898 25268 12242
rect 25424 12170 25452 12407
rect 25412 12164 25464 12170
rect 25412 12106 25464 12112
rect 25228 11892 25280 11898
rect 25228 11834 25280 11840
rect 25228 11552 25280 11558
rect 25228 11494 25280 11500
rect 24950 11248 25006 11257
rect 24950 11183 25006 11192
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24688 10810 24716 11086
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 24400 10464 24452 10470
rect 24400 10406 24452 10412
rect 24412 10266 24440 10406
rect 24766 10296 24822 10305
rect 24400 10260 24452 10266
rect 24766 10231 24822 10240
rect 24400 10202 24452 10208
rect 24216 10124 24268 10130
rect 24216 10066 24268 10072
rect 24228 9722 24256 10066
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24216 9716 24268 9722
rect 24216 9658 24268 9664
rect 24780 9178 24808 10231
rect 24964 9722 24992 11183
rect 25136 11076 25188 11082
rect 25136 11018 25188 11024
rect 25148 10742 25176 11018
rect 25136 10736 25188 10742
rect 25136 10678 25188 10684
rect 25240 10169 25268 11494
rect 25226 10160 25282 10169
rect 25226 10095 25282 10104
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 24124 9172 24176 9178
rect 24124 9114 24176 9120
rect 24768 9172 24820 9178
rect 24768 9114 24820 9120
rect 23480 8628 23532 8634
rect 23480 8570 23532 8576
rect 22468 8560 22520 8566
rect 22468 8502 22520 8508
rect 23020 8560 23072 8566
rect 23020 8502 23072 8508
rect 23112 8560 23164 8566
rect 23112 8502 23164 8508
rect 21732 8356 21784 8362
rect 21732 8298 21784 8304
rect 21548 8016 21600 8022
rect 21548 7958 21600 7964
rect 19248 7948 19300 7954
rect 19248 7890 19300 7896
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 19260 7478 19288 7890
rect 19524 7880 19576 7886
rect 19524 7822 19576 7828
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 19248 7472 19300 7478
rect 19248 7414 19300 7420
rect 19536 6934 19564 7822
rect 21192 7546 21220 7822
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 19812 7274 19840 7482
rect 21560 7478 21588 7958
rect 21744 7886 21772 8298
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21548 7472 21600 7478
rect 21548 7414 21600 7420
rect 21560 7274 21588 7414
rect 19800 7268 19852 7274
rect 19800 7210 19852 7216
rect 21548 7268 21600 7274
rect 21548 7210 21600 7216
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19524 6928 19576 6934
rect 19524 6870 19576 6876
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19260 6458 19288 6802
rect 20088 6662 20116 7142
rect 21560 6798 21588 7210
rect 21744 6934 21772 7822
rect 21732 6928 21784 6934
rect 21732 6870 21784 6876
rect 21548 6792 21600 6798
rect 21548 6734 21600 6740
rect 20076 6656 20128 6662
rect 20076 6598 20128 6604
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 20088 6322 20116 6598
rect 20076 6316 20128 6322
rect 20076 6258 20128 6264
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19246 82 19302 480
rect 18984 54 19302 82
rect 22480 82 22508 8502
rect 22652 7744 22704 7750
rect 22652 7686 22704 7692
rect 22664 7256 22692 7686
rect 23124 7546 23152 8502
rect 24136 8498 24164 9114
rect 25044 9036 25096 9042
rect 25044 8978 25096 8984
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24216 8560 24268 8566
rect 24216 8502 24268 8508
rect 24124 8492 24176 8498
rect 24124 8434 24176 8440
rect 24228 8362 24256 8502
rect 24308 8492 24360 8498
rect 24308 8434 24360 8440
rect 24216 8356 24268 8362
rect 24216 8298 24268 8304
rect 23940 8016 23992 8022
rect 23940 7958 23992 7964
rect 23112 7540 23164 7546
rect 23112 7482 23164 7488
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 22744 7268 22796 7274
rect 22664 7228 22744 7256
rect 22664 6866 22692 7228
rect 22744 7210 22796 7216
rect 22652 6860 22704 6866
rect 22652 6802 22704 6808
rect 22664 6458 22692 6802
rect 23124 6458 23152 7482
rect 23296 7200 23348 7206
rect 23296 7142 23348 7148
rect 23308 6934 23336 7142
rect 23296 6928 23348 6934
rect 23296 6870 23348 6876
rect 22652 6452 22704 6458
rect 22652 6394 22704 6400
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 23492 5914 23520 7482
rect 23952 7478 23980 7958
rect 24124 7880 24176 7886
rect 24124 7822 24176 7828
rect 24136 7546 24164 7822
rect 24320 7800 24348 8434
rect 25056 8294 25084 8978
rect 27618 8800 27674 8809
rect 27618 8735 27674 8744
rect 27632 8634 27660 8735
rect 27620 8628 27672 8634
rect 27620 8570 27672 8576
rect 24400 8288 24452 8294
rect 24400 8230 24452 8236
rect 25044 8288 25096 8294
rect 25044 8230 25096 8236
rect 25136 8288 25188 8294
rect 25136 8230 25188 8236
rect 24412 7886 24440 8230
rect 24400 7880 24452 7886
rect 24400 7822 24452 7828
rect 24228 7772 24348 7800
rect 24676 7812 24728 7818
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 23940 7472 23992 7478
rect 23940 7414 23992 7420
rect 23952 7206 23980 7414
rect 24228 7410 24256 7772
rect 24676 7754 24728 7760
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24688 7478 24716 7754
rect 24676 7472 24728 7478
rect 24676 7414 24728 7420
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 23940 7200 23992 7206
rect 23940 7142 23992 7148
rect 24228 6882 24256 7346
rect 25056 7002 25084 8230
rect 25148 7857 25176 8230
rect 25410 7984 25466 7993
rect 25410 7919 25466 7928
rect 25134 7848 25190 7857
rect 25134 7783 25190 7792
rect 25424 7546 25452 7919
rect 27618 7712 27674 7721
rect 27618 7647 27674 7656
rect 27632 7546 27660 7647
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 27620 7540 27672 7546
rect 27620 7482 27672 7488
rect 25044 6996 25096 7002
rect 25044 6938 25096 6944
rect 24676 6928 24728 6934
rect 24228 6854 24348 6882
rect 24676 6870 24728 6876
rect 25226 6896 25282 6905
rect 24320 6798 24348 6854
rect 24216 6792 24268 6798
rect 24216 6734 24268 6740
rect 24308 6792 24360 6798
rect 24308 6734 24360 6740
rect 23480 5908 23532 5914
rect 23480 5850 23532 5856
rect 24228 5574 24256 6734
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24688 6322 24716 6870
rect 25226 6831 25282 6840
rect 25240 6458 25268 6831
rect 25964 6724 26016 6730
rect 25964 6666 26016 6672
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 24676 6316 24728 6322
rect 24676 6258 24728 6264
rect 24582 6216 24638 6225
rect 24582 6151 24638 6160
rect 24596 5642 24624 6151
rect 24676 5772 24728 5778
rect 24676 5714 24728 5720
rect 24584 5636 24636 5642
rect 24584 5578 24636 5584
rect 24216 5568 24268 5574
rect 24216 5510 24268 5516
rect 24228 2650 24256 5510
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 5370 24716 5714
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 24398 5264 24454 5273
rect 24398 5199 24454 5208
rect 24412 4758 24440 5199
rect 24400 4752 24452 4758
rect 24400 4694 24452 4700
rect 24584 4684 24636 4690
rect 24636 4644 24716 4672
rect 24584 4626 24636 4632
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24688 4282 24716 4644
rect 24676 4276 24728 4282
rect 24676 4218 24728 4224
rect 24490 4040 24546 4049
rect 24490 3975 24546 3984
rect 24504 3670 24532 3975
rect 24492 3664 24544 3670
rect 24492 3606 24544 3612
rect 24584 3596 24636 3602
rect 24636 3556 24716 3584
rect 24584 3538 24636 3544
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24688 3194 24716 3556
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 24216 2644 24268 2650
rect 24216 2586 24268 2592
rect 25136 2508 25188 2514
rect 25136 2450 25188 2456
rect 25148 2310 25176 2450
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 25148 2009 25176 2246
rect 25134 2000 25190 2009
rect 25134 1935 25190 1944
rect 22742 82 22798 480
rect 22480 54 22798 82
rect 25976 82 26004 6666
rect 27618 6624 27674 6633
rect 27618 6559 27674 6568
rect 27632 6458 27660 6559
rect 27620 6452 27672 6458
rect 27620 6394 27672 6400
rect 27620 5772 27672 5778
rect 27620 5714 27672 5720
rect 27632 5681 27660 5714
rect 27618 5672 27674 5681
rect 27618 5607 27674 5616
rect 27618 4584 27674 4593
rect 27618 4519 27674 4528
rect 27632 4282 27660 4519
rect 27620 4276 27672 4282
rect 27620 4218 27672 4224
rect 27618 3496 27674 3505
rect 27618 3431 27674 3440
rect 27632 3194 27660 3431
rect 27620 3188 27672 3194
rect 27620 3130 27672 3136
rect 27618 2272 27674 2281
rect 27618 2207 27674 2216
rect 27632 513 27660 2207
rect 27618 504 27674 513
rect 26238 82 26294 480
rect 27618 439 27674 448
rect 25976 54 26294 82
rect 19246 0 19302 54
rect 22742 0 22798 54
rect 26238 0 26294 54
<< via2 >>
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 9494 21392 9550 21448
rect 9126 20440 9182 20496
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 8850 13368 8906 13424
rect 7562 10648 7618 10704
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10782 14320 10838 14376
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 9954 5208 10010 5264
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 13634 22480 13690 22536
rect 13266 13812 13268 13832
rect 13268 13812 13320 13832
rect 13320 13812 13322 13832
rect 13266 13776 13322 13812
rect 13450 13776 13506 13832
rect 10874 3984 10930 4040
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 14186 12144 14242 12200
rect 11886 2488 11942 2544
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 15382 14320 15438 14376
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14278 7928 14334 7984
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14462 7792 14518 7848
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 17038 23840 17094 23896
rect 16026 6840 16082 6896
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 16302 6160 16358 6216
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 17130 20476 17132 20496
rect 17132 20476 17184 20496
rect 17184 20476 17186 20496
rect 17130 20440 17186 20476
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 21454 22480 21510 22536
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 23386 21392 23442 21448
rect 17406 12144 17462 12200
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 23110 13368 23166 13424
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 20350 10648 20406 10704
rect 18326 2352 18382 2408
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 25134 25744 25190 25800
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 26146 26832 26202 26888
rect 25778 25064 25834 25120
rect 25502 24520 25558 24576
rect 24030 23840 24086 23896
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24766 22616 24822 22672
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24766 14592 24822 14648
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 25778 21664 25834 21720
rect 25778 20576 25834 20632
rect 26054 19488 26110 19544
rect 27618 19080 27674 19136
rect 25410 17448 25466 17504
rect 27618 17040 27674 17096
rect 27618 15952 27674 16008
rect 25410 14184 25466 14240
rect 25410 12416 25466 12472
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24950 11192 25006 11248
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24766 10240 24822 10296
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 25226 10104 25282 10160
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 27618 8744 27674 8800
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 25410 7928 25466 7984
rect 25134 7792 25190 7848
rect 27618 7656 27674 7712
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 25226 6840 25282 6896
rect 24582 6160 24638 6216
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24398 5208 24454 5264
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24490 3984 24546 4040
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 25134 1944 25190 2000
rect 27618 6568 27674 6624
rect 27618 5616 27674 5672
rect 27618 4528 27674 4584
rect 27618 3440 27674 3496
rect 27618 2216 27674 2272
rect 27618 448 27674 504
<< metal3 >>
rect 27520 27344 28000 27464
rect 26141 26890 26207 26893
rect 27662 26890 27722 27344
rect 26141 26888 27722 26890
rect 26141 26832 26146 26888
rect 26202 26832 27722 26888
rect 26141 26830 27722 26832
rect 26141 26827 26207 26830
rect 27520 26256 28000 26376
rect 25129 25802 25195 25805
rect 27662 25802 27722 26256
rect 25129 25800 27722 25802
rect 25129 25744 25134 25800
rect 25190 25744 27722 25800
rect 25129 25742 27722 25744
rect 25129 25739 25195 25742
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 27520 25304 28000 25424
rect 25773 25122 25839 25125
rect 27662 25122 27722 25304
rect 25773 25120 27722 25122
rect 25773 25064 25778 25120
rect 25834 25064 27722 25120
rect 25773 25062 27722 25064
rect 25773 25059 25839 25062
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 25497 24578 25563 24581
rect 25497 24576 27722 24578
rect 25497 24520 25502 24576
rect 25558 24520 27722 24576
rect 25497 24518 27722 24520
rect 25497 24515 25563 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 27662 24336 27722 24518
rect 27520 24216 28000 24336
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 17033 23898 17099 23901
rect 24025 23898 24091 23901
rect 17033 23896 24091 23898
rect 17033 23840 17038 23896
rect 17094 23840 24030 23896
rect 24086 23840 24091 23896
rect 17033 23838 24091 23840
rect 17033 23835 17099 23838
rect 24025 23835 24091 23838
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 27520 23128 28000 23248
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 24761 22674 24827 22677
rect 27662 22674 27722 23128
rect 24761 22672 27722 22674
rect 24761 22616 24766 22672
rect 24822 22616 27722 22672
rect 24761 22614 27722 22616
rect 24761 22611 24827 22614
rect 13629 22538 13695 22541
rect 21449 22538 21515 22541
rect 13629 22536 21515 22538
rect 13629 22480 13634 22536
rect 13690 22480 21454 22536
rect 21510 22480 21515 22536
rect 13629 22478 21515 22480
rect 13629 22475 13695 22478
rect 21449 22475 21515 22478
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 27520 22176 28000 22296
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 25773 21722 25839 21725
rect 27662 21722 27722 22176
rect 25773 21720 27722 21722
rect 25773 21664 25778 21720
rect 25834 21664 27722 21720
rect 25773 21662 27722 21664
rect 25773 21659 25839 21662
rect 9489 21450 9555 21453
rect 23381 21450 23447 21453
rect 9489 21448 23447 21450
rect 9489 21392 9494 21448
rect 9550 21392 23386 21448
rect 23442 21392 23447 21448
rect 9489 21390 23447 21392
rect 9489 21387 9555 21390
rect 23381 21387 23447 21390
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 27520 21088 28000 21208
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 25773 20634 25839 20637
rect 27662 20634 27722 21088
rect 25773 20632 27722 20634
rect 25773 20576 25778 20632
rect 25834 20576 27722 20632
rect 25773 20574 27722 20576
rect 25773 20571 25839 20574
rect 9121 20498 9187 20501
rect 17125 20498 17191 20501
rect 9121 20496 17191 20498
rect 9121 20440 9126 20496
rect 9182 20440 17130 20496
rect 17186 20440 17191 20496
rect 9121 20438 17191 20440
rect 9121 20435 9187 20438
rect 17125 20435 17191 20438
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 27520 20000 28000 20120
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 26049 19546 26115 19549
rect 27662 19546 27722 20000
rect 26049 19544 27722 19546
rect 26049 19488 26054 19544
rect 26110 19488 27722 19544
rect 26049 19486 27722 19488
rect 26049 19483 26115 19486
rect 27520 19136 28000 19168
rect 27520 19080 27618 19136
rect 27674 19080 28000 19136
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 27520 19048 28000 19080
rect 19610 19007 19930 19008
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 27520 17960 28000 18080
rect 19610 17919 19930 17920
rect 25405 17506 25471 17509
rect 27662 17506 27722 17960
rect 25405 17504 27722 17506
rect 25405 17448 25410 17504
rect 25466 17448 27722 17504
rect 25405 17446 27722 17448
rect 25405 17443 25471 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 27520 17096 28000 17128
rect 27520 17040 27618 17096
rect 27674 17040 28000 17096
rect 27520 17008 28000 17040
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 27520 16008 28000 16040
rect 27520 15952 27618 16008
rect 27674 15952 28000 16008
rect 27520 15920 28000 15952
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 27520 14832 28000 14952
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 24761 14650 24827 14653
rect 27662 14650 27722 14832
rect 24761 14648 27722 14650
rect 24761 14592 24766 14648
rect 24822 14592 27722 14648
rect 24761 14590 27722 14592
rect 24761 14587 24827 14590
rect 10777 14378 10843 14381
rect 15377 14378 15443 14381
rect 10777 14376 15443 14378
rect 10777 14320 10782 14376
rect 10838 14320 15382 14376
rect 15438 14320 15443 14376
rect 10777 14318 15443 14320
rect 10777 14315 10843 14318
rect 15377 14315 15443 14318
rect 25405 14242 25471 14245
rect 27654 14242 27660 14244
rect 25405 14240 27660 14242
rect 25405 14184 25410 14240
rect 25466 14184 27660 14240
rect 25405 14182 27660 14184
rect 25405 14179 25471 14182
rect 27654 14180 27660 14182
rect 27724 14180 27730 14244
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 27520 13972 28000 14000
rect 27520 13908 27660 13972
rect 27724 13908 28000 13972
rect 27520 13880 28000 13908
rect 13261 13834 13327 13837
rect 13445 13834 13511 13837
rect 13261 13832 13511 13834
rect 13261 13776 13266 13832
rect 13322 13776 13450 13832
rect 13506 13776 13511 13832
rect 13261 13774 13511 13776
rect 13261 13771 13327 13774
rect 13445 13771 13511 13774
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 8845 13426 8911 13429
rect 23105 13426 23171 13429
rect 8845 13424 23171 13426
rect 8845 13368 8850 13424
rect 8906 13368 23110 13424
rect 23166 13368 23171 13424
rect 8845 13366 23171 13368
rect 8845 13363 8911 13366
rect 23105 13363 23171 13366
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 27520 12792 28000 12912
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 25405 12474 25471 12477
rect 27662 12474 27722 12792
rect 25405 12472 27722 12474
rect 25405 12416 25410 12472
rect 25466 12416 27722 12472
rect 25405 12414 27722 12416
rect 25405 12411 25471 12414
rect 14181 12202 14247 12205
rect 17401 12202 17467 12205
rect 14181 12200 17467 12202
rect 14181 12144 14186 12200
rect 14242 12144 17406 12200
rect 17462 12144 17467 12200
rect 14181 12142 17467 12144
rect 14181 12139 14247 12142
rect 17401 12139 17467 12142
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 27520 11704 28000 11824
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 24945 11250 25011 11253
rect 27662 11250 27722 11704
rect 24945 11248 27722 11250
rect 24945 11192 24950 11248
rect 25006 11192 27722 11248
rect 24945 11190 27722 11192
rect 24945 11187 25011 11190
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 27520 10752 28000 10872
rect 7557 10706 7623 10709
rect 20345 10706 20411 10709
rect 7557 10704 20411 10706
rect 7557 10648 7562 10704
rect 7618 10648 20350 10704
rect 20406 10648 20411 10704
rect 7557 10646 20411 10648
rect 7557 10643 7623 10646
rect 20345 10643 20411 10646
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 24761 10298 24827 10301
rect 27662 10298 27722 10752
rect 24761 10296 27722 10298
rect 24761 10240 24766 10296
rect 24822 10240 27722 10296
rect 24761 10238 27722 10240
rect 24761 10235 24827 10238
rect 25221 10162 25287 10165
rect 25221 10160 27722 10162
rect 25221 10104 25226 10160
rect 25282 10104 27722 10160
rect 25221 10102 27722 10104
rect 25221 10099 25287 10102
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 27662 9784 27722 10102
rect 24277 9759 24597 9760
rect 27520 9664 28000 9784
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 27520 8800 28000 8832
rect 27520 8744 27618 8800
rect 27674 8744 28000 8800
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 27520 8712 28000 8744
rect 24277 8671 24597 8672
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 14273 7986 14339 7989
rect 25405 7986 25471 7989
rect 14273 7984 25471 7986
rect 14273 7928 14278 7984
rect 14334 7928 25410 7984
rect 25466 7928 25471 7984
rect 14273 7926 25471 7928
rect 14273 7923 14339 7926
rect 25405 7923 25471 7926
rect 14457 7850 14523 7853
rect 25129 7850 25195 7853
rect 14457 7848 25195 7850
rect 14457 7792 14462 7848
rect 14518 7792 25134 7848
rect 25190 7792 25195 7848
rect 14457 7790 25195 7792
rect 14457 7787 14523 7790
rect 25129 7787 25195 7790
rect 27520 7712 28000 7744
rect 27520 7656 27618 7712
rect 27674 7656 28000 7712
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 27520 7624 28000 7656
rect 24277 7583 24597 7584
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 16021 6898 16087 6901
rect 25221 6898 25287 6901
rect 16021 6896 25287 6898
rect 16021 6840 16026 6896
rect 16082 6840 25226 6896
rect 25282 6840 25287 6896
rect 16021 6838 25287 6840
rect 16021 6835 16087 6838
rect 25221 6835 25287 6838
rect 27520 6624 28000 6656
rect 27520 6568 27618 6624
rect 27674 6568 28000 6624
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 27520 6536 28000 6568
rect 24277 6495 24597 6496
rect 16297 6218 16363 6221
rect 24577 6218 24643 6221
rect 16297 6216 24643 6218
rect 16297 6160 16302 6216
rect 16358 6160 24582 6216
rect 24638 6160 24643 6216
rect 16297 6158 24643 6160
rect 16297 6155 16363 6158
rect 24577 6155 24643 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 27520 5672 28000 5704
rect 27520 5616 27618 5672
rect 27674 5616 28000 5672
rect 27520 5584 28000 5616
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 9949 5266 10015 5269
rect 24393 5266 24459 5269
rect 9949 5264 24459 5266
rect 9949 5208 9954 5264
rect 10010 5208 24398 5264
rect 24454 5208 24459 5264
rect 9949 5206 24459 5208
rect 9949 5203 10015 5206
rect 24393 5203 24459 5206
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 27520 4584 28000 4616
rect 27520 4528 27618 4584
rect 27674 4528 28000 4584
rect 27520 4496 28000 4528
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 10869 4042 10935 4045
rect 24485 4042 24551 4045
rect 10869 4040 24551 4042
rect 10869 3984 10874 4040
rect 10930 3984 24490 4040
rect 24546 3984 24551 4040
rect 10869 3982 24551 3984
rect 10869 3979 10935 3982
rect 24485 3979 24551 3982
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 27520 3496 28000 3528
rect 27520 3440 27618 3496
rect 27674 3440 28000 3496
rect 27520 3408 28000 3440
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 11881 2546 11947 2549
rect 27520 2548 28000 2576
rect 27470 2546 27476 2548
rect 11881 2544 27476 2546
rect 11881 2488 11886 2544
rect 11942 2488 27476 2544
rect 11881 2486 27476 2488
rect 11881 2483 11947 2486
rect 27470 2484 27476 2486
rect 27540 2484 27660 2548
rect 27724 2484 28000 2548
rect 27520 2456 28000 2484
rect 18321 2410 18387 2413
rect 18321 2408 27354 2410
rect 18321 2352 18326 2408
rect 18382 2352 27354 2408
rect 18321 2350 27354 2352
rect 18321 2347 18387 2350
rect 27294 2274 27354 2350
rect 27613 2274 27679 2277
rect 27294 2272 27679 2274
rect 27294 2216 27618 2272
rect 27674 2216 27679 2272
rect 27294 2214 27679 2216
rect 27613 2211 27679 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 25129 2002 25195 2005
rect 25129 2000 27722 2002
rect 25129 1944 25134 2000
rect 25190 1944 27722 2000
rect 25129 1942 27722 1944
rect 25129 1939 25195 1942
rect 27662 1488 27722 1942
rect 27520 1368 28000 1488
rect 27520 504 28000 536
rect 27520 448 27618 504
rect 27674 448 28000 504
rect 27520 416 28000 448
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 27660 14180 27724 14244
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 27660 13908 27724 13972
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 27476 2484 27540 2548
rect 27660 2484 27724 2548
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 27659 14244 27725 14245
rect 27659 14180 27660 14244
rect 27724 14180 27725 14244
rect 27659 14179 27725 14180
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 27662 13973 27722 14179
rect 27659 13972 27725 13973
rect 27659 13908 27660 13972
rect 27724 13908 27725 13972
rect 27659 13907 27725 13908
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 27475 2548 27541 2549
rect 27475 2484 27476 2548
rect 27540 2484 27541 2548
rect 27475 2483 27541 2484
rect 27659 2548 27725 2549
rect 27659 2484 27660 2548
rect 27724 2484 27725 2548
rect 27659 2483 27725 2484
rect 27478 2410 27538 2483
rect 27662 2410 27722 2483
rect 27478 2350 27722 2410
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_110 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11224 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_114
timestamp 1586364061
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_262
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_253
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_0_274
timestamp 1586364061
transform 1 0 26312 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_258
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_270
timestamp 1586364061
transform 1 0 25944 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_253
timestamp 1586364061
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_258
timestamp 1586364061
transform 1 0 24840 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_270
timestamp 1586364061
transform 1 0 25944 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18216 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_188
timestamp 1586364061
transform 1 0 18400 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_200
timestamp 1586364061
transform 1 0 19504 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_212
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_224
timestamp 1586364061
transform 1 0 21712 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 774 592
use scs8hd_decap_8  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_253
timestamp 1586364061
transform 1 0 24380 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_164
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_3  FILLER_7_172
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_177
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _208_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18124 0 1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_187
timestamp 1586364061
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_181
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_188
timestamp 1586364061
transform 1 0 18400 0 1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_199
timestamp 1586364061
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_199
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_211
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_211
timestamp 1586364061
transform 1 0 20516 0 1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 22540 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_223
timestamp 1586364061
transform 1 0 21620 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_231
timestamp 1586364061
transform 1 0 22356 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_235
timestamp 1586364061
transform 1 0 22724 0 1 5984
box -38 -48 590 592
use scs8hd_inv_8  _189_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use scs8hd_conb_1  _221_
timestamp 1586364061
transform 1 0 23460 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_246
timestamp 1586364061
transform 1 0 23736 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_241
timestamp 1586364061
transform 1 0 23276 0 1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24104 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_252
timestamp 1586364061
transform 1 0 24288 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_258
timestamp 1586364061
transform 1 0 24840 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_254
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_258
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_270
timestamp 1586364061
transform 1 0 25944 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_274
timestamp 1586364061
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_265
timestamp 1586364061
transform 1 0 25484 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_151
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 16008 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_158
timestamp 1586364061
transform 1 0 15640 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_161
timestamp 1586364061
transform 1 0 15916 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 17572 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_171
timestamp 1586364061
transform 1 0 16836 0 -1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_188
timestamp 1586364061
transform 1 0 18400 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_192
timestamp 1586364061
transform 1 0 18768 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_196
timestamp 1586364061
transform 1 0 19136 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_200
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_204
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_208
timestamp 1586364061
transform 1 0 20240 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_8  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_8  _188_
timestamp 1586364061
transform 1 0 22540 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22080 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_223
timestamp 1586364061
transform 1 0 21620 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_226
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_230
timestamp 1586364061
transform 1 0 22264 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_242
timestamp 1586364061
transform 1 0 23368 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_12  FILLER_8_259
timestamp 1586364061
transform 1 0 24932 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_271
timestamp 1586364061
transform 1 0 26036 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_nor2_4  _145_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_158
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_162
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_180
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_197
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_210
timestamp 1586364061
transform 1 0 20424 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21712 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_235
timestamp 1586364061
transform 1 0 22724 0 1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23828 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_241
timestamp 1586364061
transform 1 0 23276 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_262
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25392 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_273
timestamp 1586364061
transform 1 0 26220 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15732 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 15456 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_158
timestamp 1586364061
transform 1 0 15640 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_170
timestamp 1586364061
transform 1 0 16744 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_174
timestamp 1586364061
transform 1 0 17112 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_189
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_193
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 866 592
use scs8hd_fill_2  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 20240 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_210
timestamp 1586364061
transform 1 0 20424 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_10_223
timestamp 1586364061
transform 1 0 21620 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_235
timestamp 1586364061
transform 1 0 22724 0 -1 8160
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 -1 8160
box -38 -48 866 592
use scs8hd_fill_2  FILLER_10_247
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_258
timestamp 1586364061
transform 1 0 24840 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_270
timestamp 1586364061
transform 1 0 25944 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_274
timestamp 1586364061
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 13156 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_133
timestamp 1586364061
transform 1 0 13340 0 1 8160
box -38 -48 590 592
use scs8hd_buf_1  _132_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13892 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_142
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_146
timestamp 1586364061
transform 1 0 14536 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_150
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_11_162
timestamp 1586364061
transform 1 0 16008 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_177
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_181
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 20056 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_199
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_205
timestamp 1586364061
transform 1 0 19964 0 1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21252 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_217
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_221
timestamp 1586364061
transform 1 0 21436 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21620 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_225
timestamp 1586364061
transform 1 0 21804 0 1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23828 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_236
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_240
timestamp 1586364061
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_258
timestamp 1586364061
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_262
timestamp 1586364061
transform 1 0 25208 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_273
timestamp 1586364061
transform 1 0 26220 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_inv_8  _185_
timestamp 1586364061
transform 1 0 13156 0 -1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14904 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_140
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_148
timestamp 1586364061
transform 1 0 14720 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_152
timestamp 1586364061
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use scs8hd_conb_1  _219_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_157
timestamp 1586364061
transform 1 0 15548 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_161
timestamp 1586364061
transform 1 0 15916 0 -1 9248
box -38 -48 1142 592
use scs8hd_or2_4  _099_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 17204 0 -1 9248
box -38 -48 682 592
use scs8hd_fill_2  FILLER_12_173
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_182
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_8  _187_
timestamp 1586364061
transform 1 0 19228 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  FILLER_12_194
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_8  _186_
timestamp 1586364061
transform 1 0 22724 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24012 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_244
timestamp 1586364061
transform 1 0 23552 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_248
timestamp 1586364061
transform 1 0 23920 0 -1 9248
box -38 -48 130 592
use scs8hd_buf_2  _234_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24564 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_259
timestamp 1586364061
transform 1 0 24932 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_271
timestamp 1586364061
transform 1 0 26036 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13156 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_129
timestamp 1586364061
transform 1 0 12972 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_143
timestamp 1586364061
transform 1 0 14260 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_139
timestamp 1586364061
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_142
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_146
timestamp 1586364061
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14904 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_163
timestamp 1586364061
transform 1 0 16100 0 1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_8  _137_
timestamp 1586364061
transform 1 0 17020 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 774 592
use scs8hd_decap_4  FILLER_14_168
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_172
timestamp 1586364061
transform 1 0 16928 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_182
timestamp 1586364061
transform 1 0 17848 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 18216 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_192
timestamp 1586364061
transform 1 0 18768 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_188
timestamp 1586364061
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 18584 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 18676 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18952 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_207
timestamp 1586364061
transform 1 0 20148 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_200
timestamp 1586364061
transform 1 0 19504 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_204
timestamp 1586364061
transform 1 0 19872 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_14_210
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_211
timestamp 1586364061
transform 1 0 20516 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20332 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20700 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_219
timestamp 1586364061
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use scs8hd_conb_1  _220_
timestamp 1586364061
transform 1 0 21344 0 -1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22356 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22724 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_226
timestamp 1586364061
transform 1 0 21896 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_230
timestamp 1586364061
transform 1 0 22264 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_233
timestamp 1586364061
transform 1 0 22540 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_223
timestamp 1586364061
transform 1 0 21620 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_228
timestamp 1586364061
transform 1 0 22080 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_8  _192_
timestamp 1586364061
transform 1 0 23920 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 23920 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_237
timestamp 1586364061
transform 1 0 22908 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_243
timestamp 1586364061
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_240
timestamp 1586364061
transform 1 0 23184 0 -1 10336
box -38 -48 774 592
use scs8hd_buf_2  _233_
timestamp 1586364061
transform 1 0 24564 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24932 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_250
timestamp 1586364061
transform 1 0 24104 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_259
timestamp 1586364061
transform 1 0 24932 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_257
timestamp 1586364061
transform 1 0 24748 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_261
timestamp 1586364061
transform 1 0 25116 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_263
timestamp 1586364061
transform 1 0 25300 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_13_275
timestamp 1586364061
transform 1 0 26404 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_273
timestamp 1586364061
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_101
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_113
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_15_121
timestamp 1586364061
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12880 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_139
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use scs8hd_or4_4  _166_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_158
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_162
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 18400 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19688 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_201
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_204
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_221
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21896 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 21620 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_225
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_235
timestamp 1586364061
transform 1 0 22724 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 22908 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23920 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23276 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_239
timestamp 1586364061
transform 1 0 23092 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_243
timestamp 1586364061
transform 1 0 23460 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24288 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_250
timestamp 1586364061
transform 1 0 24104 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25484 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_263
timestamp 1586364061
transform 1 0 25300 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_267
timestamp 1586364061
transform 1 0 25668 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_275
timestamp 1586364061
transform 1 0 26404 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 590 592
use scs8hd_inv_8  _101_
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_12  FILLER_16_108
timestamp 1586364061
transform 1 0 11040 0 -1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_120
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 13156 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_133
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__D
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_143
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_147
timestamp 1586364061
transform 1 0 14628 0 -1 11424
box -38 -48 406 592
use scs8hd_inv_8  _184_
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 314 592
use scs8hd_nand2_4  _138_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 16928 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_168
timestamp 1586364061
transform 1 0 16560 0 -1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_183
timestamp 1586364061
transform 1 0 17940 0 -1 11424
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_194
timestamp 1586364061
transform 1 0 18952 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_199
timestamp 1586364061
transform 1 0 19412 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 22724 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_228
timestamp 1586364061
transform 1 0 22080 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_234
timestamp 1586364061
transform 1 0 22632 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_246
timestamp 1586364061
transform 1 0 23736 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24472 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_17_94
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use scs8hd_nand2_4  _108_
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use scs8hd_or2_4  _102_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_111
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_17_119
timestamp 1586364061
transform 1 0 12052 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_130
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_134
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 406 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 866 592
use scs8hd_decap_4  FILLER_17_149
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 406 592
use scs8hd_inv_8  _121_
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_153
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_156
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_160
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 18492 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__D
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_187
timestamp 1586364061
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_191
timestamp 1586364061
transform 1 0 18676 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 20056 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 19872 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_195
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_199
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_203
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_215
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 774 592
use scs8hd_conb_1  _213_
timestamp 1586364061
transform 1 0 22540 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21712 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22080 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_223
timestamp 1586364061
transform 1 0 21620 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_226
timestamp 1586364061
transform 1 0 21896 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_230
timestamp 1586364061
transform 1 0 22264 0 1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_236
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_248
timestamp 1586364061
transform 1 0 23920 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 24104 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_252
timestamp 1586364061
transform 1 0 24288 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_259
timestamp 1586364061
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 25484 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_263
timestamp 1586364061
transform 1 0 25300 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_267
timestamp 1586364061
transform 1 0 25668 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_275
timestamp 1586364061
transform 1 0 26404 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_8  _173_
timestamp 1586364061
transform 1 0 10396 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_97
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_100
timestamp 1586364061
transform 1 0 10304 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_110
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_1  _098_
timestamp 1586364061
transform 1 0 12144 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_114
timestamp 1586364061
transform 1 0 11592 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_18_123
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 13156 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_127
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_134
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_138
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__143__D
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__D
timestamp 1586364061
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _140_
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__C
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _146_
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__D
timestamp 1586364061
transform 1 0 17020 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_167
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_171
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_184
timestamp 1586364061
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_188
timestamp 1586364061
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_192
timestamp 1586364061
transform 1 0 18768 0 -1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21068 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21436 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_219
timestamp 1586364061
transform 1 0 21252 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_18_223
timestamp 1586364061
transform 1 0 21620 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_235
timestamp 1586364061
transform 1 0 22724 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 23644 0 -1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_18_243
timestamp 1586364061
transform 1 0 23460 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _232_
timestamp 1586364061
transform 1 0 25208 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_18_254
timestamp 1586364061
transform 1 0 24472 0 -1 12512
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_266
timestamp 1586364061
transform 1 0 25576 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_274
timestamp 1586364061
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_94
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_107
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_1  _109_
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_111
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_115
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_115
timestamp 1586364061
transform 1 0 11684 0 -1 13600
box -38 -48 774 592
use scs8hd_or4_4  _118_
timestamp 1586364061
transform 1 0 13432 0 -1 13600
box -38 -48 866 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 12972 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_138
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_126
timestamp 1586364061
transform 1 0 12696 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_130
timestamp 1586364061
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use scs8hd_or4_4  _143_
timestamp 1586364061
transform 1 0 14536 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 14536 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 14904 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_142
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_143
timestamp 1586364061
transform 1 0 14260 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_148
timestamp 1586364061
transform 1 0 14720 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_152
timestamp 1586364061
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_157
timestamp 1586364061
transform 1 0 15548 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_155
timestamp 1586364061
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 15732 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_1  _129_
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_161
timestamp 1586364061
transform 1 0 15916 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_163
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__D
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use scs8hd_or4_4  _134_
timestamp 1586364061
transform 1 0 17020 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_186
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_182
timestamp 1586364061
transform 1 0 17848 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_193
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 18768 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 18400 0 -1 13600
box -38 -48 222 592
use scs8hd_or4_4  _149_
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use scs8hd_buf_1  _139_
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 20056 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_199
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_204
timestamp 1586364061
transform 1 0 19872 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_194
timestamp 1586364061
transform 1 0 18952 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20976 0 1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_212
timestamp 1586364061
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22632 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_227
timestamp 1586364061
transform 1 0 21988 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_226
timestamp 1586364061
transform 1 0 21896 0 -1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_236
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_243
timestamp 1586364061
transform 1 0 23460 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_247
timestamp 1586364061
transform 1 0 23828 0 -1 13600
box -38 -48 406 592
use scs8hd_conb_1  _214_
timestamp 1586364061
transform 1 0 25208 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_254
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_258
timestamp 1586364061
transform 1 0 24840 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_260
timestamp 1586364061
transform 1 0 25024 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_265
timestamp 1586364061
transform 1 0 25484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_272
timestamp 1586364061
transform 1 0 26128 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_90
timestamp 1586364061
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_105
timestamp 1586364061
transform 1 0 10764 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 590 592
use scs8hd_decap_4  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 406 592
use scs8hd_or4_4  _115_
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_127
timestamp 1586364061
transform 1 0 12788 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_130
timestamp 1586364061
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_143
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_151
timestamp 1586364061
transform 1 0 14996 0 1 13600
box -38 -48 222 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 15364 0 1 13600
box -38 -48 314 592
use scs8hd_or4_4  _157_
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__D
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_158
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_162
timestamp 1586364061
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_or4_4  _160_
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__160__D
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_buf_1  _114_
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__C
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_204
timestamp 1586364061
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 21436 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_213
timestamp 1586364061
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_217
timestamp 1586364061
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_230
timestamp 1586364061
transform 1 0 22264 0 1 13600
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_238
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 406 592
use scs8hd_buf_2  _231_
timestamp 1586364061
transform 1 0 25208 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 24656 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_254
timestamp 1586364061
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_258
timestamp 1586364061
transform 1 0 24840 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 25760 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_266
timestamp 1586364061
transform 1 0 25576 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_270
timestamp 1586364061
transform 1 0 25944 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_276
timestamp 1586364061
transform 1 0 26496 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_6  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10212 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_101
timestamp 1586364061
transform 1 0 10396 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_107
timestamp 1586364061
transform 1 0 10948 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 774 592
use scs8hd_or4_4  _104_
timestamp 1586364061
transform 1 0 13340 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__D
timestamp 1586364061
transform 1 0 13156 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_125
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__C
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_142
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_146
timestamp 1586364061
transform 1 0 14536 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_150
timestamp 1586364061
transform 1 0 14904 0 -1 14688
box -38 -48 130 592
use scs8hd_inv_8  _095_
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 314 592
use scs8hd_or4_4  _153_
timestamp 1586364061
transform 1 0 17112 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__D
timestamp 1586364061
transform 1 0 16928 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_168
timestamp 1586364061
transform 1 0 16560 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 18124 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 18492 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18860 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_183
timestamp 1586364061
transform 1 0 17940 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_187
timestamp 1586364061
transform 1 0 18308 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_191
timestamp 1586364061
transform 1 0 18676 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_8  _198_
timestamp 1586364061
transform 1 0 19228 0 -1 14688
box -38 -48 866 592
use scs8hd_fill_2  FILLER_22_195
timestamp 1586364061
transform 1 0 19044 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21252 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22448 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_228
timestamp 1586364061
transform 1 0 22080 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_234
timestamp 1586364061
transform 1 0 22632 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 22816 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_6  FILLER_22_245
timestamp 1586364061
transform 1 0 23644 0 -1 14688
box -38 -48 590 592
use scs8hd_buf_2  _230_
timestamp 1586364061
transform 1 0 24564 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_253
timestamp 1586364061
transform 1 0 24380 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_259
timestamp 1586364061
transform 1 0 24932 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_271
timestamp 1586364061
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 8648 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_91
timestamp 1586364061
transform 1 0 9476 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_95
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _217_
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_or4_4  _110_
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 12880 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_126
timestamp 1586364061
transform 1 0 12696 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_130
timestamp 1586364061
transform 1 0 13064 0 1 14688
box -38 -48 222 592
use scs8hd_or4_4  _123_
timestamp 1586364061
transform 1 0 14996 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_143
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_160
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_164
timestamp 1586364061
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _152_
timestamp 1586364061
transform 1 0 16560 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 17020 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_or4_4  _163_
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_193
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19872 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19688 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_201
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 20884 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_213
timestamp 1586364061
transform 1 0 20700 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_217
timestamp 1586364061
transform 1 0 21068 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_221
timestamp 1586364061
transform 1 0 21436 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24012 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_236
timestamp 1586364061
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_240
timestamp 1586364061
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25208 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_260
timestamp 1586364061
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_264
timestamp 1586364061
transform 1 0 25392 0 1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_23_276
timestamp 1586364061
transform 1 0 26496 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_96
timestamp 1586364061
transform 1 0 9936 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 10120 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_100
timestamp 1586364061
transform 1 0 10304 0 -1 15776
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 12512 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_123
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 130 592
use scs8hd_or4_4  _126_
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__D
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_126
timestamp 1586364061
transform 1 0 12696 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_131
timestamp 1586364061
transform 1 0 13156 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_144
timestamp 1586364061
transform 1 0 14352 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_150
timestamp 1586364061
transform 1 0 14904 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 15640 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 15456 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_161
timestamp 1586364061
transform 1 0 15916 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_165
timestamp 1586364061
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 17020 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 16468 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 16836 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_169
timestamp 1586364061
transform 1 0 16652 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_176
timestamp 1586364061
transform 1 0 17296 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18768 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 18400 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_180
timestamp 1586364061
transform 1 0 17664 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_186
timestamp 1586364061
transform 1 0 18216 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_203
timestamp 1586364061
transform 1 0 19780 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_207
timestamp 1586364061
transform 1 0 20148 0 -1 15776
box -38 -48 590 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_213
timestamp 1586364061
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 22448 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_224
timestamp 1586364061
transform 1 0 21712 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_229
timestamp 1586364061
transform 1 0 22172 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 23828 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_243
timestamp 1586364061
transform 1 0 23460 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_249
timestamp 1586364061
transform 1 0 24012 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_12  FILLER_24_260
timestamp 1586364061
transform 1 0 25024 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_272
timestamp 1586364061
transform 1 0 26128 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_25_82
timestamp 1586364061
transform 1 0 8648 0 1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_87
timestamp 1586364061
transform 1 0 9108 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_91
timestamp 1586364061
transform 1 0 9476 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_104
timestamp 1586364061
transform 1 0 10672 0 1 15776
box -38 -48 774 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 12512 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_133
timestamp 1586364061
transform 1 0 13340 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_137
timestamp 1586364061
transform 1 0 13708 0 1 15776
box -38 -48 222 592
use scs8hd_inv_8  _183_
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_150
timestamp 1586364061
transform 1 0 14904 0 1 15776
box -38 -48 406 592
use scs8hd_nor3_4  _168_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_156
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_193
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19964 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19780 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_197
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_201
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 20976 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_214
timestamp 1586364061
transform 1 0 20792 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_218
timestamp 1586364061
transform 1 0 21160 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21528 0 1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21988 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22356 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_225
timestamp 1586364061
transform 1 0 21804 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_229
timestamp 1586364061
transform 1 0 22172 0 1 15776
box -38 -48 222 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 23828 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 23276 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_240
timestamp 1586364061
transform 1 0 23184 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_243
timestamp 1586364061
transform 1 0 23460 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_256
timestamp 1586364061
transform 1 0 24656 0 1 15776
box -38 -48 774 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 25392 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 25944 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_268
timestamp 1586364061
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_272
timestamp 1586364061
transform 1 0 26128 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_276
timestamp 1586364061
transform 1 0 26496 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 8464 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 590 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 9844 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_91
timestamp 1586364061
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_95
timestamp 1586364061
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_104
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_108
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_108
timestamp 1586364061
transform 1 0 11040 0 1 16864
box -38 -48 406 592
use scs8hd_inv_8  _172_
timestamp 1586364061
transform 1 0 11408 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_121
timestamp 1586364061
transform 1 0 12236 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12696 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12696 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_125
timestamp 1586364061
transform 1 0 12604 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_128
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_26_138
timestamp 1586364061
transform 1 0 13800 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_137
timestamp 1586364061
transform 1 0 13708 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14444 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_143
timestamp 1586364061
transform 1 0 14260 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_147
timestamp 1586364061
transform 1 0 14628 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_141
timestamp 1586364061
transform 1 0 14076 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_158
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_154
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_157
timestamp 1586364061
transform 1 0 15548 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_164
timestamp 1586364061
transform 1 0 16192 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_161
timestamp 1586364061
transform 1 0 15916 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 16008 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use scs8hd_nor3_4  _169_
timestamp 1586364061
transform 1 0 16008 0 1 16864
box -38 -48 1234 592
use scs8hd_nor3_4  _171_
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 18400 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_180
timestamp 1586364061
transform 1 0 17664 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_186
timestamp 1586364061
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use scs8hd_conb_1  _216_
timestamp 1586364061
transform 1 0 19780 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_197
timestamp 1586364061
transform 1 0 19228 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_6  FILLER_26_207
timestamp 1586364061
transform 1 0 20148 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_195
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_199
timestamp 1586364061
transform 1 0 19412 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_206
timestamp 1586364061
transform 1 0 20056 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 20792 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 20608 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_213
timestamp 1586364061
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_210
timestamp 1586364061
transform 1 0 20424 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_227
timestamp 1586364061
transform 1 0 21988 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_223
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_26_224
timestamp 1586364061
transform 1 0 21712 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22080 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 22080 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_230
timestamp 1586364061
transform 1 0 22264 0 1 16864
box -38 -48 314 592
use scs8hd_decap_6  FILLER_26_235
timestamp 1586364061
transform 1 0 22724 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_3  FILLER_26_230
timestamp 1586364061
transform 1 0 22264 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22540 0 -1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 16864
box -38 -48 314 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 23276 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_236
timestamp 1586364061
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _215_
timestamp 1586364061
transform 1 0 24840 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 25208 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24288 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_250
timestamp 1586364061
transform 1 0 24104 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_254
timestamp 1586364061
transform 1 0 24472 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_261
timestamp 1586364061
transform 1 0 25116 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_254
timestamp 1586364061
transform 1 0 24472 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_258
timestamp 1586364061
transform 1 0 24840 0 1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 25760 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_273
timestamp 1586364061
transform 1 0 26220 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_266
timestamp 1586364061
transform 1 0 25576 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_270
timestamp 1586364061
transform 1 0 25944 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_27_276
timestamp 1586364061
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_85
timestamp 1586364061
transform 1 0 8924 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_91
timestamp 1586364061
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_104
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_8  _175_
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_4  FILLER_28_121
timestamp 1586364061
transform 1 0 12236 0 -1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12696 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13248 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_125
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_128
timestamp 1586364061
transform 1 0 12880 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14720 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_150
timestamp 1586364061
transform 1 0 14904 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_8  _182_
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 16284 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_163
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use scs8hd_nor3_4  _170_
timestamp 1586364061
transform 1 0 16836 0 -1 17952
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 16652 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_167
timestamp 1586364061
transform 1 0 16468 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18860 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_184
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_188
timestamp 1586364061
transform 1 0 18400 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_192
timestamp 1586364061
transform 1 0 18768 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21068 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_210
timestamp 1586364061
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_220
timestamp 1586364061
transform 1 0 21344 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 22080 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21528 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21896 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_224
timestamp 1586364061
transform 1 0 21712 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23828 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 23644 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_8  FILLER_28_256
timestamp 1586364061
transform 1 0 24656 0 -1 17952
box -38 -48 774 592
use scs8hd_conb_1  _209_
timestamp 1586364061
transform 1 0 25392 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_267
timestamp 1586364061
transform 1 0 25668 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_80
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_29_92
timestamp 1586364061
transform 1 0 9568 0 1 17952
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10304 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_111
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_115
timestamp 1586364061
transform 1 0 11684 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_119
timestamp 1586364061
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_127
timestamp 1586364061
transform 1 0 12788 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14720 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14536 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_140
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_144
timestamp 1586364061
transform 1 0 14352 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 16284 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_157
timestamp 1586364061
transform 1 0 15548 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_161
timestamp 1586364061
transform 1 0 15916 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_168
timestamp 1586364061
transform 1 0 16560 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_173
timestamp 1586364061
transform 1 0 17020 0 1 17952
box -38 -48 774 592
use scs8hd_inv_8  _204_
timestamp 1586364061
transform 1 0 18400 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 18216 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_181
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_197
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_201
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_205
timestamp 1586364061
transform 1 0 19964 0 1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 20608 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_209
timestamp 1586364061
transform 1 0 20332 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_221
timestamp 1586364061
transform 1 0 21436 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 22080 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21712 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_226
timestamp 1586364061
transform 1 0 21896 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_230
timestamp 1586364061
transform 1 0 22264 0 1 17952
box -38 -48 314 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_236
timestamp 1586364061
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_240
timestamp 1586364061
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use scs8hd_buf_2  _228_
timestamp 1586364061
transform 1 0 25208 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 24656 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_254
timestamp 1586364061
transform 1 0 24472 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_258
timestamp 1586364061
transform 1 0 24840 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 25760 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_266
timestamp 1586364061
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_270
timestamp 1586364061
transform 1 0 25944 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_276
timestamp 1586364061
transform 1 0 26496 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11132 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10304 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_99
timestamp 1586364061
transform 1 0 10212 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_108
timestamp 1586364061
transform 1 0 11040 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_118
timestamp 1586364061
transform 1 0 11960 0 -1 19040
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 13800 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_135
timestamp 1586364061
transform 1 0 13524 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_140
timestamp 1586364061
transform 1 0 13984 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_152
timestamp 1586364061
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 16284 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_163
timestamp 1586364061
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_167
timestamp 1586364061
transform 1 0 16468 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_30_179
timestamp 1586364061
transform 1 0 17572 0 -1 19040
box -38 -48 222 592
use scs8hd_conb_1  _211_
timestamp 1586364061
transform 1 0 17756 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18768 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18216 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_184
timestamp 1586364061
transform 1 0 18032 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_188
timestamp 1586364061
transform 1 0 18400 0 -1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_201
timestamp 1586364061
transform 1 0 19596 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_205
timestamp 1586364061
transform 1 0 19964 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21068 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_213
timestamp 1586364061
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_220
timestamp 1586364061
transform 1 0 21344 0 -1 19040
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 22080 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21804 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_224
timestamp 1586364061
transform 1 0 21712 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_247
timestamp 1586364061
transform 1 0 23828 0 -1 19040
box -38 -48 130 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 24564 0 -1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24288 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_250
timestamp 1586364061
transform 1 0 24104 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_254
timestamp 1586364061
transform 1 0 24472 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_259
timestamp 1586364061
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_271
timestamp 1586364061
transform 1 0 26036 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_80
timestamp 1586364061
transform 1 0 8464 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_84
timestamp 1586364061
transform 1 0 8832 0 1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_31_92
timestamp 1586364061
transform 1 0 9568 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_95
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use scs8hd_inv_8  _174_
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_99
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 12604 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 12972 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_127
timestamp 1586364061
transform 1 0 12788 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_131
timestamp 1586364061
transform 1 0 13156 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 14904 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_152
timestamp 1586364061
transform 1 0 15088 0 1 19040
box -38 -48 222 592
use scs8hd_inv_8  _181_
timestamp 1586364061
transform 1 0 15640 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 15272 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_156
timestamp 1586364061
transform 1 0 15456 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_167
timestamp 1586364061
transform 1 0 16468 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_173
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_177
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_195
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_199
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _164_
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 21160 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_212
timestamp 1586364061
transform 1 0 20608 0 1 19040
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 22356 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_229
timestamp 1586364061
transform 1 0 22172 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_233
timestamp 1586364061
transform 1 0 22540 0 1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23920 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_237
timestamp 1586364061
transform 1 0 22908 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_240
timestamp 1586364061
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25484 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25944 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_268
timestamp 1586364061
transform 1 0 25760 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_272
timestamp 1586364061
transform 1 0 26128 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_276
timestamp 1586364061
transform 1 0 26496 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_conb_1  _222_
timestamp 1586364061
transform 1 0 11224 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_102
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 774 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 12512 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_113
timestamp 1586364061
transform 1 0 11500 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_32_121
timestamp 1586364061
transform 1 0 12236 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13524 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_133
timestamp 1586364061
transform 1 0 13340 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_137
timestamp 1586364061
transform 1 0 13708 0 -1 20128
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 590 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_163
timestamp 1586364061
transform 1 0 16100 0 -1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 17204 0 -1 20128
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_32_167
timestamp 1586364061
transform 1 0 16468 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_32_186
timestamp 1586364061
transform 1 0 18216 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_8  _206_
timestamp 1586364061
transform 1 0 19228 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_3  FILLER_32_194
timestamp 1586364061
transform 1 0 18952 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_206
timestamp 1586364061
transform 1 0 20056 0 -1 20128
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 21344 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_219
timestamp 1586364061
transform 1 0 21252 0 -1 20128
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21804 0 -1 20128
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_32_222
timestamp 1586364061
transform 1 0 21528 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23736 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23276 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_236
timestamp 1586364061
transform 1 0 22816 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_240
timestamp 1586364061
transform 1 0 23184 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_32_243
timestamp 1586364061
transform 1 0 23460 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24840 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_255
timestamp 1586364061
transform 1 0 24564 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_32_260
timestamp 1586364061
transform 1 0 25024 0 -1 20128
box -38 -48 314 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_266
timestamp 1586364061
transform 1 0 25576 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_274
timestamp 1586364061
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_33_82
timestamp 1586364061
transform 1 0 8648 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 9844 0 1 20128
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 8924 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_87
timestamp 1586364061
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_91
timestamp 1586364061
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_104
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_108
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_104
timestamp 1586364061
transform 1 0 10672 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_108
timestamp 1586364061
transform 1 0 11040 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use scs8hd_decap_6  FILLER_34_120
timestamp 1586364061
transform 1 0 12144 0 -1 21216
box -38 -48 590 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 12696 0 1 20128
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12696 0 -1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 13708 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_137
timestamp 1586364061
transform 1 0 13708 0 -1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14260 0 1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14076 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13892 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_139
timestamp 1586364061
transform 1 0 13892 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_154
timestamp 1586364061
transform 1 0 15272 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_158
timestamp 1586364061
transform 1 0 15640 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_165
timestamp 1586364061
transform 1 0 16284 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_173
timestamp 1586364061
transform 1 0 17020 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_177
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_169
timestamp 1586364061
transform 1 0 16652 0 -1 21216
box -38 -48 406 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 18768 0 1 20128
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18768 0 -1 21216
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18584 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_181
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 590 592
use scs8hd_decap_8  FILLER_34_182
timestamp 1586364061
transform 1 0 17848 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_195
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_199
timestamp 1586364061
transform 1 0 19412 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_203
timestamp 1586364061
transform 1 0 19780 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_207
timestamp 1586364061
transform 1 0 20148 0 -1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_212
timestamp 1586364061
transform 1 0 20608 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_213
timestamp 1586364061
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_34_221
timestamp 1586364061
transform 1 0 21436 0 -1 21216
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21528 0 -1 21216
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21528 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22356 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_224
timestamp 1586364061
transform 1 0 21712 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_228
timestamp 1586364061
transform 1 0 22080 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_233
timestamp 1586364061
transform 1 0 22540 0 -1 21216
box -38 -48 774 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23276 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_236
timestamp 1586364061
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_240
timestamp 1586364061
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_254
timestamp 1586364061
transform 1 0 24472 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_260
timestamp 1586364061
transform 1 0 25024 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_250
timestamp 1586364061
transform 1 0 24104 0 -1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_265
timestamp 1586364061
transform 1 0 25484 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_34_267
timestamp 1586364061
transform 1 0 25668 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4324 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_38
timestamp 1586364061
transform 1 0 4600 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_42
timestamp 1586364061
transform 1 0 4968 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_54
timestamp 1586364061
transform 1 0 6072 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_60
timestamp 1586364061
transform 1 0 6624 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_inv_8  _177_
timestamp 1586364061
transform 1 0 8556 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_78
timestamp 1586364061
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_90
timestamp 1586364061
transform 1 0 9384 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_35_109
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11316 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_113
timestamp 1586364061
transform 1 0 11500 0 1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_35_121
timestamp 1586364061
transform 1 0 12236 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13432 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 12880 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_127
timestamp 1586364061
transform 1 0 12788 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_130
timestamp 1586364061
transform 1 0 13064 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_145
timestamp 1586364061
transform 1 0 14444 0 1 21216
box -38 -48 774 592
use scs8hd_conb_1  _225_
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_153
timestamp 1586364061
transform 1 0 15180 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_158
timestamp 1586364061
transform 1 0 15640 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_162
timestamp 1586364061
transform 1 0 16008 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_175
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_179
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_35_192
timestamp 1586364061
transform 1 0 18768 0 1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19964 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19780 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_195
timestamp 1586364061
transform 1 0 19044 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_199
timestamp 1586364061
transform 1 0 19412 0 1 21216
box -38 -48 406 592
use scs8hd_decap_8  FILLER_35_214
timestamp 1586364061
transform 1 0 20792 0 1 21216
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21712 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21528 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_235
timestamp 1586364061
transform 1 0 22724 0 1 21216
box -38 -48 222 592
use scs8hd_inv_8  _197_
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 22908 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_239
timestamp 1586364061
transform 1 0 23092 0 1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_254
timestamp 1586364061
transform 1 0 24472 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_258
timestamp 1586364061
transform 1 0 24840 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_265
timestamp 1586364061
transform 1 0 25484 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_86
timestamp 1586364061
transform 1 0 9016 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_89
timestamp 1586364061
transform 1 0 9292 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_97
timestamp 1586364061
transform 1 0 10028 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_107
timestamp 1586364061
transform 1 0 10948 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_111
timestamp 1586364061
transform 1 0 11316 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_123
timestamp 1586364061
transform 1 0 12420 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_8  _179_
timestamp 1586364061
transform 1 0 13340 0 -1 22304
box -38 -48 866 592
use scs8hd_fill_2  FILLER_36_131
timestamp 1586364061
transform 1 0 13156 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_142
timestamp 1586364061
transform 1 0 14168 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  FILLER_36_150
timestamp 1586364061
transform 1 0 14904 0 -1 22304
box -38 -48 314 592
use scs8hd_inv_8  _180_
timestamp 1586364061
transform 1 0 15548 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 17112 0 -1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 18308 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_185
timestamp 1586364061
transform 1 0 18124 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_189
timestamp 1586364061
transform 1 0 18492 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 22304
box -38 -48 866 592
use scs8hd_fill_2  FILLER_36_206
timestamp 1586364061
transform 1 0 20056 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_210
timestamp 1586364061
transform 1 0 20424 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_8  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 22632 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21712 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22448 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_223
timestamp 1586364061
transform 1 0 21620 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_226
timestamp 1586364061
transform 1 0 21896 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_230
timestamp 1586364061
transform 1 0 22264 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23644 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24012 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_243
timestamp 1586364061
transform 1 0 23460 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_247
timestamp 1586364061
transform 1 0 23828 0 -1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_258
timestamp 1586364061
transform 1 0 24840 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_270
timestamp 1586364061
transform 1 0 25944 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_274
timestamp 1586364061
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8280 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 406 592
use scs8hd_decap_4  FILLER_37_80
timestamp 1586364061
transform 1 0 8464 0 1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9108 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_84
timestamp 1586364061
transform 1 0 8832 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_96
timestamp 1586364061
transform 1 0 9936 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_100
timestamp 1586364061
transform 1 0 10304 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_113
timestamp 1586364061
transform 1 0 11500 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_117
timestamp 1586364061
transform 1 0 11868 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_126
timestamp 1586364061
transform 1 0 12696 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_130
timestamp 1586364061
transform 1 0 13064 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_134
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13892 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_148
timestamp 1586364061
transform 1 0 14720 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_152
timestamp 1586364061
transform 1 0 15088 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_156
timestamp 1586364061
transform 1 0 15456 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_160
timestamp 1586364061
transform 1 0 15824 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_175
timestamp 1586364061
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_179
timestamp 1586364061
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_193
timestamp 1586364061
transform 1 0 18860 0 1 22304
box -38 -48 222 592
use scs8hd_inv_8  _199_
timestamp 1586364061
transform 1 0 19596 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 19412 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 19044 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_197
timestamp 1586364061
transform 1 0 19228 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21436 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_210
timestamp 1586364061
transform 1 0 20424 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_214
timestamp 1586364061
transform 1 0 20792 0 1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_37_217
timestamp 1586364061
transform 1 0 21068 0 1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_223
timestamp 1586364061
transform 1 0 21620 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_236
timestamp 1586364061
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_240
timestamp 1586364061
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_254
timestamp 1586364061
transform 1 0 24472 0 1 22304
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_265
timestamp 1586364061
transform 1 0 25484 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_273
timestamp 1586364061
transform 1 0 26220 0 1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8280 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_76
timestamp 1586364061
transform 1 0 8096 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_81
timestamp 1586364061
transform 1 0 8556 0 -1 23392
box -38 -48 774 592
use scs8hd_conb_1  _223_
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_38_89
timestamp 1586364061
transform 1 0 9292 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_6  FILLER_38_96
timestamp 1586364061
transform 1 0 9936 0 -1 23392
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 10488 0 -1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_113
timestamp 1586364061
transform 1 0 11500 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_8  FILLER_38_124
timestamp 1586364061
transform 1 0 12512 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_151
timestamp 1586364061
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_163
timestamp 1586364061
transform 1 0 16100 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17112 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17572 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_168
timestamp 1586364061
transform 1 0 16560 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_38_177
timestamp 1586364061
transform 1 0 17388 0 -1 23392
box -38 -48 222 592
use scs8hd_inv_8  _205_
timestamp 1586364061
transform 1 0 18124 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_4  FILLER_38_181
timestamp 1586364061
transform 1 0 17756 0 -1 23392
box -38 -48 406 592
use scs8hd_buf_2  _240_
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19136 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_194
timestamp 1586364061
transform 1 0 18952 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_198
timestamp 1586364061
transform 1 0 19320 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_38_206
timestamp 1586364061
transform 1 0 20056 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_218
timestamp 1586364061
transform 1 0 21160 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22080 0 -1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_38_226
timestamp 1586364061
transform 1 0 21896 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_38_237
timestamp 1586364061
transform 1 0 22908 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_254
timestamp 1586364061
transform 1 0 24472 0 -1 23392
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_265
timestamp 1586364061
transform 1 0 25484 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_38_273
timestamp 1586364061
transform 1 0 26220 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3220 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_39_22
timestamp 1586364061
transform 1 0 3128 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_26
timestamp 1586364061
transform 1 0 3496 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3680 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_30
timestamp 1586364061
transform 1 0 3864 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5336 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_42
timestamp 1586364061
transform 1 0 4968 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_49
timestamp 1586364061
transform 1 0 5612 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6348 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7360 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_60
timestamp 1586364061
transform 1 0 6624 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_71
timestamp 1586364061
transform 1 0 7636 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_75
timestamp 1586364061
transform 1 0 8004 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_79
timestamp 1586364061
transform 1 0 8372 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_83
timestamp 1586364061
transform 1 0 8740 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_72
timestamp 1586364061
transform 1 0 7728 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9476 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8924 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9936 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_87
timestamp 1586364061
transform 1 0 9108 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_94
timestamp 1586364061
transform 1 0 9752 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_84
timestamp 1586364061
transform 1 0 8832 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_8  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_8  _176_
timestamp 1586364061
transform 1 0 10488 0 1 23392
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10488 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10304 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_101
timestamp 1586364061
transform 1 0 10396 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_111
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_115
timestamp 1586364061
transform 1 0 11684 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_121
timestamp 1586364061
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_116
timestamp 1586364061
transform 1 0 11776 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_3  FILLER_40_124
timestamp 1586364061
transform 1 0 12512 0 -1 24480
box -38 -48 314 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 13708 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _242_
timestamp 1586364061
transform 1 0 12788 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 12604 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 13156 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 13708 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_129
timestamp 1586364061
transform 1 0 12972 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_133
timestamp 1586364061
transform 1 0 13340 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_131
timestamp 1586364061
transform 1 0 13156 0 -1 24480
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13892 0 -1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14260 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_141
timestamp 1586364061
transform 1 0 14076 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_145
timestamp 1586364061
transform 1 0 14444 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_142
timestamp 1586364061
transform 1 0 14168 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_3  FILLER_40_150
timestamp 1586364061
transform 1 0 14904 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_8  _178_
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 15824 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_158
timestamp 1586364061
transform 1 0 15640 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_162
timestamp 1586364061
transform 1 0 16008 0 1 23392
box -38 -48 590 592
use scs8hd_decap_8  FILLER_40_163
timestamp 1586364061
transform 1 0 16100 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_2  _237_
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 16652 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_168
timestamp 1586364061
transform 1 0 16560 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_174
timestamp 1586364061
transform 1 0 17112 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_8  _207_
timestamp 1586364061
transform 1 0 18124 0 1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_182
timestamp 1586364061
transform 1 0 17848 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_186
timestamp 1586364061
transform 1 0 18216 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19688 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_194
timestamp 1586364061
transform 1 0 18952 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_198
timestamp 1586364061
transform 1 0 19320 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_200
timestamp 1586364061
transform 1 0 19504 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_204
timestamp 1586364061
transform 1 0 19872 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 21252 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 20884 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_211
timestamp 1586364061
transform 1 0 20516 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_217
timestamp 1586364061
transform 1 0 21068 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_212
timestamp 1586364061
transform 1 0 20608 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_219
timestamp 1586364061
transform 1 0 21252 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_223
timestamp 1586364061
transform 1 0 21620 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_227
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_39_235
timestamp 1586364061
transform 1 0 22724 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_231
timestamp 1586364061
transform 1 0 22356 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 866 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 23644 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_240
timestamp 1586364061
transform 1 0 23184 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_243
timestamp 1586364061
transform 1 0 23460 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_249
timestamp 1586364061
transform 1 0 24012 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_2  _235_
timestamp 1586364061
transform 1 0 25208 0 1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24748 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_254
timestamp 1586364061
transform 1 0 24472 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_260
timestamp 1586364061
transform 1 0 25024 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 25760 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_266
timestamp 1586364061
transform 1 0 25576 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_270
timestamp 1586364061
transform 1 0 25944 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_276
timestamp 1586364061
transform 1 0 26496 0 1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_40_272
timestamp 1586364061
transform 1 0 26128 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9476 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9936 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_90
timestamp 1586364061
transform 1 0 9384 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_94
timestamp 1586364061
transform 1 0 9752 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_conb_1  _224_
timestamp 1586364061
transform 1 0 13708 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_126
timestamp 1586364061
transform 1 0 12696 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_130
timestamp 1586364061
transform 1 0 13064 0 1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_41_136
timestamp 1586364061
transform 1 0 13616 0 1 24480
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14720 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_140
timestamp 1586364061
transform 1 0 13984 0 1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_41_151
timestamp 1586364061
transform 1 0 14996 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15824 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15180 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16284 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_155
timestamp 1586364061
transform 1 0 15364 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_163
timestamp 1586364061
transform 1 0 16100 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_167
timestamp 1586364061
transform 1 0 16468 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_174
timestamp 1586364061
transform 1 0 17112 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_178
timestamp 1586364061
transform 1 0 17480 0 1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_193
timestamp 1586364061
transform 1 0 18860 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_205
timestamp 1586364061
transform 1 0 19964 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_217
timestamp 1586364061
transform 1 0 21068 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_229
timestamp 1586364061
transform 1 0 22172 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_41_241
timestamp 1586364061
transform 1 0 23276 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_253
timestamp 1586364061
transform 1 0 24380 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_258
timestamp 1586364061
transform 1 0 24840 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_262
timestamp 1586364061
transform 1 0 25208 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_41_266
timestamp 1586364061
transform 1 0 25576 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  FILLER_41_274
timestamp 1586364061
transform 1 0 26312 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_6  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_258
timestamp 1586364061
transform 1 0 24840 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_270
timestamp 1586364061
transform 1 0 25944 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_1  FILLER_42_276
timestamp 1586364061
transform 1 0 26496 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
<< labels >>
rlabel metal2 s 5262 0 5318 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 8758 0 8814 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 12254 0 12310 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 15750 0 15806 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 19246 0 19302 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 22742 0 22798 480 6 address[5]
port 5 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 chanx_right_in[0]
port 6 nsew default input
rlabel metal3 s 27520 2456 28000 2576 6 chanx_right_in[1]
port 7 nsew default input
rlabel metal3 s 27520 3408 28000 3528 6 chanx_right_in[2]
port 8 nsew default input
rlabel metal3 s 27520 4496 28000 4616 6 chanx_right_in[3]
port 9 nsew default input
rlabel metal3 s 27520 5584 28000 5704 6 chanx_right_in[4]
port 10 nsew default input
rlabel metal3 s 27520 6536 28000 6656 6 chanx_right_in[5]
port 11 nsew default input
rlabel metal3 s 27520 7624 28000 7744 6 chanx_right_in[6]
port 12 nsew default input
rlabel metal3 s 27520 8712 28000 8832 6 chanx_right_in[7]
port 13 nsew default input
rlabel metal3 s 27520 9664 28000 9784 6 chanx_right_in[8]
port 14 nsew default input
rlabel metal3 s 27520 10752 28000 10872 6 chanx_right_out[0]
port 15 nsew default tristate
rlabel metal3 s 27520 11704 28000 11824 6 chanx_right_out[1]
port 16 nsew default tristate
rlabel metal3 s 27520 12792 28000 12912 6 chanx_right_out[2]
port 17 nsew default tristate
rlabel metal3 s 27520 13880 28000 14000 6 chanx_right_out[3]
port 18 nsew default tristate
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_out[4]
port 19 nsew default tristate
rlabel metal3 s 27520 15920 28000 16040 6 chanx_right_out[5]
port 20 nsew default tristate
rlabel metal3 s 27520 17008 28000 17128 6 chanx_right_out[6]
port 21 nsew default tristate
rlabel metal3 s 27520 17960 28000 18080 6 chanx_right_out[7]
port 22 nsew default tristate
rlabel metal3 s 27520 19048 28000 19168 6 chanx_right_out[8]
port 23 nsew default tristate
rlabel metal2 s 8758 27520 8814 28000 6 chany_top_in[0]
port 24 nsew default input
rlabel metal2 s 9770 27520 9826 28000 6 chany_top_in[1]
port 25 nsew default input
rlabel metal2 s 10782 27520 10838 28000 6 chany_top_in[2]
port 26 nsew default input
rlabel metal2 s 11794 27520 11850 28000 6 chany_top_in[3]
port 27 nsew default input
rlabel metal2 s 12898 27520 12954 28000 6 chany_top_in[4]
port 28 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_in[5]
port 29 nsew default input
rlabel metal2 s 14922 27520 14978 28000 6 chany_top_in[6]
port 30 nsew default input
rlabel metal2 s 15934 27520 15990 28000 6 chany_top_in[7]
port 31 nsew default input
rlabel metal2 s 17038 27520 17094 28000 6 chany_top_in[8]
port 32 nsew default input
rlabel metal2 s 18050 27520 18106 28000 6 chany_top_out[0]
port 33 nsew default tristate
rlabel metal2 s 19062 27520 19118 28000 6 chany_top_out[1]
port 34 nsew default tristate
rlabel metal2 s 20074 27520 20130 28000 6 chany_top_out[2]
port 35 nsew default tristate
rlabel metal2 s 21178 27520 21234 28000 6 chany_top_out[3]
port 36 nsew default tristate
rlabel metal2 s 22190 27520 22246 28000 6 chany_top_out[4]
port 37 nsew default tristate
rlabel metal2 s 23202 27520 23258 28000 6 chany_top_out[5]
port 38 nsew default tristate
rlabel metal2 s 24214 27520 24270 28000 6 chany_top_out[6]
port 39 nsew default tristate
rlabel metal2 s 25318 27520 25374 28000 6 chany_top_out[7]
port 40 nsew default tristate
rlabel metal2 s 26330 27520 26386 28000 6 chany_top_out[8]
port 41 nsew default tristate
rlabel metal2 s 26238 0 26294 480 6 data_in
port 42 nsew default input
rlabel metal2 s 1766 0 1822 480 6 enable
port 43 nsew default input
rlabel metal3 s 27520 25304 28000 25424 6 right_bottom_grid_pin_11_
port 44 nsew default input
rlabel metal3 s 27520 26256 28000 26376 6 right_bottom_grid_pin_13_
port 45 nsew default input
rlabel metal3 s 27520 27344 28000 27464 6 right_bottom_grid_pin_15_
port 46 nsew default input
rlabel metal3 s 27520 20000 28000 20120 6 right_bottom_grid_pin_1_
port 47 nsew default input
rlabel metal3 s 27520 21088 28000 21208 6 right_bottom_grid_pin_3_
port 48 nsew default input
rlabel metal3 s 27520 22176 28000 22296 6 right_bottom_grid_pin_5_
port 49 nsew default input
rlabel metal3 s 27520 23128 28000 23248 6 right_bottom_grid_pin_7_
port 50 nsew default input
rlabel metal3 s 27520 24216 28000 24336 6 right_bottom_grid_pin_9_
port 51 nsew default input
rlabel metal3 s 27520 416 28000 536 6 right_top_grid_pin_10_
port 52 nsew default input
rlabel metal2 s 5630 27520 5686 28000 6 top_left_grid_pin_11_
port 53 nsew default input
rlabel metal2 s 6642 27520 6698 28000 6 top_left_grid_pin_13_
port 54 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 top_left_grid_pin_15_
port 55 nsew default input
rlabel metal2 s 478 27520 534 28000 6 top_left_grid_pin_1_
port 56 nsew default input
rlabel metal2 s 1490 27520 1546 28000 6 top_left_grid_pin_3_
port 57 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 top_left_grid_pin_5_
port 58 nsew default input
rlabel metal2 s 3514 27520 3570 28000 6 top_left_grid_pin_7_
port 59 nsew default input
rlabel metal2 s 4618 27520 4674 28000 6 top_left_grid_pin_9_
port 60 nsew default input
rlabel metal2 s 27342 27520 27398 28000 6 top_right_grid_pin_11_
port 61 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 62 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 63 nsew default input
<< end >>
