magic
tech sky130A
magscale 1 2
timestamp 1608156043
<< obsli1 >>
rect 1104 2159 21620 20145
<< obsm1 >>
rect 14 1300 22526 21956
<< metal2 >>
rect 294 22000 350 22800
rect 846 22000 902 22800
rect 1398 22000 1454 22800
rect 1950 22000 2006 22800
rect 2502 22000 2558 22800
rect 3054 22000 3110 22800
rect 3606 22000 3662 22800
rect 4158 22000 4214 22800
rect 4710 22000 4766 22800
rect 5262 22000 5318 22800
rect 5814 22000 5870 22800
rect 6366 22000 6422 22800
rect 6918 22000 6974 22800
rect 7470 22000 7526 22800
rect 8022 22000 8078 22800
rect 8574 22000 8630 22800
rect 9126 22000 9182 22800
rect 9678 22000 9734 22800
rect 10230 22000 10286 22800
rect 10782 22000 10838 22800
rect 11334 22000 11390 22800
rect 11978 22000 12034 22800
rect 12530 22000 12586 22800
rect 13082 22000 13138 22800
rect 13634 22000 13690 22800
rect 14186 22000 14242 22800
rect 14738 22000 14794 22800
rect 15290 22000 15346 22800
rect 15842 22000 15898 22800
rect 16394 22000 16450 22800
rect 16946 22000 17002 22800
rect 17498 22000 17554 22800
rect 18050 22000 18106 22800
rect 18602 22000 18658 22800
rect 19154 22000 19210 22800
rect 19706 22000 19762 22800
rect 20258 22000 20314 22800
rect 20810 22000 20866 22800
rect 21362 22000 21418 22800
rect 21914 22000 21970 22800
rect 22466 22000 22522 22800
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 1950 0 2006 800
rect 2502 0 2558 800
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4158 0 4214 800
rect 4710 0 4766 800
rect 5262 0 5318 800
rect 5814 0 5870 800
rect 6366 0 6422 800
rect 6918 0 6974 800
rect 7470 0 7526 800
rect 8022 0 8078 800
rect 8574 0 8630 800
rect 9126 0 9182 800
rect 9678 0 9734 800
rect 10230 0 10286 800
rect 10782 0 10838 800
rect 11334 0 11390 800
rect 11978 0 12034 800
rect 12530 0 12586 800
rect 13082 0 13138 800
rect 13634 0 13690 800
rect 14186 0 14242 800
rect 14738 0 14794 800
rect 15290 0 15346 800
rect 15842 0 15898 800
rect 16394 0 16450 800
rect 16946 0 17002 800
rect 17498 0 17554 800
rect 18050 0 18106 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21914 0 21970 800
rect 22466 0 22522 800
<< obsm2 >>
rect 20 21944 238 22545
rect 406 21944 790 22545
rect 958 21944 1342 22545
rect 1510 21944 1894 22545
rect 2062 21944 2446 22545
rect 2614 21944 2998 22545
rect 3166 21944 3550 22545
rect 3718 21944 4102 22545
rect 4270 21944 4654 22545
rect 4822 21944 5206 22545
rect 5374 21944 5758 22545
rect 5926 21944 6310 22545
rect 6478 21944 6862 22545
rect 7030 21944 7414 22545
rect 7582 21944 7966 22545
rect 8134 21944 8518 22545
rect 8686 21944 9070 22545
rect 9238 21944 9622 22545
rect 9790 21944 10174 22545
rect 10342 21944 10726 22545
rect 10894 21944 11278 22545
rect 11446 21944 11922 22545
rect 12090 21944 12474 22545
rect 12642 21944 13026 22545
rect 13194 21944 13578 22545
rect 13746 21944 14130 22545
rect 14298 21944 14682 22545
rect 14850 21944 15234 22545
rect 15402 21944 15786 22545
rect 15954 21944 16338 22545
rect 16506 21944 16890 22545
rect 17058 21944 17442 22545
rect 17610 21944 17994 22545
rect 18162 21944 18546 22545
rect 18714 21944 19098 22545
rect 19266 21944 19650 22545
rect 19818 21944 20202 22545
rect 20370 21944 20754 22545
rect 20922 21944 21306 22545
rect 21474 21944 21858 22545
rect 22026 21944 22410 22545
rect 20 856 22520 21944
rect 20 167 238 856
rect 406 167 790 856
rect 958 167 1342 856
rect 1510 167 1894 856
rect 2062 167 2446 856
rect 2614 167 2998 856
rect 3166 167 3550 856
rect 3718 167 4102 856
rect 4270 167 4654 856
rect 4822 167 5206 856
rect 5374 167 5758 856
rect 5926 167 6310 856
rect 6478 167 6862 856
rect 7030 167 7414 856
rect 7582 167 7966 856
rect 8134 167 8518 856
rect 8686 167 9070 856
rect 9238 167 9622 856
rect 9790 167 10174 856
rect 10342 167 10726 856
rect 10894 167 11278 856
rect 11446 167 11922 856
rect 12090 167 12474 856
rect 12642 167 13026 856
rect 13194 167 13578 856
rect 13746 167 14130 856
rect 14298 167 14682 856
rect 14850 167 15234 856
rect 15402 167 15786 856
rect 15954 167 16338 856
rect 16506 167 16890 856
rect 17058 167 17442 856
rect 17610 167 17994 856
rect 18162 167 18546 856
rect 18714 167 19098 856
rect 19266 167 19650 856
rect 19818 167 20202 856
rect 20370 167 20754 856
rect 20922 167 21306 856
rect 21474 167 21858 856
rect 22026 167 22410 856
<< metal3 >>
rect 22000 22448 22800 22568
rect 22000 22040 22800 22160
rect 22000 21496 22800 21616
rect 22000 21088 22800 21208
rect 22000 20544 22800 20664
rect 22000 20136 22800 20256
rect 22000 19728 22800 19848
rect 22000 19184 22800 19304
rect 22000 18776 22800 18896
rect 22000 18232 22800 18352
rect 22000 17824 22800 17944
rect 0 17144 800 17264
rect 22000 17280 22800 17400
rect 22000 16872 22800 16992
rect 22000 16464 22800 16584
rect 22000 15920 22800 16040
rect 22000 15512 22800 15632
rect 22000 14968 22800 15088
rect 22000 14560 22800 14680
rect 22000 14016 22800 14136
rect 22000 13608 22800 13728
rect 22000 13200 22800 13320
rect 22000 12656 22800 12776
rect 22000 12248 22800 12368
rect 22000 11704 22800 11824
rect 22000 11296 22800 11416
rect 22000 10752 22800 10872
rect 22000 10344 22800 10464
rect 22000 9936 22800 10056
rect 22000 9392 22800 9512
rect 22000 8984 22800 9104
rect 22000 8440 22800 8560
rect 22000 8032 22800 8152
rect 22000 7488 22800 7608
rect 22000 7080 22800 7200
rect 22000 6672 22800 6792
rect 22000 6128 22800 6248
rect 0 5720 800 5840
rect 22000 5720 22800 5840
rect 22000 5176 22800 5296
rect 22000 4768 22800 4888
rect 22000 4224 22800 4344
rect 22000 3816 22800 3936
rect 22000 3408 22800 3528
rect 22000 2864 22800 2984
rect 22000 2456 22800 2576
rect 22000 1912 22800 2032
rect 22000 1504 22800 1624
rect 22000 960 22800 1080
rect 22000 552 22800 672
rect 22000 144 22800 264
<< obsm3 >>
rect 800 22368 21920 22541
rect 800 22240 22000 22368
rect 800 21960 21920 22240
rect 800 21696 22000 21960
rect 800 21416 21920 21696
rect 800 21288 22000 21416
rect 800 21008 21920 21288
rect 800 20744 22000 21008
rect 800 20464 21920 20744
rect 800 20336 22000 20464
rect 800 20056 21920 20336
rect 800 19928 22000 20056
rect 800 19648 21920 19928
rect 800 19384 22000 19648
rect 800 19104 21920 19384
rect 800 18976 22000 19104
rect 800 18696 21920 18976
rect 800 18432 22000 18696
rect 800 18152 21920 18432
rect 800 18024 22000 18152
rect 800 17744 21920 18024
rect 800 17480 22000 17744
rect 800 17344 21920 17480
rect 880 17200 21920 17344
rect 880 17072 22000 17200
rect 880 17064 21920 17072
rect 800 16792 21920 17064
rect 800 16664 22000 16792
rect 800 16384 21920 16664
rect 800 16120 22000 16384
rect 800 15840 21920 16120
rect 800 15712 22000 15840
rect 800 15432 21920 15712
rect 800 15168 22000 15432
rect 800 14888 21920 15168
rect 800 14760 22000 14888
rect 800 14480 21920 14760
rect 800 14216 22000 14480
rect 800 13936 21920 14216
rect 800 13808 22000 13936
rect 800 13528 21920 13808
rect 800 13400 22000 13528
rect 800 13120 21920 13400
rect 800 12856 22000 13120
rect 800 12576 21920 12856
rect 800 12448 22000 12576
rect 800 12168 21920 12448
rect 800 11904 22000 12168
rect 800 11624 21920 11904
rect 800 11496 22000 11624
rect 800 11216 21920 11496
rect 800 10952 22000 11216
rect 800 10672 21920 10952
rect 800 10544 22000 10672
rect 800 10264 21920 10544
rect 800 10136 22000 10264
rect 800 9856 21920 10136
rect 800 9592 22000 9856
rect 800 9312 21920 9592
rect 800 9184 22000 9312
rect 800 8904 21920 9184
rect 800 8640 22000 8904
rect 800 8360 21920 8640
rect 800 8232 22000 8360
rect 800 7952 21920 8232
rect 800 7688 22000 7952
rect 800 7408 21920 7688
rect 800 7280 22000 7408
rect 800 7000 21920 7280
rect 800 6872 22000 7000
rect 800 6592 21920 6872
rect 800 6328 22000 6592
rect 800 6048 21920 6328
rect 800 5920 22000 6048
rect 880 5640 21920 5920
rect 800 5376 22000 5640
rect 800 5096 21920 5376
rect 800 4968 22000 5096
rect 800 4688 21920 4968
rect 800 4424 22000 4688
rect 800 4144 21920 4424
rect 800 4016 22000 4144
rect 800 3736 21920 4016
rect 800 3608 22000 3736
rect 800 3328 21920 3608
rect 800 3064 22000 3328
rect 800 2784 21920 3064
rect 800 2656 22000 2784
rect 800 2376 21920 2656
rect 800 2112 22000 2376
rect 800 1832 21920 2112
rect 800 1704 22000 1832
rect 800 1424 21920 1704
rect 800 1160 22000 1424
rect 800 880 21920 1160
rect 800 752 22000 880
rect 800 472 21920 752
rect 800 344 22000 472
rect 800 171 21920 344
<< metal4 >>
rect 4376 2128 4696 20176
rect 7808 2128 8128 20176
<< obsm4 >>
rect 11240 1531 19261 20176
<< labels >>
rlabel metal2 s 294 0 350 800 6 bottom_left_grid_pin_1_
port 1 nsew default input
rlabel metal3 s 0 5720 800 5840 6 ccff_head
port 2 nsew default input
rlabel metal3 s 0 17144 800 17264 6 ccff_tail
port 3 nsew default output
rlabel metal3 s 22000 3816 22800 3936 6 chanx_right_in[0]
port 4 nsew default input
rlabel metal3 s 22000 8440 22800 8560 6 chanx_right_in[10]
port 5 nsew default input
rlabel metal3 s 22000 8984 22800 9104 6 chanx_right_in[11]
port 6 nsew default input
rlabel metal3 s 22000 9392 22800 9512 6 chanx_right_in[12]
port 7 nsew default input
rlabel metal3 s 22000 9936 22800 10056 6 chanx_right_in[13]
port 8 nsew default input
rlabel metal3 s 22000 10344 22800 10464 6 chanx_right_in[14]
port 9 nsew default input
rlabel metal3 s 22000 10752 22800 10872 6 chanx_right_in[15]
port 10 nsew default input
rlabel metal3 s 22000 11296 22800 11416 6 chanx_right_in[16]
port 11 nsew default input
rlabel metal3 s 22000 11704 22800 11824 6 chanx_right_in[17]
port 12 nsew default input
rlabel metal3 s 22000 12248 22800 12368 6 chanx_right_in[18]
port 13 nsew default input
rlabel metal3 s 22000 12656 22800 12776 6 chanx_right_in[19]
port 14 nsew default input
rlabel metal3 s 22000 4224 22800 4344 6 chanx_right_in[1]
port 15 nsew default input
rlabel metal3 s 22000 4768 22800 4888 6 chanx_right_in[2]
port 16 nsew default input
rlabel metal3 s 22000 5176 22800 5296 6 chanx_right_in[3]
port 17 nsew default input
rlabel metal3 s 22000 5720 22800 5840 6 chanx_right_in[4]
port 18 nsew default input
rlabel metal3 s 22000 6128 22800 6248 6 chanx_right_in[5]
port 19 nsew default input
rlabel metal3 s 22000 6672 22800 6792 6 chanx_right_in[6]
port 20 nsew default input
rlabel metal3 s 22000 7080 22800 7200 6 chanx_right_in[7]
port 21 nsew default input
rlabel metal3 s 22000 7488 22800 7608 6 chanx_right_in[8]
port 22 nsew default input
rlabel metal3 s 22000 8032 22800 8152 6 chanx_right_in[9]
port 23 nsew default input
rlabel metal3 s 22000 13200 22800 13320 6 chanx_right_out[0]
port 24 nsew default output
rlabel metal3 s 22000 17824 22800 17944 6 chanx_right_out[10]
port 25 nsew default output
rlabel metal3 s 22000 18232 22800 18352 6 chanx_right_out[11]
port 26 nsew default output
rlabel metal3 s 22000 18776 22800 18896 6 chanx_right_out[12]
port 27 nsew default output
rlabel metal3 s 22000 19184 22800 19304 6 chanx_right_out[13]
port 28 nsew default output
rlabel metal3 s 22000 19728 22800 19848 6 chanx_right_out[14]
port 29 nsew default output
rlabel metal3 s 22000 20136 22800 20256 6 chanx_right_out[15]
port 30 nsew default output
rlabel metal3 s 22000 20544 22800 20664 6 chanx_right_out[16]
port 31 nsew default output
rlabel metal3 s 22000 21088 22800 21208 6 chanx_right_out[17]
port 32 nsew default output
rlabel metal3 s 22000 21496 22800 21616 6 chanx_right_out[18]
port 33 nsew default output
rlabel metal3 s 22000 22040 22800 22160 6 chanx_right_out[19]
port 34 nsew default output
rlabel metal3 s 22000 13608 22800 13728 6 chanx_right_out[1]
port 35 nsew default output
rlabel metal3 s 22000 14016 22800 14136 6 chanx_right_out[2]
port 36 nsew default output
rlabel metal3 s 22000 14560 22800 14680 6 chanx_right_out[3]
port 37 nsew default output
rlabel metal3 s 22000 14968 22800 15088 6 chanx_right_out[4]
port 38 nsew default output
rlabel metal3 s 22000 15512 22800 15632 6 chanx_right_out[5]
port 39 nsew default output
rlabel metal3 s 22000 15920 22800 16040 6 chanx_right_out[6]
port 40 nsew default output
rlabel metal3 s 22000 16464 22800 16584 6 chanx_right_out[7]
port 41 nsew default output
rlabel metal3 s 22000 16872 22800 16992 6 chanx_right_out[8]
port 42 nsew default output
rlabel metal3 s 22000 17280 22800 17400 6 chanx_right_out[9]
port 43 nsew default output
rlabel metal2 s 846 0 902 800 6 chany_bottom_in[0]
port 44 nsew default input
rlabel metal2 s 6366 0 6422 800 6 chany_bottom_in[10]
port 45 nsew default input
rlabel metal2 s 6918 0 6974 800 6 chany_bottom_in[11]
port 46 nsew default input
rlabel metal2 s 7470 0 7526 800 6 chany_bottom_in[12]
port 47 nsew default input
rlabel metal2 s 8022 0 8078 800 6 chany_bottom_in[13]
port 48 nsew default input
rlabel metal2 s 8574 0 8630 800 6 chany_bottom_in[14]
port 49 nsew default input
rlabel metal2 s 9126 0 9182 800 6 chany_bottom_in[15]
port 50 nsew default input
rlabel metal2 s 9678 0 9734 800 6 chany_bottom_in[16]
port 51 nsew default input
rlabel metal2 s 10230 0 10286 800 6 chany_bottom_in[17]
port 52 nsew default input
rlabel metal2 s 10782 0 10838 800 6 chany_bottom_in[18]
port 53 nsew default input
rlabel metal2 s 11334 0 11390 800 6 chany_bottom_in[19]
port 54 nsew default input
rlabel metal2 s 1398 0 1454 800 6 chany_bottom_in[1]
port 55 nsew default input
rlabel metal2 s 1950 0 2006 800 6 chany_bottom_in[2]
port 56 nsew default input
rlabel metal2 s 2502 0 2558 800 6 chany_bottom_in[3]
port 57 nsew default input
rlabel metal2 s 3054 0 3110 800 6 chany_bottom_in[4]
port 58 nsew default input
rlabel metal2 s 3606 0 3662 800 6 chany_bottom_in[5]
port 59 nsew default input
rlabel metal2 s 4158 0 4214 800 6 chany_bottom_in[6]
port 60 nsew default input
rlabel metal2 s 4710 0 4766 800 6 chany_bottom_in[7]
port 61 nsew default input
rlabel metal2 s 5262 0 5318 800 6 chany_bottom_in[8]
port 62 nsew default input
rlabel metal2 s 5814 0 5870 800 6 chany_bottom_in[9]
port 63 nsew default input
rlabel metal2 s 11978 0 12034 800 6 chany_bottom_out[0]
port 64 nsew default output
rlabel metal2 s 17498 0 17554 800 6 chany_bottom_out[10]
port 65 nsew default output
rlabel metal2 s 18050 0 18106 800 6 chany_bottom_out[11]
port 66 nsew default output
rlabel metal2 s 18602 0 18658 800 6 chany_bottom_out[12]
port 67 nsew default output
rlabel metal2 s 19154 0 19210 800 6 chany_bottom_out[13]
port 68 nsew default output
rlabel metal2 s 19706 0 19762 800 6 chany_bottom_out[14]
port 69 nsew default output
rlabel metal2 s 20258 0 20314 800 6 chany_bottom_out[15]
port 70 nsew default output
rlabel metal2 s 20810 0 20866 800 6 chany_bottom_out[16]
port 71 nsew default output
rlabel metal2 s 21362 0 21418 800 6 chany_bottom_out[17]
port 72 nsew default output
rlabel metal2 s 21914 0 21970 800 6 chany_bottom_out[18]
port 73 nsew default output
rlabel metal2 s 22466 0 22522 800 6 chany_bottom_out[19]
port 74 nsew default output
rlabel metal2 s 12530 0 12586 800 6 chany_bottom_out[1]
port 75 nsew default output
rlabel metal2 s 13082 0 13138 800 6 chany_bottom_out[2]
port 76 nsew default output
rlabel metal2 s 13634 0 13690 800 6 chany_bottom_out[3]
port 77 nsew default output
rlabel metal2 s 14186 0 14242 800 6 chany_bottom_out[4]
port 78 nsew default output
rlabel metal2 s 14738 0 14794 800 6 chany_bottom_out[5]
port 79 nsew default output
rlabel metal2 s 15290 0 15346 800 6 chany_bottom_out[6]
port 80 nsew default output
rlabel metal2 s 15842 0 15898 800 6 chany_bottom_out[7]
port 81 nsew default output
rlabel metal2 s 16394 0 16450 800 6 chany_bottom_out[8]
port 82 nsew default output
rlabel metal2 s 16946 0 17002 800 6 chany_bottom_out[9]
port 83 nsew default output
rlabel metal2 s 846 22000 902 22800 6 chany_top_in[0]
port 84 nsew default input
rlabel metal2 s 6366 22000 6422 22800 6 chany_top_in[10]
port 85 nsew default input
rlabel metal2 s 6918 22000 6974 22800 6 chany_top_in[11]
port 86 nsew default input
rlabel metal2 s 7470 22000 7526 22800 6 chany_top_in[12]
port 87 nsew default input
rlabel metal2 s 8022 22000 8078 22800 6 chany_top_in[13]
port 88 nsew default input
rlabel metal2 s 8574 22000 8630 22800 6 chany_top_in[14]
port 89 nsew default input
rlabel metal2 s 9126 22000 9182 22800 6 chany_top_in[15]
port 90 nsew default input
rlabel metal2 s 9678 22000 9734 22800 6 chany_top_in[16]
port 91 nsew default input
rlabel metal2 s 10230 22000 10286 22800 6 chany_top_in[17]
port 92 nsew default input
rlabel metal2 s 10782 22000 10838 22800 6 chany_top_in[18]
port 93 nsew default input
rlabel metal2 s 11334 22000 11390 22800 6 chany_top_in[19]
port 94 nsew default input
rlabel metal2 s 1398 22000 1454 22800 6 chany_top_in[1]
port 95 nsew default input
rlabel metal2 s 1950 22000 2006 22800 6 chany_top_in[2]
port 96 nsew default input
rlabel metal2 s 2502 22000 2558 22800 6 chany_top_in[3]
port 97 nsew default input
rlabel metal2 s 3054 22000 3110 22800 6 chany_top_in[4]
port 98 nsew default input
rlabel metal2 s 3606 22000 3662 22800 6 chany_top_in[5]
port 99 nsew default input
rlabel metal2 s 4158 22000 4214 22800 6 chany_top_in[6]
port 100 nsew default input
rlabel metal2 s 4710 22000 4766 22800 6 chany_top_in[7]
port 101 nsew default input
rlabel metal2 s 5262 22000 5318 22800 6 chany_top_in[8]
port 102 nsew default input
rlabel metal2 s 5814 22000 5870 22800 6 chany_top_in[9]
port 103 nsew default input
rlabel metal2 s 11978 22000 12034 22800 6 chany_top_out[0]
port 104 nsew default output
rlabel metal2 s 17498 22000 17554 22800 6 chany_top_out[10]
port 105 nsew default output
rlabel metal2 s 18050 22000 18106 22800 6 chany_top_out[11]
port 106 nsew default output
rlabel metal2 s 18602 22000 18658 22800 6 chany_top_out[12]
port 107 nsew default output
rlabel metal2 s 19154 22000 19210 22800 6 chany_top_out[13]
port 108 nsew default output
rlabel metal2 s 19706 22000 19762 22800 6 chany_top_out[14]
port 109 nsew default output
rlabel metal2 s 20258 22000 20314 22800 6 chany_top_out[15]
port 110 nsew default output
rlabel metal2 s 20810 22000 20866 22800 6 chany_top_out[16]
port 111 nsew default output
rlabel metal2 s 21362 22000 21418 22800 6 chany_top_out[17]
port 112 nsew default output
rlabel metal2 s 21914 22000 21970 22800 6 chany_top_out[18]
port 113 nsew default output
rlabel metal2 s 22466 22000 22522 22800 6 chany_top_out[19]
port 114 nsew default output
rlabel metal2 s 12530 22000 12586 22800 6 chany_top_out[1]
port 115 nsew default output
rlabel metal2 s 13082 22000 13138 22800 6 chany_top_out[2]
port 116 nsew default output
rlabel metal2 s 13634 22000 13690 22800 6 chany_top_out[3]
port 117 nsew default output
rlabel metal2 s 14186 22000 14242 22800 6 chany_top_out[4]
port 118 nsew default output
rlabel metal2 s 14738 22000 14794 22800 6 chany_top_out[5]
port 119 nsew default output
rlabel metal2 s 15290 22000 15346 22800 6 chany_top_out[6]
port 120 nsew default output
rlabel metal2 s 15842 22000 15898 22800 6 chany_top_out[7]
port 121 nsew default output
rlabel metal2 s 16394 22000 16450 22800 6 chany_top_out[8]
port 122 nsew default output
rlabel metal2 s 16946 22000 17002 22800 6 chany_top_out[9]
port 123 nsew default output
rlabel metal3 s 22000 22448 22800 22568 6 prog_clk_0_E_in
port 124 nsew default input
rlabel metal3 s 22000 144 22800 264 6 right_bottom_grid_pin_34_
port 125 nsew default input
rlabel metal3 s 22000 552 22800 672 6 right_bottom_grid_pin_35_
port 126 nsew default input
rlabel metal3 s 22000 960 22800 1080 6 right_bottom_grid_pin_36_
port 127 nsew default input
rlabel metal3 s 22000 1504 22800 1624 6 right_bottom_grid_pin_37_
port 128 nsew default input
rlabel metal3 s 22000 1912 22800 2032 6 right_bottom_grid_pin_38_
port 129 nsew default input
rlabel metal3 s 22000 2456 22800 2576 6 right_bottom_grid_pin_39_
port 130 nsew default input
rlabel metal3 s 22000 2864 22800 2984 6 right_bottom_grid_pin_40_
port 131 nsew default input
rlabel metal3 s 22000 3408 22800 3528 6 right_bottom_grid_pin_41_
port 132 nsew default input
rlabel metal2 s 294 22000 350 22800 6 top_left_grid_pin_1_
port 133 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 134 nsew power input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 135 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 22800 22800
string LEFview TRUE
<< end >>
