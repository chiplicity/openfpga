magic
tech sky130A
magscale 1 2
timestamp 1608764939
<< checkpaint >>
rect -1260 -1260 18260 21260
<< locali >>
rect 8309 14807 8343 14909
rect 11345 14331 11379 14501
rect 4997 12223 5031 12393
rect 4629 11203 4663 11305
rect 2731 10217 2823 10251
rect 2789 9979 2823 10217
rect 2697 7259 2731 7361
rect 10517 6647 10551 6817
rect 8125 5015 8159 5117
rect 12265 5015 12299 5321
<< viali >>
rect 3065 17289 3099 17323
rect 4997 17289 5031 17323
rect 5549 17289 5583 17323
rect 6101 17289 6135 17323
rect 9965 17289 9999 17323
rect 1777 17221 1811 17255
rect 3617 17221 3651 17255
rect 7113 17221 7147 17255
rect 10701 17221 10735 17255
rect 8217 17153 8251 17187
rect 9229 17153 9263 17187
rect 11345 17153 11379 17187
rect 13185 17153 13219 17187
rect 14105 17153 14139 17187
rect 15117 17153 15151 17187
rect 1593 17085 1627 17119
rect 2881 17085 2915 17119
rect 3433 17085 3467 17119
rect 4813 17085 4847 17119
rect 5365 17085 5399 17119
rect 5917 17085 5951 17119
rect 6929 17085 6963 17119
rect 8033 17085 8067 17119
rect 9781 17085 9815 17119
rect 11069 17085 11103 17119
rect 8125 17017 8159 17051
rect 14197 17017 14231 17051
rect 7665 16949 7699 16983
rect 8677 16949 8711 16983
rect 9045 16949 9079 16983
rect 9137 16949 9171 16983
rect 11161 16949 11195 16983
rect 12633 16949 12667 16983
rect 13001 16949 13035 16983
rect 13093 16949 13127 16983
rect 1777 16745 1811 16779
rect 2329 16745 2363 16779
rect 4537 16745 4571 16779
rect 6745 16745 6779 16779
rect 8401 16745 8435 16779
rect 10149 16745 10183 16779
rect 11069 16745 11103 16779
rect 11529 16745 11563 16779
rect 13737 16745 13771 16779
rect 3157 16677 3191 16711
rect 5632 16677 5666 16711
rect 7266 16677 7300 16711
rect 1593 16609 1627 16643
rect 2145 16609 2179 16643
rect 2881 16609 2915 16643
rect 4353 16609 4387 16643
rect 7021 16609 7055 16643
rect 8677 16609 8711 16643
rect 10057 16609 10091 16643
rect 11437 16609 11471 16643
rect 12624 16609 12658 16643
rect 14197 16609 14231 16643
rect 14565 16609 14599 16643
rect 5365 16541 5399 16575
rect 10333 16541 10367 16575
rect 11713 16541 11747 16575
rect 12357 16541 12391 16575
rect 14933 16541 14967 16575
rect 8861 16405 8895 16439
rect 9689 16405 9723 16439
rect 2513 16201 2547 16235
rect 3617 16201 3651 16235
rect 4169 16201 4203 16235
rect 5365 16201 5399 16235
rect 8033 16201 8067 16235
rect 12449 16201 12483 16235
rect 3065 16133 3099 16167
rect 1777 16065 1811 16099
rect 6377 16065 6411 16099
rect 7481 16065 7515 16099
rect 13001 16065 13035 16099
rect 1593 15997 1627 16031
rect 2329 15997 2363 16031
rect 2881 15997 2915 16031
rect 3433 15997 3467 16031
rect 3985 15997 4019 16031
rect 5181 15997 5215 16031
rect 7849 15997 7883 16031
rect 8401 15997 8435 16031
rect 8668 15997 8702 16031
rect 10057 15997 10091 16031
rect 10324 15997 10358 16031
rect 13461 15997 13495 16031
rect 6101 15929 6135 15963
rect 13706 15929 13740 15963
rect 5733 15861 5767 15895
rect 6193 15861 6227 15895
rect 6837 15861 6871 15895
rect 7205 15861 7239 15895
rect 7297 15861 7331 15895
rect 9781 15861 9815 15895
rect 11437 15861 11471 15895
rect 11713 15861 11747 15895
rect 12817 15861 12851 15895
rect 12909 15861 12943 15895
rect 14841 15861 14875 15895
rect 15117 15861 15151 15895
rect 2421 15657 2455 15691
rect 6561 15657 6595 15691
rect 7021 15657 7055 15691
rect 7481 15657 7515 15691
rect 8033 15657 8067 15691
rect 10149 15657 10183 15691
rect 13645 15657 13679 15691
rect 13921 15657 13955 15691
rect 1777 15589 1811 15623
rect 3433 15589 3467 15623
rect 4988 15589 5022 15623
rect 8401 15589 8435 15623
rect 8493 15589 8527 15623
rect 12532 15589 12566 15623
rect 14381 15589 14415 15623
rect 1501 15521 1535 15555
rect 2237 15521 2271 15555
rect 3341 15521 3375 15555
rect 4721 15521 4755 15555
rect 6377 15521 6411 15555
rect 7389 15521 7423 15555
rect 9045 15521 9079 15555
rect 10057 15521 10091 15555
rect 11069 15521 11103 15555
rect 14289 15521 14323 15555
rect 3525 15453 3559 15487
rect 7573 15453 7607 15487
rect 8585 15453 8619 15487
rect 10241 15453 10275 15487
rect 11161 15453 11195 15487
rect 11345 15453 11379 15487
rect 12265 15453 12299 15487
rect 14473 15453 14507 15487
rect 6101 15385 6135 15419
rect 9229 15385 9263 15419
rect 9689 15385 9723 15419
rect 2973 15317 3007 15351
rect 10701 15317 10735 15351
rect 4077 15113 4111 15147
rect 4353 15113 4387 15147
rect 6377 15113 6411 15147
rect 7481 15113 7515 15147
rect 9873 15113 9907 15147
rect 10149 15113 10183 15147
rect 12449 15113 12483 15147
rect 14473 15113 14507 15147
rect 11161 15045 11195 15079
rect 13461 15045 13495 15079
rect 2329 14977 2363 15011
rect 4905 14977 4939 15011
rect 5917 14977 5951 15011
rect 8033 14977 8067 15011
rect 10609 14977 10643 15011
rect 10701 14977 10735 15011
rect 11713 14977 11747 15011
rect 12909 14977 12943 15011
rect 13001 14977 13035 15011
rect 13921 14977 13955 15011
rect 14105 14977 14139 15011
rect 14933 14977 14967 15011
rect 15025 14977 15059 15011
rect 2697 14909 2731 14943
rect 2964 14909 2998 14943
rect 4813 14909 4847 14943
rect 6561 14909 6595 14943
rect 7849 14909 7883 14943
rect 8309 14909 8343 14943
rect 8493 14909 8527 14943
rect 10517 14909 10551 14943
rect 11529 14909 11563 14943
rect 12817 14909 12851 14943
rect 2053 14841 2087 14875
rect 7021 14841 7055 14875
rect 8760 14841 8794 14875
rect 11621 14841 11655 14875
rect 13829 14841 13863 14875
rect 1685 14773 1719 14807
rect 2145 14773 2179 14807
rect 4721 14773 4755 14807
rect 5365 14773 5399 14807
rect 5733 14773 5767 14807
rect 5825 14773 5859 14807
rect 7941 14773 7975 14807
rect 8309 14773 8343 14807
rect 14841 14773 14875 14807
rect 2881 14569 2915 14603
rect 5825 14569 5859 14603
rect 6285 14569 6319 14603
rect 7573 14569 7607 14603
rect 8585 14569 8619 14603
rect 3433 14501 3467 14535
rect 4414 14501 4448 14535
rect 9045 14501 9079 14535
rect 11345 14501 11379 14535
rect 11796 14501 11830 14535
rect 14013 14501 14047 14535
rect 1501 14433 1535 14467
rect 1768 14433 1802 14467
rect 3157 14433 3191 14467
rect 6193 14433 6227 14467
rect 7941 14433 7975 14467
rect 8953 14433 8987 14467
rect 10140 14433 10174 14467
rect 4169 14365 4203 14399
rect 6377 14365 6411 14399
rect 8033 14365 8067 14399
rect 8217 14365 8251 14399
rect 9137 14365 9171 14399
rect 9873 14365 9907 14399
rect 11529 14365 11563 14399
rect 13921 14365 13955 14399
rect 14197 14365 14231 14399
rect 5549 14297 5583 14331
rect 11253 14297 11287 14331
rect 11345 14297 11379 14331
rect 12909 14229 12943 14263
rect 1961 14025 1995 14059
rect 2973 14025 3007 14059
rect 3985 14025 4019 14059
rect 5549 14025 5583 14059
rect 11253 14025 11287 14059
rect 14887 14025 14921 14059
rect 10425 13957 10459 13991
rect 10701 13957 10735 13991
rect 14473 13957 14507 13991
rect 2605 13889 2639 13923
rect 3433 13889 3467 13923
rect 3525 13889 3559 13923
rect 4537 13889 4571 13923
rect 4997 13889 5031 13923
rect 6009 13889 6043 13923
rect 6193 13889 6227 13923
rect 6837 13889 6871 13923
rect 11805 13889 11839 13923
rect 2329 13821 2363 13855
rect 4445 13821 4479 13855
rect 5917 13821 5951 13855
rect 7093 13821 7127 13855
rect 9045 13821 9079 13855
rect 10885 13821 10919 13855
rect 11713 13821 11747 13855
rect 13093 13821 13127 13855
rect 14816 13821 14850 13855
rect 3341 13753 3375 13787
rect 4353 13753 4387 13787
rect 9312 13753 9346 13787
rect 13360 13753 13394 13787
rect 2421 13685 2455 13719
rect 8217 13685 8251 13719
rect 11621 13685 11655 13719
rect 2697 13481 2731 13515
rect 5089 13481 5123 13515
rect 6009 13481 6043 13515
rect 8953 13481 8987 13515
rect 9321 13481 9355 13515
rect 11713 13481 11747 13515
rect 11989 13481 12023 13515
rect 14013 13481 14047 13515
rect 3065 13413 3099 13447
rect 6101 13413 6135 13447
rect 12357 13413 12391 13447
rect 14473 13413 14507 13447
rect 2053 13345 2087 13379
rect 4997 13345 5031 13379
rect 7481 13345 7515 13379
rect 7840 13345 7874 13379
rect 9505 13345 9539 13379
rect 10333 13345 10367 13379
rect 10600 13345 10634 13379
rect 13369 13345 13403 13379
rect 14381 13345 14415 13379
rect 2145 13277 2179 13311
rect 2237 13277 2271 13311
rect 3157 13277 3191 13311
rect 3249 13277 3283 13311
rect 5273 13277 5307 13311
rect 6285 13277 6319 13311
rect 7573 13277 7607 13311
rect 12449 13277 12483 13311
rect 12541 13277 12575 13311
rect 13461 13277 13495 13311
rect 13553 13277 13587 13311
rect 14565 13277 14599 13311
rect 1685 13209 1719 13243
rect 7297 13209 7331 13243
rect 13001 13209 13035 13243
rect 4629 13141 4663 13175
rect 5641 13141 5675 13175
rect 2145 12937 2179 12971
rect 4537 12937 4571 12971
rect 5365 12937 5399 12971
rect 10885 12937 10919 12971
rect 12449 12937 12483 12971
rect 1593 12801 1627 12835
rect 2605 12801 2639 12835
rect 2789 12801 2823 12835
rect 5825 12801 5859 12835
rect 6009 12801 6043 12835
rect 7389 12801 7423 12835
rect 10425 12801 10459 12835
rect 11529 12801 11563 12835
rect 13001 12801 13035 12835
rect 14381 12801 14415 12835
rect 14565 12801 14599 12835
rect 1409 12733 1443 12767
rect 3157 12733 3191 12767
rect 3413 12733 3447 12767
rect 6561 12733 6595 12767
rect 7297 12733 7331 12767
rect 8033 12733 8067 12767
rect 10241 12733 10275 12767
rect 10333 12733 10367 12767
rect 12909 12733 12943 12767
rect 2513 12665 2547 12699
rect 5733 12665 5767 12699
rect 8300 12665 8334 12699
rect 11253 12665 11287 12699
rect 14289 12665 14323 12699
rect 6377 12597 6411 12631
rect 6837 12597 6871 12631
rect 7205 12597 7239 12631
rect 9413 12597 9447 12631
rect 9873 12597 9907 12631
rect 11345 12597 11379 12631
rect 12817 12597 12851 12631
rect 13921 12597 13955 12631
rect 3341 12393 3375 12427
rect 4537 12393 4571 12427
rect 4997 12393 5031 12427
rect 6469 12393 6503 12427
rect 8125 12393 8159 12427
rect 9689 12393 9723 12427
rect 12541 12393 12575 12427
rect 13185 12393 13219 12427
rect 13553 12393 13587 12427
rect 14197 12393 14231 12427
rect 14565 12393 14599 12427
rect 2228 12257 2262 12291
rect 3893 12257 3927 12291
rect 4445 12257 4479 12291
rect 6990 12325 7024 12359
rect 11130 12325 11164 12359
rect 13645 12325 13679 12359
rect 14657 12325 14691 12359
rect 5089 12257 5123 12291
rect 5356 12257 5390 12291
rect 8861 12257 8895 12291
rect 10057 12257 10091 12291
rect 1961 12189 1995 12223
rect 4721 12189 4755 12223
rect 4997 12189 5031 12223
rect 6745 12189 6779 12223
rect 8217 12189 8251 12223
rect 8953 12189 8987 12223
rect 9045 12189 9079 12223
rect 10149 12189 10183 12223
rect 10333 12189 10367 12223
rect 10885 12189 10919 12223
rect 13737 12189 13771 12223
rect 14749 12189 14783 12223
rect 3709 12121 3743 12155
rect 8493 12121 8527 12155
rect 4077 12053 4111 12087
rect 12265 12053 12299 12087
rect 1869 11849 1903 11883
rect 4261 11849 4295 11883
rect 5733 11849 5767 11883
rect 7757 11849 7791 11883
rect 8677 11849 8711 11883
rect 9689 11849 9723 11883
rect 10701 11849 10735 11883
rect 2513 11713 2547 11747
rect 2881 11713 2915 11747
rect 5273 11713 5307 11747
rect 6285 11713 6319 11747
rect 7481 11713 7515 11747
rect 8401 11713 8435 11747
rect 9229 11713 9263 11747
rect 10241 11713 10275 11747
rect 11161 11713 11195 11747
rect 11253 11713 11287 11747
rect 13185 11713 13219 11747
rect 15117 11713 15151 11747
rect 3148 11645 3182 11679
rect 6193 11645 6227 11679
rect 7297 11645 7331 11679
rect 10149 11645 10183 11679
rect 13001 11645 13035 11679
rect 14841 11645 14875 11679
rect 2237 11577 2271 11611
rect 6101 11577 6135 11611
rect 8125 11577 8159 11611
rect 9137 11577 9171 11611
rect 10057 11577 10091 11611
rect 11069 11577 11103 11611
rect 2329 11509 2363 11543
rect 4629 11509 4663 11543
rect 4997 11509 5031 11543
rect 5089 11509 5123 11543
rect 6929 11509 6963 11543
rect 7389 11509 7423 11543
rect 8217 11509 8251 11543
rect 9045 11509 9079 11543
rect 2789 11305 2823 11339
rect 4629 11305 4663 11339
rect 4813 11305 4847 11339
rect 5181 11305 5215 11339
rect 7205 11305 7239 11339
rect 7573 11305 7607 11339
rect 8585 11305 8619 11339
rect 10425 11305 10459 11339
rect 13093 11305 13127 11339
rect 1676 11237 1710 11271
rect 5273 11237 5307 11271
rect 10793 11237 10827 11271
rect 1409 11169 1443 11203
rect 3065 11169 3099 11203
rect 4077 11169 4111 11203
rect 4629 11169 4663 11203
rect 5825 11169 5859 11203
rect 6092 11169 6126 11203
rect 7941 11169 7975 11203
rect 8953 11169 8987 11203
rect 9045 11169 9079 11203
rect 10333 11169 10367 11203
rect 11713 11169 11747 11203
rect 11980 11169 12014 11203
rect 3249 11101 3283 11135
rect 4261 11101 4295 11135
rect 5457 11101 5491 11135
rect 8033 11101 8067 11135
rect 8217 11101 8251 11135
rect 9229 11101 9263 11135
rect 10885 11101 10919 11135
rect 10977 11101 11011 11135
rect 10149 10965 10183 10999
rect 2237 10761 2271 10795
rect 5641 10761 5675 10795
rect 9045 10761 9079 10795
rect 12081 10761 12115 10795
rect 9689 10693 9723 10727
rect 2881 10625 2915 10659
rect 3893 10625 3927 10659
rect 6101 10625 6135 10659
rect 7205 10625 7239 10659
rect 10333 10625 10367 10659
rect 12633 10625 12667 10659
rect 14841 10625 14875 10659
rect 1501 10557 1535 10591
rect 1777 10557 1811 10591
rect 3617 10557 3651 10591
rect 4261 10557 4295 10591
rect 5917 10557 5951 10591
rect 7665 10557 7699 10591
rect 7932 10557 7966 10591
rect 10701 10557 10735 10591
rect 10968 10557 11002 10591
rect 12900 10557 12934 10591
rect 14749 10557 14783 10591
rect 4528 10489 4562 10523
rect 10057 10489 10091 10523
rect 2605 10421 2639 10455
rect 2697 10421 2731 10455
rect 3249 10421 3283 10455
rect 3709 10421 3743 10455
rect 10149 10421 10183 10455
rect 14013 10421 14047 10455
rect 14289 10421 14323 10455
rect 14657 10421 14691 10455
rect 2237 10217 2271 10251
rect 2697 10217 2731 10251
rect 2881 10217 2915 10251
rect 7113 10217 7147 10251
rect 8769 10217 8803 10251
rect 11345 10217 11379 10251
rect 13829 10217 13863 10251
rect 14381 10217 14415 10251
rect 2329 10149 2363 10183
rect 2513 10013 2547 10047
rect 4905 10149 4939 10183
rect 5978 10149 6012 10183
rect 9137 10149 9171 10183
rect 3249 10081 3283 10115
rect 4813 10081 4847 10115
rect 5733 10081 5767 10115
rect 8309 10081 8343 10115
rect 10221 10081 10255 10115
rect 12357 10081 12391 10115
rect 13737 10081 13771 10115
rect 3341 10013 3375 10047
rect 3433 10013 3467 10047
rect 5089 10013 5123 10047
rect 8401 10013 8435 10047
rect 8585 10013 8619 10047
rect 9229 10013 9263 10047
rect 9321 10013 9355 10047
rect 9965 10013 9999 10047
rect 12449 10013 12483 10047
rect 12633 10013 12667 10047
rect 14013 10013 14047 10047
rect 2789 9945 2823 9979
rect 1869 9877 1903 9911
rect 4445 9877 4479 9911
rect 7941 9877 7975 9911
rect 11989 9877 12023 9911
rect 13369 9877 13403 9911
rect 1777 9605 1811 9639
rect 5457 9605 5491 9639
rect 8769 9605 8803 9639
rect 9321 9605 9355 9639
rect 10149 9605 10183 9639
rect 11345 9605 11379 9639
rect 12449 9605 12483 9639
rect 13461 9605 13495 9639
rect 2421 9537 2455 9571
rect 5089 9537 5123 9571
rect 6561 9537 6595 9571
rect 9873 9537 9907 9571
rect 10701 9537 10735 9571
rect 11989 9537 12023 9571
rect 13093 9537 13127 9571
rect 14013 9537 14047 9571
rect 2145 9469 2179 9503
rect 2789 9469 2823 9503
rect 5641 9469 5675 9503
rect 6285 9469 6319 9503
rect 9781 9469 9815 9503
rect 10609 9469 10643 9503
rect 11713 9469 11747 9503
rect 13829 9469 13863 9503
rect 2237 9401 2271 9435
rect 3056 9401 3090 9435
rect 4905 9401 4939 9435
rect 7481 9401 7515 9435
rect 11805 9401 11839 9435
rect 13921 9401 13955 9435
rect 4169 9333 4203 9367
rect 4445 9333 4479 9367
rect 4813 9333 4847 9367
rect 5917 9333 5951 9367
rect 6377 9333 6411 9367
rect 9689 9333 9723 9367
rect 10517 9333 10551 9367
rect 12817 9333 12851 9367
rect 12909 9333 12943 9367
rect 3525 9129 3559 9163
rect 4077 9129 4111 9163
rect 6377 9129 6411 9163
rect 8493 9129 8527 9163
rect 8861 9129 8895 9163
rect 9689 9129 9723 9163
rect 12449 9129 12483 9163
rect 13921 9129 13955 9163
rect 5242 9061 5276 9095
rect 10057 9061 10091 9095
rect 12909 9061 12943 9095
rect 1409 8993 1443 9027
rect 1685 8993 1719 9027
rect 2145 8993 2179 9027
rect 2412 8993 2446 9027
rect 4537 8993 4571 9027
rect 6920 8993 6954 9027
rect 10968 8993 11002 9027
rect 12817 8993 12851 9027
rect 13829 8993 13863 9027
rect 4997 8925 5031 8959
rect 6653 8925 6687 8959
rect 8953 8925 8987 8959
rect 9137 8925 9171 8959
rect 10149 8925 10183 8959
rect 10241 8925 10275 8959
rect 10701 8925 10735 8959
rect 13093 8925 13127 8959
rect 14013 8925 14047 8959
rect 8033 8857 8067 8891
rect 12081 8857 12115 8891
rect 13461 8857 13495 8891
rect 5733 8585 5767 8619
rect 8585 8585 8619 8619
rect 14197 8585 14231 8619
rect 2789 8517 2823 8551
rect 8309 8517 8343 8551
rect 9689 8517 9723 8551
rect 2421 8449 2455 8483
rect 3341 8449 3375 8483
rect 4353 8449 4387 8483
rect 5457 8449 5491 8483
rect 6193 8449 6227 8483
rect 6377 8449 6411 8483
rect 6929 8449 6963 8483
rect 9137 8449 9171 8483
rect 9965 8449 9999 8483
rect 11621 8449 11655 8483
rect 2145 8381 2179 8415
rect 3249 8381 3283 8415
rect 4169 8381 4203 8415
rect 5181 8381 5215 8415
rect 7196 8381 7230 8415
rect 9873 8381 9907 8415
rect 12817 8381 12851 8415
rect 2237 8313 2271 8347
rect 3157 8313 3191 8347
rect 5273 8313 5307 8347
rect 6101 8313 6135 8347
rect 9045 8313 9079 8347
rect 10232 8313 10266 8347
rect 13084 8313 13118 8347
rect 1777 8245 1811 8279
rect 3801 8245 3835 8279
rect 4261 8245 4295 8279
rect 4813 8245 4847 8279
rect 8953 8245 8987 8279
rect 11345 8245 11379 8279
rect 2973 8041 3007 8075
rect 3341 8041 3375 8075
rect 4169 8041 4203 8075
rect 4537 8041 4571 8075
rect 6561 8041 6595 8075
rect 6837 8041 6871 8075
rect 8585 8041 8619 8075
rect 10057 8041 10091 8075
rect 10701 8041 10735 8075
rect 12173 8041 12207 8075
rect 12725 8041 12759 8075
rect 2513 7973 2547 8007
rect 3433 7973 3467 8007
rect 10149 7973 10183 8007
rect 11161 7973 11195 8007
rect 13185 7973 13219 8007
rect 1501 7905 1535 7939
rect 2237 7905 2271 7939
rect 4629 7905 4663 7939
rect 5448 7905 5482 7939
rect 7205 7905 7239 7939
rect 8953 7905 8987 7939
rect 11069 7905 11103 7939
rect 12081 7905 12115 7939
rect 13093 7905 13127 7939
rect 1685 7837 1719 7871
rect 3525 7837 3559 7871
rect 4813 7837 4847 7871
rect 5181 7837 5215 7871
rect 7297 7837 7331 7871
rect 7389 7837 7423 7871
rect 9045 7837 9079 7871
rect 9137 7837 9171 7871
rect 10241 7837 10275 7871
rect 11253 7837 11287 7871
rect 12265 7837 12299 7871
rect 13277 7837 13311 7871
rect 11713 7769 11747 7803
rect 9689 7701 9723 7735
rect 4537 7497 4571 7531
rect 5549 7497 5583 7531
rect 6837 7497 6871 7531
rect 10057 7497 10091 7531
rect 11069 7497 11103 7531
rect 4261 7429 4295 7463
rect 9689 7429 9723 7463
rect 2513 7361 2547 7395
rect 2697 7361 2731 7395
rect 5089 7361 5123 7395
rect 6193 7361 6227 7395
rect 7389 7361 7423 7395
rect 10609 7361 10643 7395
rect 11713 7361 11747 7395
rect 13093 7361 13127 7395
rect 2237 7293 2271 7327
rect 2881 7293 2915 7327
rect 6009 7293 6043 7327
rect 8033 7293 8067 7327
rect 8309 7293 8343 7327
rect 10517 7293 10551 7327
rect 11437 7293 11471 7327
rect 12909 7293 12943 7327
rect 2697 7225 2731 7259
rect 3126 7225 3160 7259
rect 4905 7225 4939 7259
rect 7297 7225 7331 7259
rect 8576 7225 8610 7259
rect 1869 7157 1903 7191
rect 2329 7157 2363 7191
rect 4997 7157 5031 7191
rect 5917 7157 5951 7191
rect 7205 7157 7239 7191
rect 7849 7157 7883 7191
rect 10425 7157 10459 7191
rect 11529 7157 11563 7191
rect 12449 7157 12483 7191
rect 12817 7157 12851 7191
rect 3065 6953 3099 6987
rect 4813 6953 4847 6987
rect 9137 6953 9171 6987
rect 9689 6953 9723 6987
rect 12633 6953 12667 6987
rect 5181 6885 5215 6919
rect 10057 6885 10091 6919
rect 11520 6885 11554 6919
rect 1952 6817 1986 6851
rect 4721 6817 4755 6851
rect 5273 6817 5307 6851
rect 6009 6817 6043 6851
rect 7113 6817 7147 6851
rect 7757 6817 7791 6851
rect 8024 6817 8058 6851
rect 10149 6817 10183 6851
rect 10517 6817 10551 6851
rect 10885 6817 10919 6851
rect 11253 6817 11287 6851
rect 13277 6817 13311 6851
rect 13369 6817 13403 6851
rect 1685 6749 1719 6783
rect 5365 6749 5399 6783
rect 7205 6749 7239 6783
rect 7389 6749 7423 6783
rect 10241 6749 10275 6783
rect 13461 6749 13495 6783
rect 4537 6613 4571 6647
rect 6193 6613 6227 6647
rect 6745 6613 6779 6647
rect 10517 6613 10551 6647
rect 10701 6613 10735 6647
rect 12909 6613 12943 6647
rect 3065 6409 3099 6443
rect 4537 6409 4571 6443
rect 8493 6409 8527 6443
rect 11345 6409 11379 6443
rect 8217 6341 8251 6375
rect 10885 6341 10919 6375
rect 3893 6273 3927 6307
rect 5089 6273 5123 6307
rect 6193 6273 6227 6307
rect 6377 6273 6411 6307
rect 9137 6273 9171 6307
rect 9505 6273 9539 6307
rect 11897 6273 11931 6307
rect 12449 6273 12483 6307
rect 1685 6205 1719 6239
rect 6101 6205 6135 6239
rect 6837 6205 6871 6239
rect 9772 6205 9806 6239
rect 11805 6205 11839 6239
rect 1952 6137 1986 6171
rect 3709 6137 3743 6171
rect 4997 6137 5031 6171
rect 7104 6137 7138 6171
rect 8953 6137 8987 6171
rect 11713 6137 11747 6171
rect 3341 6069 3375 6103
rect 3801 6069 3835 6103
rect 4905 6069 4939 6103
rect 5733 6069 5767 6103
rect 8861 6069 8895 6103
rect 4077 5865 4111 5899
rect 4445 5865 4479 5899
rect 4537 5865 4571 5899
rect 6929 5865 6963 5899
rect 1685 5797 1719 5831
rect 2513 5797 2547 5831
rect 5540 5797 5574 5831
rect 14749 5797 14783 5831
rect 1409 5729 1443 5763
rect 3433 5729 3467 5763
rect 5273 5729 5307 5763
rect 7757 5729 7791 5763
rect 7849 5729 7883 5763
rect 8401 5729 8435 5763
rect 8953 5729 8987 5763
rect 10333 5729 10367 5763
rect 13369 5729 13403 5763
rect 14473 5729 14507 5763
rect 2605 5661 2639 5695
rect 2697 5661 2731 5695
rect 4629 5661 4663 5695
rect 8033 5661 8067 5695
rect 10425 5661 10459 5695
rect 10609 5661 10643 5695
rect 13461 5661 13495 5695
rect 13645 5661 13679 5695
rect 8585 5593 8619 5627
rect 13001 5593 13035 5627
rect 2145 5525 2179 5559
rect 3617 5525 3651 5559
rect 6653 5525 6687 5559
rect 7389 5525 7423 5559
rect 9137 5525 9171 5559
rect 9965 5525 9999 5559
rect 5273 5321 5307 5355
rect 9689 5321 9723 5355
rect 12081 5321 12115 5355
rect 12265 5321 12299 5355
rect 13829 5321 13863 5355
rect 2605 5185 2639 5219
rect 2697 5185 2731 5219
rect 6377 5185 6411 5219
rect 6837 5185 6871 5219
rect 7941 5185 7975 5219
rect 1593 5117 1627 5151
rect 3157 5117 3191 5151
rect 3893 5117 3927 5151
rect 4149 5117 4183 5151
rect 6101 5117 6135 5151
rect 7665 5117 7699 5151
rect 8125 5117 8159 5151
rect 8309 5117 8343 5151
rect 9965 5117 9999 5151
rect 10701 5117 10735 5151
rect 6193 5049 6227 5083
rect 8576 5049 8610 5083
rect 10946 5049 10980 5083
rect 14749 5185 14783 5219
rect 12449 5117 12483 5151
rect 14565 5117 14599 5151
rect 12694 5049 12728 5083
rect 1777 4981 1811 5015
rect 2145 4981 2179 5015
rect 2513 4981 2547 5015
rect 3341 4981 3375 5015
rect 5733 4981 5767 5015
rect 7297 4981 7331 5015
rect 7757 4981 7791 5015
rect 8125 4981 8159 5015
rect 10149 4981 10183 5015
rect 12265 4981 12299 5015
rect 14105 4981 14139 5015
rect 14473 4981 14507 5015
rect 1869 4777 1903 4811
rect 2329 4777 2363 4811
rect 2881 4777 2915 4811
rect 3249 4777 3283 4811
rect 7573 4777 7607 4811
rect 8953 4777 8987 4811
rect 13921 4777 13955 4811
rect 14565 4777 14599 4811
rect 2237 4709 2271 4743
rect 6092 4709 6126 4743
rect 8033 4709 8067 4743
rect 9045 4709 9079 4743
rect 10508 4709 10542 4743
rect 14657 4709 14691 4743
rect 3341 4641 3375 4675
rect 4077 4641 4111 4675
rect 4629 4641 4663 4675
rect 5181 4641 5215 4675
rect 5825 4641 5859 4675
rect 7941 4641 7975 4675
rect 9689 4641 9723 4675
rect 12808 4641 12842 4675
rect 2421 4573 2455 4607
rect 3525 4573 3559 4607
rect 8217 4573 8251 4607
rect 9229 4573 9263 4607
rect 10241 4573 10275 4607
rect 12541 4573 12575 4607
rect 14749 4573 14783 4607
rect 5365 4505 5399 4539
rect 9873 4505 9907 4539
rect 11621 4505 11655 4539
rect 4261 4437 4295 4471
rect 4813 4437 4847 4471
rect 7205 4437 7239 4471
rect 8585 4437 8619 4471
rect 14197 4437 14231 4471
rect 4353 4233 4387 4267
rect 9229 4233 9263 4267
rect 9505 4233 9539 4267
rect 9781 4233 9815 4267
rect 1685 4097 1719 4131
rect 5273 4097 5307 4131
rect 6193 4097 6227 4131
rect 6377 4097 6411 4131
rect 10425 4097 10459 4131
rect 11989 4097 12023 4131
rect 13093 4097 13127 4131
rect 14013 4097 14047 4131
rect 14473 4097 14507 4131
rect 1501 4029 1535 4063
rect 2237 4029 2271 4063
rect 2513 4029 2547 4063
rect 2973 4029 3007 4063
rect 6101 4029 6135 4063
rect 6837 4029 6871 4063
rect 7849 4029 7883 4063
rect 9689 4029 9723 4063
rect 10793 4029 10827 4063
rect 13921 4029 13955 4063
rect 3240 3961 3274 3995
rect 5089 3961 5123 3995
rect 8116 3961 8150 3995
rect 13829 3961 13863 3995
rect 4721 3893 4755 3927
rect 5181 3893 5215 3927
rect 5733 3893 5767 3927
rect 7021 3893 7055 3927
rect 10149 3893 10183 3927
rect 10241 3893 10275 3927
rect 10977 3893 11011 3927
rect 11345 3893 11379 3927
rect 11713 3893 11747 3927
rect 11805 3893 11839 3927
rect 12449 3893 12483 3927
rect 12817 3893 12851 3927
rect 12909 3893 12943 3927
rect 13461 3893 13495 3927
rect 9045 3689 9079 3723
rect 10333 3689 10367 3723
rect 11437 3689 11471 3723
rect 11805 3689 11839 3723
rect 12909 3689 12943 3723
rect 13921 3689 13955 3723
rect 2228 3621 2262 3655
rect 6736 3621 6770 3655
rect 13829 3621 13863 3655
rect 1409 3553 1443 3587
rect 1961 3553 1995 3587
rect 3893 3553 3927 3587
rect 4620 3553 4654 3587
rect 8953 3553 8987 3587
rect 12817 3553 12851 3587
rect 4353 3485 4387 3519
rect 6469 3485 6503 3519
rect 9229 3485 9263 3519
rect 10425 3485 10459 3519
rect 10609 3485 10643 3519
rect 11897 3485 11931 3519
rect 12081 3485 12115 3519
rect 13093 3485 13127 3519
rect 14013 3485 14047 3519
rect 3709 3417 3743 3451
rect 5733 3417 5767 3451
rect 12449 3417 12483 3451
rect 1593 3349 1627 3383
rect 3341 3349 3375 3383
rect 7849 3349 7883 3383
rect 8585 3349 8619 3383
rect 9965 3349 9999 3383
rect 13461 3349 13495 3383
rect 2237 3145 2271 3179
rect 5733 3145 5767 3179
rect 9321 3145 9355 3179
rect 10977 3145 11011 3179
rect 11345 3145 11379 3179
rect 14289 3145 14323 3179
rect 1685 3009 1719 3043
rect 2697 3009 2731 3043
rect 2881 3009 2915 3043
rect 3801 3009 3835 3043
rect 4905 3009 4939 3043
rect 6377 3009 6411 3043
rect 7389 3009 7423 3043
rect 7941 3009 7975 3043
rect 9597 3009 9631 3043
rect 11897 3009 11931 3043
rect 12449 3009 12483 3043
rect 12909 3009 12943 3043
rect 1501 2941 1535 2975
rect 4629 2941 4663 2975
rect 8208 2941 8242 2975
rect 14841 2941 14875 2975
rect 2605 2873 2639 2907
rect 3617 2873 3651 2907
rect 7205 2873 7239 2907
rect 7297 2873 7331 2907
rect 9864 2873 9898 2907
rect 11713 2873 11747 2907
rect 13176 2873 13210 2907
rect 15117 2873 15151 2907
rect 3249 2805 3283 2839
rect 3709 2805 3743 2839
rect 4261 2805 4295 2839
rect 4721 2805 4755 2839
rect 5273 2805 5307 2839
rect 6101 2805 6135 2839
rect 6193 2805 6227 2839
rect 6837 2805 6871 2839
rect 11805 2805 11839 2839
rect 4353 2601 4387 2635
rect 4813 2601 4847 2635
rect 5457 2601 5491 2635
rect 5917 2601 5951 2635
rect 7113 2601 7147 2635
rect 8033 2601 8067 2635
rect 8677 2601 8711 2635
rect 9781 2601 9815 2635
rect 10241 2601 10275 2635
rect 12081 2601 12115 2635
rect 12633 2601 12667 2635
rect 13093 2601 13127 2635
rect 13829 2601 13863 2635
rect 14381 2601 14415 2635
rect 4721 2533 4755 2567
rect 9045 2533 9079 2567
rect 10149 2533 10183 2567
rect 11345 2533 11379 2567
rect 1501 2465 1535 2499
rect 2053 2465 2087 2499
rect 2320 2465 2354 2499
rect 5825 2465 5859 2499
rect 6929 2465 6963 2499
rect 8125 2465 8159 2499
rect 11253 2465 11287 2499
rect 11897 2465 11931 2499
rect 13001 2465 13035 2499
rect 13645 2465 13679 2499
rect 14197 2465 14231 2499
rect 14749 2465 14783 2499
rect 4997 2397 5031 2431
rect 6101 2397 6135 2431
rect 8217 2397 8251 2431
rect 9137 2397 9171 2431
rect 9321 2397 9355 2431
rect 10425 2397 10459 2431
rect 11529 2397 11563 2431
rect 13185 2397 13219 2431
rect 7665 2329 7699 2363
rect 10885 2329 10919 2363
rect 1685 2261 1719 2295
rect 3433 2261 3467 2295
rect 14933 2261 14967 2295
<< metal1 >>
rect 4062 17960 4068 18012
rect 4120 18000 4126 18012
rect 14090 18000 14096 18012
rect 4120 17972 14096 18000
rect 4120 17960 4126 17972
rect 14090 17960 14096 17972
rect 14148 17960 14154 18012
rect 8938 17620 8944 17672
rect 8996 17660 9002 17672
rect 9490 17660 9496 17672
rect 8996 17632 9496 17660
rect 8996 17620 9002 17632
rect 9490 17620 9496 17632
rect 9548 17620 9554 17672
rect 5350 17552 5356 17604
rect 5408 17592 5414 17604
rect 11514 17592 11520 17604
rect 5408 17564 11520 17592
rect 5408 17552 5414 17564
rect 11514 17552 11520 17564
rect 11572 17552 11578 17604
rect 198 17484 204 17536
rect 256 17524 262 17536
rect 14182 17524 14188 17536
rect 256 17496 14188 17524
rect 256 17484 262 17496
rect 14182 17484 14188 17496
rect 14240 17484 14246 17536
rect 1104 17434 15824 17456
rect 1104 17382 3447 17434
rect 3499 17382 3511 17434
rect 3563 17382 3575 17434
rect 3627 17382 3639 17434
rect 3691 17382 8378 17434
rect 8430 17382 8442 17434
rect 8494 17382 8506 17434
rect 8558 17382 8570 17434
rect 8622 17382 13308 17434
rect 13360 17382 13372 17434
rect 13424 17382 13436 17434
rect 13488 17382 13500 17434
rect 13552 17382 15824 17434
rect 1104 17360 15824 17382
rect 2774 17280 2780 17332
rect 2832 17320 2838 17332
rect 3053 17323 3111 17329
rect 3053 17320 3065 17323
rect 2832 17292 3065 17320
rect 2832 17280 2838 17292
rect 3053 17289 3065 17292
rect 3099 17289 3111 17323
rect 3053 17283 3111 17289
rect 4614 17280 4620 17332
rect 4672 17320 4678 17332
rect 4985 17323 5043 17329
rect 4985 17320 4997 17323
rect 4672 17292 4997 17320
rect 4672 17280 4678 17292
rect 4985 17289 4997 17292
rect 5031 17289 5043 17323
rect 4985 17283 5043 17289
rect 5074 17280 5080 17332
rect 5132 17320 5138 17332
rect 5537 17323 5595 17329
rect 5537 17320 5549 17323
rect 5132 17292 5549 17320
rect 5132 17280 5138 17292
rect 5537 17289 5549 17292
rect 5583 17289 5595 17323
rect 5537 17283 5595 17289
rect 5626 17280 5632 17332
rect 5684 17320 5690 17332
rect 6089 17323 6147 17329
rect 6089 17320 6101 17323
rect 5684 17292 6101 17320
rect 5684 17280 5690 17292
rect 6089 17289 6101 17292
rect 6135 17289 6147 17323
rect 6089 17283 6147 17289
rect 7834 17280 7840 17332
rect 7892 17320 7898 17332
rect 9953 17323 10011 17329
rect 9953 17320 9965 17323
rect 7892 17292 9965 17320
rect 7892 17280 7898 17292
rect 9953 17289 9965 17292
rect 9999 17289 10011 17323
rect 12710 17320 12716 17332
rect 9953 17283 10011 17289
rect 10060 17292 12716 17320
rect 1765 17255 1823 17261
rect 1765 17221 1777 17255
rect 1811 17252 1823 17255
rect 2866 17252 2872 17264
rect 1811 17224 2872 17252
rect 1811 17221 1823 17224
rect 1765 17215 1823 17221
rect 2866 17212 2872 17224
rect 2924 17212 2930 17264
rect 2958 17212 2964 17264
rect 3016 17252 3022 17264
rect 3605 17255 3663 17261
rect 3605 17252 3617 17255
rect 3016 17224 3617 17252
rect 3016 17212 3022 17224
rect 3605 17221 3617 17224
rect 3651 17221 3663 17255
rect 3605 17215 3663 17221
rect 5810 17212 5816 17264
rect 5868 17252 5874 17264
rect 7101 17255 7159 17261
rect 7101 17252 7113 17255
rect 5868 17224 7113 17252
rect 5868 17212 5874 17224
rect 7101 17221 7113 17224
rect 7147 17221 7159 17255
rect 10060 17252 10088 17292
rect 12710 17280 12716 17292
rect 12768 17280 12774 17332
rect 7101 17215 7159 17221
rect 8036 17224 10088 17252
rect 10689 17255 10747 17261
rect 1578 17116 1584 17128
rect 1539 17088 1584 17116
rect 1578 17076 1584 17088
rect 1636 17076 1642 17128
rect 2869 17119 2927 17125
rect 2869 17085 2881 17119
rect 2915 17085 2927 17119
rect 2869 17079 2927 17085
rect 3421 17119 3479 17125
rect 3421 17085 3433 17119
rect 3467 17116 3479 17119
rect 3878 17116 3884 17128
rect 3467 17088 3884 17116
rect 3467 17085 3479 17088
rect 3421 17079 3479 17085
rect 2884 17048 2912 17079
rect 3878 17076 3884 17088
rect 3936 17076 3942 17128
rect 4801 17119 4859 17125
rect 4801 17085 4813 17119
rect 4847 17085 4859 17119
rect 5350 17116 5356 17128
rect 5311 17088 5356 17116
rect 4801 17079 4859 17085
rect 4154 17048 4160 17060
rect 2884 17020 4160 17048
rect 4154 17008 4160 17020
rect 4212 17008 4218 17060
rect 4816 17048 4844 17079
rect 5350 17076 5356 17088
rect 5408 17076 5414 17128
rect 5905 17119 5963 17125
rect 5905 17085 5917 17119
rect 5951 17116 5963 17119
rect 6822 17116 6828 17128
rect 5951 17088 6828 17116
rect 5951 17085 5963 17088
rect 5905 17079 5963 17085
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 8036 17125 8064 17224
rect 10689 17221 10701 17255
rect 10735 17252 10747 17255
rect 13722 17252 13728 17264
rect 10735 17224 13728 17252
rect 10735 17221 10747 17224
rect 10689 17215 10747 17221
rect 13722 17212 13728 17224
rect 13780 17212 13786 17264
rect 8205 17187 8263 17193
rect 8205 17153 8217 17187
rect 8251 17153 8263 17187
rect 8205 17147 8263 17153
rect 6917 17119 6975 17125
rect 6917 17085 6929 17119
rect 6963 17085 6975 17119
rect 6917 17079 6975 17085
rect 8021 17119 8079 17125
rect 8021 17085 8033 17119
rect 8067 17085 8079 17119
rect 8220 17116 8248 17147
rect 8386 17144 8392 17196
rect 8444 17184 8450 17196
rect 9217 17187 9275 17193
rect 9217 17184 9229 17187
rect 8444 17156 9229 17184
rect 8444 17144 8450 17156
rect 9217 17153 9229 17156
rect 9263 17153 9275 17187
rect 11238 17184 11244 17196
rect 9217 17147 9275 17153
rect 9324 17156 11244 17184
rect 9324 17116 9352 17156
rect 11238 17144 11244 17156
rect 11296 17144 11302 17196
rect 11333 17187 11391 17193
rect 11333 17153 11345 17187
rect 11379 17184 11391 17187
rect 11606 17184 11612 17196
rect 11379 17156 11612 17184
rect 11379 17153 11391 17156
rect 11333 17147 11391 17153
rect 11606 17144 11612 17156
rect 11664 17144 11670 17196
rect 13170 17184 13176 17196
rect 13131 17156 13176 17184
rect 13170 17144 13176 17156
rect 13228 17144 13234 17196
rect 14090 17184 14096 17196
rect 14051 17156 14096 17184
rect 14090 17144 14096 17156
rect 14148 17144 14154 17196
rect 15102 17184 15108 17196
rect 15063 17156 15108 17184
rect 15102 17144 15108 17156
rect 15160 17144 15166 17196
rect 8220 17088 9352 17116
rect 9769 17119 9827 17125
rect 8021 17079 8079 17085
rect 9769 17085 9781 17119
rect 9815 17116 9827 17119
rect 10226 17116 10232 17128
rect 9815 17088 10232 17116
rect 9815 17085 9827 17088
rect 9769 17079 9827 17085
rect 6546 17048 6552 17060
rect 4816 17020 6552 17048
rect 6546 17008 6552 17020
rect 6604 17008 6610 17060
rect 6932 17048 6960 17079
rect 10226 17076 10232 17088
rect 10284 17076 10290 17128
rect 11057 17119 11115 17125
rect 11057 17085 11069 17119
rect 11103 17116 11115 17119
rect 12434 17116 12440 17128
rect 11103 17088 12440 17116
rect 11103 17085 11115 17088
rect 11057 17079 11115 17085
rect 12434 17076 12440 17088
rect 12492 17076 12498 17128
rect 8113 17051 8171 17057
rect 6932 17020 8064 17048
rect 2866 16940 2872 16992
rect 2924 16980 2930 16992
rect 7653 16983 7711 16989
rect 7653 16980 7665 16983
rect 2924 16952 7665 16980
rect 2924 16940 2930 16952
rect 7653 16949 7665 16952
rect 7699 16949 7711 16983
rect 8036 16980 8064 17020
rect 8113 17017 8125 17051
rect 8159 17048 8171 17051
rect 14185 17051 14243 17057
rect 8159 17020 12664 17048
rect 8159 17017 8171 17020
rect 8113 17011 8171 17017
rect 8294 16980 8300 16992
rect 8036 16952 8300 16980
rect 7653 16943 7711 16949
rect 8294 16940 8300 16952
rect 8352 16940 8358 16992
rect 8662 16980 8668 16992
rect 8623 16952 8668 16980
rect 8662 16940 8668 16952
rect 8720 16940 8726 16992
rect 9030 16980 9036 16992
rect 8991 16952 9036 16980
rect 9030 16940 9036 16952
rect 9088 16940 9094 16992
rect 9122 16940 9128 16992
rect 9180 16980 9186 16992
rect 9180 16952 9225 16980
rect 9180 16940 9186 16952
rect 11146 16940 11152 16992
rect 11204 16980 11210 16992
rect 12636 16989 12664 17020
rect 14185 17017 14197 17051
rect 14231 17048 14243 17051
rect 15010 17048 15016 17060
rect 14231 17020 15016 17048
rect 14231 17017 14243 17020
rect 14185 17011 14243 17017
rect 15010 17008 15016 17020
rect 15068 17008 15074 17060
rect 12621 16983 12679 16989
rect 11204 16952 11249 16980
rect 11204 16940 11210 16952
rect 12621 16949 12633 16983
rect 12667 16949 12679 16983
rect 12986 16980 12992 16992
rect 12947 16952 12992 16980
rect 12621 16943 12679 16949
rect 12986 16940 12992 16952
rect 13044 16940 13050 16992
rect 13081 16983 13139 16989
rect 13081 16949 13093 16983
rect 13127 16980 13139 16983
rect 13906 16980 13912 16992
rect 13127 16952 13912 16980
rect 13127 16949 13139 16952
rect 13081 16943 13139 16949
rect 13906 16940 13912 16952
rect 13964 16940 13970 16992
rect 1104 16890 15824 16912
rect 1104 16838 5912 16890
rect 5964 16838 5976 16890
rect 6028 16838 6040 16890
rect 6092 16838 6104 16890
rect 6156 16838 10843 16890
rect 10895 16838 10907 16890
rect 10959 16838 10971 16890
rect 11023 16838 11035 16890
rect 11087 16838 15824 16890
rect 1104 16816 15824 16838
rect 934 16736 940 16788
rect 992 16776 998 16788
rect 1765 16779 1823 16785
rect 1765 16776 1777 16779
rect 992 16748 1777 16776
rect 992 16736 998 16748
rect 1765 16745 1777 16748
rect 1811 16745 1823 16779
rect 1765 16739 1823 16745
rect 2317 16779 2375 16785
rect 2317 16745 2329 16779
rect 2363 16745 2375 16779
rect 2317 16739 2375 16745
rect 1394 16668 1400 16720
rect 1452 16708 1458 16720
rect 2332 16708 2360 16739
rect 4246 16736 4252 16788
rect 4304 16776 4310 16788
rect 4525 16779 4583 16785
rect 4525 16776 4537 16779
rect 4304 16748 4537 16776
rect 4304 16736 4310 16748
rect 4525 16745 4537 16748
rect 4571 16745 4583 16779
rect 4525 16739 4583 16745
rect 6733 16779 6791 16785
rect 6733 16745 6745 16779
rect 6779 16745 6791 16779
rect 8386 16776 8392 16788
rect 8347 16748 8392 16776
rect 6733 16739 6791 16745
rect 3142 16708 3148 16720
rect 1452 16680 2360 16708
rect 3103 16680 3148 16708
rect 1452 16668 1458 16680
rect 3142 16668 3148 16680
rect 3200 16668 3206 16720
rect 5620 16711 5678 16717
rect 5620 16677 5632 16711
rect 5666 16708 5678 16711
rect 5718 16708 5724 16720
rect 5666 16680 5724 16708
rect 5666 16677 5678 16680
rect 5620 16671 5678 16677
rect 5718 16668 5724 16680
rect 5776 16668 5782 16720
rect 6362 16668 6368 16720
rect 6420 16708 6426 16720
rect 6748 16708 6776 16739
rect 8386 16736 8392 16748
rect 8444 16736 8450 16788
rect 8662 16736 8668 16788
rect 8720 16776 8726 16788
rect 10137 16779 10195 16785
rect 10137 16776 10149 16779
rect 8720 16748 10149 16776
rect 8720 16736 8726 16748
rect 10137 16745 10149 16748
rect 10183 16745 10195 16779
rect 10137 16739 10195 16745
rect 11057 16779 11115 16785
rect 11057 16745 11069 16779
rect 11103 16776 11115 16779
rect 11146 16776 11152 16788
rect 11103 16748 11152 16776
rect 11103 16745 11115 16748
rect 11057 16739 11115 16745
rect 11146 16736 11152 16748
rect 11204 16736 11210 16788
rect 11517 16779 11575 16785
rect 11517 16745 11529 16779
rect 11563 16776 11575 16779
rect 12618 16776 12624 16788
rect 11563 16748 12624 16776
rect 11563 16745 11575 16748
rect 11517 16739 11575 16745
rect 12618 16736 12624 16748
rect 12676 16776 12682 16788
rect 13078 16776 13084 16788
rect 12676 16748 13084 16776
rect 12676 16736 12682 16748
rect 13078 16736 13084 16748
rect 13136 16736 13142 16788
rect 13170 16736 13176 16788
rect 13228 16776 13234 16788
rect 13725 16779 13783 16785
rect 13725 16776 13737 16779
rect 13228 16748 13737 16776
rect 13228 16736 13234 16748
rect 13725 16745 13737 16748
rect 13771 16745 13783 16779
rect 13725 16739 13783 16745
rect 7254 16711 7312 16717
rect 7254 16708 7266 16711
rect 6420 16680 7266 16708
rect 6420 16668 6426 16680
rect 7254 16677 7266 16680
rect 7300 16677 7312 16711
rect 7254 16671 7312 16677
rect 8294 16668 8300 16720
rect 8352 16708 8358 16720
rect 9490 16708 9496 16720
rect 8352 16680 9496 16708
rect 8352 16668 8358 16680
rect 9490 16668 9496 16680
rect 9548 16668 9554 16720
rect 11790 16708 11796 16720
rect 9968 16680 11796 16708
rect 1581 16643 1639 16649
rect 1581 16609 1593 16643
rect 1627 16640 1639 16643
rect 1670 16640 1676 16652
rect 1627 16612 1676 16640
rect 1627 16609 1639 16612
rect 1581 16603 1639 16609
rect 1670 16600 1676 16612
rect 1728 16600 1734 16652
rect 2133 16643 2191 16649
rect 2133 16609 2145 16643
rect 2179 16640 2191 16643
rect 2498 16640 2504 16652
rect 2179 16612 2504 16640
rect 2179 16609 2191 16612
rect 2133 16603 2191 16609
rect 2498 16600 2504 16612
rect 2556 16600 2562 16652
rect 2866 16640 2872 16652
rect 2827 16612 2872 16640
rect 2866 16600 2872 16612
rect 2924 16600 2930 16652
rect 4341 16643 4399 16649
rect 4341 16609 4353 16643
rect 4387 16640 4399 16643
rect 6730 16640 6736 16652
rect 4387 16612 6736 16640
rect 4387 16609 4399 16612
rect 4341 16603 4399 16609
rect 6730 16600 6736 16612
rect 6788 16600 6794 16652
rect 7009 16643 7067 16649
rect 7009 16640 7021 16643
rect 6840 16612 7021 16640
rect 5353 16575 5411 16581
rect 5353 16541 5365 16575
rect 5399 16541 5411 16575
rect 5353 16535 5411 16541
rect 5368 16448 5396 16535
rect 5350 16436 5356 16448
rect 5263 16408 5356 16436
rect 5350 16396 5356 16408
rect 5408 16436 5414 16448
rect 6840 16436 6868 16612
rect 7009 16609 7021 16612
rect 7055 16609 7067 16643
rect 7009 16603 7067 16609
rect 8665 16643 8723 16649
rect 8665 16609 8677 16643
rect 8711 16640 8723 16643
rect 9968 16640 9996 16680
rect 11790 16668 11796 16680
rect 11848 16668 11854 16720
rect 8711 16612 9996 16640
rect 10045 16643 10103 16649
rect 8711 16609 8723 16612
rect 8665 16603 8723 16609
rect 10045 16609 10057 16643
rect 10091 16609 10103 16643
rect 11422 16640 11428 16652
rect 11383 16612 11428 16640
rect 10045 16603 10103 16609
rect 8110 16532 8116 16584
rect 8168 16572 8174 16584
rect 8168 16544 9536 16572
rect 8168 16532 8174 16544
rect 8018 16464 8024 16516
rect 8076 16504 8082 16516
rect 8938 16504 8944 16516
rect 8076 16476 8944 16504
rect 8076 16464 8082 16476
rect 8938 16464 8944 16476
rect 8996 16464 9002 16516
rect 9508 16504 9536 16544
rect 9582 16532 9588 16584
rect 9640 16572 9646 16584
rect 10060 16572 10088 16603
rect 11422 16600 11428 16612
rect 11480 16600 11486 16652
rect 12612 16643 12670 16649
rect 12612 16609 12624 16643
rect 12658 16640 12670 16643
rect 13998 16640 14004 16652
rect 12658 16612 14004 16640
rect 12658 16609 12670 16612
rect 12612 16603 12670 16609
rect 13998 16600 14004 16612
rect 14056 16600 14062 16652
rect 14182 16640 14188 16652
rect 14143 16612 14188 16640
rect 14182 16600 14188 16612
rect 14240 16600 14246 16652
rect 14553 16643 14611 16649
rect 14553 16609 14565 16643
rect 14599 16640 14611 16643
rect 14826 16640 14832 16652
rect 14599 16612 14832 16640
rect 14599 16609 14611 16612
rect 14553 16603 14611 16609
rect 14826 16600 14832 16612
rect 14884 16600 14890 16652
rect 9640 16544 10088 16572
rect 10321 16575 10379 16581
rect 9640 16532 9646 16544
rect 10321 16541 10333 16575
rect 10367 16572 10379 16575
rect 11698 16572 11704 16584
rect 10367 16544 11704 16572
rect 10367 16541 10379 16544
rect 10321 16535 10379 16541
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 11974 16532 11980 16584
rect 12032 16572 12038 16584
rect 12345 16575 12403 16581
rect 12345 16572 12357 16575
rect 12032 16544 12357 16572
rect 12032 16532 12038 16544
rect 12345 16541 12357 16544
rect 12391 16541 12403 16575
rect 12345 16535 12403 16541
rect 14921 16575 14979 16581
rect 14921 16541 14933 16575
rect 14967 16572 14979 16575
rect 15010 16572 15016 16584
rect 14967 16544 15016 16572
rect 14967 16541 14979 16544
rect 14921 16535 14979 16541
rect 15010 16532 15016 16544
rect 15068 16532 15074 16584
rect 11330 16504 11336 16516
rect 9508 16476 11336 16504
rect 11330 16464 11336 16476
rect 11388 16464 11394 16516
rect 5408 16408 6868 16436
rect 5408 16396 5414 16408
rect 7650 16396 7656 16448
rect 7708 16436 7714 16448
rect 8849 16439 8907 16445
rect 8849 16436 8861 16439
rect 7708 16408 8861 16436
rect 7708 16396 7714 16408
rect 8849 16405 8861 16408
rect 8895 16405 8907 16439
rect 8849 16399 8907 16405
rect 9677 16439 9735 16445
rect 9677 16405 9689 16439
rect 9723 16436 9735 16439
rect 9766 16436 9772 16448
rect 9723 16408 9772 16436
rect 9723 16405 9735 16408
rect 9677 16399 9735 16405
rect 9766 16396 9772 16408
rect 9824 16396 9830 16448
rect 10594 16396 10600 16448
rect 10652 16436 10658 16448
rect 15194 16436 15200 16448
rect 10652 16408 15200 16436
rect 10652 16396 10658 16408
rect 15194 16396 15200 16408
rect 15252 16436 15258 16448
rect 15930 16436 15936 16448
rect 15252 16408 15936 16436
rect 15252 16396 15258 16408
rect 15930 16396 15936 16408
rect 15988 16396 15994 16448
rect 1104 16346 15824 16368
rect 1104 16294 3447 16346
rect 3499 16294 3511 16346
rect 3563 16294 3575 16346
rect 3627 16294 3639 16346
rect 3691 16294 8378 16346
rect 8430 16294 8442 16346
rect 8494 16294 8506 16346
rect 8558 16294 8570 16346
rect 8622 16294 13308 16346
rect 13360 16294 13372 16346
rect 13424 16294 13436 16346
rect 13488 16294 13500 16346
rect 13552 16294 15824 16346
rect 1104 16272 15824 16294
rect 1854 16192 1860 16244
rect 1912 16232 1918 16244
rect 2501 16235 2559 16241
rect 2501 16232 2513 16235
rect 1912 16204 2513 16232
rect 1912 16192 1918 16204
rect 2501 16201 2513 16204
rect 2547 16201 2559 16235
rect 2501 16195 2559 16201
rect 3326 16192 3332 16244
rect 3384 16232 3390 16244
rect 3605 16235 3663 16241
rect 3605 16232 3617 16235
rect 3384 16204 3617 16232
rect 3384 16192 3390 16204
rect 3605 16201 3617 16204
rect 3651 16201 3663 16235
rect 3605 16195 3663 16201
rect 3786 16192 3792 16244
rect 3844 16232 3850 16244
rect 4157 16235 4215 16241
rect 4157 16232 4169 16235
rect 3844 16204 4169 16232
rect 3844 16192 3850 16204
rect 4157 16201 4169 16204
rect 4203 16201 4215 16235
rect 4157 16195 4215 16201
rect 5353 16235 5411 16241
rect 5353 16201 5365 16235
rect 5399 16232 5411 16235
rect 6270 16232 6276 16244
rect 5399 16204 6276 16232
rect 5399 16201 5411 16204
rect 5353 16195 5411 16201
rect 6270 16192 6276 16204
rect 6328 16192 6334 16244
rect 7006 16192 7012 16244
rect 7064 16232 7070 16244
rect 8021 16235 8079 16241
rect 8021 16232 8033 16235
rect 7064 16204 8033 16232
rect 7064 16192 7070 16204
rect 8021 16201 8033 16204
rect 8067 16201 8079 16235
rect 8021 16195 8079 16201
rect 9030 16192 9036 16244
rect 9088 16232 9094 16244
rect 11422 16232 11428 16244
rect 9088 16204 11428 16232
rect 9088 16192 9094 16204
rect 11422 16192 11428 16204
rect 11480 16192 11486 16244
rect 12434 16192 12440 16244
rect 12492 16232 12498 16244
rect 12492 16204 12537 16232
rect 12492 16192 12498 16204
rect 2222 16124 2228 16176
rect 2280 16164 2286 16176
rect 3053 16167 3111 16173
rect 3053 16164 3065 16167
rect 2280 16136 3065 16164
rect 2280 16124 2286 16136
rect 3053 16133 3065 16136
rect 3099 16133 3111 16167
rect 3053 16127 3111 16133
rect 6454 16124 6460 16176
rect 6512 16164 6518 16176
rect 8110 16164 8116 16176
rect 6512 16136 8116 16164
rect 6512 16124 6518 16136
rect 8110 16124 8116 16136
rect 8168 16124 8174 16176
rect 1762 16096 1768 16108
rect 1723 16068 1768 16096
rect 1762 16056 1768 16068
rect 1820 16056 1826 16108
rect 5534 16096 5540 16108
rect 3252 16068 5540 16096
rect 1581 16031 1639 16037
rect 1581 15997 1593 16031
rect 1627 16028 1639 16031
rect 2314 16028 2320 16040
rect 1627 16000 2176 16028
rect 2275 16000 2320 16028
rect 1627 15997 1639 16000
rect 1581 15991 1639 15997
rect 2148 15960 2176 16000
rect 2314 15988 2320 16000
rect 2372 15988 2378 16040
rect 2869 16031 2927 16037
rect 2869 15997 2881 16031
rect 2915 16028 2927 16031
rect 3252 16028 3280 16068
rect 5534 16056 5540 16068
rect 5592 16056 5598 16108
rect 6362 16096 6368 16108
rect 6323 16068 6368 16096
rect 6362 16056 6368 16068
rect 6420 16056 6426 16108
rect 7469 16099 7527 16105
rect 7469 16065 7481 16099
rect 7515 16096 7527 16099
rect 7650 16096 7656 16108
rect 7515 16068 7656 16096
rect 7515 16065 7527 16068
rect 7469 16059 7527 16065
rect 7650 16056 7656 16068
rect 7708 16056 7714 16108
rect 11698 16056 11704 16108
rect 11756 16096 11762 16108
rect 12989 16099 13047 16105
rect 12989 16096 13001 16099
rect 11756 16068 13001 16096
rect 11756 16056 11762 16068
rect 12989 16065 13001 16068
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 2915 16000 3280 16028
rect 2915 15997 2927 16000
rect 2869 15991 2927 15997
rect 3326 15988 3332 16040
rect 3384 16028 3390 16040
rect 3421 16031 3479 16037
rect 3421 16028 3433 16031
rect 3384 16000 3433 16028
rect 3384 15988 3390 16000
rect 3421 15997 3433 16000
rect 3467 15997 3479 16031
rect 3421 15991 3479 15997
rect 3786 15988 3792 16040
rect 3844 16028 3850 16040
rect 3973 16031 4031 16037
rect 3973 16028 3985 16031
rect 3844 16000 3985 16028
rect 3844 15988 3850 16000
rect 3973 15997 3985 16000
rect 4019 15997 4031 16031
rect 5166 16028 5172 16040
rect 5127 16000 5172 16028
rect 3973 15991 4031 15997
rect 5166 15988 5172 16000
rect 5224 15988 5230 16040
rect 7834 16028 7840 16040
rect 7795 16000 7840 16028
rect 7834 15988 7840 16000
rect 7892 15988 7898 16040
rect 8386 16028 8392 16040
rect 8347 16000 8392 16028
rect 8386 15988 8392 16000
rect 8444 15988 8450 16040
rect 8662 16037 8668 16040
rect 8656 16028 8668 16037
rect 8623 16000 8668 16028
rect 8656 15991 8668 16000
rect 8662 15988 8668 15991
rect 8720 15988 8726 16040
rect 9122 15988 9128 16040
rect 9180 16028 9186 16040
rect 10045 16031 10103 16037
rect 10045 16028 10057 16031
rect 9180 16000 10057 16028
rect 9180 15988 9186 16000
rect 10045 15997 10057 16000
rect 10091 15997 10103 16031
rect 10312 16031 10370 16037
rect 10312 16028 10324 16031
rect 10045 15991 10103 15997
rect 10244 16000 10324 16028
rect 2774 15960 2780 15972
rect 2148 15932 2780 15960
rect 2774 15920 2780 15932
rect 2832 15920 2838 15972
rect 6089 15963 6147 15969
rect 2976 15932 5764 15960
rect 2590 15852 2596 15904
rect 2648 15892 2654 15904
rect 2976 15892 3004 15932
rect 5736 15901 5764 15932
rect 6089 15929 6101 15963
rect 6135 15960 6147 15963
rect 9582 15960 9588 15972
rect 6135 15932 9588 15960
rect 6135 15929 6147 15932
rect 6089 15923 6147 15929
rect 9582 15920 9588 15932
rect 9640 15920 9646 15972
rect 10134 15960 10140 15972
rect 9692 15932 10140 15960
rect 2648 15864 3004 15892
rect 5721 15895 5779 15901
rect 2648 15852 2654 15864
rect 5721 15861 5733 15895
rect 5767 15861 5779 15895
rect 5721 15855 5779 15861
rect 6181 15895 6239 15901
rect 6181 15861 6193 15895
rect 6227 15892 6239 15895
rect 6825 15895 6883 15901
rect 6825 15892 6837 15895
rect 6227 15864 6837 15892
rect 6227 15861 6239 15864
rect 6181 15855 6239 15861
rect 6825 15861 6837 15864
rect 6871 15861 6883 15895
rect 6825 15855 6883 15861
rect 7006 15852 7012 15904
rect 7064 15892 7070 15904
rect 7193 15895 7251 15901
rect 7193 15892 7205 15895
rect 7064 15864 7205 15892
rect 7064 15852 7070 15864
rect 7193 15861 7205 15864
rect 7239 15861 7251 15895
rect 7193 15855 7251 15861
rect 7282 15852 7288 15904
rect 7340 15892 7346 15904
rect 7340 15864 7385 15892
rect 7340 15852 7346 15864
rect 8386 15852 8392 15904
rect 8444 15892 8450 15904
rect 9692 15892 9720 15932
rect 10134 15920 10140 15932
rect 10192 15920 10198 15972
rect 8444 15864 9720 15892
rect 9769 15895 9827 15901
rect 8444 15852 8450 15864
rect 9769 15861 9781 15895
rect 9815 15892 9827 15895
rect 10244 15892 10272 16000
rect 10312 15997 10324 16000
rect 10358 16028 10370 16031
rect 11716 16028 11744 16056
rect 10358 16000 11744 16028
rect 10358 15997 10370 16000
rect 10312 15991 10370 15997
rect 11974 15988 11980 16040
rect 12032 16028 12038 16040
rect 13449 16031 13507 16037
rect 13449 16028 13461 16031
rect 12032 16000 13461 16028
rect 12032 15988 12038 16000
rect 13449 15997 13461 16000
rect 13495 15997 13507 16031
rect 13449 15991 13507 15997
rect 11238 15920 11244 15972
rect 11296 15960 11302 15972
rect 13538 15960 13544 15972
rect 11296 15932 13544 15960
rect 11296 15920 11302 15932
rect 13538 15920 13544 15932
rect 13596 15960 13602 15972
rect 13694 15963 13752 15969
rect 13694 15960 13706 15963
rect 13596 15932 13706 15960
rect 13596 15920 13602 15932
rect 13694 15929 13706 15932
rect 13740 15929 13752 15963
rect 15286 15960 15292 15972
rect 13694 15923 13752 15929
rect 13832 15932 15292 15960
rect 9815 15864 10272 15892
rect 11425 15895 11483 15901
rect 9815 15861 9827 15864
rect 9769 15855 9827 15861
rect 11425 15861 11437 15895
rect 11471 15892 11483 15895
rect 11606 15892 11612 15904
rect 11471 15864 11612 15892
rect 11471 15861 11483 15864
rect 11425 15855 11483 15861
rect 11606 15852 11612 15864
rect 11664 15852 11670 15904
rect 11701 15895 11759 15901
rect 11701 15861 11713 15895
rect 11747 15892 11759 15895
rect 12805 15895 12863 15901
rect 12805 15892 12817 15895
rect 11747 15864 12817 15892
rect 11747 15861 11759 15864
rect 11701 15855 11759 15861
rect 12805 15861 12817 15864
rect 12851 15861 12863 15895
rect 12805 15855 12863 15861
rect 12897 15895 12955 15901
rect 12897 15861 12909 15895
rect 12943 15892 12955 15895
rect 13832 15892 13860 15932
rect 15286 15920 15292 15932
rect 15344 15960 15350 15972
rect 16390 15960 16396 15972
rect 15344 15932 16396 15960
rect 15344 15920 15350 15932
rect 16390 15920 16396 15932
rect 16448 15920 16454 15972
rect 14826 15892 14832 15904
rect 12943 15864 13860 15892
rect 14787 15864 14832 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 14826 15852 14832 15864
rect 14884 15852 14890 15904
rect 14918 15852 14924 15904
rect 14976 15892 14982 15904
rect 15105 15895 15163 15901
rect 15105 15892 15117 15895
rect 14976 15864 15117 15892
rect 14976 15852 14982 15864
rect 15105 15861 15117 15864
rect 15151 15861 15163 15895
rect 15105 15855 15163 15861
rect 1104 15802 15824 15824
rect 1104 15750 5912 15802
rect 5964 15750 5976 15802
rect 6028 15750 6040 15802
rect 6092 15750 6104 15802
rect 6156 15750 10843 15802
rect 10895 15750 10907 15802
rect 10959 15750 10971 15802
rect 11023 15750 11035 15802
rect 11087 15750 15824 15802
rect 1104 15728 15824 15750
rect 566 15648 572 15700
rect 624 15688 630 15700
rect 2409 15691 2467 15697
rect 2409 15688 2421 15691
rect 624 15660 2421 15688
rect 624 15648 630 15660
rect 2409 15657 2421 15660
rect 2455 15657 2467 15691
rect 2409 15651 2467 15657
rect 6549 15691 6607 15697
rect 6549 15657 6561 15691
rect 6595 15688 6607 15691
rect 6638 15688 6644 15700
rect 6595 15660 6644 15688
rect 6595 15657 6607 15660
rect 6549 15651 6607 15657
rect 6638 15648 6644 15660
rect 6696 15648 6702 15700
rect 7006 15688 7012 15700
rect 6967 15660 7012 15688
rect 7006 15648 7012 15660
rect 7064 15648 7070 15700
rect 7466 15688 7472 15700
rect 7379 15660 7472 15688
rect 7466 15648 7472 15660
rect 7524 15688 7530 15700
rect 7926 15688 7932 15700
rect 7524 15660 7932 15688
rect 7524 15648 7530 15660
rect 7926 15648 7932 15660
rect 7984 15648 7990 15700
rect 8021 15691 8079 15697
rect 8021 15657 8033 15691
rect 8067 15688 8079 15691
rect 10137 15691 10195 15697
rect 10137 15688 10149 15691
rect 8067 15660 10149 15688
rect 8067 15657 8079 15660
rect 8021 15651 8079 15657
rect 10137 15657 10149 15660
rect 10183 15657 10195 15691
rect 10137 15651 10195 15657
rect 10226 15648 10232 15700
rect 10284 15688 10290 15700
rect 11238 15688 11244 15700
rect 10284 15660 11244 15688
rect 10284 15648 10290 15660
rect 11238 15648 11244 15660
rect 11296 15648 11302 15700
rect 12802 15688 12808 15700
rect 11900 15660 12808 15688
rect 1762 15620 1768 15632
rect 1723 15592 1768 15620
rect 1762 15580 1768 15592
rect 1820 15580 1826 15632
rect 2590 15620 2596 15632
rect 2148 15592 2596 15620
rect 1489 15555 1547 15561
rect 1489 15521 1501 15555
rect 1535 15552 1547 15555
rect 2148 15552 2176 15592
rect 2590 15580 2596 15592
rect 2648 15580 2654 15632
rect 3421 15623 3479 15629
rect 3421 15589 3433 15623
rect 3467 15620 3479 15623
rect 3970 15620 3976 15632
rect 3467 15592 3976 15620
rect 3467 15589 3479 15592
rect 3421 15583 3479 15589
rect 3970 15580 3976 15592
rect 4028 15580 4034 15632
rect 4976 15623 5034 15629
rect 4976 15589 4988 15623
rect 5022 15620 5034 15623
rect 8386 15620 8392 15632
rect 5022 15592 7512 15620
rect 8347 15592 8392 15620
rect 5022 15589 5034 15592
rect 4976 15583 5034 15589
rect 1535 15524 2176 15552
rect 2225 15555 2283 15561
rect 1535 15521 1547 15524
rect 1489 15515 1547 15521
rect 2225 15521 2237 15555
rect 2271 15552 2283 15555
rect 3234 15552 3240 15564
rect 2271 15524 3240 15552
rect 2271 15521 2283 15524
rect 2225 15515 2283 15521
rect 3234 15512 3240 15524
rect 3292 15512 3298 15564
rect 3329 15555 3387 15561
rect 3329 15521 3341 15555
rect 3375 15552 3387 15555
rect 4338 15552 4344 15564
rect 3375 15524 4344 15552
rect 3375 15521 3387 15524
rect 3329 15515 3387 15521
rect 4338 15512 4344 15524
rect 4396 15512 4402 15564
rect 4709 15555 4767 15561
rect 4709 15521 4721 15555
rect 4755 15552 4767 15555
rect 5350 15552 5356 15564
rect 4755 15524 5356 15552
rect 4755 15521 4767 15524
rect 4709 15515 4767 15521
rect 5350 15512 5356 15524
rect 5408 15512 5414 15564
rect 6362 15552 6368 15564
rect 6323 15524 6368 15552
rect 6362 15512 6368 15524
rect 6420 15512 6426 15564
rect 6546 15512 6552 15564
rect 6604 15552 6610 15564
rect 7190 15552 7196 15564
rect 6604 15524 7196 15552
rect 6604 15512 6610 15524
rect 7190 15512 7196 15524
rect 7248 15552 7254 15564
rect 7377 15555 7435 15561
rect 7377 15552 7389 15555
rect 7248 15524 7389 15552
rect 7248 15512 7254 15524
rect 7377 15521 7389 15524
rect 7423 15521 7435 15555
rect 7484 15552 7512 15592
rect 8386 15580 8392 15592
rect 8444 15580 8450 15632
rect 8481 15623 8539 15629
rect 8481 15589 8493 15623
rect 8527 15620 8539 15623
rect 11900 15620 11928 15660
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 13170 15688 13176 15700
rect 13004 15660 13176 15688
rect 8527 15592 11928 15620
rect 12520 15623 12578 15629
rect 8527 15589 8539 15592
rect 8481 15583 8539 15589
rect 12520 15589 12532 15623
rect 12566 15620 12578 15623
rect 13004 15620 13032 15660
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 13538 15648 13544 15700
rect 13596 15688 13602 15700
rect 13633 15691 13691 15697
rect 13633 15688 13645 15691
rect 13596 15660 13645 15688
rect 13596 15648 13602 15660
rect 13633 15657 13645 15660
rect 13679 15657 13691 15691
rect 13906 15688 13912 15700
rect 13867 15660 13912 15688
rect 13633 15651 13691 15657
rect 13906 15648 13912 15660
rect 13964 15648 13970 15700
rect 15102 15648 15108 15700
rect 15160 15688 15166 15700
rect 16758 15688 16764 15700
rect 15160 15660 16764 15688
rect 15160 15648 15166 15660
rect 16758 15648 16764 15660
rect 16816 15648 16822 15700
rect 12566 15592 13032 15620
rect 12566 15589 12578 15592
rect 12520 15583 12578 15589
rect 13078 15580 13084 15632
rect 13136 15620 13142 15632
rect 14369 15623 14427 15629
rect 14369 15620 14381 15623
rect 13136 15592 14381 15620
rect 13136 15580 13142 15592
rect 14369 15589 14381 15592
rect 14415 15589 14427 15623
rect 14369 15583 14427 15589
rect 7484 15524 7604 15552
rect 7377 15515 7435 15521
rect 2774 15444 2780 15496
rect 2832 15444 2838 15496
rect 2958 15444 2964 15496
rect 3016 15484 3022 15496
rect 7576 15493 7604 15524
rect 8110 15512 8116 15564
rect 8168 15552 8174 15564
rect 8846 15552 8852 15564
rect 8168 15524 8852 15552
rect 8168 15512 8174 15524
rect 8846 15512 8852 15524
rect 8904 15512 8910 15564
rect 9030 15552 9036 15564
rect 8991 15524 9036 15552
rect 9030 15512 9036 15524
rect 9088 15552 9094 15564
rect 9306 15552 9312 15564
rect 9088 15524 9312 15552
rect 9088 15512 9094 15524
rect 9306 15512 9312 15524
rect 9364 15512 9370 15564
rect 10042 15552 10048 15564
rect 10003 15524 10048 15552
rect 10042 15512 10048 15524
rect 10100 15512 10106 15564
rect 10134 15512 10140 15564
rect 10192 15552 10198 15564
rect 10962 15552 10968 15564
rect 10192 15524 10968 15552
rect 10192 15512 10198 15524
rect 10962 15512 10968 15524
rect 11020 15512 11026 15564
rect 11057 15555 11115 15561
rect 11057 15521 11069 15555
rect 11103 15552 11115 15555
rect 11514 15552 11520 15564
rect 11103 15524 11520 15552
rect 11103 15521 11115 15524
rect 11057 15515 11115 15521
rect 11514 15512 11520 15524
rect 11572 15512 11578 15564
rect 14274 15552 14280 15564
rect 14235 15524 14280 15552
rect 14274 15512 14280 15524
rect 14332 15512 14338 15564
rect 3513 15487 3571 15493
rect 3513 15484 3525 15487
rect 3016 15456 3525 15484
rect 3016 15444 3022 15456
rect 3513 15453 3525 15456
rect 3559 15453 3571 15487
rect 3513 15447 3571 15453
rect 7561 15487 7619 15493
rect 7561 15453 7573 15487
rect 7607 15484 7619 15487
rect 8018 15484 8024 15496
rect 7607 15456 8024 15484
rect 7607 15453 7619 15456
rect 7561 15447 7619 15453
rect 8018 15444 8024 15456
rect 8076 15484 8082 15496
rect 8573 15487 8631 15493
rect 8573 15484 8585 15487
rect 8076 15456 8585 15484
rect 8076 15444 8082 15456
rect 8573 15453 8585 15456
rect 8619 15453 8631 15487
rect 10229 15487 10287 15493
rect 10229 15484 10241 15487
rect 8573 15447 8631 15453
rect 8680 15456 10241 15484
rect 2792 15416 2820 15444
rect 2792 15388 3096 15416
rect 2774 15308 2780 15360
rect 2832 15348 2838 15360
rect 2961 15351 3019 15357
rect 2961 15348 2973 15351
rect 2832 15320 2973 15348
rect 2832 15308 2838 15320
rect 2961 15317 2973 15320
rect 3007 15317 3019 15351
rect 3068 15348 3096 15388
rect 5718 15376 5724 15428
rect 5776 15416 5782 15428
rect 6089 15419 6147 15425
rect 6089 15416 6101 15419
rect 5776 15388 6101 15416
rect 5776 15376 5782 15388
rect 6089 15385 6101 15388
rect 6135 15416 6147 15419
rect 7650 15416 7656 15428
rect 6135 15388 7656 15416
rect 6135 15385 6147 15388
rect 6089 15379 6147 15385
rect 7650 15376 7656 15388
rect 7708 15416 7714 15428
rect 8680 15416 8708 15456
rect 10229 15453 10241 15456
rect 10275 15453 10287 15487
rect 10229 15447 10287 15453
rect 10410 15444 10416 15496
rect 10468 15484 10474 15496
rect 11149 15487 11207 15493
rect 11149 15484 11161 15487
rect 10468 15456 11161 15484
rect 10468 15444 10474 15456
rect 11149 15453 11161 15456
rect 11195 15453 11207 15487
rect 11149 15447 11207 15453
rect 11333 15487 11391 15493
rect 11333 15453 11345 15487
rect 11379 15484 11391 15487
rect 11698 15484 11704 15496
rect 11379 15456 11704 15484
rect 11379 15453 11391 15456
rect 11333 15447 11391 15453
rect 11698 15444 11704 15456
rect 11756 15444 11762 15496
rect 11974 15444 11980 15496
rect 12032 15484 12038 15496
rect 12158 15484 12164 15496
rect 12032 15456 12164 15484
rect 12032 15444 12038 15456
rect 12158 15444 12164 15456
rect 12216 15484 12222 15496
rect 12253 15487 12311 15493
rect 12253 15484 12265 15487
rect 12216 15456 12265 15484
rect 12216 15444 12222 15456
rect 12253 15453 12265 15456
rect 12299 15453 12311 15487
rect 12253 15447 12311 15453
rect 13998 15444 14004 15496
rect 14056 15484 14062 15496
rect 14461 15487 14519 15493
rect 14461 15484 14473 15487
rect 14056 15456 14473 15484
rect 14056 15444 14062 15456
rect 14461 15453 14473 15456
rect 14507 15484 14519 15487
rect 14550 15484 14556 15496
rect 14507 15456 14556 15484
rect 14507 15453 14519 15456
rect 14461 15447 14519 15453
rect 14550 15444 14556 15456
rect 14608 15444 14614 15496
rect 7708 15388 8708 15416
rect 7708 15376 7714 15388
rect 8754 15376 8760 15428
rect 8812 15416 8818 15428
rect 9217 15419 9275 15425
rect 9217 15416 9229 15419
rect 8812 15388 9229 15416
rect 8812 15376 8818 15388
rect 9217 15385 9229 15388
rect 9263 15385 9275 15419
rect 9217 15379 9275 15385
rect 9582 15376 9588 15428
rect 9640 15416 9646 15428
rect 9677 15419 9735 15425
rect 9677 15416 9689 15419
rect 9640 15388 9689 15416
rect 9640 15376 9646 15388
rect 9677 15385 9689 15388
rect 9723 15385 9735 15419
rect 9677 15379 9735 15385
rect 9968 15388 12296 15416
rect 9968 15348 9996 15388
rect 12268 15360 12296 15388
rect 3068 15320 9996 15348
rect 10689 15351 10747 15357
rect 2961 15311 3019 15317
rect 10689 15317 10701 15351
rect 10735 15348 10747 15351
rect 11514 15348 11520 15360
rect 10735 15320 11520 15348
rect 10735 15317 10747 15320
rect 10689 15311 10747 15317
rect 11514 15308 11520 15320
rect 11572 15308 11578 15360
rect 12250 15308 12256 15360
rect 12308 15308 12314 15360
rect 1104 15258 15824 15280
rect 1104 15206 3447 15258
rect 3499 15206 3511 15258
rect 3563 15206 3575 15258
rect 3627 15206 3639 15258
rect 3691 15206 8378 15258
rect 8430 15206 8442 15258
rect 8494 15206 8506 15258
rect 8558 15206 8570 15258
rect 8622 15206 13308 15258
rect 13360 15206 13372 15258
rect 13424 15206 13436 15258
rect 13488 15206 13500 15258
rect 13552 15206 15824 15258
rect 1104 15184 15824 15206
rect 4062 15144 4068 15156
rect 2516 15116 4068 15144
rect 2317 15011 2375 15017
rect 2317 14977 2329 15011
rect 2363 15008 2375 15011
rect 2516 15008 2544 15116
rect 4062 15104 4068 15116
rect 4120 15104 4126 15156
rect 4338 15144 4344 15156
rect 4299 15116 4344 15144
rect 4338 15104 4344 15116
rect 4396 15104 4402 15156
rect 5350 15104 5356 15156
rect 5408 15144 5414 15156
rect 6365 15147 6423 15153
rect 6365 15144 6377 15147
rect 5408 15116 6377 15144
rect 5408 15104 5414 15116
rect 6365 15113 6377 15116
rect 6411 15113 6423 15147
rect 6365 15107 6423 15113
rect 7282 15104 7288 15156
rect 7340 15144 7346 15156
rect 7469 15147 7527 15153
rect 7469 15144 7481 15147
rect 7340 15116 7481 15144
rect 7340 15104 7346 15116
rect 7469 15113 7481 15116
rect 7515 15113 7527 15147
rect 7469 15107 7527 15113
rect 8018 15104 8024 15156
rect 8076 15144 8082 15156
rect 9861 15147 9919 15153
rect 9861 15144 9873 15147
rect 8076 15116 9873 15144
rect 8076 15104 8082 15116
rect 9861 15113 9873 15116
rect 9907 15113 9919 15147
rect 9861 15107 9919 15113
rect 9876 15076 9904 15107
rect 10042 15104 10048 15156
rect 10100 15144 10106 15156
rect 10137 15147 10195 15153
rect 10137 15144 10149 15147
rect 10100 15116 10149 15144
rect 10100 15104 10106 15116
rect 10137 15113 10149 15116
rect 10183 15113 10195 15147
rect 10137 15107 10195 15113
rect 10226 15104 10232 15156
rect 10284 15144 10290 15156
rect 10284 15116 11928 15144
rect 10284 15104 10290 15116
rect 11149 15079 11207 15085
rect 9876 15048 10732 15076
rect 2363 14980 2544 15008
rect 2363 14977 2375 14980
rect 2317 14971 2375 14977
rect 4522 14968 4528 15020
rect 4580 15008 4586 15020
rect 4893 15011 4951 15017
rect 4893 15008 4905 15011
rect 4580 14980 4905 15008
rect 4580 14968 4586 14980
rect 4893 14977 4905 14980
rect 4939 14977 4951 15011
rect 4893 14971 4951 14977
rect 5626 14968 5632 15020
rect 5684 15008 5690 15020
rect 5905 15011 5963 15017
rect 5905 15008 5917 15011
rect 5684 14980 5917 15008
rect 5684 14968 5690 14980
rect 5905 14977 5917 14980
rect 5951 14977 5963 15011
rect 7742 15008 7748 15020
rect 5905 14971 5963 14977
rect 7300 14980 7748 15008
rect 1486 14900 1492 14952
rect 1544 14940 1550 14952
rect 2958 14949 2964 14952
rect 2685 14943 2743 14949
rect 2685 14940 2697 14943
rect 1544 14912 2697 14940
rect 1544 14900 1550 14912
rect 2685 14909 2697 14912
rect 2731 14940 2743 14943
rect 2731 14912 2912 14940
rect 2731 14909 2743 14912
rect 2685 14903 2743 14909
rect 2041 14875 2099 14881
rect 2041 14841 2053 14875
rect 2087 14872 2099 14875
rect 2774 14872 2780 14884
rect 2087 14844 2780 14872
rect 2087 14841 2099 14844
rect 2041 14835 2099 14841
rect 2774 14832 2780 14844
rect 2832 14832 2838 14884
rect 2884 14872 2912 14912
rect 2952 14903 2964 14949
rect 3016 14940 3022 14952
rect 4798 14940 4804 14952
rect 3016 14912 3052 14940
rect 4759 14912 4804 14940
rect 2958 14900 2964 14903
rect 3016 14900 3022 14912
rect 4798 14900 4804 14912
rect 4856 14900 4862 14952
rect 6546 14940 6552 14952
rect 6507 14912 6552 14940
rect 6546 14900 6552 14912
rect 6604 14900 6610 14952
rect 7300 14940 7328 14980
rect 7742 14968 7748 14980
rect 7800 14968 7806 15020
rect 8018 15008 8024 15020
rect 7979 14980 8024 15008
rect 8018 14968 8024 14980
rect 8076 14968 8082 15020
rect 9674 14968 9680 15020
rect 9732 15008 9738 15020
rect 10134 15008 10140 15020
rect 9732 14980 10140 15008
rect 9732 14968 9738 14980
rect 10134 14968 10140 14980
rect 10192 14968 10198 15020
rect 10594 15008 10600 15020
rect 10555 14980 10600 15008
rect 10594 14968 10600 14980
rect 10652 14968 10658 15020
rect 10704 15017 10732 15048
rect 11149 15045 11161 15079
rect 11195 15076 11207 15079
rect 11900 15076 11928 15116
rect 12250 15104 12256 15156
rect 12308 15144 12314 15156
rect 12437 15147 12495 15153
rect 12437 15144 12449 15147
rect 12308 15116 12449 15144
rect 12308 15104 12314 15116
rect 12437 15113 12449 15116
rect 12483 15113 12495 15147
rect 12437 15107 12495 15113
rect 12986 15104 12992 15156
rect 13044 15144 13050 15156
rect 14461 15147 14519 15153
rect 14461 15144 14473 15147
rect 13044 15116 14473 15144
rect 13044 15104 13050 15116
rect 14461 15113 14473 15116
rect 14507 15113 14519 15147
rect 14461 15107 14519 15113
rect 14550 15104 14556 15156
rect 14608 15144 14614 15156
rect 14608 15116 15056 15144
rect 14608 15104 14614 15116
rect 13449 15079 13507 15085
rect 11195 15048 11836 15076
rect 11900 15048 13216 15076
rect 11195 15045 11207 15048
rect 11149 15039 11207 15045
rect 10689 15011 10747 15017
rect 10689 14977 10701 15011
rect 10735 14977 10747 15011
rect 10689 14971 10747 14977
rect 11606 14968 11612 15020
rect 11664 15008 11670 15020
rect 11701 15011 11759 15017
rect 11701 15008 11713 15011
rect 11664 14980 11713 15008
rect 11664 14968 11670 14980
rect 11701 14977 11713 14980
rect 11747 14977 11759 15011
rect 11808 15008 11836 15048
rect 12897 15011 12955 15017
rect 12897 15008 12909 15011
rect 11808 14980 12909 15008
rect 11701 14971 11759 14977
rect 12897 14977 12909 14980
rect 12943 14977 12955 15011
rect 12897 14971 12955 14977
rect 12986 14968 12992 15020
rect 13044 15008 13050 15020
rect 13188 15008 13216 15048
rect 13449 15045 13461 15079
rect 13495 15076 13507 15079
rect 13495 15048 14964 15076
rect 13495 15045 13507 15048
rect 13449 15039 13507 15045
rect 13909 15011 13967 15017
rect 13909 15008 13921 15011
rect 13044 14980 13089 15008
rect 13188 14980 13921 15008
rect 13044 14968 13050 14980
rect 13909 14977 13921 14980
rect 13955 14977 13967 15011
rect 14090 15008 14096 15020
rect 14051 14980 14096 15008
rect 13909 14971 13967 14977
rect 14090 14968 14096 14980
rect 14148 14968 14154 15020
rect 14936 15017 14964 15048
rect 15028 15017 15056 15116
rect 14921 15011 14979 15017
rect 14921 14977 14933 15011
rect 14967 14977 14979 15011
rect 14921 14971 14979 14977
rect 15013 15011 15071 15017
rect 15013 14977 15025 15011
rect 15059 14977 15071 15011
rect 15013 14971 15071 14977
rect 6932 14912 7328 14940
rect 5442 14872 5448 14884
rect 2884 14844 5448 14872
rect 5442 14832 5448 14844
rect 5500 14832 5506 14884
rect 5534 14832 5540 14884
rect 5592 14872 5598 14884
rect 6932 14872 6960 14912
rect 7374 14900 7380 14952
rect 7432 14940 7438 14952
rect 7837 14943 7895 14949
rect 7837 14940 7849 14943
rect 7432 14912 7849 14940
rect 7432 14900 7438 14912
rect 7837 14909 7849 14912
rect 7883 14940 7895 14943
rect 8297 14943 8355 14949
rect 8297 14940 8309 14943
rect 7883 14912 8309 14940
rect 7883 14909 7895 14912
rect 7837 14903 7895 14909
rect 8297 14909 8309 14912
rect 8343 14909 8355 14943
rect 8297 14903 8355 14909
rect 8481 14943 8539 14949
rect 8481 14909 8493 14943
rect 8527 14940 8539 14943
rect 8570 14940 8576 14952
rect 8527 14912 8576 14940
rect 8527 14909 8539 14912
rect 8481 14903 8539 14909
rect 8570 14900 8576 14912
rect 8628 14900 8634 14952
rect 10505 14943 10563 14949
rect 10505 14940 10517 14943
rect 8680 14912 10517 14940
rect 5592 14844 6960 14872
rect 7009 14875 7067 14881
rect 5592 14832 5598 14844
rect 7009 14841 7021 14875
rect 7055 14872 7067 14875
rect 8680 14872 8708 14912
rect 10505 14909 10517 14912
rect 10551 14909 10563 14943
rect 11514 14940 11520 14952
rect 11475 14912 11520 14940
rect 10505 14903 10563 14909
rect 11514 14900 11520 14912
rect 11572 14900 11578 14952
rect 12805 14943 12863 14949
rect 12805 14909 12817 14943
rect 12851 14940 12863 14943
rect 13722 14940 13728 14952
rect 12851 14912 13728 14940
rect 12851 14909 12863 14912
rect 12805 14903 12863 14909
rect 13722 14900 13728 14912
rect 13780 14900 13786 14952
rect 7055 14844 8708 14872
rect 8748 14875 8806 14881
rect 7055 14841 7067 14844
rect 7009 14835 7067 14841
rect 8748 14841 8760 14875
rect 8794 14872 8806 14875
rect 8938 14872 8944 14884
rect 8794 14844 8944 14872
rect 8794 14841 8806 14844
rect 8748 14835 8806 14841
rect 8938 14832 8944 14844
rect 8996 14832 9002 14884
rect 9766 14832 9772 14884
rect 9824 14872 9830 14884
rect 11609 14875 11667 14881
rect 11609 14872 11621 14875
rect 9824 14844 11621 14872
rect 9824 14832 9830 14844
rect 11609 14841 11621 14844
rect 11655 14841 11667 14875
rect 13817 14875 13875 14881
rect 13817 14872 13829 14875
rect 11609 14835 11667 14841
rect 12912 14844 13829 14872
rect 1394 14764 1400 14816
rect 1452 14804 1458 14816
rect 1673 14807 1731 14813
rect 1673 14804 1685 14807
rect 1452 14776 1685 14804
rect 1452 14764 1458 14776
rect 1673 14773 1685 14776
rect 1719 14773 1731 14807
rect 1673 14767 1731 14773
rect 1946 14764 1952 14816
rect 2004 14804 2010 14816
rect 2133 14807 2191 14813
rect 2133 14804 2145 14807
rect 2004 14776 2145 14804
rect 2004 14764 2010 14776
rect 2133 14773 2145 14776
rect 2179 14773 2191 14807
rect 4706 14804 4712 14816
rect 4667 14776 4712 14804
rect 2133 14767 2191 14773
rect 4706 14764 4712 14776
rect 4764 14764 4770 14816
rect 5350 14804 5356 14816
rect 5311 14776 5356 14804
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 5718 14804 5724 14816
rect 5679 14776 5724 14804
rect 5718 14764 5724 14776
rect 5776 14764 5782 14816
rect 5810 14764 5816 14816
rect 5868 14804 5874 14816
rect 5868 14776 5913 14804
rect 5868 14764 5874 14776
rect 7926 14764 7932 14816
rect 7984 14804 7990 14816
rect 8297 14807 8355 14813
rect 7984 14776 8029 14804
rect 7984 14764 7990 14776
rect 8297 14773 8309 14807
rect 8343 14804 8355 14807
rect 9582 14804 9588 14816
rect 8343 14776 9588 14804
rect 8343 14773 8355 14776
rect 8297 14767 8355 14773
rect 9582 14764 9588 14776
rect 9640 14764 9646 14816
rect 10042 14764 10048 14816
rect 10100 14804 10106 14816
rect 10318 14804 10324 14816
rect 10100 14776 10324 14804
rect 10100 14764 10106 14776
rect 10318 14764 10324 14776
rect 10376 14804 10382 14816
rect 12912 14804 12940 14844
rect 13817 14841 13829 14844
rect 13863 14841 13875 14875
rect 13817 14835 13875 14841
rect 10376 14776 12940 14804
rect 10376 14764 10382 14776
rect 13262 14764 13268 14816
rect 13320 14804 13326 14816
rect 14829 14807 14887 14813
rect 14829 14804 14841 14807
rect 13320 14776 14841 14804
rect 13320 14764 13326 14776
rect 14829 14773 14841 14776
rect 14875 14773 14887 14807
rect 14829 14767 14887 14773
rect 1104 14714 15824 14736
rect 1104 14662 5912 14714
rect 5964 14662 5976 14714
rect 6028 14662 6040 14714
rect 6092 14662 6104 14714
rect 6156 14662 10843 14714
rect 10895 14662 10907 14714
rect 10959 14662 10971 14714
rect 11023 14662 11035 14714
rect 11087 14662 15824 14714
rect 1104 14640 15824 14662
rect 2869 14603 2927 14609
rect 2869 14569 2881 14603
rect 2915 14600 2927 14603
rect 2958 14600 2964 14612
rect 2915 14572 2964 14600
rect 2915 14569 2927 14572
rect 2869 14563 2927 14569
rect 2958 14560 2964 14572
rect 3016 14560 3022 14612
rect 5718 14560 5724 14612
rect 5776 14600 5782 14612
rect 5813 14603 5871 14609
rect 5813 14600 5825 14603
rect 5776 14572 5825 14600
rect 5776 14560 5782 14572
rect 5813 14569 5825 14572
rect 5859 14569 5871 14603
rect 6270 14600 6276 14612
rect 6231 14572 6276 14600
rect 5813 14563 5871 14569
rect 6270 14560 6276 14572
rect 6328 14600 6334 14612
rect 7374 14600 7380 14612
rect 6328 14572 7380 14600
rect 6328 14560 6334 14572
rect 7374 14560 7380 14572
rect 7432 14560 7438 14612
rect 7561 14603 7619 14609
rect 7561 14569 7573 14603
rect 7607 14600 7619 14603
rect 7926 14600 7932 14612
rect 7607 14572 7932 14600
rect 7607 14569 7619 14572
rect 7561 14563 7619 14569
rect 7926 14560 7932 14572
rect 7984 14560 7990 14612
rect 8573 14603 8631 14609
rect 8573 14569 8585 14603
rect 8619 14569 8631 14603
rect 8573 14563 8631 14569
rect 3418 14532 3424 14544
rect 3379 14504 3424 14532
rect 3418 14492 3424 14504
rect 3476 14492 3482 14544
rect 4062 14492 4068 14544
rect 4120 14532 4126 14544
rect 4402 14535 4460 14541
rect 4402 14532 4414 14535
rect 4120 14504 4414 14532
rect 4120 14492 4126 14504
rect 4402 14501 4414 14504
rect 4448 14501 4460 14535
rect 8588 14532 8616 14563
rect 8754 14560 8760 14612
rect 8812 14600 8818 14612
rect 14642 14600 14648 14612
rect 8812 14572 14648 14600
rect 8812 14560 8818 14572
rect 14642 14560 14648 14572
rect 14700 14560 14706 14612
rect 4402 14495 4460 14501
rect 5828 14504 8616 14532
rect 9033 14535 9091 14541
rect 1486 14464 1492 14476
rect 1447 14436 1492 14464
rect 1486 14424 1492 14436
rect 1544 14424 1550 14476
rect 1756 14467 1814 14473
rect 1756 14433 1768 14467
rect 1802 14464 1814 14467
rect 2682 14464 2688 14476
rect 1802 14436 2688 14464
rect 1802 14433 1814 14436
rect 1756 14427 1814 14433
rect 2682 14424 2688 14436
rect 2740 14424 2746 14476
rect 3145 14467 3203 14473
rect 3145 14433 3157 14467
rect 3191 14464 3203 14467
rect 5828 14464 5856 14504
rect 9033 14501 9045 14535
rect 9079 14532 9091 14535
rect 10594 14532 10600 14544
rect 9079 14504 10600 14532
rect 9079 14501 9091 14504
rect 9033 14495 9091 14501
rect 10594 14492 10600 14504
rect 10652 14492 10658 14544
rect 11333 14535 11391 14541
rect 11333 14501 11345 14535
rect 11379 14532 11391 14535
rect 11784 14535 11842 14541
rect 11784 14532 11796 14535
rect 11379 14504 11796 14532
rect 11379 14501 11391 14504
rect 11333 14495 11391 14501
rect 11784 14501 11796 14504
rect 11830 14532 11842 14535
rect 12986 14532 12992 14544
rect 11830 14504 12992 14532
rect 11830 14501 11842 14504
rect 11784 14495 11842 14501
rect 12986 14492 12992 14504
rect 13044 14492 13050 14544
rect 13998 14532 14004 14544
rect 13959 14504 14004 14532
rect 13998 14492 14004 14504
rect 14056 14492 14062 14544
rect 3191 14436 5856 14464
rect 6181 14467 6239 14473
rect 3191 14433 3203 14436
rect 3145 14427 3203 14433
rect 6181 14433 6193 14467
rect 6227 14464 6239 14467
rect 7006 14464 7012 14476
rect 6227 14436 7012 14464
rect 6227 14433 6239 14436
rect 6181 14427 6239 14433
rect 7006 14424 7012 14436
rect 7064 14464 7070 14476
rect 7466 14464 7472 14476
rect 7064 14436 7472 14464
rect 7064 14424 7070 14436
rect 7466 14424 7472 14436
rect 7524 14424 7530 14476
rect 7929 14467 7987 14473
rect 7929 14433 7941 14467
rect 7975 14464 7987 14467
rect 8110 14464 8116 14476
rect 7975 14436 8116 14464
rect 7975 14433 7987 14436
rect 7929 14427 7987 14433
rect 8110 14424 8116 14436
rect 8168 14424 8174 14476
rect 8941 14467 8999 14473
rect 8941 14433 8953 14467
rect 8987 14464 8999 14467
rect 9950 14464 9956 14476
rect 8987 14436 9956 14464
rect 8987 14433 8999 14436
rect 8941 14427 8999 14433
rect 9950 14424 9956 14436
rect 10008 14424 10014 14476
rect 10128 14467 10186 14473
rect 10128 14433 10140 14467
rect 10174 14464 10186 14467
rect 11606 14464 11612 14476
rect 10174 14436 11612 14464
rect 10174 14433 10186 14436
rect 10128 14427 10186 14433
rect 11606 14424 11612 14436
rect 11664 14424 11670 14476
rect 4154 14396 4160 14408
rect 4115 14368 4160 14396
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 6365 14399 6423 14405
rect 6365 14365 6377 14399
rect 6411 14365 6423 14399
rect 6365 14359 6423 14365
rect 8021 14399 8079 14405
rect 8021 14365 8033 14399
rect 8067 14365 8079 14399
rect 8021 14359 8079 14365
rect 8205 14399 8263 14405
rect 8205 14365 8217 14399
rect 8251 14365 8263 14399
rect 8205 14359 8263 14365
rect 5537 14331 5595 14337
rect 5537 14297 5549 14331
rect 5583 14328 5595 14331
rect 6178 14328 6184 14340
rect 5583 14300 6184 14328
rect 5583 14297 5595 14300
rect 5537 14291 5595 14297
rect 6178 14288 6184 14300
rect 6236 14328 6242 14340
rect 6380 14328 6408 14359
rect 6236 14300 6408 14328
rect 6236 14288 6242 14300
rect 3234 14220 3240 14272
rect 3292 14260 3298 14272
rect 4338 14260 4344 14272
rect 3292 14232 4344 14260
rect 3292 14220 3298 14232
rect 4338 14220 4344 14232
rect 4396 14260 4402 14272
rect 5718 14260 5724 14272
rect 4396 14232 5724 14260
rect 4396 14220 4402 14232
rect 5718 14220 5724 14232
rect 5776 14260 5782 14272
rect 8036 14260 8064 14359
rect 8220 14328 8248 14359
rect 9122 14356 9128 14408
rect 9180 14396 9186 14408
rect 9861 14399 9919 14405
rect 9180 14368 9225 14396
rect 9180 14356 9186 14368
rect 9861 14365 9873 14399
rect 9907 14365 9919 14399
rect 11517 14399 11575 14405
rect 11517 14396 11529 14399
rect 9861 14359 9919 14365
rect 10888 14368 11529 14396
rect 8938 14328 8944 14340
rect 8220 14300 8944 14328
rect 8938 14288 8944 14300
rect 8996 14288 9002 14340
rect 9030 14288 9036 14340
rect 9088 14328 9094 14340
rect 9876 14328 9904 14359
rect 9088 14300 9904 14328
rect 9088 14288 9094 14300
rect 5776 14232 8064 14260
rect 9876 14260 9904 14300
rect 10502 14260 10508 14272
rect 9876 14232 10508 14260
rect 5776 14220 5782 14232
rect 10502 14220 10508 14232
rect 10560 14260 10566 14272
rect 10888 14260 10916 14368
rect 11517 14365 11529 14368
rect 11563 14365 11575 14399
rect 11517 14359 11575 14365
rect 13722 14356 13728 14408
rect 13780 14396 13786 14408
rect 13909 14399 13967 14405
rect 13909 14396 13921 14399
rect 13780 14368 13921 14396
rect 13780 14356 13786 14368
rect 13909 14365 13921 14368
rect 13955 14365 13967 14399
rect 13909 14359 13967 14365
rect 14185 14399 14243 14405
rect 14185 14365 14197 14399
rect 14231 14365 14243 14399
rect 14185 14359 14243 14365
rect 11241 14331 11299 14337
rect 11241 14297 11253 14331
rect 11287 14328 11299 14331
rect 11333 14331 11391 14337
rect 11333 14328 11345 14331
rect 11287 14300 11345 14328
rect 11287 14297 11299 14300
rect 11241 14291 11299 14297
rect 11333 14297 11345 14300
rect 11379 14297 11391 14331
rect 14200 14328 14228 14359
rect 11333 14291 11391 14297
rect 12728 14300 14228 14328
rect 10560 14232 10916 14260
rect 10560 14220 10566 14232
rect 10962 14220 10968 14272
rect 11020 14260 11026 14272
rect 12728 14260 12756 14300
rect 11020 14232 12756 14260
rect 12897 14263 12955 14269
rect 11020 14220 11026 14232
rect 12897 14229 12909 14263
rect 12943 14260 12955 14263
rect 12986 14260 12992 14272
rect 12943 14232 12992 14260
rect 12943 14229 12955 14232
rect 12897 14223 12955 14229
rect 12986 14220 12992 14232
rect 13044 14260 13050 14272
rect 14090 14260 14096 14272
rect 13044 14232 14096 14260
rect 13044 14220 13050 14232
rect 14090 14220 14096 14232
rect 14148 14220 14154 14272
rect 1104 14170 15824 14192
rect 1104 14118 3447 14170
rect 3499 14118 3511 14170
rect 3563 14118 3575 14170
rect 3627 14118 3639 14170
rect 3691 14118 8378 14170
rect 8430 14118 8442 14170
rect 8494 14118 8506 14170
rect 8558 14118 8570 14170
rect 8622 14118 13308 14170
rect 13360 14118 13372 14170
rect 13424 14118 13436 14170
rect 13488 14118 13500 14170
rect 13552 14118 15824 14170
rect 1104 14096 15824 14118
rect 1946 14056 1952 14068
rect 1907 14028 1952 14056
rect 1946 14016 1952 14028
rect 2004 14016 2010 14068
rect 2961 14059 3019 14065
rect 2961 14025 2973 14059
rect 3007 14025 3019 14059
rect 3970 14056 3976 14068
rect 3931 14028 3976 14056
rect 2961 14019 3019 14025
rect 2976 13988 3004 14019
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 4154 14016 4160 14068
rect 4212 14056 4218 14068
rect 5074 14056 5080 14068
rect 4212 14028 5080 14056
rect 4212 14016 4218 14028
rect 5074 14016 5080 14028
rect 5132 14056 5138 14068
rect 5537 14059 5595 14065
rect 5132 14028 5488 14056
rect 5132 14016 5138 14028
rect 5460 14000 5488 14028
rect 5537 14025 5549 14059
rect 5583 14056 5595 14059
rect 5810 14056 5816 14068
rect 5583 14028 5816 14056
rect 5583 14025 5595 14028
rect 5537 14019 5595 14025
rect 5810 14016 5816 14028
rect 5868 14016 5874 14068
rect 5902 14016 5908 14068
rect 5960 14056 5966 14068
rect 9674 14056 9680 14068
rect 5960 14028 9680 14056
rect 5960 14016 5966 14028
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 9950 14016 9956 14068
rect 10008 14056 10014 14068
rect 11241 14059 11299 14065
rect 11241 14056 11253 14059
rect 10008 14028 11253 14056
rect 10008 14016 10014 14028
rect 11241 14025 11253 14028
rect 11287 14025 11299 14059
rect 11241 14019 11299 14025
rect 13998 14016 14004 14068
rect 14056 14056 14062 14068
rect 14875 14059 14933 14065
rect 14875 14056 14887 14059
rect 14056 14028 14887 14056
rect 14056 14016 14062 14028
rect 14875 14025 14887 14028
rect 14921 14025 14933 14059
rect 14875 14019 14933 14025
rect 5258 13988 5264 14000
rect 2516 13960 3004 13988
rect 3436 13960 5264 13988
rect 2317 13855 2375 13861
rect 2317 13821 2329 13855
rect 2363 13852 2375 13855
rect 2516 13852 2544 13960
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13920 2651 13923
rect 2958 13920 2964 13932
rect 2639 13892 2964 13920
rect 2639 13889 2651 13892
rect 2593 13883 2651 13889
rect 2958 13880 2964 13892
rect 3016 13880 3022 13932
rect 3436 13929 3464 13960
rect 5258 13948 5264 13960
rect 5316 13948 5322 14000
rect 5442 13948 5448 14000
rect 5500 13988 5506 14000
rect 10413 13991 10471 13997
rect 10413 13988 10425 13991
rect 5500 13960 6868 13988
rect 5500 13948 5506 13960
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13889 3479 13923
rect 3421 13883 3479 13889
rect 3513 13923 3571 13929
rect 3513 13889 3525 13923
rect 3559 13920 3571 13923
rect 4522 13920 4528 13932
rect 3559 13892 4528 13920
rect 3559 13889 3571 13892
rect 3513 13883 3571 13889
rect 2363 13824 2544 13852
rect 2363 13821 2375 13824
rect 2317 13815 2375 13821
rect 2682 13812 2688 13864
rect 2740 13852 2746 13864
rect 3234 13852 3240 13864
rect 2740 13824 3240 13852
rect 2740 13812 2746 13824
rect 3234 13812 3240 13824
rect 3292 13852 3298 13864
rect 3528 13852 3556 13883
rect 4522 13880 4528 13892
rect 4580 13880 4586 13932
rect 4706 13880 4712 13932
rect 4764 13920 4770 13932
rect 4985 13923 5043 13929
rect 4985 13920 4997 13923
rect 4764 13892 4997 13920
rect 4764 13880 4770 13892
rect 4985 13889 4997 13892
rect 5031 13889 5043 13923
rect 4985 13883 5043 13889
rect 5718 13880 5724 13932
rect 5776 13920 5782 13932
rect 5997 13923 6055 13929
rect 5997 13920 6009 13923
rect 5776 13892 6009 13920
rect 5776 13880 5782 13892
rect 5997 13889 6009 13892
rect 6043 13889 6055 13923
rect 6178 13920 6184 13932
rect 6139 13892 6184 13920
rect 5997 13883 6055 13889
rect 6178 13880 6184 13892
rect 6236 13920 6242 13932
rect 6840 13929 6868 13960
rect 10060 13960 10425 13988
rect 6825 13923 6883 13929
rect 6236 13892 6776 13920
rect 6236 13880 6242 13892
rect 3292 13824 3556 13852
rect 4433 13855 4491 13861
rect 3292 13812 3298 13824
rect 4433 13821 4445 13855
rect 4479 13852 4491 13855
rect 4890 13852 4896 13864
rect 4479 13824 4896 13852
rect 4479 13821 4491 13824
rect 4433 13815 4491 13821
rect 4890 13812 4896 13824
rect 4948 13852 4954 13864
rect 5810 13852 5816 13864
rect 4948 13824 5816 13852
rect 4948 13812 4954 13824
rect 5810 13812 5816 13824
rect 5868 13812 5874 13864
rect 5905 13855 5963 13861
rect 5905 13821 5917 13855
rect 5951 13852 5963 13855
rect 6748 13852 6776 13892
rect 6825 13889 6837 13923
rect 6871 13889 6883 13923
rect 6825 13883 6883 13889
rect 7081 13855 7139 13861
rect 7081 13852 7093 13855
rect 5951 13824 6500 13852
rect 6748 13824 7093 13852
rect 5951 13821 5963 13824
rect 5905 13815 5963 13821
rect 3326 13784 3332 13796
rect 3287 13756 3332 13784
rect 3326 13744 3332 13756
rect 3384 13744 3390 13796
rect 4341 13787 4399 13793
rect 4341 13753 4353 13787
rect 4387 13784 4399 13787
rect 4706 13784 4712 13796
rect 4387 13756 4712 13784
rect 4387 13753 4399 13756
rect 4341 13747 4399 13753
rect 4706 13744 4712 13756
rect 4764 13784 4770 13796
rect 6362 13784 6368 13796
rect 4764 13756 6368 13784
rect 4764 13744 4770 13756
rect 6362 13744 6368 13756
rect 6420 13744 6426 13796
rect 6472 13784 6500 13824
rect 7081 13821 7093 13824
rect 7127 13821 7139 13855
rect 7081 13815 7139 13821
rect 8662 13812 8668 13864
rect 8720 13852 8726 13864
rect 9030 13852 9036 13864
rect 8720 13824 9036 13852
rect 8720 13812 8726 13824
rect 9030 13812 9036 13824
rect 9088 13812 9094 13864
rect 9122 13812 9128 13864
rect 9180 13852 9186 13864
rect 10060 13852 10088 13960
rect 10413 13957 10425 13960
rect 10459 13957 10471 13991
rect 10413 13951 10471 13957
rect 10502 13948 10508 14000
rect 10560 13988 10566 14000
rect 10689 13991 10747 13997
rect 10689 13988 10701 13991
rect 10560 13960 10701 13988
rect 10560 13948 10566 13960
rect 10689 13957 10701 13960
rect 10735 13988 10747 13991
rect 12158 13988 12164 14000
rect 10735 13960 12164 13988
rect 10735 13957 10747 13960
rect 10689 13951 10747 13957
rect 12158 13948 12164 13960
rect 12216 13988 12222 14000
rect 14461 13991 14519 13997
rect 12216 13960 13124 13988
rect 12216 13948 12222 13960
rect 11606 13920 11612 13932
rect 9180 13824 10088 13852
rect 10152 13892 11612 13920
rect 9180 13812 9186 13824
rect 7190 13784 7196 13796
rect 6472 13756 7196 13784
rect 7190 13744 7196 13756
rect 7248 13784 7254 13796
rect 8110 13784 8116 13796
rect 7248 13756 8116 13784
rect 7248 13744 7254 13756
rect 8110 13744 8116 13756
rect 8168 13744 8174 13796
rect 9300 13787 9358 13793
rect 9300 13753 9312 13787
rect 9346 13784 9358 13787
rect 10152 13784 10180 13892
rect 11606 13880 11612 13892
rect 11664 13920 11670 13932
rect 11793 13923 11851 13929
rect 11793 13920 11805 13923
rect 11664 13892 11805 13920
rect 11664 13880 11670 13892
rect 11793 13889 11805 13892
rect 11839 13889 11851 13923
rect 13096 13920 13124 13960
rect 14461 13957 14473 13991
rect 14507 13988 14519 13991
rect 14550 13988 14556 14000
rect 14507 13960 14556 13988
rect 14507 13957 14519 13960
rect 14461 13951 14519 13957
rect 14550 13948 14556 13960
rect 14608 13948 14614 14000
rect 13096 13892 13216 13920
rect 11793 13883 11851 13889
rect 10226 13812 10232 13864
rect 10284 13852 10290 13864
rect 10873 13855 10931 13861
rect 10873 13852 10885 13855
rect 10284 13824 10885 13852
rect 10284 13812 10290 13824
rect 10873 13821 10885 13824
rect 10919 13821 10931 13855
rect 10873 13815 10931 13821
rect 11701 13855 11759 13861
rect 11701 13821 11713 13855
rect 11747 13852 11759 13855
rect 12434 13852 12440 13864
rect 11747 13824 12440 13852
rect 11747 13821 11759 13824
rect 11701 13815 11759 13821
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 13081 13855 13139 13861
rect 13081 13821 13093 13855
rect 13127 13852 13139 13855
rect 13188 13852 13216 13892
rect 13127 13824 13216 13852
rect 14804 13855 14862 13861
rect 13127 13821 13139 13824
rect 13081 13815 13139 13821
rect 14804 13821 14816 13855
rect 14850 13852 14862 13855
rect 15010 13852 15016 13864
rect 14850 13824 15016 13852
rect 14850 13821 14862 13824
rect 14804 13815 14862 13821
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 9346 13756 10180 13784
rect 9346 13753 9358 13756
rect 9300 13747 9358 13753
rect 12986 13744 12992 13796
rect 13044 13784 13050 13796
rect 13348 13787 13406 13793
rect 13348 13784 13360 13787
rect 13044 13756 13360 13784
rect 13044 13744 13050 13756
rect 13348 13753 13360 13756
rect 13394 13784 13406 13787
rect 13538 13784 13544 13796
rect 13394 13756 13544 13784
rect 13394 13753 13406 13756
rect 13348 13747 13406 13753
rect 13538 13744 13544 13756
rect 13596 13744 13602 13796
rect 14642 13744 14648 13796
rect 14700 13784 14706 13796
rect 15562 13784 15568 13796
rect 14700 13756 15568 13784
rect 14700 13744 14706 13756
rect 15562 13744 15568 13756
rect 15620 13744 15626 13796
rect 2406 13676 2412 13728
rect 2464 13716 2470 13728
rect 2464 13688 2509 13716
rect 2464 13676 2470 13688
rect 7466 13676 7472 13728
rect 7524 13716 7530 13728
rect 8205 13719 8263 13725
rect 8205 13716 8217 13719
rect 7524 13688 8217 13716
rect 7524 13676 7530 13688
rect 8205 13685 8217 13688
rect 8251 13685 8263 13719
rect 8205 13679 8263 13685
rect 11609 13719 11667 13725
rect 11609 13685 11621 13719
rect 11655 13716 11667 13719
rect 11974 13716 11980 13728
rect 11655 13688 11980 13716
rect 11655 13685 11667 13688
rect 11609 13679 11667 13685
rect 11974 13676 11980 13688
rect 12032 13676 12038 13728
rect 1104 13626 15824 13648
rect 1104 13574 5912 13626
rect 5964 13574 5976 13626
rect 6028 13574 6040 13626
rect 6092 13574 6104 13626
rect 6156 13574 10843 13626
rect 10895 13574 10907 13626
rect 10959 13574 10971 13626
rect 11023 13574 11035 13626
rect 11087 13574 15824 13626
rect 1104 13552 15824 13574
rect 2406 13472 2412 13524
rect 2464 13512 2470 13524
rect 2685 13515 2743 13521
rect 2685 13512 2697 13515
rect 2464 13484 2697 13512
rect 2464 13472 2470 13484
rect 2685 13481 2697 13484
rect 2731 13481 2743 13515
rect 2685 13475 2743 13481
rect 5077 13515 5135 13521
rect 5077 13481 5089 13515
rect 5123 13512 5135 13515
rect 5350 13512 5356 13524
rect 5123 13484 5356 13512
rect 5123 13481 5135 13484
rect 5077 13475 5135 13481
rect 5350 13472 5356 13484
rect 5408 13472 5414 13524
rect 5997 13515 6055 13521
rect 5997 13481 6009 13515
rect 6043 13512 6055 13515
rect 6454 13512 6460 13524
rect 6043 13484 6460 13512
rect 6043 13481 6055 13484
rect 5997 13475 6055 13481
rect 6454 13472 6460 13484
rect 6512 13472 6518 13524
rect 8938 13512 8944 13524
rect 8899 13484 8944 13512
rect 8938 13472 8944 13484
rect 8996 13472 9002 13524
rect 9309 13515 9367 13521
rect 9309 13481 9321 13515
rect 9355 13512 9367 13515
rect 10226 13512 10232 13524
rect 9355 13484 10232 13512
rect 9355 13481 9367 13484
rect 9309 13475 9367 13481
rect 10226 13472 10232 13484
rect 10284 13472 10290 13524
rect 11606 13472 11612 13524
rect 11664 13512 11670 13524
rect 11701 13515 11759 13521
rect 11701 13512 11713 13515
rect 11664 13484 11713 13512
rect 11664 13472 11670 13484
rect 11701 13481 11713 13484
rect 11747 13481 11759 13515
rect 11974 13512 11980 13524
rect 11935 13484 11980 13512
rect 11701 13475 11759 13481
rect 11974 13472 11980 13484
rect 12032 13472 12038 13524
rect 14001 13515 14059 13521
rect 12084 13484 13492 13512
rect 2314 13404 2320 13456
rect 2372 13444 2378 13456
rect 3053 13447 3111 13453
rect 3053 13444 3065 13447
rect 2372 13416 3065 13444
rect 2372 13404 2378 13416
rect 3053 13413 3065 13416
rect 3099 13413 3111 13447
rect 3053 13407 3111 13413
rect 3878 13404 3884 13456
rect 3936 13444 3942 13456
rect 6089 13447 6147 13453
rect 6089 13444 6101 13447
rect 3936 13416 6101 13444
rect 3936 13404 3942 13416
rect 6089 13413 6101 13416
rect 6135 13413 6147 13447
rect 6089 13407 6147 13413
rect 7392 13416 9536 13444
rect 1762 13336 1768 13388
rect 1820 13376 1826 13388
rect 2041 13379 2099 13385
rect 2041 13376 2053 13379
rect 1820 13348 2053 13376
rect 1820 13336 1826 13348
rect 2041 13345 2053 13348
rect 2087 13345 2099 13379
rect 2041 13339 2099 13345
rect 4985 13379 5043 13385
rect 4985 13345 4997 13379
rect 5031 13376 5043 13379
rect 5350 13376 5356 13388
rect 5031 13348 5356 13376
rect 5031 13345 5043 13348
rect 4985 13339 5043 13345
rect 5350 13336 5356 13348
rect 5408 13336 5414 13388
rect 2130 13308 2136 13320
rect 2091 13280 2136 13308
rect 2130 13268 2136 13280
rect 2188 13268 2194 13320
rect 2222 13268 2228 13320
rect 2280 13308 2286 13320
rect 3142 13308 3148 13320
rect 2280 13280 2325 13308
rect 3103 13280 3148 13308
rect 2280 13268 2286 13280
rect 3142 13268 3148 13280
rect 3200 13268 3206 13320
rect 3234 13268 3240 13320
rect 3292 13308 3298 13320
rect 5261 13311 5319 13317
rect 3292 13280 3337 13308
rect 3292 13268 3298 13280
rect 5261 13277 5273 13311
rect 5307 13308 5319 13311
rect 5718 13308 5724 13320
rect 5307 13280 5724 13308
rect 5307 13277 5319 13280
rect 5261 13271 5319 13277
rect 5718 13268 5724 13280
rect 5776 13268 5782 13320
rect 6270 13308 6276 13320
rect 6231 13280 6276 13308
rect 6270 13268 6276 13280
rect 6328 13268 6334 13320
rect 1673 13243 1731 13249
rect 1673 13209 1685 13243
rect 1719 13240 1731 13243
rect 5534 13240 5540 13252
rect 1719 13212 5540 13240
rect 1719 13209 1731 13212
rect 1673 13203 1731 13209
rect 5534 13200 5540 13212
rect 5592 13200 5598 13252
rect 6638 13200 6644 13252
rect 6696 13240 6702 13252
rect 7285 13243 7343 13249
rect 7285 13240 7297 13243
rect 6696 13212 7297 13240
rect 6696 13200 6702 13212
rect 7285 13209 7297 13212
rect 7331 13240 7343 13243
rect 7392 13240 7420 13416
rect 7469 13379 7527 13385
rect 7469 13345 7481 13379
rect 7515 13376 7527 13379
rect 7650 13376 7656 13388
rect 7515 13348 7656 13376
rect 7515 13345 7527 13348
rect 7469 13339 7527 13345
rect 7650 13336 7656 13348
rect 7708 13336 7714 13388
rect 7828 13379 7886 13385
rect 7828 13345 7840 13379
rect 7874 13376 7886 13379
rect 9122 13376 9128 13388
rect 7874 13348 9128 13376
rect 7874 13345 7886 13348
rect 7828 13339 7886 13345
rect 9122 13336 9128 13348
rect 9180 13336 9186 13388
rect 9508 13385 9536 13416
rect 9582 13404 9588 13456
rect 9640 13444 9646 13456
rect 12084 13444 12112 13484
rect 9640 13416 12112 13444
rect 12345 13447 12403 13453
rect 9640 13404 9646 13416
rect 12345 13413 12357 13447
rect 12391 13444 12403 13447
rect 12526 13444 12532 13456
rect 12391 13416 12532 13444
rect 12391 13413 12403 13416
rect 12345 13407 12403 13413
rect 12526 13404 12532 13416
rect 12584 13404 12590 13456
rect 13464 13444 13492 13484
rect 14001 13481 14013 13515
rect 14047 13512 14059 13515
rect 14274 13512 14280 13524
rect 14047 13484 14280 13512
rect 14047 13481 14059 13484
rect 14001 13475 14059 13481
rect 14274 13472 14280 13484
rect 14332 13472 14338 13524
rect 14461 13447 14519 13453
rect 14461 13444 14473 13447
rect 13464 13416 14473 13444
rect 14461 13413 14473 13416
rect 14507 13413 14519 13447
rect 14461 13407 14519 13413
rect 9493 13379 9551 13385
rect 9493 13345 9505 13379
rect 9539 13345 9551 13379
rect 9493 13339 9551 13345
rect 10321 13379 10379 13385
rect 10321 13345 10333 13379
rect 10367 13376 10379 13379
rect 10410 13376 10416 13388
rect 10367 13348 10416 13376
rect 10367 13345 10379 13348
rect 10321 13339 10379 13345
rect 10410 13336 10416 13348
rect 10468 13336 10474 13388
rect 10588 13379 10646 13385
rect 10588 13345 10600 13379
rect 10634 13376 10646 13379
rect 10870 13376 10876 13388
rect 10634 13348 10876 13376
rect 10634 13345 10646 13348
rect 10588 13339 10646 13345
rect 10870 13336 10876 13348
rect 10928 13376 10934 13388
rect 12250 13376 12256 13388
rect 10928 13348 12256 13376
rect 10928 13336 10934 13348
rect 12250 13336 12256 13348
rect 12308 13376 12314 13388
rect 12308 13348 12572 13376
rect 12308 13336 12314 13348
rect 12544 13317 12572 13348
rect 12986 13336 12992 13388
rect 13044 13376 13050 13388
rect 13357 13379 13415 13385
rect 13357 13376 13369 13379
rect 13044 13348 13369 13376
rect 13044 13336 13050 13348
rect 13357 13345 13369 13348
rect 13403 13345 13415 13379
rect 13357 13339 13415 13345
rect 13722 13336 13728 13388
rect 13780 13376 13786 13388
rect 14369 13379 14427 13385
rect 14369 13376 14381 13379
rect 13780 13348 14381 13376
rect 13780 13336 13786 13348
rect 14369 13345 14381 13348
rect 14415 13345 14427 13379
rect 14369 13339 14427 13345
rect 7561 13311 7619 13317
rect 7561 13277 7573 13311
rect 7607 13277 7619 13311
rect 7561 13271 7619 13277
rect 12437 13311 12495 13317
rect 12437 13277 12449 13311
rect 12483 13277 12495 13311
rect 12437 13271 12495 13277
rect 12529 13311 12587 13317
rect 12529 13277 12541 13311
rect 12575 13277 12587 13311
rect 12529 13271 12587 13277
rect 13449 13311 13507 13317
rect 13449 13277 13461 13311
rect 13495 13277 13507 13311
rect 13449 13271 13507 13277
rect 7331 13212 7420 13240
rect 7331 13209 7343 13212
rect 7285 13203 7343 13209
rect 1578 13132 1584 13184
rect 1636 13172 1642 13184
rect 3970 13172 3976 13184
rect 1636 13144 3976 13172
rect 1636 13132 1642 13144
rect 3970 13132 3976 13144
rect 4028 13132 4034 13184
rect 4614 13172 4620 13184
rect 4575 13144 4620 13172
rect 4614 13132 4620 13144
rect 4672 13132 4678 13184
rect 5629 13175 5687 13181
rect 5629 13141 5641 13175
rect 5675 13172 5687 13175
rect 5810 13172 5816 13184
rect 5675 13144 5816 13172
rect 5675 13141 5687 13144
rect 5629 13135 5687 13141
rect 5810 13132 5816 13144
rect 5868 13132 5874 13184
rect 7576 13172 7604 13271
rect 9030 13172 9036 13184
rect 7576 13144 9036 13172
rect 9030 13132 9036 13144
rect 9088 13132 9094 13184
rect 12452 13172 12480 13271
rect 12989 13243 13047 13249
rect 12989 13209 13001 13243
rect 13035 13240 13047 13243
rect 13078 13240 13084 13252
rect 13035 13212 13084 13240
rect 13035 13209 13047 13212
rect 12989 13203 13047 13209
rect 13078 13200 13084 13212
rect 13136 13200 13142 13252
rect 13464 13240 13492 13271
rect 13538 13268 13544 13320
rect 13596 13308 13602 13320
rect 14553 13311 14611 13317
rect 14553 13308 14565 13311
rect 13596 13280 14565 13308
rect 13596 13268 13602 13280
rect 14553 13277 14565 13280
rect 14599 13277 14611 13311
rect 14553 13271 14611 13277
rect 13998 13240 14004 13252
rect 13464 13212 14004 13240
rect 13998 13200 14004 13212
rect 14056 13200 14062 13252
rect 14642 13172 14648 13184
rect 12452 13144 14648 13172
rect 14642 13132 14648 13144
rect 14700 13132 14706 13184
rect 1104 13082 15824 13104
rect 1104 13030 3447 13082
rect 3499 13030 3511 13082
rect 3563 13030 3575 13082
rect 3627 13030 3639 13082
rect 3691 13030 8378 13082
rect 8430 13030 8442 13082
rect 8494 13030 8506 13082
rect 8558 13030 8570 13082
rect 8622 13030 13308 13082
rect 13360 13030 13372 13082
rect 13424 13030 13436 13082
rect 13488 13030 13500 13082
rect 13552 13030 15824 13082
rect 1104 13008 15824 13030
rect 2133 12971 2191 12977
rect 2133 12937 2145 12971
rect 2179 12968 2191 12971
rect 3142 12968 3148 12980
rect 2179 12940 3148 12968
rect 2179 12937 2191 12940
rect 2133 12931 2191 12937
rect 3142 12928 3148 12940
rect 3200 12928 3206 12980
rect 3786 12928 3792 12980
rect 3844 12968 3850 12980
rect 4062 12968 4068 12980
rect 3844 12940 4068 12968
rect 3844 12928 3850 12940
rect 4062 12928 4068 12940
rect 4120 12928 4126 12980
rect 4522 12968 4528 12980
rect 4483 12940 4528 12968
rect 4522 12928 4528 12940
rect 4580 12928 4586 12980
rect 5350 12968 5356 12980
rect 5311 12940 5356 12968
rect 5350 12928 5356 12940
rect 5408 12928 5414 12980
rect 10594 12928 10600 12980
rect 10652 12968 10658 12980
rect 10873 12971 10931 12977
rect 10873 12968 10885 12971
rect 10652 12940 10885 12968
rect 10652 12928 10658 12940
rect 10873 12937 10885 12940
rect 10919 12937 10931 12971
rect 10873 12931 10931 12937
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 12492 12940 12537 12968
rect 12492 12928 12498 12940
rect 12710 12928 12716 12980
rect 12768 12968 12774 12980
rect 13170 12968 13176 12980
rect 12768 12940 13176 12968
rect 12768 12928 12774 12940
rect 13170 12928 13176 12940
rect 13228 12928 13234 12980
rect 5902 12860 5908 12912
rect 5960 12900 5966 12912
rect 5960 12872 6040 12900
rect 5960 12860 5966 12872
rect 1578 12832 1584 12844
rect 1539 12804 1584 12832
rect 1578 12792 1584 12804
rect 1636 12792 1642 12844
rect 1670 12792 1676 12844
rect 1728 12832 1734 12844
rect 2593 12835 2651 12841
rect 2593 12832 2605 12835
rect 1728 12804 2605 12832
rect 1728 12792 1734 12804
rect 2593 12801 2605 12804
rect 2639 12801 2651 12835
rect 2593 12795 2651 12801
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12832 2835 12835
rect 5810 12832 5816 12844
rect 2823 12804 3280 12832
rect 5771 12804 5816 12832
rect 2823 12801 2835 12804
rect 2777 12795 2835 12801
rect 3252 12776 3280 12804
rect 5810 12792 5816 12804
rect 5868 12792 5874 12844
rect 6012 12841 6040 12872
rect 6730 12860 6736 12912
rect 6788 12900 6794 12912
rect 7926 12900 7932 12912
rect 6788 12872 7932 12900
rect 6788 12860 6794 12872
rect 7926 12860 7932 12872
rect 7984 12860 7990 12912
rect 9140 12872 11376 12900
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12832 6055 12835
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 6043 12804 7389 12832
rect 6043 12801 6055 12804
rect 5997 12795 6055 12801
rect 7377 12801 7389 12804
rect 7423 12832 7435 12835
rect 7466 12832 7472 12844
rect 7423 12804 7472 12832
rect 7423 12801 7435 12804
rect 7377 12795 7435 12801
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 1394 12764 1400 12776
rect 1355 12736 1400 12764
rect 1394 12724 1400 12736
rect 1452 12724 1458 12776
rect 2866 12724 2872 12776
rect 2924 12764 2930 12776
rect 3145 12767 3203 12773
rect 3145 12764 3157 12767
rect 2924 12736 3157 12764
rect 2924 12724 2930 12736
rect 3145 12733 3157 12736
rect 3191 12733 3203 12767
rect 3145 12727 3203 12733
rect 3234 12724 3240 12776
rect 3292 12764 3298 12776
rect 3401 12767 3459 12773
rect 3401 12764 3413 12767
rect 3292 12736 3413 12764
rect 3292 12724 3298 12736
rect 3401 12733 3413 12736
rect 3447 12733 3459 12767
rect 6362 12764 6368 12776
rect 3401 12727 3459 12733
rect 5644 12736 6368 12764
rect 2501 12699 2559 12705
rect 2501 12665 2513 12699
rect 2547 12696 2559 12699
rect 5644 12696 5672 12736
rect 6362 12724 6368 12736
rect 6420 12724 6426 12776
rect 6549 12767 6607 12773
rect 6549 12733 6561 12767
rect 6595 12764 6607 12767
rect 6638 12764 6644 12776
rect 6595 12736 6644 12764
rect 6595 12733 6607 12736
rect 6549 12727 6607 12733
rect 6638 12724 6644 12736
rect 6696 12724 6702 12776
rect 6822 12724 6828 12776
rect 6880 12724 6886 12776
rect 7190 12724 7196 12776
rect 7248 12764 7254 12776
rect 7285 12767 7343 12773
rect 7285 12764 7297 12767
rect 7248 12736 7297 12764
rect 7248 12724 7254 12736
rect 7285 12733 7297 12736
rect 7331 12733 7343 12767
rect 8018 12764 8024 12776
rect 7979 12736 8024 12764
rect 7285 12727 7343 12733
rect 8018 12724 8024 12736
rect 8076 12724 8082 12776
rect 9030 12764 9036 12776
rect 8128 12736 9036 12764
rect 2547 12668 5672 12696
rect 5721 12699 5779 12705
rect 2547 12665 2559 12668
rect 2501 12659 2559 12665
rect 5721 12665 5733 12699
rect 5767 12696 5779 12699
rect 6840 12696 6868 12724
rect 8128 12696 8156 12736
rect 9030 12724 9036 12736
rect 9088 12724 9094 12776
rect 8294 12705 8300 12708
rect 5767 12668 8156 12696
rect 5767 12665 5779 12668
rect 5721 12659 5779 12665
rect 8288 12659 8300 12705
rect 8352 12696 8358 12708
rect 8352 12668 8388 12696
rect 8294 12656 8300 12659
rect 8352 12656 8358 12668
rect 4246 12588 4252 12640
rect 4304 12628 4310 12640
rect 6365 12631 6423 12637
rect 6365 12628 6377 12631
rect 4304 12600 6377 12628
rect 4304 12588 4310 12600
rect 6365 12597 6377 12600
rect 6411 12628 6423 12631
rect 6546 12628 6552 12640
rect 6411 12600 6552 12628
rect 6411 12597 6423 12600
rect 6365 12591 6423 12597
rect 6546 12588 6552 12600
rect 6604 12588 6610 12640
rect 6822 12628 6828 12640
rect 6783 12600 6828 12628
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 7193 12631 7251 12637
rect 7193 12597 7205 12631
rect 7239 12628 7251 12631
rect 7834 12628 7840 12640
rect 7239 12600 7840 12628
rect 7239 12597 7251 12600
rect 7193 12591 7251 12597
rect 7834 12588 7840 12600
rect 7892 12628 7898 12640
rect 9140 12628 9168 12872
rect 10410 12832 10416 12844
rect 10371 12804 10416 12832
rect 10410 12792 10416 12804
rect 10468 12832 10474 12844
rect 10870 12832 10876 12844
rect 10468 12804 10876 12832
rect 10468 12792 10474 12804
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 9490 12724 9496 12776
rect 9548 12764 9554 12776
rect 10229 12767 10287 12773
rect 10229 12764 10241 12767
rect 9548 12736 10241 12764
rect 9548 12724 9554 12736
rect 10229 12733 10241 12736
rect 10275 12733 10287 12767
rect 10229 12727 10287 12733
rect 10318 12724 10324 12776
rect 10376 12764 10382 12776
rect 10376 12736 10421 12764
rect 10376 12724 10382 12736
rect 11241 12699 11299 12705
rect 11241 12696 11253 12699
rect 9876 12668 11253 12696
rect 7892 12600 9168 12628
rect 9401 12631 9459 12637
rect 7892 12588 7898 12600
rect 9401 12597 9413 12631
rect 9447 12628 9459 12631
rect 9766 12628 9772 12640
rect 9447 12600 9772 12628
rect 9447 12597 9459 12600
rect 9401 12591 9459 12597
rect 9766 12588 9772 12600
rect 9824 12588 9830 12640
rect 9876 12637 9904 12668
rect 11241 12665 11253 12668
rect 11287 12665 11299 12699
rect 11348 12696 11376 12872
rect 12802 12860 12808 12912
rect 12860 12900 12866 12912
rect 12860 12872 13308 12900
rect 12860 12860 12866 12872
rect 13280 12844 13308 12872
rect 11517 12835 11575 12841
rect 11517 12801 11529 12835
rect 11563 12832 11575 12835
rect 11606 12832 11612 12844
rect 11563 12804 11612 12832
rect 11563 12801 11575 12804
rect 11517 12795 11575 12801
rect 11606 12792 11612 12804
rect 11664 12792 11670 12844
rect 12250 12792 12256 12844
rect 12308 12832 12314 12844
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 12308 12804 13001 12832
rect 12308 12792 12314 12804
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 13262 12792 13268 12844
rect 13320 12832 13326 12844
rect 14369 12835 14427 12841
rect 14369 12832 14381 12835
rect 13320 12804 14381 12832
rect 13320 12792 13326 12804
rect 14369 12801 14381 12804
rect 14415 12801 14427 12835
rect 14550 12832 14556 12844
rect 14511 12804 14556 12832
rect 14369 12795 14427 12801
rect 14550 12792 14556 12804
rect 14608 12792 14614 12844
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 12897 12767 12955 12773
rect 12897 12764 12909 12767
rect 12492 12736 12909 12764
rect 12492 12724 12498 12736
rect 12897 12733 12909 12736
rect 12943 12764 12955 12767
rect 13814 12764 13820 12776
rect 12943 12736 13820 12764
rect 12943 12733 12955 12736
rect 12897 12727 12955 12733
rect 13814 12724 13820 12736
rect 13872 12724 13878 12776
rect 14277 12699 14335 12705
rect 14277 12696 14289 12699
rect 11348 12668 14289 12696
rect 11241 12659 11299 12665
rect 14277 12665 14289 12668
rect 14323 12696 14335 12699
rect 14550 12696 14556 12708
rect 14323 12668 14556 12696
rect 14323 12665 14335 12668
rect 14277 12659 14335 12665
rect 14550 12656 14556 12668
rect 14608 12656 14614 12708
rect 9861 12631 9919 12637
rect 9861 12597 9873 12631
rect 9907 12597 9919 12631
rect 11330 12628 11336 12640
rect 11291 12600 11336 12628
rect 9861 12591 9919 12597
rect 11330 12588 11336 12600
rect 11388 12588 11394 12640
rect 11790 12588 11796 12640
rect 11848 12628 11854 12640
rect 12250 12628 12256 12640
rect 11848 12600 12256 12628
rect 11848 12588 11854 12600
rect 12250 12588 12256 12600
rect 12308 12628 12314 12640
rect 12805 12631 12863 12637
rect 12805 12628 12817 12631
rect 12308 12600 12817 12628
rect 12308 12588 12314 12600
rect 12805 12597 12817 12600
rect 12851 12597 12863 12631
rect 13906 12628 13912 12640
rect 13867 12600 13912 12628
rect 12805 12591 12863 12597
rect 13906 12588 13912 12600
rect 13964 12588 13970 12640
rect 1104 12538 15824 12560
rect 1104 12486 5912 12538
rect 5964 12486 5976 12538
rect 6028 12486 6040 12538
rect 6092 12486 6104 12538
rect 6156 12486 10843 12538
rect 10895 12486 10907 12538
rect 10959 12486 10971 12538
rect 11023 12486 11035 12538
rect 11087 12486 15824 12538
rect 1104 12464 15824 12486
rect 3234 12384 3240 12436
rect 3292 12424 3298 12436
rect 3329 12427 3387 12433
rect 3329 12424 3341 12427
rect 3292 12396 3341 12424
rect 3292 12384 3298 12396
rect 3329 12393 3341 12396
rect 3375 12393 3387 12427
rect 3329 12387 3387 12393
rect 4525 12427 4583 12433
rect 4525 12393 4537 12427
rect 4571 12424 4583 12427
rect 4614 12424 4620 12436
rect 4571 12396 4620 12424
rect 4571 12393 4583 12396
rect 4525 12387 4583 12393
rect 4614 12384 4620 12396
rect 4672 12384 4678 12436
rect 4985 12427 5043 12433
rect 4985 12393 4997 12427
rect 5031 12424 5043 12427
rect 5031 12396 5672 12424
rect 5031 12393 5043 12396
rect 4985 12387 5043 12393
rect 5644 12356 5672 12396
rect 5718 12384 5724 12436
rect 5776 12424 5782 12436
rect 6270 12424 6276 12436
rect 5776 12396 6276 12424
rect 5776 12384 5782 12396
rect 6270 12384 6276 12396
rect 6328 12424 6334 12436
rect 6457 12427 6515 12433
rect 6457 12424 6469 12427
rect 6328 12396 6469 12424
rect 6328 12384 6334 12396
rect 6457 12393 6469 12396
rect 6503 12393 6515 12427
rect 8113 12427 8171 12433
rect 8113 12424 8125 12427
rect 6457 12387 6515 12393
rect 7116 12396 8125 12424
rect 6472 12356 6500 12387
rect 6978 12359 7036 12365
rect 6978 12356 6990 12359
rect 5644 12328 6408 12356
rect 6472 12328 6990 12356
rect 2222 12297 2228 12300
rect 2216 12288 2228 12297
rect 2183 12260 2228 12288
rect 2216 12251 2228 12260
rect 2222 12248 2228 12251
rect 2280 12248 2286 12300
rect 3881 12291 3939 12297
rect 3881 12257 3893 12291
rect 3927 12288 3939 12291
rect 4246 12288 4252 12300
rect 3927 12260 4252 12288
rect 3927 12257 3939 12260
rect 3881 12251 3939 12257
rect 4246 12248 4252 12260
rect 4304 12248 4310 12300
rect 4430 12288 4436 12300
rect 4391 12260 4436 12288
rect 4430 12248 4436 12260
rect 4488 12248 4494 12300
rect 5074 12288 5080 12300
rect 5035 12260 5080 12288
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 5344 12291 5402 12297
rect 5344 12257 5356 12291
rect 5390 12288 5402 12291
rect 5810 12288 5816 12300
rect 5390 12260 5816 12288
rect 5390 12257 5402 12260
rect 5344 12251 5402 12257
rect 5810 12248 5816 12260
rect 5868 12248 5874 12300
rect 6380 12288 6408 12328
rect 6978 12325 6990 12328
rect 7024 12325 7036 12359
rect 6978 12319 7036 12325
rect 7116 12288 7144 12396
rect 8113 12393 8125 12396
rect 8159 12424 8171 12427
rect 8294 12424 8300 12436
rect 8159 12396 8300 12424
rect 8159 12393 8171 12396
rect 8113 12387 8171 12393
rect 8294 12384 8300 12396
rect 8352 12384 8358 12436
rect 9677 12427 9735 12433
rect 9677 12393 9689 12427
rect 9723 12393 9735 12427
rect 11330 12424 11336 12436
rect 9677 12387 9735 12393
rect 10152 12396 11336 12424
rect 7190 12316 7196 12368
rect 7248 12356 7254 12368
rect 7558 12356 7564 12368
rect 7248 12328 7564 12356
rect 7248 12316 7254 12328
rect 7558 12316 7564 12328
rect 7616 12316 7622 12368
rect 9692 12356 9720 12387
rect 10152 12356 10180 12396
rect 11330 12384 11336 12396
rect 11388 12384 11394 12436
rect 12526 12424 12532 12436
rect 12487 12396 12532 12424
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 13170 12424 13176 12436
rect 13131 12396 13176 12424
rect 13170 12384 13176 12396
rect 13228 12384 13234 12436
rect 13541 12427 13599 12433
rect 13541 12393 13553 12427
rect 13587 12424 13599 12427
rect 14185 12427 14243 12433
rect 14185 12424 14197 12427
rect 13587 12396 14197 12424
rect 13587 12393 13599 12396
rect 13541 12387 13599 12393
rect 14185 12393 14197 12396
rect 14231 12393 14243 12427
rect 14185 12387 14243 12393
rect 14553 12427 14611 12433
rect 14553 12393 14565 12427
rect 14599 12424 14611 12427
rect 14918 12424 14924 12436
rect 14599 12396 14924 12424
rect 14599 12393 14611 12396
rect 14553 12387 14611 12393
rect 14918 12384 14924 12396
rect 14976 12384 14982 12436
rect 9692 12328 10180 12356
rect 10962 12316 10968 12368
rect 11020 12356 11026 12368
rect 11118 12359 11176 12365
rect 11118 12356 11130 12359
rect 11020 12328 11130 12356
rect 11020 12316 11026 12328
rect 11118 12325 11130 12328
rect 11164 12325 11176 12359
rect 11118 12319 11176 12325
rect 13633 12359 13691 12365
rect 13633 12325 13645 12359
rect 13679 12356 13691 12359
rect 13906 12356 13912 12368
rect 13679 12328 13912 12356
rect 13679 12325 13691 12328
rect 13633 12319 13691 12325
rect 13906 12316 13912 12328
rect 13964 12316 13970 12368
rect 14645 12359 14703 12365
rect 14645 12325 14657 12359
rect 14691 12356 14703 12359
rect 14734 12356 14740 12368
rect 14691 12328 14740 12356
rect 14691 12325 14703 12328
rect 14645 12319 14703 12325
rect 14734 12316 14740 12328
rect 14792 12356 14798 12368
rect 14792 12328 14964 12356
rect 14792 12316 14798 12328
rect 14936 12300 14964 12328
rect 6380 12260 7144 12288
rect 8662 12248 8668 12300
rect 8720 12288 8726 12300
rect 8849 12291 8907 12297
rect 8849 12288 8861 12291
rect 8720 12260 8861 12288
rect 8720 12248 8726 12260
rect 8849 12257 8861 12260
rect 8895 12257 8907 12291
rect 8849 12251 8907 12257
rect 10045 12291 10103 12297
rect 10045 12257 10057 12291
rect 10091 12288 10103 12291
rect 10686 12288 10692 12300
rect 10091 12260 10692 12288
rect 10091 12257 10103 12260
rect 10045 12251 10103 12257
rect 10686 12248 10692 12260
rect 10744 12248 10750 12300
rect 12342 12288 12348 12300
rect 10796 12260 12348 12288
rect 1949 12223 2007 12229
rect 1949 12189 1961 12223
rect 1995 12189 2007 12223
rect 1949 12183 2007 12189
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12220 4767 12223
rect 4985 12223 5043 12229
rect 4985 12220 4997 12223
rect 4755 12192 4997 12220
rect 4755 12189 4767 12192
rect 4709 12183 4767 12189
rect 4985 12189 4997 12192
rect 5031 12189 5043 12223
rect 6730 12220 6736 12232
rect 6691 12192 6736 12220
rect 4985 12183 5043 12189
rect 1394 12044 1400 12096
rect 1452 12084 1458 12096
rect 1964 12084 1992 12183
rect 6730 12180 6736 12192
rect 6788 12180 6794 12232
rect 8202 12220 8208 12232
rect 8163 12192 8208 12220
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 8938 12220 8944 12232
rect 8899 12192 8944 12220
rect 8938 12180 8944 12192
rect 8996 12180 9002 12232
rect 9033 12223 9091 12229
rect 9033 12189 9045 12223
rect 9079 12189 9091 12223
rect 9033 12183 9091 12189
rect 3697 12155 3755 12161
rect 3697 12121 3709 12155
rect 3743 12152 3755 12155
rect 4246 12152 4252 12164
rect 3743 12124 4252 12152
rect 3743 12121 3755 12124
rect 3697 12115 3755 12121
rect 2866 12084 2872 12096
rect 1452 12056 2872 12084
rect 1452 12044 1458 12056
rect 2866 12044 2872 12056
rect 2924 12084 2930 12096
rect 3712 12084 3740 12115
rect 4246 12112 4252 12124
rect 4304 12112 4310 12164
rect 8481 12155 8539 12161
rect 8481 12152 8493 12155
rect 7668 12124 8493 12152
rect 2924 12056 3740 12084
rect 2924 12044 2930 12056
rect 3786 12044 3792 12096
rect 3844 12084 3850 12096
rect 4065 12087 4123 12093
rect 4065 12084 4077 12087
rect 3844 12056 4077 12084
rect 3844 12044 3850 12056
rect 4065 12053 4077 12056
rect 4111 12053 4123 12087
rect 4065 12047 4123 12053
rect 5258 12044 5264 12096
rect 5316 12084 5322 12096
rect 7668 12084 7696 12124
rect 8481 12121 8493 12124
rect 8527 12121 8539 12155
rect 8481 12115 8539 12121
rect 8846 12112 8852 12164
rect 8904 12152 8910 12164
rect 9048 12152 9076 12183
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 9732 12192 10149 12220
rect 9732 12180 9738 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12220 10379 12223
rect 10410 12220 10416 12232
rect 10367 12192 10416 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 10796 12152 10824 12260
rect 12342 12248 12348 12260
rect 12400 12248 12406 12300
rect 13078 12248 13084 12300
rect 13136 12248 13142 12300
rect 14458 12248 14464 12300
rect 14516 12288 14522 12300
rect 14516 12260 14780 12288
rect 14516 12248 14522 12260
rect 10870 12180 10876 12232
rect 10928 12220 10934 12232
rect 13096 12220 13124 12248
rect 14752 12229 14780 12260
rect 14918 12248 14924 12300
rect 14976 12248 14982 12300
rect 13725 12223 13783 12229
rect 13725 12220 13737 12223
rect 10928 12192 10973 12220
rect 13096 12192 13737 12220
rect 10928 12180 10934 12192
rect 13725 12189 13737 12192
rect 13771 12189 13783 12223
rect 13725 12183 13783 12189
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12189 14795 12223
rect 14737 12183 14795 12189
rect 8904 12124 9076 12152
rect 9140 12124 10824 12152
rect 8904 12112 8910 12124
rect 5316 12056 7696 12084
rect 5316 12044 5322 12056
rect 7926 12044 7932 12096
rect 7984 12084 7990 12096
rect 9140 12084 9168 12124
rect 7984 12056 9168 12084
rect 7984 12044 7990 12056
rect 10410 12044 10416 12096
rect 10468 12084 10474 12096
rect 12253 12087 12311 12093
rect 12253 12084 12265 12087
rect 10468 12056 12265 12084
rect 10468 12044 10474 12056
rect 12253 12053 12265 12056
rect 12299 12053 12311 12087
rect 12253 12047 12311 12053
rect 1104 11994 15824 12016
rect 1104 11942 3447 11994
rect 3499 11942 3511 11994
rect 3563 11942 3575 11994
rect 3627 11942 3639 11994
rect 3691 11942 8378 11994
rect 8430 11942 8442 11994
rect 8494 11942 8506 11994
rect 8558 11942 8570 11994
rect 8622 11942 13308 11994
rect 13360 11942 13372 11994
rect 13424 11942 13436 11994
rect 13488 11942 13500 11994
rect 13552 11942 15824 11994
rect 1104 11920 15824 11942
rect 1857 11883 1915 11889
rect 1857 11849 1869 11883
rect 1903 11880 1915 11883
rect 2130 11880 2136 11892
rect 1903 11852 2136 11880
rect 1903 11849 1915 11852
rect 1857 11843 1915 11849
rect 2130 11840 2136 11852
rect 2188 11840 2194 11892
rect 4249 11883 4307 11889
rect 4249 11880 4261 11883
rect 2700 11852 4261 11880
rect 2498 11744 2504 11756
rect 2411 11716 2504 11744
rect 2498 11704 2504 11716
rect 2556 11744 2562 11756
rect 2700 11744 2728 11852
rect 4249 11849 4261 11852
rect 4295 11849 4307 11883
rect 4249 11843 4307 11849
rect 4430 11840 4436 11892
rect 4488 11880 4494 11892
rect 5721 11883 5779 11889
rect 5721 11880 5733 11883
rect 4488 11852 5733 11880
rect 4488 11840 4494 11852
rect 5721 11849 5733 11852
rect 5767 11849 5779 11883
rect 5721 11843 5779 11849
rect 6362 11840 6368 11892
rect 6420 11880 6426 11892
rect 7745 11883 7803 11889
rect 7745 11880 7757 11883
rect 6420 11852 7757 11880
rect 6420 11840 6426 11852
rect 7745 11849 7757 11852
rect 7791 11849 7803 11883
rect 8662 11880 8668 11892
rect 8623 11852 8668 11880
rect 7745 11843 7803 11849
rect 8662 11840 8668 11852
rect 8720 11840 8726 11892
rect 9030 11840 9036 11892
rect 9088 11880 9094 11892
rect 9582 11880 9588 11892
rect 9088 11852 9588 11880
rect 9088 11840 9094 11852
rect 9582 11840 9588 11852
rect 9640 11840 9646 11892
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 10686 11880 10692 11892
rect 9732 11852 9777 11880
rect 10647 11852 10692 11880
rect 9732 11840 9738 11852
rect 10686 11840 10692 11852
rect 10744 11840 10750 11892
rect 14918 11812 14924 11824
rect 7300 11784 14924 11812
rect 2866 11744 2872 11756
rect 2556 11716 2728 11744
rect 2827 11716 2872 11744
rect 2556 11704 2562 11716
rect 2866 11704 2872 11716
rect 2924 11704 2930 11756
rect 4890 11704 4896 11756
rect 4948 11744 4954 11756
rect 5166 11744 5172 11756
rect 4948 11716 5172 11744
rect 4948 11704 4954 11716
rect 5166 11704 5172 11716
rect 5224 11704 5230 11756
rect 5261 11747 5319 11753
rect 5261 11713 5273 11747
rect 5307 11744 5319 11747
rect 5442 11744 5448 11756
rect 5307 11716 5448 11744
rect 5307 11713 5319 11716
rect 5261 11707 5319 11713
rect 3142 11685 3148 11688
rect 3136 11676 3148 11685
rect 3055 11648 3148 11676
rect 3136 11639 3148 11648
rect 3200 11676 3206 11688
rect 5276 11676 5304 11707
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 6270 11744 6276 11756
rect 6231 11716 6276 11744
rect 6270 11704 6276 11716
rect 6328 11704 6334 11756
rect 7300 11744 7328 11784
rect 14918 11772 14924 11784
rect 14976 11772 14982 11824
rect 7466 11744 7472 11756
rect 7208 11716 7328 11744
rect 7427 11716 7472 11744
rect 3200 11648 5304 11676
rect 6181 11679 6239 11685
rect 3142 11636 3148 11639
rect 3200 11636 3206 11648
rect 6181 11645 6193 11679
rect 6227 11676 6239 11679
rect 6822 11676 6828 11688
rect 6227 11648 6828 11676
rect 6227 11645 6239 11648
rect 6181 11639 6239 11645
rect 6822 11636 6828 11648
rect 6880 11636 6886 11688
rect 7208 11676 7236 11716
rect 7466 11704 7472 11716
rect 7524 11704 7530 11756
rect 8389 11747 8447 11753
rect 8389 11713 8401 11747
rect 8435 11744 8447 11747
rect 9214 11744 9220 11756
rect 8435 11716 9220 11744
rect 8435 11713 8447 11716
rect 8389 11707 8447 11713
rect 9214 11704 9220 11716
rect 9272 11704 9278 11756
rect 9766 11704 9772 11756
rect 9824 11744 9830 11756
rect 10229 11747 10287 11753
rect 10229 11744 10241 11747
rect 9824 11716 10241 11744
rect 9824 11704 9830 11716
rect 10229 11713 10241 11716
rect 10275 11744 10287 11747
rect 10686 11744 10692 11756
rect 10275 11716 10692 11744
rect 10275 11713 10287 11716
rect 10229 11707 10287 11713
rect 10686 11704 10692 11716
rect 10744 11744 10750 11756
rect 10962 11744 10968 11756
rect 10744 11716 10968 11744
rect 10744 11704 10750 11716
rect 10962 11704 10968 11716
rect 11020 11704 11026 11756
rect 11146 11744 11152 11756
rect 11107 11716 11152 11744
rect 11146 11704 11152 11716
rect 11204 11704 11210 11756
rect 11241 11747 11299 11753
rect 11241 11713 11253 11747
rect 11287 11713 11299 11747
rect 11241 11707 11299 11713
rect 7116 11648 7236 11676
rect 7285 11679 7343 11685
rect 2225 11611 2283 11617
rect 2225 11577 2237 11611
rect 2271 11608 2283 11611
rect 2774 11608 2780 11620
rect 2271 11580 2780 11608
rect 2271 11577 2283 11580
rect 2225 11571 2283 11577
rect 2774 11568 2780 11580
rect 2832 11568 2838 11620
rect 3234 11568 3240 11620
rect 3292 11608 3298 11620
rect 5626 11608 5632 11620
rect 3292 11580 5632 11608
rect 3292 11568 3298 11580
rect 5626 11568 5632 11580
rect 5684 11568 5690 11620
rect 6089 11611 6147 11617
rect 6089 11577 6101 11611
rect 6135 11608 6147 11611
rect 6135 11580 6960 11608
rect 6135 11577 6147 11580
rect 6089 11571 6147 11577
rect 2314 11500 2320 11552
rect 2372 11540 2378 11552
rect 4614 11540 4620 11552
rect 2372 11512 2417 11540
rect 4575 11512 4620 11540
rect 2372 11500 2378 11512
rect 4614 11500 4620 11512
rect 4672 11500 4678 11552
rect 4890 11500 4896 11552
rect 4948 11540 4954 11552
rect 4985 11543 5043 11549
rect 4985 11540 4997 11543
rect 4948 11512 4997 11540
rect 4948 11500 4954 11512
rect 4985 11509 4997 11512
rect 5031 11509 5043 11543
rect 4985 11503 5043 11509
rect 5077 11543 5135 11549
rect 5077 11509 5089 11543
rect 5123 11540 5135 11543
rect 6454 11540 6460 11552
rect 5123 11512 6460 11540
rect 5123 11509 5135 11512
rect 5077 11503 5135 11509
rect 6454 11500 6460 11512
rect 6512 11500 6518 11552
rect 6932 11549 6960 11580
rect 6917 11543 6975 11549
rect 6917 11509 6929 11543
rect 6963 11509 6975 11543
rect 7116 11540 7144 11648
rect 7285 11645 7297 11679
rect 7331 11676 7343 11679
rect 8202 11676 8208 11688
rect 7331 11648 8208 11676
rect 7331 11645 7343 11648
rect 7285 11639 7343 11645
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 9950 11636 9956 11688
rect 10008 11676 10014 11688
rect 10137 11679 10195 11685
rect 10137 11676 10149 11679
rect 10008 11648 10149 11676
rect 10008 11636 10014 11648
rect 10137 11645 10149 11648
rect 10183 11676 10195 11679
rect 10410 11676 10416 11688
rect 10183 11648 10416 11676
rect 10183 11645 10195 11648
rect 10137 11639 10195 11645
rect 10410 11636 10416 11648
rect 10468 11636 10474 11688
rect 10980 11676 11008 11704
rect 11256 11676 11284 11707
rect 11514 11704 11520 11756
rect 11572 11744 11578 11756
rect 13173 11747 13231 11753
rect 13173 11744 13185 11747
rect 11572 11716 13185 11744
rect 11572 11704 11578 11716
rect 13173 11713 13185 11716
rect 13219 11713 13231 11747
rect 15102 11744 15108 11756
rect 15063 11716 15108 11744
rect 13173 11707 13231 11713
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 10980 11648 11284 11676
rect 12989 11679 13047 11685
rect 12989 11645 13001 11679
rect 13035 11676 13047 11679
rect 14642 11676 14648 11688
rect 13035 11648 14648 11676
rect 13035 11645 13047 11648
rect 12989 11639 13047 11645
rect 14642 11636 14648 11648
rect 14700 11676 14706 11688
rect 14829 11679 14887 11685
rect 14829 11676 14841 11679
rect 14700 11648 14841 11676
rect 14700 11636 14706 11648
rect 14829 11645 14841 11648
rect 14875 11645 14887 11679
rect 14829 11639 14887 11645
rect 7190 11568 7196 11620
rect 7248 11608 7254 11620
rect 8113 11611 8171 11617
rect 8113 11608 8125 11611
rect 7248 11580 8125 11608
rect 7248 11568 7254 11580
rect 8113 11577 8125 11580
rect 8159 11577 8171 11611
rect 8113 11571 8171 11577
rect 8294 11568 8300 11620
rect 8352 11608 8358 11620
rect 9125 11611 9183 11617
rect 9125 11608 9137 11611
rect 8352 11580 9137 11608
rect 8352 11568 8358 11580
rect 9125 11577 9137 11580
rect 9171 11577 9183 11611
rect 9125 11571 9183 11577
rect 9858 11568 9864 11620
rect 9916 11608 9922 11620
rect 10045 11611 10103 11617
rect 10045 11608 10057 11611
rect 9916 11580 10057 11608
rect 9916 11568 9922 11580
rect 10045 11577 10057 11580
rect 10091 11577 10103 11611
rect 10045 11571 10103 11577
rect 11054 11568 11060 11620
rect 11112 11608 11118 11620
rect 11112 11580 11157 11608
rect 11112 11568 11118 11580
rect 13078 11568 13084 11620
rect 13136 11608 13142 11620
rect 13998 11608 14004 11620
rect 13136 11580 14004 11608
rect 13136 11568 13142 11580
rect 13998 11568 14004 11580
rect 14056 11568 14062 11620
rect 7377 11543 7435 11549
rect 7377 11540 7389 11543
rect 7116 11512 7389 11540
rect 6917 11503 6975 11509
rect 7377 11509 7389 11512
rect 7423 11509 7435 11543
rect 7377 11503 7435 11509
rect 8205 11543 8263 11549
rect 8205 11509 8217 11543
rect 8251 11540 8263 11543
rect 8662 11540 8668 11552
rect 8251 11512 8668 11540
rect 8251 11509 8263 11512
rect 8205 11503 8263 11509
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 9033 11543 9091 11549
rect 9033 11509 9045 11543
rect 9079 11540 9091 11543
rect 9490 11540 9496 11552
rect 9079 11512 9496 11540
rect 9079 11509 9091 11512
rect 9033 11503 9091 11509
rect 9490 11500 9496 11512
rect 9548 11540 9554 11552
rect 13906 11540 13912 11552
rect 9548 11512 13912 11540
rect 9548 11500 9554 11512
rect 13906 11500 13912 11512
rect 13964 11500 13970 11552
rect 1104 11450 15824 11472
rect 1104 11398 5912 11450
rect 5964 11398 5976 11450
rect 6028 11398 6040 11450
rect 6092 11398 6104 11450
rect 6156 11398 10843 11450
rect 10895 11398 10907 11450
rect 10959 11398 10971 11450
rect 11023 11398 11035 11450
rect 11087 11398 15824 11450
rect 1104 11376 15824 11398
rect 2222 11296 2228 11348
rect 2280 11336 2286 11348
rect 2777 11339 2835 11345
rect 2777 11336 2789 11339
rect 2280 11308 2789 11336
rect 2280 11296 2286 11308
rect 2777 11305 2789 11308
rect 2823 11305 2835 11339
rect 2777 11299 2835 11305
rect 4617 11339 4675 11345
rect 4617 11305 4629 11339
rect 4663 11336 4675 11339
rect 4801 11339 4859 11345
rect 4801 11336 4813 11339
rect 4663 11308 4813 11336
rect 4663 11305 4675 11308
rect 4617 11299 4675 11305
rect 4801 11305 4813 11308
rect 4847 11305 4859 11339
rect 4801 11299 4859 11305
rect 5169 11339 5227 11345
rect 5169 11305 5181 11339
rect 5215 11336 5227 11339
rect 5718 11336 5724 11348
rect 5215 11308 5724 11336
rect 5215 11305 5227 11308
rect 5169 11299 5227 11305
rect 5718 11296 5724 11308
rect 5776 11296 5782 11348
rect 6270 11336 6276 11348
rect 5828 11308 6276 11336
rect 1664 11271 1722 11277
rect 1664 11237 1676 11271
rect 1710 11268 1722 11271
rect 2498 11268 2504 11280
rect 1710 11240 2504 11268
rect 1710 11237 1722 11240
rect 1664 11231 1722 11237
rect 2498 11228 2504 11240
rect 2556 11228 2562 11280
rect 5258 11268 5264 11280
rect 3068 11240 4752 11268
rect 5219 11240 5264 11268
rect 1394 11200 1400 11212
rect 1355 11172 1400 11200
rect 1394 11160 1400 11172
rect 1452 11160 1458 11212
rect 3068 11209 3096 11240
rect 3053 11203 3111 11209
rect 3053 11169 3065 11203
rect 3099 11169 3111 11203
rect 3053 11163 3111 11169
rect 4065 11203 4123 11209
rect 4065 11169 4077 11203
rect 4111 11200 4123 11203
rect 4617 11203 4675 11209
rect 4617 11200 4629 11203
rect 4111 11172 4629 11200
rect 4111 11169 4123 11172
rect 4065 11163 4123 11169
rect 4617 11169 4629 11172
rect 4663 11169 4675 11203
rect 4617 11163 4675 11169
rect 2866 11092 2872 11144
rect 2924 11132 2930 11144
rect 3237 11135 3295 11141
rect 3237 11132 3249 11135
rect 2924 11104 3249 11132
rect 2924 11092 2930 11104
rect 3237 11101 3249 11104
rect 3283 11101 3295 11135
rect 3237 11095 3295 11101
rect 4249 11135 4307 11141
rect 4249 11101 4261 11135
rect 4295 11101 4307 11135
rect 4249 11095 4307 11101
rect 3234 10956 3240 11008
rect 3292 10996 3298 11008
rect 4264 10996 4292 11095
rect 4724 11064 4752 11240
rect 5258 11228 5264 11240
rect 5316 11228 5322 11280
rect 5828 11209 5856 11308
rect 6270 11296 6276 11308
rect 6328 11336 6334 11348
rect 6730 11336 6736 11348
rect 6328 11308 6736 11336
rect 6328 11296 6334 11308
rect 6730 11296 6736 11308
rect 6788 11296 6794 11348
rect 7193 11339 7251 11345
rect 7193 11305 7205 11339
rect 7239 11305 7251 11339
rect 7193 11299 7251 11305
rect 7561 11339 7619 11345
rect 7561 11305 7573 11339
rect 7607 11336 7619 11339
rect 8294 11336 8300 11348
rect 7607 11308 8300 11336
rect 7607 11305 7619 11308
rect 7561 11299 7619 11305
rect 6178 11268 6184 11280
rect 6012 11240 6184 11268
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11169 5871 11203
rect 6012 11200 6040 11240
rect 6178 11228 6184 11240
rect 6236 11268 6242 11280
rect 7208 11268 7236 11299
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 8573 11339 8631 11345
rect 8573 11305 8585 11339
rect 8619 11336 8631 11339
rect 8938 11336 8944 11348
rect 8619 11308 8944 11336
rect 8619 11305 8631 11308
rect 8573 11299 8631 11305
rect 8938 11296 8944 11308
rect 8996 11296 9002 11348
rect 9030 11296 9036 11348
rect 9088 11336 9094 11348
rect 9306 11336 9312 11348
rect 9088 11308 9312 11336
rect 9088 11296 9094 11308
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 10318 11296 10324 11348
rect 10376 11336 10382 11348
rect 10413 11339 10471 11345
rect 10413 11336 10425 11339
rect 10376 11308 10425 11336
rect 10376 11296 10382 11308
rect 10413 11305 10425 11308
rect 10459 11305 10471 11339
rect 10413 11299 10471 11305
rect 11238 11296 11244 11348
rect 11296 11336 11302 11348
rect 13081 11339 13139 11345
rect 13081 11336 13093 11339
rect 11296 11308 13093 11336
rect 11296 11296 11302 11308
rect 13081 11305 13093 11308
rect 13127 11305 13139 11339
rect 13081 11299 13139 11305
rect 8846 11268 8852 11280
rect 6236 11240 7236 11268
rect 7852 11240 8852 11268
rect 6236 11228 6242 11240
rect 5813 11163 5871 11169
rect 5920 11172 6040 11200
rect 6080 11203 6138 11209
rect 5445 11135 5503 11141
rect 5445 11101 5457 11135
rect 5491 11132 5503 11135
rect 5920 11132 5948 11172
rect 6080 11169 6092 11203
rect 6126 11200 6138 11203
rect 6454 11200 6460 11212
rect 6126 11172 6460 11200
rect 6126 11169 6138 11172
rect 6080 11163 6138 11169
rect 6454 11160 6460 11172
rect 6512 11200 6518 11212
rect 7852 11200 7880 11240
rect 8846 11228 8852 11240
rect 8904 11228 8910 11280
rect 10134 11228 10140 11280
rect 10192 11268 10198 11280
rect 10781 11271 10839 11277
rect 10781 11268 10793 11271
rect 10192 11240 10793 11268
rect 10192 11228 10198 11240
rect 10781 11237 10793 11240
rect 10827 11237 10839 11271
rect 10781 11231 10839 11237
rect 6512 11172 7880 11200
rect 6512 11160 6518 11172
rect 7926 11160 7932 11212
rect 7984 11200 7990 11212
rect 8938 11200 8944 11212
rect 7984 11172 8029 11200
rect 8899 11172 8944 11200
rect 7984 11160 7990 11172
rect 8938 11160 8944 11172
rect 8996 11160 9002 11212
rect 9033 11203 9091 11209
rect 9033 11169 9045 11203
rect 9079 11200 9091 11203
rect 9079 11172 10088 11200
rect 9079 11169 9091 11172
rect 9033 11163 9091 11169
rect 5491 11104 5948 11132
rect 5491 11101 5503 11104
rect 5445 11095 5503 11101
rect 6914 11092 6920 11144
rect 6972 11132 6978 11144
rect 7944 11132 7972 11160
rect 6972 11104 7972 11132
rect 6972 11092 6978 11104
rect 8018 11092 8024 11144
rect 8076 11132 8082 11144
rect 8205 11135 8263 11141
rect 8076 11104 8121 11132
rect 8076 11092 8082 11104
rect 8205 11101 8217 11135
rect 8251 11101 8263 11135
rect 9214 11132 9220 11144
rect 9175 11104 9220 11132
rect 8205 11095 8263 11101
rect 8220 11064 8248 11095
rect 9214 11092 9220 11104
rect 9272 11092 9278 11144
rect 10060 11132 10088 11172
rect 10226 11160 10232 11212
rect 10284 11200 10290 11212
rect 10321 11203 10379 11209
rect 10321 11200 10333 11203
rect 10284 11172 10333 11200
rect 10284 11160 10290 11172
rect 10321 11169 10333 11172
rect 10367 11169 10379 11203
rect 10321 11163 10379 11169
rect 10686 11160 10692 11212
rect 10744 11200 10750 11212
rect 11698 11200 11704 11212
rect 10744 11172 11008 11200
rect 10744 11160 10750 11172
rect 10134 11132 10140 11144
rect 10060 11104 10140 11132
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 10870 11132 10876 11144
rect 10831 11104 10876 11132
rect 10870 11092 10876 11104
rect 10928 11092 10934 11144
rect 10980 11141 11008 11172
rect 11072 11172 11704 11200
rect 10965 11135 11023 11141
rect 10965 11101 10977 11135
rect 11011 11101 11023 11135
rect 10965 11095 11023 11101
rect 9306 11064 9312 11076
rect 4724 11036 5856 11064
rect 3292 10968 4292 10996
rect 3292 10956 3298 10968
rect 4798 10956 4804 11008
rect 4856 10996 4862 11008
rect 5074 10996 5080 11008
rect 4856 10968 5080 10996
rect 4856 10956 4862 10968
rect 5074 10956 5080 10968
rect 5132 10956 5138 11008
rect 5828 10996 5856 11036
rect 6748 11036 8156 11064
rect 8220 11036 9312 11064
rect 6748 10996 6776 11036
rect 5828 10968 6776 10996
rect 7006 10956 7012 11008
rect 7064 10996 7070 11008
rect 7558 10996 7564 11008
rect 7064 10968 7564 10996
rect 7064 10956 7070 10968
rect 7558 10956 7564 10968
rect 7616 10956 7622 11008
rect 8128 10996 8156 11036
rect 9306 11024 9312 11036
rect 9364 11024 9370 11076
rect 11072 11064 11100 11172
rect 11698 11160 11704 11172
rect 11756 11160 11762 11212
rect 11968 11203 12026 11209
rect 11968 11169 11980 11203
rect 12014 11200 12026 11203
rect 12526 11200 12532 11212
rect 12014 11172 12532 11200
rect 12014 11169 12026 11172
rect 11968 11163 12026 11169
rect 12526 11160 12532 11172
rect 12584 11160 12590 11212
rect 10520 11036 11100 11064
rect 10520 11008 10548 11036
rect 9582 10996 9588 11008
rect 8128 10968 9588 10996
rect 9582 10956 9588 10968
rect 9640 10956 9646 11008
rect 10137 10999 10195 11005
rect 10137 10965 10149 10999
rect 10183 10996 10195 10999
rect 10502 10996 10508 11008
rect 10183 10968 10508 10996
rect 10183 10965 10195 10968
rect 10137 10959 10195 10965
rect 10502 10956 10508 10968
rect 10560 10956 10566 11008
rect 1104 10906 15824 10928
rect 1104 10854 3447 10906
rect 3499 10854 3511 10906
rect 3563 10854 3575 10906
rect 3627 10854 3639 10906
rect 3691 10854 8378 10906
rect 8430 10854 8442 10906
rect 8494 10854 8506 10906
rect 8558 10854 8570 10906
rect 8622 10854 13308 10906
rect 13360 10854 13372 10906
rect 13424 10854 13436 10906
rect 13488 10854 13500 10906
rect 13552 10854 15824 10906
rect 1104 10832 15824 10854
rect 2225 10795 2283 10801
rect 2225 10761 2237 10795
rect 2271 10792 2283 10795
rect 2314 10792 2320 10804
rect 2271 10764 2320 10792
rect 2271 10761 2283 10764
rect 2225 10755 2283 10761
rect 2314 10752 2320 10764
rect 2372 10752 2378 10804
rect 3804 10764 5212 10792
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10656 2927 10659
rect 3142 10656 3148 10668
rect 2915 10628 3148 10656
rect 2915 10625 2927 10628
rect 2869 10619 2927 10625
rect 3142 10616 3148 10628
rect 3200 10656 3206 10668
rect 3418 10656 3424 10668
rect 3200 10628 3424 10656
rect 3200 10616 3206 10628
rect 3418 10616 3424 10628
rect 3476 10616 3482 10668
rect 1489 10591 1547 10597
rect 1489 10557 1501 10591
rect 1535 10557 1547 10591
rect 1489 10551 1547 10557
rect 1765 10591 1823 10597
rect 1765 10557 1777 10591
rect 1811 10588 1823 10591
rect 2958 10588 2964 10600
rect 1811 10560 2964 10588
rect 1811 10557 1823 10560
rect 1765 10551 1823 10557
rect 1504 10520 1532 10551
rect 2958 10548 2964 10560
rect 3016 10548 3022 10600
rect 3605 10591 3663 10597
rect 3605 10557 3617 10591
rect 3651 10588 3663 10591
rect 3804 10588 3832 10764
rect 5184 10724 5212 10764
rect 5442 10752 5448 10804
rect 5500 10792 5506 10804
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 5500 10764 5641 10792
rect 5500 10752 5506 10764
rect 5629 10761 5641 10764
rect 5675 10761 5687 10795
rect 5629 10755 5687 10761
rect 6730 10752 6736 10804
rect 6788 10792 6794 10804
rect 8018 10792 8024 10804
rect 6788 10764 8024 10792
rect 6788 10752 6794 10764
rect 8018 10752 8024 10764
rect 8076 10752 8082 10804
rect 8846 10752 8852 10804
rect 8904 10792 8910 10804
rect 9033 10795 9091 10801
rect 9033 10792 9045 10795
rect 8904 10764 9045 10792
rect 8904 10752 8910 10764
rect 9033 10761 9045 10764
rect 9079 10761 9091 10795
rect 9033 10755 9091 10761
rect 10686 10752 10692 10804
rect 10744 10792 10750 10804
rect 12069 10795 12127 10801
rect 12069 10792 12081 10795
rect 10744 10764 12081 10792
rect 10744 10752 10750 10764
rect 12069 10761 12081 10764
rect 12115 10761 12127 10795
rect 12069 10755 12127 10761
rect 7282 10724 7288 10736
rect 5184 10696 7288 10724
rect 7282 10684 7288 10696
rect 7340 10724 7346 10736
rect 7558 10724 7564 10736
rect 7340 10696 7564 10724
rect 7340 10684 7346 10696
rect 7558 10684 7564 10696
rect 7616 10684 7622 10736
rect 9582 10684 9588 10736
rect 9640 10724 9646 10736
rect 9677 10727 9735 10733
rect 9677 10724 9689 10727
rect 9640 10696 9689 10724
rect 9640 10684 9646 10696
rect 9677 10693 9689 10696
rect 9723 10693 9735 10727
rect 9677 10687 9735 10693
rect 3881 10659 3939 10665
rect 3881 10625 3893 10659
rect 3927 10625 3939 10659
rect 3881 10619 3939 10625
rect 3651 10560 3832 10588
rect 3651 10557 3663 10560
rect 3605 10551 3663 10557
rect 3786 10520 3792 10532
rect 1504 10492 3792 10520
rect 3786 10480 3792 10492
rect 3844 10480 3850 10532
rect 3896 10520 3924 10619
rect 5626 10616 5632 10668
rect 5684 10656 5690 10668
rect 6089 10659 6147 10665
rect 6089 10656 6101 10659
rect 5684 10628 6101 10656
rect 5684 10616 5690 10628
rect 6089 10625 6101 10628
rect 6135 10625 6147 10659
rect 7190 10656 7196 10668
rect 7151 10628 7196 10656
rect 6089 10619 6147 10625
rect 7190 10616 7196 10628
rect 7248 10616 7254 10668
rect 10042 10616 10048 10668
rect 10100 10656 10106 10668
rect 10226 10656 10232 10668
rect 10100 10628 10232 10656
rect 10100 10616 10106 10628
rect 10226 10616 10232 10628
rect 10284 10616 10290 10668
rect 10321 10659 10379 10665
rect 10321 10625 10333 10659
rect 10367 10656 10379 10659
rect 10367 10628 10824 10656
rect 10367 10625 10379 10628
rect 10321 10619 10379 10625
rect 4246 10588 4252 10600
rect 4159 10560 4252 10588
rect 4246 10548 4252 10560
rect 4304 10588 4310 10600
rect 5442 10588 5448 10600
rect 4304 10560 5448 10588
rect 4304 10548 4310 10560
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 5534 10548 5540 10600
rect 5592 10588 5598 10600
rect 5905 10591 5963 10597
rect 5905 10588 5917 10591
rect 5592 10560 5917 10588
rect 5592 10548 5598 10560
rect 5905 10557 5917 10560
rect 5951 10557 5963 10591
rect 5905 10551 5963 10557
rect 7653 10591 7711 10597
rect 7653 10557 7665 10591
rect 7699 10557 7711 10591
rect 7653 10551 7711 10557
rect 4522 10529 4528 10532
rect 4516 10520 4528 10529
rect 3896 10492 4528 10520
rect 4516 10483 4528 10492
rect 4522 10480 4528 10483
rect 4580 10480 4586 10532
rect 7190 10520 7196 10532
rect 4632 10492 7196 10520
rect 2590 10452 2596 10464
rect 2551 10424 2596 10452
rect 2590 10412 2596 10424
rect 2648 10412 2654 10464
rect 2685 10455 2743 10461
rect 2685 10421 2697 10455
rect 2731 10452 2743 10455
rect 3237 10455 3295 10461
rect 3237 10452 3249 10455
rect 2731 10424 3249 10452
rect 2731 10421 2743 10424
rect 2685 10415 2743 10421
rect 3237 10421 3249 10424
rect 3283 10421 3295 10455
rect 3237 10415 3295 10421
rect 3697 10455 3755 10461
rect 3697 10421 3709 10455
rect 3743 10452 3755 10455
rect 4338 10452 4344 10464
rect 3743 10424 4344 10452
rect 3743 10421 3755 10424
rect 3697 10415 3755 10421
rect 4338 10412 4344 10424
rect 4396 10452 4402 10464
rect 4632 10452 4660 10492
rect 7190 10480 7196 10492
rect 7248 10480 7254 10532
rect 7668 10520 7696 10551
rect 7742 10548 7748 10600
rect 7800 10588 7806 10600
rect 7920 10591 7978 10597
rect 7920 10588 7932 10591
rect 7800 10560 7932 10588
rect 7800 10548 7806 10560
rect 7920 10557 7932 10560
rect 7966 10588 7978 10591
rect 9214 10588 9220 10600
rect 7966 10560 9220 10588
rect 7966 10557 7978 10560
rect 7920 10551 7978 10557
rect 9214 10548 9220 10560
rect 9272 10548 9278 10600
rect 9766 10588 9772 10600
rect 9315 10560 9772 10588
rect 9315 10520 9343 10560
rect 9766 10548 9772 10560
rect 9824 10588 9830 10600
rect 10502 10588 10508 10600
rect 9824 10560 10508 10588
rect 9824 10548 9830 10560
rect 10502 10548 10508 10560
rect 10560 10588 10566 10600
rect 10689 10591 10747 10597
rect 10689 10588 10701 10591
rect 10560 10560 10701 10588
rect 10560 10548 10566 10560
rect 10689 10557 10701 10560
rect 10735 10557 10747 10591
rect 10796 10588 10824 10628
rect 11698 10616 11704 10668
rect 11756 10656 11762 10668
rect 12621 10659 12679 10665
rect 12621 10656 12633 10659
rect 11756 10628 12633 10656
rect 11756 10616 11762 10628
rect 12621 10625 12633 10628
rect 12667 10625 12679 10659
rect 12621 10619 12679 10625
rect 13998 10616 14004 10668
rect 14056 10656 14062 10668
rect 14829 10659 14887 10665
rect 14829 10656 14841 10659
rect 14056 10628 14841 10656
rect 14056 10616 14062 10628
rect 14829 10625 14841 10628
rect 14875 10625 14887 10659
rect 14829 10619 14887 10625
rect 10956 10591 11014 10597
rect 10956 10588 10968 10591
rect 10796 10560 10968 10588
rect 10689 10551 10747 10557
rect 10956 10557 10968 10560
rect 11002 10588 11014 10591
rect 11238 10588 11244 10600
rect 11002 10560 11244 10588
rect 11002 10557 11014 10560
rect 10956 10551 11014 10557
rect 11238 10548 11244 10560
rect 11296 10548 11302 10600
rect 12888 10591 12946 10597
rect 12888 10557 12900 10591
rect 12934 10588 12946 10591
rect 14016 10588 14044 10616
rect 12934 10560 14044 10588
rect 14737 10591 14795 10597
rect 12934 10557 12946 10560
rect 12888 10551 12946 10557
rect 14737 10557 14749 10591
rect 14783 10588 14795 10591
rect 15102 10588 15108 10600
rect 14783 10560 15108 10588
rect 14783 10557 14795 10560
rect 14737 10551 14795 10557
rect 15102 10548 15108 10560
rect 15160 10548 15166 10600
rect 7668 10492 9343 10520
rect 10045 10523 10103 10529
rect 10045 10489 10057 10523
rect 10091 10520 10103 10523
rect 11882 10520 11888 10532
rect 10091 10492 11888 10520
rect 10091 10489 10103 10492
rect 10045 10483 10103 10489
rect 11882 10480 11888 10492
rect 11940 10480 11946 10532
rect 4396 10424 4660 10452
rect 4396 10412 4402 10424
rect 4706 10412 4712 10464
rect 4764 10452 4770 10464
rect 5166 10452 5172 10464
rect 4764 10424 5172 10452
rect 4764 10412 4770 10424
rect 5166 10412 5172 10424
rect 5224 10412 5230 10464
rect 10137 10455 10195 10461
rect 10137 10421 10149 10455
rect 10183 10452 10195 10455
rect 11330 10452 11336 10464
rect 10183 10424 11336 10452
rect 10183 10421 10195 10424
rect 10137 10415 10195 10421
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 12526 10412 12532 10464
rect 12584 10452 12590 10464
rect 14001 10455 14059 10461
rect 14001 10452 14013 10455
rect 12584 10424 14013 10452
rect 12584 10412 12590 10424
rect 14001 10421 14013 10424
rect 14047 10421 14059 10455
rect 14274 10452 14280 10464
rect 14235 10424 14280 10452
rect 14001 10415 14059 10421
rect 14274 10412 14280 10424
rect 14332 10412 14338 10464
rect 14366 10412 14372 10464
rect 14424 10452 14430 10464
rect 14645 10455 14703 10461
rect 14645 10452 14657 10455
rect 14424 10424 14657 10452
rect 14424 10412 14430 10424
rect 14645 10421 14657 10424
rect 14691 10421 14703 10455
rect 14645 10415 14703 10421
rect 1104 10362 15824 10384
rect 1104 10310 5912 10362
rect 5964 10310 5976 10362
rect 6028 10310 6040 10362
rect 6092 10310 6104 10362
rect 6156 10310 10843 10362
rect 10895 10310 10907 10362
rect 10959 10310 10971 10362
rect 11023 10310 11035 10362
rect 11087 10310 15824 10362
rect 1104 10288 15824 10310
rect 2225 10251 2283 10257
rect 2225 10217 2237 10251
rect 2271 10248 2283 10251
rect 2685 10251 2743 10257
rect 2685 10248 2697 10251
rect 2271 10220 2697 10248
rect 2271 10217 2283 10220
rect 2225 10211 2283 10217
rect 2685 10217 2697 10220
rect 2731 10217 2743 10251
rect 2685 10211 2743 10217
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 2869 10251 2927 10257
rect 2869 10248 2881 10251
rect 2832 10220 2881 10248
rect 2832 10208 2838 10220
rect 2869 10217 2881 10220
rect 2915 10217 2927 10251
rect 2869 10211 2927 10217
rect 4522 10208 4528 10260
rect 4580 10248 4586 10260
rect 7101 10251 7159 10257
rect 7101 10248 7113 10251
rect 4580 10220 7113 10248
rect 4580 10208 4586 10220
rect 7101 10217 7113 10220
rect 7147 10217 7159 10251
rect 7101 10211 7159 10217
rect 8757 10251 8815 10257
rect 8757 10217 8769 10251
rect 8803 10248 8815 10251
rect 8938 10248 8944 10260
rect 8803 10220 8944 10248
rect 8803 10217 8815 10220
rect 8757 10211 8815 10217
rect 8938 10208 8944 10220
rect 8996 10208 9002 10260
rect 9214 10208 9220 10260
rect 9272 10248 9278 10260
rect 11333 10251 11391 10257
rect 11333 10248 11345 10251
rect 9272 10220 11345 10248
rect 9272 10208 9278 10220
rect 11333 10217 11345 10220
rect 11379 10217 11391 10251
rect 11333 10211 11391 10217
rect 11606 10208 11612 10260
rect 11664 10248 11670 10260
rect 13630 10248 13636 10260
rect 11664 10220 13636 10248
rect 11664 10208 11670 10220
rect 13630 10208 13636 10220
rect 13688 10248 13694 10260
rect 13817 10251 13875 10257
rect 13817 10248 13829 10251
rect 13688 10220 13829 10248
rect 13688 10208 13694 10220
rect 13817 10217 13829 10220
rect 13863 10217 13875 10251
rect 14366 10248 14372 10260
rect 14327 10220 14372 10248
rect 13817 10211 13875 10217
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 2314 10180 2320 10192
rect 2275 10152 2320 10180
rect 2314 10140 2320 10152
rect 2372 10140 2378 10192
rect 4893 10183 4951 10189
rect 4893 10149 4905 10183
rect 4939 10180 4951 10183
rect 5074 10180 5080 10192
rect 4939 10152 5080 10180
rect 4939 10149 4951 10152
rect 4893 10143 4951 10149
rect 5074 10140 5080 10152
rect 5132 10180 5138 10192
rect 5350 10180 5356 10192
rect 5132 10152 5356 10180
rect 5132 10140 5138 10152
rect 5350 10140 5356 10152
rect 5408 10140 5414 10192
rect 5810 10140 5816 10192
rect 5868 10180 5874 10192
rect 5966 10183 6024 10189
rect 5966 10180 5978 10183
rect 5868 10152 5978 10180
rect 5868 10140 5874 10152
rect 5966 10149 5978 10152
rect 6012 10149 6024 10183
rect 5966 10143 6024 10149
rect 7006 10140 7012 10192
rect 7064 10180 7070 10192
rect 9125 10183 9183 10189
rect 7064 10152 9076 10180
rect 7064 10140 7070 10152
rect 3237 10115 3295 10121
rect 3237 10081 3249 10115
rect 3283 10112 3295 10115
rect 3878 10112 3884 10124
rect 3283 10084 3884 10112
rect 3283 10081 3295 10084
rect 3237 10075 3295 10081
rect 3878 10072 3884 10084
rect 3936 10112 3942 10124
rect 4798 10112 4804 10124
rect 3936 10084 4660 10112
rect 4759 10084 4804 10112
rect 3936 10072 3942 10084
rect 2501 10047 2559 10053
rect 2501 10013 2513 10047
rect 2547 10044 2559 10047
rect 3142 10044 3148 10056
rect 2547 10016 3148 10044
rect 2547 10013 2559 10016
rect 2501 10007 2559 10013
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 3326 10044 3332 10056
rect 3287 10016 3332 10044
rect 3326 10004 3332 10016
rect 3384 10004 3390 10056
rect 3418 10004 3424 10056
rect 3476 10044 3482 10056
rect 3476 10016 3521 10044
rect 3476 10004 3482 10016
rect 2777 9979 2835 9985
rect 2777 9945 2789 9979
rect 2823 9976 2835 9979
rect 4522 9976 4528 9988
rect 2823 9948 4528 9976
rect 2823 9945 2835 9948
rect 2777 9939 2835 9945
rect 4522 9936 4528 9948
rect 4580 9936 4586 9988
rect 1854 9908 1860 9920
rect 1815 9880 1860 9908
rect 1854 9868 1860 9880
rect 1912 9868 1918 9920
rect 4338 9868 4344 9920
rect 4396 9908 4402 9920
rect 4433 9911 4491 9917
rect 4433 9908 4445 9911
rect 4396 9880 4445 9908
rect 4396 9868 4402 9880
rect 4433 9877 4445 9880
rect 4479 9877 4491 9911
rect 4632 9908 4660 10084
rect 4798 10072 4804 10084
rect 4856 10072 4862 10124
rect 5442 10072 5448 10124
rect 5500 10112 5506 10124
rect 5721 10115 5779 10121
rect 5721 10112 5733 10115
rect 5500 10084 5733 10112
rect 5500 10072 5506 10084
rect 5721 10081 5733 10084
rect 5767 10112 5779 10115
rect 6270 10112 6276 10124
rect 5767 10084 6276 10112
rect 5767 10081 5779 10084
rect 5721 10075 5779 10081
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 8297 10115 8355 10121
rect 8297 10081 8309 10115
rect 8343 10112 8355 10115
rect 8662 10112 8668 10124
rect 8343 10084 8668 10112
rect 8343 10081 8355 10084
rect 8297 10075 8355 10081
rect 8662 10072 8668 10084
rect 8720 10072 8726 10124
rect 5074 10044 5080 10056
rect 5035 10016 5080 10044
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 8573 10047 8631 10053
rect 8573 10013 8585 10047
rect 8619 10044 8631 10047
rect 8846 10044 8852 10056
rect 8619 10016 8852 10044
rect 8619 10013 8631 10016
rect 8573 10007 8631 10013
rect 8404 9976 8432 10007
rect 8846 10004 8852 10016
rect 8904 10004 8910 10056
rect 8754 9976 8760 9988
rect 8404 9948 8760 9976
rect 8754 9936 8760 9948
rect 8812 9936 8818 9988
rect 9048 9976 9076 10152
rect 9125 10149 9137 10183
rect 9171 10180 9183 10183
rect 9398 10180 9404 10192
rect 9171 10152 9404 10180
rect 9171 10149 9183 10152
rect 9125 10143 9183 10149
rect 9398 10140 9404 10152
rect 9456 10140 9462 10192
rect 9674 10140 9680 10192
rect 9732 10180 9738 10192
rect 9732 10152 10456 10180
rect 9732 10140 9738 10152
rect 9858 10112 9864 10124
rect 9324 10084 9864 10112
rect 9324 10056 9352 10084
rect 9858 10072 9864 10084
rect 9916 10112 9922 10124
rect 10209 10115 10267 10121
rect 10209 10112 10221 10115
rect 9916 10084 10221 10112
rect 9916 10072 9922 10084
rect 10209 10081 10221 10084
rect 10255 10081 10267 10115
rect 10428 10112 10456 10152
rect 10502 10140 10508 10192
rect 10560 10180 10566 10192
rect 15102 10180 15108 10192
rect 10560 10152 15108 10180
rect 10560 10140 10566 10152
rect 15102 10140 15108 10152
rect 15160 10140 15166 10192
rect 12158 10112 12164 10124
rect 10428 10084 12164 10112
rect 10209 10075 10267 10081
rect 12158 10072 12164 10084
rect 12216 10112 12222 10124
rect 12345 10115 12403 10121
rect 12345 10112 12357 10115
rect 12216 10084 12357 10112
rect 12216 10072 12222 10084
rect 12345 10081 12357 10084
rect 12391 10081 12403 10115
rect 12345 10075 12403 10081
rect 13725 10115 13783 10121
rect 13725 10081 13737 10115
rect 13771 10112 13783 10115
rect 14090 10112 14096 10124
rect 13771 10084 14096 10112
rect 13771 10081 13783 10084
rect 13725 10075 13783 10081
rect 14090 10072 14096 10084
rect 14148 10072 14154 10124
rect 9122 10004 9128 10056
rect 9180 10044 9186 10056
rect 9217 10047 9275 10053
rect 9217 10044 9229 10047
rect 9180 10016 9229 10044
rect 9180 10004 9186 10016
rect 9217 10013 9229 10016
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 9306 10004 9312 10056
rect 9364 10044 9370 10056
rect 9364 10016 9409 10044
rect 9364 10004 9370 10016
rect 9766 10004 9772 10056
rect 9824 10044 9830 10056
rect 9953 10047 10011 10053
rect 9953 10044 9965 10047
rect 9824 10016 9965 10044
rect 9824 10004 9830 10016
rect 9953 10013 9965 10016
rect 9999 10013 10011 10047
rect 9953 10007 10011 10013
rect 12437 10047 12495 10053
rect 12437 10013 12449 10047
rect 12483 10013 12495 10047
rect 12437 10007 12495 10013
rect 12621 10047 12679 10053
rect 12621 10013 12633 10047
rect 12667 10013 12679 10047
rect 12621 10007 12679 10013
rect 9048 9948 9996 9976
rect 7466 9908 7472 9920
rect 4632 9880 7472 9908
rect 4433 9871 4491 9877
rect 7466 9868 7472 9880
rect 7524 9868 7530 9920
rect 7929 9911 7987 9917
rect 7929 9877 7941 9911
rect 7975 9908 7987 9911
rect 9766 9908 9772 9920
rect 7975 9880 9772 9908
rect 7975 9877 7987 9880
rect 7929 9871 7987 9877
rect 9766 9868 9772 9880
rect 9824 9868 9830 9920
rect 9968 9908 9996 9948
rect 11606 9908 11612 9920
rect 9968 9880 11612 9908
rect 11606 9868 11612 9880
rect 11664 9868 11670 9920
rect 11698 9868 11704 9920
rect 11756 9908 11762 9920
rect 11977 9911 12035 9917
rect 11977 9908 11989 9911
rect 11756 9880 11989 9908
rect 11756 9868 11762 9880
rect 11977 9877 11989 9880
rect 12023 9877 12035 9911
rect 12452 9908 12480 10007
rect 12636 9976 12664 10007
rect 12802 10004 12808 10056
rect 12860 10044 12866 10056
rect 12986 10044 12992 10056
rect 12860 10016 12992 10044
rect 12860 10004 12866 10016
rect 12986 10004 12992 10016
rect 13044 10004 13050 10056
rect 13998 10044 14004 10056
rect 13959 10016 14004 10044
rect 13998 10004 14004 10016
rect 14056 10004 14062 10056
rect 14016 9976 14044 10004
rect 12636 9948 14044 9976
rect 12618 9908 12624 9920
rect 12452 9880 12624 9908
rect 11977 9871 12035 9877
rect 12618 9868 12624 9880
rect 12676 9868 12682 9920
rect 12894 9868 12900 9920
rect 12952 9908 12958 9920
rect 13078 9908 13084 9920
rect 12952 9880 13084 9908
rect 12952 9868 12958 9880
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 13357 9911 13415 9917
rect 13357 9877 13369 9911
rect 13403 9908 13415 9911
rect 14366 9908 14372 9920
rect 13403 9880 14372 9908
rect 13403 9877 13415 9880
rect 13357 9871 13415 9877
rect 14366 9868 14372 9880
rect 14424 9868 14430 9920
rect 1104 9818 15824 9840
rect 1104 9766 3447 9818
rect 3499 9766 3511 9818
rect 3563 9766 3575 9818
rect 3627 9766 3639 9818
rect 3691 9766 8378 9818
rect 8430 9766 8442 9818
rect 8494 9766 8506 9818
rect 8558 9766 8570 9818
rect 8622 9766 13308 9818
rect 13360 9766 13372 9818
rect 13424 9766 13436 9818
rect 13488 9766 13500 9818
rect 13552 9766 15824 9818
rect 1104 9744 15824 9766
rect 3142 9664 3148 9716
rect 3200 9704 3206 9716
rect 7098 9704 7104 9716
rect 3200 9676 7104 9704
rect 3200 9664 3206 9676
rect 7098 9664 7104 9676
rect 7156 9704 7162 9716
rect 7834 9704 7840 9716
rect 7156 9676 7840 9704
rect 7156 9664 7162 9676
rect 7834 9664 7840 9676
rect 7892 9664 7898 9716
rect 9232 9676 10272 9704
rect 1762 9636 1768 9648
rect 1723 9608 1768 9636
rect 1762 9596 1768 9608
rect 1820 9596 1826 9648
rect 3878 9596 3884 9648
rect 3936 9636 3942 9648
rect 5445 9639 5503 9645
rect 5445 9636 5457 9639
rect 3936 9608 5457 9636
rect 3936 9596 3942 9608
rect 5445 9605 5457 9608
rect 5491 9605 5503 9639
rect 5445 9599 5503 9605
rect 7650 9596 7656 9648
rect 7708 9636 7714 9648
rect 8018 9636 8024 9648
rect 7708 9608 8024 9636
rect 7708 9596 7714 9608
rect 8018 9596 8024 9608
rect 8076 9636 8082 9648
rect 8757 9639 8815 9645
rect 8757 9636 8769 9639
rect 8076 9608 8769 9636
rect 8076 9596 8082 9608
rect 8757 9605 8769 9608
rect 8803 9605 8815 9639
rect 8757 9599 8815 9605
rect 8938 9596 8944 9648
rect 8996 9636 9002 9648
rect 9232 9636 9260 9676
rect 8996 9608 9260 9636
rect 9309 9639 9367 9645
rect 8996 9596 9002 9608
rect 9309 9605 9321 9639
rect 9355 9636 9367 9639
rect 10134 9636 10140 9648
rect 9355 9608 9996 9636
rect 10095 9608 10140 9636
rect 9355 9605 9367 9608
rect 9309 9599 9367 9605
rect 2409 9571 2467 9577
rect 2409 9537 2421 9571
rect 2455 9568 2467 9571
rect 2498 9568 2504 9580
rect 2455 9540 2504 9568
rect 2455 9537 2467 9540
rect 2409 9531 2467 9537
rect 2498 9528 2504 9540
rect 2556 9528 2562 9580
rect 5074 9568 5080 9580
rect 5035 9540 5080 9568
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 6549 9571 6607 9577
rect 6549 9537 6561 9571
rect 6595 9568 6607 9571
rect 7742 9568 7748 9580
rect 6595 9540 7748 9568
rect 6595 9537 6607 9540
rect 6549 9531 6607 9537
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9537 9919 9571
rect 9968 9568 9996 9608
rect 10134 9596 10140 9608
rect 10192 9596 10198 9648
rect 10244 9636 10272 9676
rect 12618 9664 12624 9716
rect 12676 9704 12682 9716
rect 12676 9676 12756 9704
rect 12676 9664 12682 9676
rect 11330 9636 11336 9648
rect 10244 9608 11192 9636
rect 11291 9608 11336 9636
rect 10318 9568 10324 9580
rect 9968 9540 10324 9568
rect 9861 9531 9919 9537
rect 1854 9460 1860 9512
rect 1912 9500 1918 9512
rect 2133 9503 2191 9509
rect 2133 9500 2145 9503
rect 1912 9472 2145 9500
rect 1912 9460 1918 9472
rect 2133 9469 2145 9472
rect 2179 9469 2191 9503
rect 2133 9463 2191 9469
rect 2774 9460 2780 9512
rect 2832 9500 2838 9512
rect 4614 9500 4620 9512
rect 2832 9472 2877 9500
rect 2976 9472 4620 9500
rect 2832 9460 2838 9472
rect 2225 9435 2283 9441
rect 2225 9401 2237 9435
rect 2271 9432 2283 9435
rect 2976 9432 3004 9472
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 4706 9460 4712 9512
rect 4764 9500 4770 9512
rect 5629 9503 5687 9509
rect 5629 9500 5641 9503
rect 4764 9472 5641 9500
rect 4764 9460 4770 9472
rect 5629 9469 5641 9472
rect 5675 9469 5687 9503
rect 5629 9463 5687 9469
rect 6273 9503 6331 9509
rect 6273 9469 6285 9503
rect 6319 9500 6331 9503
rect 8386 9500 8392 9512
rect 6319 9472 8392 9500
rect 6319 9469 6331 9472
rect 6273 9463 6331 9469
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 8846 9460 8852 9512
rect 8904 9500 8910 9512
rect 8904 9472 9536 9500
rect 8904 9460 8910 9472
rect 2271 9404 3004 9432
rect 3044 9435 3102 9441
rect 2271 9401 2283 9404
rect 2225 9395 2283 9401
rect 3044 9401 3056 9435
rect 3090 9432 3102 9435
rect 3510 9432 3516 9444
rect 3090 9404 3516 9432
rect 3090 9401 3102 9404
rect 3044 9395 3102 9401
rect 3510 9392 3516 9404
rect 3568 9392 3574 9444
rect 4893 9435 4951 9441
rect 4893 9432 4905 9435
rect 4632 9404 4905 9432
rect 4632 9376 4660 9404
rect 4893 9401 4905 9404
rect 4939 9432 4951 9435
rect 6914 9432 6920 9444
rect 4939 9404 6920 9432
rect 4939 9401 4951 9404
rect 4893 9395 4951 9401
rect 6914 9392 6920 9404
rect 6972 9392 6978 9444
rect 7469 9435 7527 9441
rect 7469 9401 7481 9435
rect 7515 9432 7527 9435
rect 9398 9432 9404 9444
rect 7515 9404 9404 9432
rect 7515 9401 7527 9404
rect 7469 9395 7527 9401
rect 9398 9392 9404 9404
rect 9456 9392 9462 9444
rect 9508 9432 9536 9472
rect 9674 9460 9680 9512
rect 9732 9500 9738 9512
rect 9769 9503 9827 9509
rect 9769 9500 9781 9503
rect 9732 9472 9781 9500
rect 9732 9460 9738 9472
rect 9769 9469 9781 9472
rect 9815 9469 9827 9503
rect 9769 9463 9827 9469
rect 9876 9432 9904 9531
rect 10318 9528 10324 9540
rect 10376 9528 10382 9580
rect 10686 9568 10692 9580
rect 10647 9540 10692 9568
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 11164 9568 11192 9608
rect 11330 9596 11336 9608
rect 11388 9596 11394 9648
rect 12437 9639 12495 9645
rect 12437 9605 12449 9639
rect 12483 9636 12495 9639
rect 12728 9636 12756 9676
rect 12483 9608 12756 9636
rect 12912 9676 14044 9704
rect 12483 9605 12495 9608
rect 12437 9599 12495 9605
rect 11790 9568 11796 9580
rect 11164 9540 11796 9568
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 11977 9571 12035 9577
rect 11977 9537 11989 9571
rect 12023 9568 12035 9571
rect 12526 9568 12532 9580
rect 12023 9540 12532 9568
rect 12023 9537 12035 9540
rect 11977 9531 12035 9537
rect 12526 9528 12532 9540
rect 12584 9568 12590 9580
rect 12912 9568 12940 9676
rect 13449 9639 13507 9645
rect 13449 9605 13461 9639
rect 13495 9605 13507 9639
rect 13449 9599 13507 9605
rect 13078 9568 13084 9580
rect 12584 9540 12940 9568
rect 13039 9540 13084 9568
rect 12584 9528 12590 9540
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 10410 9460 10416 9512
rect 10468 9500 10474 9512
rect 10597 9503 10655 9509
rect 10597 9500 10609 9503
rect 10468 9472 10609 9500
rect 10468 9460 10474 9472
rect 10597 9469 10609 9472
rect 10643 9469 10655 9503
rect 11698 9500 11704 9512
rect 11659 9472 11704 9500
rect 10597 9463 10655 9469
rect 11698 9460 11704 9472
rect 11756 9460 11762 9512
rect 11882 9460 11888 9512
rect 11940 9500 11946 9512
rect 13464 9500 13492 9599
rect 14016 9577 14044 9676
rect 14001 9571 14059 9577
rect 14001 9537 14013 9571
rect 14047 9537 14059 9571
rect 14001 9531 14059 9537
rect 11940 9472 13492 9500
rect 13817 9503 13875 9509
rect 11940 9460 11946 9472
rect 13817 9469 13829 9503
rect 13863 9500 13875 9503
rect 14274 9500 14280 9512
rect 13863 9472 14280 9500
rect 13863 9469 13875 9472
rect 13817 9463 13875 9469
rect 14274 9460 14280 9472
rect 14332 9460 14338 9512
rect 9508 9404 9904 9432
rect 11793 9435 11851 9441
rect 11793 9401 11805 9435
rect 11839 9432 11851 9435
rect 13262 9432 13268 9444
rect 11839 9404 13268 9432
rect 11839 9401 11851 9404
rect 11793 9395 11851 9401
rect 13262 9392 13268 9404
rect 13320 9392 13326 9444
rect 13909 9435 13967 9441
rect 13909 9401 13921 9435
rect 13955 9432 13967 9435
rect 14366 9432 14372 9444
rect 13955 9404 14372 9432
rect 13955 9401 13967 9404
rect 13909 9395 13967 9401
rect 14366 9392 14372 9404
rect 14424 9392 14430 9444
rect 2406 9324 2412 9376
rect 2464 9364 2470 9376
rect 3786 9364 3792 9376
rect 2464 9336 3792 9364
rect 2464 9324 2470 9336
rect 3786 9324 3792 9336
rect 3844 9364 3850 9376
rect 4157 9367 4215 9373
rect 4157 9364 4169 9367
rect 3844 9336 4169 9364
rect 3844 9324 3850 9336
rect 4157 9333 4169 9336
rect 4203 9333 4215 9367
rect 4157 9327 4215 9333
rect 4430 9324 4436 9376
rect 4488 9364 4494 9376
rect 4488 9336 4533 9364
rect 4488 9324 4494 9336
rect 4614 9324 4620 9376
rect 4672 9324 4678 9376
rect 4801 9367 4859 9373
rect 4801 9333 4813 9367
rect 4847 9364 4859 9367
rect 5166 9364 5172 9376
rect 4847 9336 5172 9364
rect 4847 9333 4859 9336
rect 4801 9327 4859 9333
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 5810 9324 5816 9376
rect 5868 9364 5874 9376
rect 5905 9367 5963 9373
rect 5905 9364 5917 9367
rect 5868 9336 5917 9364
rect 5868 9324 5874 9336
rect 5905 9333 5917 9336
rect 5951 9333 5963 9367
rect 5905 9327 5963 9333
rect 6365 9367 6423 9373
rect 6365 9333 6377 9367
rect 6411 9364 6423 9367
rect 8294 9364 8300 9376
rect 6411 9336 8300 9364
rect 6411 9333 6423 9336
rect 6365 9327 6423 9333
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 8938 9324 8944 9376
rect 8996 9364 9002 9376
rect 9122 9364 9128 9376
rect 8996 9336 9128 9364
rect 8996 9324 9002 9336
rect 9122 9324 9128 9336
rect 9180 9324 9186 9376
rect 9677 9367 9735 9373
rect 9677 9333 9689 9367
rect 9723 9364 9735 9367
rect 9858 9364 9864 9376
rect 9723 9336 9864 9364
rect 9723 9333 9735 9336
rect 9677 9327 9735 9333
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 10042 9324 10048 9376
rect 10100 9364 10106 9376
rect 10505 9367 10563 9373
rect 10505 9364 10517 9367
rect 10100 9336 10517 9364
rect 10100 9324 10106 9336
rect 10505 9333 10517 9336
rect 10551 9333 10563 9367
rect 10505 9327 10563 9333
rect 12066 9324 12072 9376
rect 12124 9364 12130 9376
rect 12805 9367 12863 9373
rect 12805 9364 12817 9367
rect 12124 9336 12817 9364
rect 12124 9324 12130 9336
rect 12805 9333 12817 9336
rect 12851 9333 12863 9367
rect 12805 9327 12863 9333
rect 12894 9324 12900 9376
rect 12952 9364 12958 9376
rect 12952 9336 12997 9364
rect 12952 9324 12958 9336
rect 1104 9274 15824 9296
rect 1104 9222 5912 9274
rect 5964 9222 5976 9274
rect 6028 9222 6040 9274
rect 6092 9222 6104 9274
rect 6156 9222 10843 9274
rect 10895 9222 10907 9274
rect 10959 9222 10971 9274
rect 11023 9222 11035 9274
rect 11087 9222 15824 9274
rect 1104 9200 15824 9222
rect 3510 9160 3516 9172
rect 3471 9132 3516 9160
rect 3510 9120 3516 9132
rect 3568 9120 3574 9172
rect 3786 9120 3792 9172
rect 3844 9160 3850 9172
rect 4065 9163 4123 9169
rect 3844 9132 4016 9160
rect 3844 9120 3850 9132
rect 2774 9092 2780 9104
rect 2148 9064 2780 9092
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 8993 1455 9027
rect 1670 9024 1676 9036
rect 1631 8996 1676 9024
rect 1397 8987 1455 8993
rect 1412 8820 1440 8987
rect 1670 8984 1676 8996
rect 1728 8984 1734 9036
rect 2148 9033 2176 9064
rect 2774 9052 2780 9064
rect 2832 9092 2838 9104
rect 3878 9092 3884 9104
rect 2832 9064 3884 9092
rect 2832 9052 2838 9064
rect 3878 9052 3884 9064
rect 3936 9052 3942 9104
rect 3988 9092 4016 9132
rect 4065 9129 4077 9163
rect 4111 9160 4123 9163
rect 4798 9160 4804 9172
rect 4111 9132 4804 9160
rect 4111 9129 4123 9132
rect 4065 9123 4123 9129
rect 4798 9120 4804 9132
rect 4856 9120 4862 9172
rect 6365 9163 6423 9169
rect 6365 9129 6377 9163
rect 6411 9160 6423 9163
rect 8481 9163 8539 9169
rect 6411 9132 6868 9160
rect 6411 9129 6423 9132
rect 6365 9123 6423 9129
rect 5230 9095 5288 9101
rect 5230 9092 5242 9095
rect 3988 9064 5242 9092
rect 5230 9061 5242 9064
rect 5276 9061 5288 9095
rect 5230 9055 5288 9061
rect 2133 9027 2191 9033
rect 2133 8993 2145 9027
rect 2179 8993 2191 9027
rect 2133 8987 2191 8993
rect 2400 9027 2458 9033
rect 2400 8993 2412 9027
rect 2446 9024 2458 9027
rect 4246 9024 4252 9036
rect 2446 8996 4252 9024
rect 2446 8993 2458 8996
rect 2400 8987 2458 8993
rect 4246 8984 4252 8996
rect 4304 8984 4310 9036
rect 4522 9024 4528 9036
rect 4483 8996 4528 9024
rect 4522 8984 4528 8996
rect 4580 8984 4586 9036
rect 6840 9024 6868 9132
rect 8481 9129 8493 9163
rect 8527 9160 8539 9163
rect 8662 9160 8668 9172
rect 8527 9132 8668 9160
rect 8527 9129 8539 9132
rect 8481 9123 8539 9129
rect 8662 9120 8668 9132
rect 8720 9120 8726 9172
rect 8849 9163 8907 9169
rect 8849 9129 8861 9163
rect 8895 9160 8907 9163
rect 9122 9160 9128 9172
rect 8895 9132 9128 9160
rect 8895 9129 8907 9132
rect 8849 9123 8907 9129
rect 9122 9120 9128 9132
rect 9180 9120 9186 9172
rect 9677 9163 9735 9169
rect 9677 9129 9689 9163
rect 9723 9160 9735 9163
rect 9858 9160 9864 9172
rect 9723 9132 9864 9160
rect 9723 9129 9735 9132
rect 9677 9123 9735 9129
rect 9858 9120 9864 9132
rect 9916 9120 9922 9172
rect 12342 9160 12348 9172
rect 9968 9132 12348 9160
rect 8294 9052 8300 9104
rect 8352 9092 8358 9104
rect 8938 9092 8944 9104
rect 8352 9064 8944 9092
rect 8352 9052 8358 9064
rect 8938 9052 8944 9064
rect 8996 9092 9002 9104
rect 9968 9092 9996 9132
rect 12342 9120 12348 9132
rect 12400 9120 12406 9172
rect 12437 9163 12495 9169
rect 12437 9129 12449 9163
rect 12483 9160 12495 9163
rect 13909 9163 13967 9169
rect 13909 9160 13921 9163
rect 12483 9132 13921 9160
rect 12483 9129 12495 9132
rect 12437 9123 12495 9129
rect 13909 9129 13921 9132
rect 13955 9129 13967 9163
rect 13909 9123 13967 9129
rect 8996 9064 9996 9092
rect 10045 9095 10103 9101
rect 8996 9052 9002 9064
rect 10045 9061 10057 9095
rect 10091 9092 10103 9095
rect 11606 9092 11612 9104
rect 10091 9064 11612 9092
rect 10091 9061 10103 9064
rect 10045 9055 10103 9061
rect 11606 9052 11612 9064
rect 11664 9052 11670 9104
rect 12897 9095 12955 9101
rect 12897 9092 12909 9095
rect 12452 9064 12909 9092
rect 12452 9036 12480 9064
rect 12897 9061 12909 9064
rect 12943 9092 12955 9095
rect 12986 9092 12992 9104
rect 12943 9064 12992 9092
rect 12943 9061 12955 9064
rect 12897 9055 12955 9061
rect 12986 9052 12992 9064
rect 13044 9052 13050 9104
rect 13630 9052 13636 9104
rect 13688 9092 13694 9104
rect 15286 9092 15292 9104
rect 13688 9064 15292 9092
rect 13688 9052 13694 9064
rect 15286 9052 15292 9064
rect 15344 9052 15350 9104
rect 6908 9027 6966 9033
rect 6908 9024 6920 9027
rect 5000 8996 6040 9024
rect 6840 8996 6920 9024
rect 3878 8916 3884 8968
rect 3936 8956 3942 8968
rect 5000 8965 5028 8996
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 3936 8928 4997 8956
rect 3936 8916 3942 8928
rect 4985 8925 4997 8928
rect 5031 8925 5043 8959
rect 6012 8956 6040 8996
rect 6908 8993 6920 8996
rect 6954 9024 6966 9027
rect 7374 9024 7380 9036
rect 6954 8996 7380 9024
rect 6954 8993 6966 8996
rect 6908 8987 6966 8993
rect 7374 8984 7380 8996
rect 7432 8984 7438 9036
rect 8386 8984 8392 9036
rect 8444 9024 8450 9036
rect 9030 9024 9036 9036
rect 8444 8996 9036 9024
rect 8444 8984 8450 8996
rect 9030 8984 9036 8996
rect 9088 9024 9094 9036
rect 10778 9024 10784 9036
rect 9088 8996 10784 9024
rect 9088 8984 9094 8996
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 10956 9027 11014 9033
rect 10956 8993 10968 9027
rect 11002 9024 11014 9027
rect 11330 9024 11336 9036
rect 11002 8996 11336 9024
rect 11002 8993 11014 8996
rect 10956 8987 11014 8993
rect 11330 8984 11336 8996
rect 11388 8984 11394 9036
rect 11514 8984 11520 9036
rect 11572 9024 11578 9036
rect 11974 9024 11980 9036
rect 11572 8996 11980 9024
rect 11572 8984 11578 8996
rect 11974 8984 11980 8996
rect 12032 8984 12038 9036
rect 12434 8984 12440 9036
rect 12492 8984 12498 9036
rect 12802 9024 12808 9036
rect 12763 8996 12808 9024
rect 12802 8984 12808 8996
rect 12860 8984 12866 9036
rect 13814 9024 13820 9036
rect 13775 8996 13820 9024
rect 13814 8984 13820 8996
rect 13872 8984 13878 9036
rect 6638 8956 6644 8968
rect 6012 8928 6644 8956
rect 4985 8919 5043 8925
rect 6638 8916 6644 8928
rect 6696 8956 6702 8968
rect 6696 8928 6789 8956
rect 6696 8916 6702 8928
rect 7834 8916 7840 8968
rect 7892 8956 7898 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 7892 8928 8953 8956
rect 7892 8916 7898 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 8021 8891 8079 8897
rect 8021 8857 8033 8891
rect 8067 8888 8079 8891
rect 9030 8888 9036 8900
rect 8067 8860 9036 8888
rect 8067 8857 8079 8860
rect 8021 8851 8079 8857
rect 9030 8848 9036 8860
rect 9088 8888 9094 8900
rect 9140 8888 9168 8919
rect 9858 8916 9864 8968
rect 9916 8956 9922 8968
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9916 8928 10149 8956
rect 9916 8916 9922 8928
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8925 10287 8959
rect 10686 8956 10692 8968
rect 10647 8928 10692 8956
rect 10229 8919 10287 8925
rect 10244 8888 10272 8919
rect 10686 8916 10692 8928
rect 10744 8916 10750 8968
rect 13078 8956 13084 8968
rect 13039 8928 13084 8956
rect 13078 8916 13084 8928
rect 13136 8916 13142 8968
rect 13998 8956 14004 8968
rect 13959 8928 14004 8956
rect 13998 8916 14004 8928
rect 14056 8916 14062 8968
rect 9088 8860 10272 8888
rect 12069 8891 12127 8897
rect 9088 8848 9094 8860
rect 12069 8857 12081 8891
rect 12115 8888 12127 8891
rect 13096 8888 13124 8916
rect 12115 8860 13124 8888
rect 12115 8857 12127 8860
rect 12069 8851 12127 8857
rect 13262 8848 13268 8900
rect 13320 8888 13326 8900
rect 13449 8891 13507 8897
rect 13449 8888 13461 8891
rect 13320 8860 13461 8888
rect 13320 8848 13326 8860
rect 13449 8857 13461 8860
rect 13495 8857 13507 8891
rect 13449 8851 13507 8857
rect 11698 8820 11704 8832
rect 1412 8792 11704 8820
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 12158 8780 12164 8832
rect 12216 8820 12222 8832
rect 13722 8820 13728 8832
rect 12216 8792 13728 8820
rect 12216 8780 12222 8792
rect 13722 8780 13728 8792
rect 13780 8780 13786 8832
rect 1104 8730 15824 8752
rect 1104 8678 3447 8730
rect 3499 8678 3511 8730
rect 3563 8678 3575 8730
rect 3627 8678 3639 8730
rect 3691 8678 8378 8730
rect 8430 8678 8442 8730
rect 8494 8678 8506 8730
rect 8558 8678 8570 8730
rect 8622 8678 13308 8730
rect 13360 8678 13372 8730
rect 13424 8678 13436 8730
rect 13488 8678 13500 8730
rect 13552 8678 15824 8730
rect 1104 8656 15824 8678
rect 4430 8616 4436 8628
rect 3804 8588 4436 8616
rect 2777 8551 2835 8557
rect 2777 8517 2789 8551
rect 2823 8517 2835 8551
rect 2777 8511 2835 8517
rect 2406 8480 2412 8492
rect 2367 8452 2412 8480
rect 2406 8440 2412 8452
rect 2464 8440 2470 8492
rect 2133 8415 2191 8421
rect 2133 8381 2145 8415
rect 2179 8412 2191 8415
rect 2792 8412 2820 8511
rect 3326 8480 3332 8492
rect 3287 8452 3332 8480
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 2179 8384 2820 8412
rect 3237 8415 3295 8421
rect 2179 8381 2191 8384
rect 2133 8375 2191 8381
rect 3237 8381 3249 8415
rect 3283 8412 3295 8415
rect 3804 8412 3832 8588
rect 4430 8576 4436 8588
rect 4488 8576 4494 8628
rect 5718 8616 5724 8628
rect 5679 8588 5724 8616
rect 5718 8576 5724 8588
rect 5776 8576 5782 8628
rect 6730 8576 6736 8628
rect 6788 8576 6794 8628
rect 8573 8619 8631 8625
rect 8573 8585 8585 8619
rect 8619 8616 8631 8619
rect 8754 8616 8760 8628
rect 8619 8588 8760 8616
rect 8619 8585 8631 8588
rect 8573 8579 8631 8585
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 10686 8616 10692 8628
rect 9968 8588 10692 8616
rect 6748 8548 6776 8576
rect 4172 8520 6776 8548
rect 8297 8551 8355 8557
rect 4172 8421 4200 8520
rect 8297 8517 8309 8551
rect 8343 8548 8355 8551
rect 8662 8548 8668 8560
rect 8343 8520 8668 8548
rect 8343 8517 8355 8520
rect 8297 8511 8355 8517
rect 8662 8508 8668 8520
rect 8720 8548 8726 8560
rect 8846 8548 8852 8560
rect 8720 8520 8852 8548
rect 8720 8508 8726 8520
rect 8846 8508 8852 8520
rect 8904 8508 8910 8560
rect 9677 8551 9735 8557
rect 8956 8520 9260 8548
rect 4246 8440 4252 8492
rect 4304 8480 4310 8492
rect 4341 8483 4399 8489
rect 4341 8480 4353 8483
rect 4304 8452 4353 8480
rect 4304 8440 4310 8452
rect 4341 8449 4353 8452
rect 4387 8480 4399 8483
rect 5074 8480 5080 8492
rect 4387 8452 5080 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 5074 8440 5080 8452
rect 5132 8480 5138 8492
rect 5442 8480 5448 8492
rect 5132 8452 5448 8480
rect 5132 8440 5138 8452
rect 5442 8440 5448 8452
rect 5500 8440 5506 8492
rect 5810 8440 5816 8492
rect 5868 8480 5874 8492
rect 6181 8483 6239 8489
rect 6181 8480 6193 8483
rect 5868 8452 6193 8480
rect 5868 8440 5874 8452
rect 6181 8449 6193 8452
rect 6227 8449 6239 8483
rect 6181 8443 6239 8449
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8480 6423 8483
rect 6454 8480 6460 8492
rect 6411 8452 6460 8480
rect 6411 8449 6423 8452
rect 6365 8443 6423 8449
rect 6454 8440 6460 8452
rect 6512 8440 6518 8492
rect 6638 8440 6644 8492
rect 6696 8480 6702 8492
rect 6917 8483 6975 8489
rect 6917 8480 6929 8483
rect 6696 8452 6929 8480
rect 6696 8440 6702 8452
rect 6917 8449 6929 8452
rect 6963 8449 6975 8483
rect 6917 8443 6975 8449
rect 7926 8440 7932 8492
rect 7984 8480 7990 8492
rect 8956 8480 8984 8520
rect 7984 8452 8984 8480
rect 7984 8440 7990 8452
rect 9030 8440 9036 8492
rect 9088 8480 9094 8492
rect 9125 8483 9183 8489
rect 9125 8480 9137 8483
rect 9088 8452 9137 8480
rect 9088 8440 9094 8452
rect 9125 8449 9137 8452
rect 9171 8449 9183 8483
rect 9125 8443 9183 8449
rect 3283 8384 3832 8412
rect 4157 8415 4215 8421
rect 3283 8381 3295 8384
rect 3237 8375 3295 8381
rect 4157 8381 4169 8415
rect 4203 8381 4215 8415
rect 4157 8375 4215 8381
rect 5169 8415 5227 8421
rect 5169 8381 5181 8415
rect 5215 8412 5227 8415
rect 6822 8412 6828 8424
rect 5215 8384 6828 8412
rect 5215 8381 5227 8384
rect 5169 8375 5227 8381
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 7184 8415 7242 8421
rect 7184 8381 7196 8415
rect 7230 8412 7242 8415
rect 9048 8412 9076 8440
rect 7230 8384 9076 8412
rect 7230 8381 7242 8384
rect 7184 8375 7242 8381
rect 2225 8347 2283 8353
rect 2225 8313 2237 8347
rect 2271 8344 2283 8347
rect 2958 8344 2964 8356
rect 2271 8316 2964 8344
rect 2271 8313 2283 8316
rect 2225 8307 2283 8313
rect 2958 8304 2964 8316
rect 3016 8304 3022 8356
rect 3145 8347 3203 8353
rect 3145 8313 3157 8347
rect 3191 8344 3203 8347
rect 4338 8344 4344 8356
rect 3191 8316 4344 8344
rect 3191 8313 3203 8316
rect 3145 8307 3203 8313
rect 4338 8304 4344 8316
rect 4396 8304 4402 8356
rect 4430 8304 4436 8356
rect 4488 8344 4494 8356
rect 5074 8344 5080 8356
rect 4488 8316 5080 8344
rect 4488 8304 4494 8316
rect 5074 8304 5080 8316
rect 5132 8304 5138 8356
rect 5261 8347 5319 8353
rect 5261 8313 5273 8347
rect 5307 8344 5319 8347
rect 5534 8344 5540 8356
rect 5307 8316 5540 8344
rect 5307 8313 5319 8316
rect 5261 8307 5319 8313
rect 5534 8304 5540 8316
rect 5592 8304 5598 8356
rect 6089 8347 6147 8353
rect 6089 8313 6101 8347
rect 6135 8344 6147 8347
rect 6362 8344 6368 8356
rect 6135 8316 6368 8344
rect 6135 8313 6147 8316
rect 6089 8307 6147 8313
rect 6362 8304 6368 8316
rect 6420 8304 6426 8356
rect 7282 8304 7288 8356
rect 7340 8344 7346 8356
rect 9033 8347 9091 8353
rect 9033 8344 9045 8347
rect 7340 8316 9045 8344
rect 7340 8304 7346 8316
rect 9033 8313 9045 8316
rect 9079 8313 9091 8347
rect 9232 8344 9260 8520
rect 9677 8517 9689 8551
rect 9723 8548 9735 8551
rect 9968 8548 9996 8588
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 10870 8576 10876 8628
rect 10928 8616 10934 8628
rect 12618 8616 12624 8628
rect 10928 8588 12624 8616
rect 10928 8576 10934 8588
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 14185 8619 14243 8625
rect 14185 8616 14197 8619
rect 14056 8588 14197 8616
rect 14056 8576 14062 8588
rect 14185 8585 14197 8588
rect 14231 8585 14243 8619
rect 14185 8579 14243 8585
rect 9723 8520 9996 8548
rect 9723 8517 9735 8520
rect 9677 8511 9735 8517
rect 9968 8489 9996 8520
rect 11238 8508 11244 8560
rect 11296 8548 11302 8560
rect 12158 8548 12164 8560
rect 11296 8520 12164 8548
rect 11296 8508 11302 8520
rect 12158 8508 12164 8520
rect 12216 8508 12222 8560
rect 9953 8483 10011 8489
rect 9953 8449 9965 8483
rect 9999 8449 10011 8483
rect 11606 8480 11612 8492
rect 11567 8452 11612 8480
rect 9953 8443 10011 8449
rect 11606 8440 11612 8452
rect 11664 8440 11670 8492
rect 9861 8415 9919 8421
rect 9861 8381 9873 8415
rect 9907 8412 9919 8415
rect 10594 8412 10600 8424
rect 9907 8384 10600 8412
rect 9907 8381 9919 8384
rect 9861 8375 9919 8381
rect 10594 8372 10600 8384
rect 10652 8372 10658 8424
rect 10686 8372 10692 8424
rect 10744 8412 10750 8424
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 10744 8384 12817 8412
rect 10744 8372 10750 8384
rect 12805 8381 12817 8384
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 10220 8347 10278 8353
rect 9232 8316 10180 8344
rect 9033 8307 9091 8313
rect 1486 8236 1492 8288
rect 1544 8276 1550 8288
rect 1765 8279 1823 8285
rect 1765 8276 1777 8279
rect 1544 8248 1777 8276
rect 1544 8236 1550 8248
rect 1765 8245 1777 8248
rect 1811 8245 1823 8279
rect 3786 8276 3792 8288
rect 3747 8248 3792 8276
rect 1765 8239 1823 8245
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 4246 8276 4252 8288
rect 4207 8248 4252 8276
rect 4246 8236 4252 8248
rect 4304 8236 4310 8288
rect 4798 8276 4804 8288
rect 4759 8248 4804 8276
rect 4798 8236 4804 8248
rect 4856 8236 4862 8288
rect 8754 8236 8760 8288
rect 8812 8276 8818 8288
rect 8941 8279 8999 8285
rect 8941 8276 8953 8279
rect 8812 8248 8953 8276
rect 8812 8236 8818 8248
rect 8941 8245 8953 8248
rect 8987 8276 8999 8279
rect 9398 8276 9404 8288
rect 8987 8248 9404 8276
rect 8987 8245 8999 8248
rect 8941 8239 8999 8245
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 10152 8276 10180 8316
rect 10220 8313 10232 8347
rect 10266 8344 10278 8347
rect 11054 8344 11060 8356
rect 10266 8316 11060 8344
rect 10266 8313 10278 8316
rect 10220 8307 10278 8313
rect 11054 8304 11060 8316
rect 11112 8304 11118 8356
rect 12526 8344 12532 8356
rect 11164 8316 12532 8344
rect 11164 8276 11192 8316
rect 12526 8304 12532 8316
rect 12584 8304 12590 8356
rect 13078 8353 13084 8356
rect 13072 8344 13084 8353
rect 12991 8316 13084 8344
rect 13072 8307 13084 8316
rect 13136 8344 13142 8356
rect 13262 8344 13268 8356
rect 13136 8316 13268 8344
rect 13078 8304 13084 8307
rect 13136 8304 13142 8316
rect 13262 8304 13268 8316
rect 13320 8304 13326 8356
rect 11330 8276 11336 8288
rect 10152 8248 11192 8276
rect 11291 8248 11336 8276
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 11606 8236 11612 8288
rect 11664 8276 11670 8288
rect 12250 8276 12256 8288
rect 11664 8248 12256 8276
rect 11664 8236 11670 8248
rect 12250 8236 12256 8248
rect 12308 8276 12314 8288
rect 12894 8276 12900 8288
rect 12308 8248 12900 8276
rect 12308 8236 12314 8248
rect 12894 8236 12900 8248
rect 12952 8236 12958 8288
rect 1104 8186 15824 8208
rect 1104 8134 5912 8186
rect 5964 8134 5976 8186
rect 6028 8134 6040 8186
rect 6092 8134 6104 8186
rect 6156 8134 10843 8186
rect 10895 8134 10907 8186
rect 10959 8134 10971 8186
rect 11023 8134 11035 8186
rect 11087 8134 15824 8186
rect 1104 8112 15824 8134
rect 2958 8072 2964 8084
rect 2919 8044 2964 8072
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 3329 8075 3387 8081
rect 3329 8041 3341 8075
rect 3375 8072 3387 8075
rect 3786 8072 3792 8084
rect 3375 8044 3792 8072
rect 3375 8041 3387 8044
rect 3329 8035 3387 8041
rect 3786 8032 3792 8044
rect 3844 8032 3850 8084
rect 4157 8075 4215 8081
rect 4157 8041 4169 8075
rect 4203 8072 4215 8075
rect 4246 8072 4252 8084
rect 4203 8044 4252 8072
rect 4203 8041 4215 8044
rect 4157 8035 4215 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 5166 8072 5172 8084
rect 4571 8044 5172 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 5442 8032 5448 8084
rect 5500 8072 5506 8084
rect 6549 8075 6607 8081
rect 6549 8072 6561 8075
rect 5500 8044 6561 8072
rect 5500 8032 5506 8044
rect 6549 8041 6561 8044
rect 6595 8041 6607 8075
rect 6549 8035 6607 8041
rect 6825 8075 6883 8081
rect 6825 8041 6837 8075
rect 6871 8072 6883 8075
rect 7282 8072 7288 8084
rect 6871 8044 7288 8072
rect 6871 8041 6883 8044
rect 6825 8035 6883 8041
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 8573 8075 8631 8081
rect 8573 8041 8585 8075
rect 8619 8072 8631 8075
rect 9674 8072 9680 8084
rect 8619 8044 9680 8072
rect 8619 8041 8631 8044
rect 8573 8035 8631 8041
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 10045 8075 10103 8081
rect 10045 8041 10057 8075
rect 10091 8072 10103 8075
rect 10318 8072 10324 8084
rect 10091 8044 10324 8072
rect 10091 8041 10103 8044
rect 10045 8035 10103 8041
rect 10318 8032 10324 8044
rect 10376 8032 10382 8084
rect 10689 8075 10747 8081
rect 10689 8041 10701 8075
rect 10735 8072 10747 8075
rect 12161 8075 12219 8081
rect 12161 8072 12173 8075
rect 10735 8044 12173 8072
rect 10735 8041 10747 8044
rect 10689 8035 10747 8041
rect 12161 8041 12173 8044
rect 12207 8041 12219 8075
rect 12161 8035 12219 8041
rect 12713 8075 12771 8081
rect 12713 8041 12725 8075
rect 12759 8072 12771 8075
rect 13814 8072 13820 8084
rect 12759 8044 13820 8072
rect 12759 8041 12771 8044
rect 12713 8035 12771 8041
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 2498 8004 2504 8016
rect 2459 7976 2504 8004
rect 2498 7964 2504 7976
rect 2556 7964 2562 8016
rect 3421 8007 3479 8013
rect 3421 7973 3433 8007
rect 3467 8004 3479 8007
rect 4338 8004 4344 8016
rect 3467 7976 4344 8004
rect 3467 7973 3479 7976
rect 3421 7967 3479 7973
rect 4338 7964 4344 7976
rect 4396 7964 4402 8016
rect 8478 8004 8484 8016
rect 4632 7976 8484 8004
rect 1486 7936 1492 7948
rect 1447 7908 1492 7936
rect 1486 7896 1492 7908
rect 1544 7896 1550 7948
rect 2225 7939 2283 7945
rect 2225 7905 2237 7939
rect 2271 7905 2283 7939
rect 2225 7899 2283 7905
rect 1670 7868 1676 7880
rect 1631 7840 1676 7868
rect 1670 7828 1676 7840
rect 1728 7828 1734 7880
rect 2240 7800 2268 7899
rect 3326 7896 3332 7948
rect 3384 7936 3390 7948
rect 3384 7908 3556 7936
rect 3384 7896 3390 7908
rect 3528 7877 3556 7908
rect 4154 7896 4160 7948
rect 4212 7936 4218 7948
rect 4632 7945 4660 7976
rect 8478 7964 8484 7976
rect 8536 7964 8542 8016
rect 9950 7964 9956 8016
rect 10008 8004 10014 8016
rect 10137 8007 10195 8013
rect 10137 8004 10149 8007
rect 10008 7976 10149 8004
rect 10008 7964 10014 7976
rect 10137 7973 10149 7976
rect 10183 7973 10195 8007
rect 10137 7967 10195 7973
rect 10778 7964 10784 8016
rect 10836 8004 10842 8016
rect 11149 8007 11207 8013
rect 11149 8004 11161 8007
rect 10836 7976 11161 8004
rect 10836 7964 10842 7976
rect 11149 7973 11161 7976
rect 11195 7973 11207 8007
rect 11149 7967 11207 7973
rect 12986 7964 12992 8016
rect 13044 8004 13050 8016
rect 13173 8007 13231 8013
rect 13173 8004 13185 8007
rect 13044 7976 13185 8004
rect 13044 7964 13050 7976
rect 13173 7973 13185 7976
rect 13219 7973 13231 8007
rect 13173 7967 13231 7973
rect 4617 7939 4675 7945
rect 4617 7936 4629 7939
rect 4212 7908 4629 7936
rect 4212 7896 4218 7908
rect 4617 7905 4629 7908
rect 4663 7905 4675 7939
rect 5436 7939 5494 7945
rect 5436 7936 5448 7939
rect 4617 7899 4675 7905
rect 5092 7908 5448 7936
rect 3513 7871 3571 7877
rect 3513 7837 3525 7871
rect 3559 7837 3571 7871
rect 3513 7831 3571 7837
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7868 4859 7871
rect 5092 7868 5120 7908
rect 5436 7905 5448 7908
rect 5482 7936 5494 7939
rect 6178 7936 6184 7948
rect 5482 7908 6184 7936
rect 5482 7905 5494 7908
rect 5436 7899 5494 7905
rect 6178 7896 6184 7908
rect 6236 7896 6242 7948
rect 7193 7939 7251 7945
rect 7193 7905 7205 7939
rect 7239 7936 7251 7939
rect 7558 7936 7564 7948
rect 7239 7908 7564 7936
rect 7239 7905 7251 7908
rect 7193 7899 7251 7905
rect 7558 7896 7564 7908
rect 7616 7936 7622 7948
rect 7742 7936 7748 7948
rect 7616 7908 7748 7936
rect 7616 7896 7622 7908
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 8846 7896 8852 7948
rect 8904 7936 8910 7948
rect 8941 7939 8999 7945
rect 8941 7936 8953 7939
rect 8904 7908 8953 7936
rect 8904 7896 8910 7908
rect 8941 7905 8953 7908
rect 8987 7905 8999 7939
rect 8941 7899 8999 7905
rect 9306 7896 9312 7948
rect 9364 7936 9370 7948
rect 11054 7936 11060 7948
rect 9364 7908 10272 7936
rect 11015 7908 11060 7936
rect 9364 7896 9370 7908
rect 4847 7840 5120 7868
rect 5169 7871 5227 7877
rect 4847 7837 4859 7840
rect 4801 7831 4859 7837
rect 5169 7837 5181 7871
rect 5215 7837 5227 7871
rect 7282 7868 7288 7880
rect 7243 7840 7288 7868
rect 5169 7831 5227 7837
rect 2240 7772 3832 7800
rect 3804 7732 3832 7772
rect 3878 7760 3884 7812
rect 3936 7800 3942 7812
rect 5184 7800 5212 7831
rect 7282 7828 7288 7840
rect 7340 7828 7346 7880
rect 7374 7828 7380 7880
rect 7432 7868 7438 7880
rect 9033 7871 9091 7877
rect 7432 7840 7477 7868
rect 7432 7828 7438 7840
rect 9033 7837 9045 7871
rect 9079 7837 9091 7871
rect 9033 7831 9091 7837
rect 3936 7772 5212 7800
rect 7300 7800 7328 7828
rect 7558 7800 7564 7812
rect 7300 7772 7564 7800
rect 3936 7760 3942 7772
rect 7558 7760 7564 7772
rect 7616 7760 7622 7812
rect 9048 7800 9076 7831
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 10244 7877 10272 7908
rect 11054 7896 11060 7908
rect 11112 7896 11118 7948
rect 11422 7896 11428 7948
rect 11480 7936 11486 7948
rect 11882 7936 11888 7948
rect 11480 7908 11888 7936
rect 11480 7896 11486 7908
rect 11882 7896 11888 7908
rect 11940 7896 11946 7948
rect 12066 7936 12072 7948
rect 12027 7908 12072 7936
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 12526 7896 12532 7948
rect 12584 7936 12590 7948
rect 12894 7936 12900 7948
rect 12584 7908 12900 7936
rect 12584 7896 12590 7908
rect 12894 7896 12900 7908
rect 12952 7936 12958 7948
rect 13081 7939 13139 7945
rect 13081 7936 13093 7939
rect 12952 7908 13093 7936
rect 12952 7896 12958 7908
rect 13081 7905 13093 7908
rect 13127 7905 13139 7939
rect 13081 7899 13139 7905
rect 10229 7871 10287 7877
rect 9180 7840 9225 7868
rect 9180 7828 9186 7840
rect 10229 7837 10241 7871
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 11241 7871 11299 7877
rect 11241 7868 11253 7871
rect 11204 7840 11253 7868
rect 11204 7828 11210 7840
rect 11241 7837 11253 7840
rect 11287 7837 11299 7871
rect 11241 7831 11299 7837
rect 11330 7828 11336 7880
rect 11388 7868 11394 7880
rect 12253 7871 12311 7877
rect 12253 7868 12265 7871
rect 11388 7840 12265 7868
rect 11388 7828 11394 7840
rect 12253 7837 12265 7840
rect 12299 7837 12311 7871
rect 13262 7868 13268 7880
rect 13223 7840 13268 7868
rect 12253 7831 12311 7837
rect 13262 7828 13268 7840
rect 13320 7828 13326 7880
rect 9048 7772 9904 7800
rect 9677 7735 9735 7741
rect 9677 7732 9689 7735
rect 3804 7704 9689 7732
rect 9677 7701 9689 7704
rect 9723 7701 9735 7735
rect 9876 7732 9904 7772
rect 9950 7760 9956 7812
rect 10008 7800 10014 7812
rect 10134 7800 10140 7812
rect 10008 7772 10140 7800
rect 10008 7760 10014 7772
rect 10134 7760 10140 7772
rect 10192 7760 10198 7812
rect 11698 7800 11704 7812
rect 11659 7772 11704 7800
rect 11698 7760 11704 7772
rect 11756 7760 11762 7812
rect 13170 7732 13176 7744
rect 9876 7704 13176 7732
rect 9677 7695 9735 7701
rect 13170 7692 13176 7704
rect 13228 7732 13234 7744
rect 15010 7732 15016 7744
rect 13228 7704 15016 7732
rect 13228 7692 13234 7704
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 1104 7642 15824 7664
rect 1104 7590 3447 7642
rect 3499 7590 3511 7642
rect 3563 7590 3575 7642
rect 3627 7590 3639 7642
rect 3691 7590 8378 7642
rect 8430 7590 8442 7642
rect 8494 7590 8506 7642
rect 8558 7590 8570 7642
rect 8622 7590 13308 7642
rect 13360 7590 13372 7642
rect 13424 7590 13436 7642
rect 13488 7590 13500 7642
rect 13552 7590 15824 7642
rect 1104 7568 15824 7590
rect 4525 7531 4583 7537
rect 4525 7528 4537 7531
rect 2792 7500 4537 7528
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 2685 7395 2743 7401
rect 2685 7392 2697 7395
rect 2547 7364 2697 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 2685 7361 2697 7364
rect 2731 7361 2743 7395
rect 2685 7355 2743 7361
rect 2225 7327 2283 7333
rect 2225 7293 2237 7327
rect 2271 7324 2283 7327
rect 2792 7324 2820 7500
rect 4525 7497 4537 7500
rect 4571 7497 4583 7531
rect 5534 7528 5540 7540
rect 5495 7500 5540 7528
rect 4525 7491 4583 7497
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 6822 7528 6828 7540
rect 6783 7500 6828 7528
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 9030 7528 9036 7540
rect 7484 7500 9036 7528
rect 4249 7463 4307 7469
rect 4249 7429 4261 7463
rect 4295 7460 4307 7463
rect 4295 7432 6224 7460
rect 4295 7429 4307 7432
rect 4249 7423 4307 7429
rect 6196 7404 6224 7432
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 5077 7395 5135 7401
rect 5077 7392 5089 7395
rect 4212 7364 5089 7392
rect 4212 7352 4218 7364
rect 5077 7361 5089 7364
rect 5123 7361 5135 7395
rect 6178 7392 6184 7404
rect 6091 7364 6184 7392
rect 5077 7355 5135 7361
rect 6178 7352 6184 7364
rect 6236 7392 6242 7404
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 6236 7364 7389 7392
rect 6236 7352 6242 7364
rect 7377 7361 7389 7364
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 2271 7296 2820 7324
rect 2271 7293 2283 7296
rect 2225 7287 2283 7293
rect 2866 7284 2872 7336
rect 2924 7324 2930 7336
rect 5997 7327 6055 7333
rect 2924 7296 2969 7324
rect 2924 7284 2930 7296
rect 5997 7293 6009 7327
rect 6043 7324 6055 7327
rect 7484 7324 7512 7500
rect 9030 7488 9036 7500
rect 9088 7488 9094 7540
rect 10045 7531 10103 7537
rect 10045 7497 10057 7531
rect 10091 7528 10103 7531
rect 10778 7528 10784 7540
rect 10091 7500 10784 7528
rect 10091 7497 10103 7500
rect 10045 7491 10103 7497
rect 10778 7488 10784 7500
rect 10836 7488 10842 7540
rect 11054 7528 11060 7540
rect 11015 7500 11060 7528
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 9677 7463 9735 7469
rect 9677 7429 9689 7463
rect 9723 7460 9735 7463
rect 10226 7460 10232 7472
rect 9723 7432 10232 7460
rect 9723 7429 9735 7432
rect 9677 7423 9735 7429
rect 10226 7420 10232 7432
rect 10284 7420 10290 7472
rect 10597 7395 10655 7401
rect 10597 7361 10609 7395
rect 10643 7392 10655 7395
rect 11606 7392 11612 7404
rect 10643 7364 11612 7392
rect 10643 7361 10655 7364
rect 10597 7355 10655 7361
rect 11606 7352 11612 7364
rect 11664 7392 11670 7404
rect 11701 7395 11759 7401
rect 11701 7392 11713 7395
rect 11664 7364 11713 7392
rect 11664 7352 11670 7364
rect 11701 7361 11713 7364
rect 11747 7392 11759 7395
rect 13081 7395 13139 7401
rect 13081 7392 13093 7395
rect 11747 7364 13093 7392
rect 11747 7361 11759 7364
rect 11701 7355 11759 7361
rect 13081 7361 13093 7364
rect 13127 7392 13139 7395
rect 13446 7392 13452 7404
rect 13127 7364 13452 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 13446 7352 13452 7364
rect 13504 7352 13510 7404
rect 8018 7324 8024 7336
rect 6043 7296 7512 7324
rect 7979 7296 8024 7324
rect 6043 7293 6055 7296
rect 5997 7287 6055 7293
rect 8018 7284 8024 7296
rect 8076 7284 8082 7336
rect 8294 7324 8300 7336
rect 8207 7296 8300 7324
rect 8294 7284 8300 7296
rect 8352 7324 8358 7336
rect 10134 7324 10140 7336
rect 8352 7296 10140 7324
rect 8352 7284 8358 7296
rect 10134 7284 10140 7296
rect 10192 7284 10198 7336
rect 10318 7284 10324 7336
rect 10376 7324 10382 7336
rect 10505 7327 10563 7333
rect 10505 7324 10517 7327
rect 10376 7296 10517 7324
rect 10376 7284 10382 7296
rect 10505 7293 10517 7296
rect 10551 7293 10563 7327
rect 10505 7287 10563 7293
rect 11425 7327 11483 7333
rect 11425 7293 11437 7327
rect 11471 7324 11483 7327
rect 11514 7324 11520 7336
rect 11471 7296 11520 7324
rect 11471 7293 11483 7296
rect 11425 7287 11483 7293
rect 11514 7284 11520 7296
rect 11572 7324 11578 7336
rect 11882 7324 11888 7336
rect 11572 7296 11888 7324
rect 11572 7284 11578 7296
rect 11882 7284 11888 7296
rect 11940 7284 11946 7336
rect 12710 7284 12716 7336
rect 12768 7324 12774 7336
rect 12897 7327 12955 7333
rect 12897 7324 12909 7327
rect 12768 7296 12909 7324
rect 12768 7284 12774 7296
rect 12897 7293 12909 7296
rect 12943 7293 12955 7327
rect 12897 7287 12955 7293
rect 2685 7259 2743 7265
rect 2685 7225 2697 7259
rect 2731 7256 2743 7259
rect 3050 7256 3056 7268
rect 2731 7228 3056 7256
rect 2731 7225 2743 7228
rect 2685 7219 2743 7225
rect 3050 7216 3056 7228
rect 3108 7265 3114 7268
rect 3108 7259 3172 7265
rect 3108 7225 3126 7259
rect 3160 7225 3172 7259
rect 4890 7256 4896 7268
rect 4851 7228 4896 7256
rect 3108 7219 3172 7225
rect 3108 7216 3114 7219
rect 4890 7216 4896 7228
rect 4948 7216 4954 7268
rect 7285 7259 7343 7265
rect 7285 7225 7297 7259
rect 7331 7256 7343 7259
rect 8564 7259 8622 7265
rect 7331 7228 8524 7256
rect 7331 7225 7343 7228
rect 7285 7219 7343 7225
rect 1394 7148 1400 7200
rect 1452 7188 1458 7200
rect 1857 7191 1915 7197
rect 1857 7188 1869 7191
rect 1452 7160 1869 7188
rect 1452 7148 1458 7160
rect 1857 7157 1869 7160
rect 1903 7157 1915 7191
rect 1857 7151 1915 7157
rect 2317 7191 2375 7197
rect 2317 7157 2329 7191
rect 2363 7188 2375 7191
rect 2866 7188 2872 7200
rect 2363 7160 2872 7188
rect 2363 7157 2375 7160
rect 2317 7151 2375 7157
rect 2866 7148 2872 7160
rect 2924 7148 2930 7200
rect 4982 7188 4988 7200
rect 4943 7160 4988 7188
rect 4982 7148 4988 7160
rect 5040 7148 5046 7200
rect 5905 7191 5963 7197
rect 5905 7157 5917 7191
rect 5951 7188 5963 7191
rect 6270 7188 6276 7200
rect 5951 7160 6276 7188
rect 5951 7157 5963 7160
rect 5905 7151 5963 7157
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 7190 7188 7196 7200
rect 7151 7160 7196 7188
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 7650 7148 7656 7200
rect 7708 7188 7714 7200
rect 7837 7191 7895 7197
rect 7837 7188 7849 7191
rect 7708 7160 7849 7188
rect 7708 7148 7714 7160
rect 7837 7157 7849 7160
rect 7883 7157 7895 7191
rect 8496 7188 8524 7228
rect 8564 7225 8576 7259
rect 8610 7256 8622 7259
rect 9306 7256 9312 7268
rect 8610 7228 9312 7256
rect 8610 7225 8622 7228
rect 8564 7219 8622 7225
rect 9306 7216 9312 7228
rect 9364 7216 9370 7268
rect 9398 7216 9404 7268
rect 9456 7256 9462 7268
rect 11698 7256 11704 7268
rect 9456 7228 11704 7256
rect 9456 7216 9462 7228
rect 11698 7216 11704 7228
rect 11756 7216 11762 7268
rect 12912 7256 12940 7287
rect 13078 7256 13084 7268
rect 12912 7228 13084 7256
rect 13078 7216 13084 7228
rect 13136 7216 13142 7268
rect 9214 7188 9220 7200
rect 8496 7160 9220 7188
rect 7837 7151 7895 7157
rect 9214 7148 9220 7160
rect 9272 7188 9278 7200
rect 9674 7188 9680 7200
rect 9272 7160 9680 7188
rect 9272 7148 9278 7160
rect 9674 7148 9680 7160
rect 9732 7188 9738 7200
rect 10413 7191 10471 7197
rect 10413 7188 10425 7191
rect 9732 7160 10425 7188
rect 9732 7148 9738 7160
rect 10413 7157 10425 7160
rect 10459 7157 10471 7191
rect 10413 7151 10471 7157
rect 10594 7148 10600 7200
rect 10652 7188 10658 7200
rect 11517 7191 11575 7197
rect 11517 7188 11529 7191
rect 10652 7160 11529 7188
rect 10652 7148 10658 7160
rect 11517 7157 11529 7160
rect 11563 7157 11575 7191
rect 11517 7151 11575 7157
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 12492 7160 12537 7188
rect 12492 7148 12498 7160
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 12805 7191 12863 7197
rect 12805 7188 12817 7191
rect 12676 7160 12817 7188
rect 12676 7148 12682 7160
rect 12805 7157 12817 7160
rect 12851 7188 12863 7191
rect 16298 7188 16304 7200
rect 12851 7160 16304 7188
rect 12851 7157 12863 7160
rect 12805 7151 12863 7157
rect 16298 7148 16304 7160
rect 16356 7148 16362 7200
rect 1104 7098 15824 7120
rect 1104 7046 5912 7098
rect 5964 7046 5976 7098
rect 6028 7046 6040 7098
rect 6092 7046 6104 7098
rect 6156 7046 10843 7098
rect 10895 7046 10907 7098
rect 10959 7046 10971 7098
rect 11023 7046 11035 7098
rect 11087 7046 15824 7098
rect 1104 7024 15824 7046
rect 3050 6984 3056 6996
rect 3011 6956 3056 6984
rect 3050 6944 3056 6956
rect 3108 6944 3114 6996
rect 4801 6987 4859 6993
rect 4801 6953 4813 6987
rect 4847 6984 4859 6987
rect 4890 6984 4896 6996
rect 4847 6956 4896 6984
rect 4847 6953 4859 6956
rect 4801 6947 4859 6953
rect 4890 6944 4896 6956
rect 4948 6944 4954 6996
rect 6270 6944 6276 6996
rect 6328 6984 6334 6996
rect 9125 6987 9183 6993
rect 6328 6956 8800 6984
rect 6328 6944 6334 6956
rect 5169 6919 5227 6925
rect 5169 6885 5181 6919
rect 5215 6916 5227 6919
rect 6822 6916 6828 6928
rect 5215 6888 6828 6916
rect 5215 6885 5227 6888
rect 5169 6879 5227 6885
rect 6822 6876 6828 6888
rect 6880 6876 6886 6928
rect 8294 6916 8300 6928
rect 7944 6888 8300 6916
rect 1940 6851 1998 6857
rect 1940 6817 1952 6851
rect 1986 6848 1998 6851
rect 4154 6848 4160 6860
rect 1986 6820 4160 6848
rect 1986 6817 1998 6820
rect 1940 6811 1998 6817
rect 4154 6808 4160 6820
rect 4212 6808 4218 6860
rect 4709 6851 4767 6857
rect 4709 6817 4721 6851
rect 4755 6817 4767 6851
rect 5258 6848 5264 6860
rect 5219 6820 5264 6848
rect 4709 6811 4767 6817
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6749 1731 6783
rect 1673 6743 1731 6749
rect 1688 6644 1716 6743
rect 4724 6712 4752 6811
rect 5258 6808 5264 6820
rect 5316 6848 5322 6860
rect 5997 6851 6055 6857
rect 5316 6820 5948 6848
rect 5316 6808 5322 6820
rect 5350 6740 5356 6792
rect 5408 6780 5414 6792
rect 5920 6780 5948 6820
rect 5997 6817 6009 6851
rect 6043 6848 6055 6851
rect 6914 6848 6920 6860
rect 6043 6820 6920 6848
rect 6043 6817 6055 6820
rect 5997 6811 6055 6817
rect 6914 6808 6920 6820
rect 6972 6808 6978 6860
rect 7098 6848 7104 6860
rect 7059 6820 7104 6848
rect 7098 6808 7104 6820
rect 7156 6808 7162 6860
rect 7745 6851 7803 6857
rect 7745 6817 7757 6851
rect 7791 6848 7803 6851
rect 7944 6848 7972 6888
rect 8294 6876 8300 6888
rect 8352 6876 8358 6928
rect 8662 6876 8668 6928
rect 8720 6876 8726 6928
rect 8772 6916 8800 6956
rect 9125 6953 9137 6987
rect 9171 6984 9183 6987
rect 9306 6984 9312 6996
rect 9171 6956 9312 6984
rect 9171 6953 9183 6956
rect 9125 6947 9183 6953
rect 9306 6944 9312 6956
rect 9364 6944 9370 6996
rect 9677 6987 9735 6993
rect 9677 6953 9689 6987
rect 9723 6984 9735 6987
rect 10318 6984 10324 6996
rect 9723 6956 10324 6984
rect 9723 6953 9735 6956
rect 9677 6947 9735 6953
rect 10318 6944 10324 6956
rect 10376 6944 10382 6996
rect 11238 6944 11244 6996
rect 11296 6984 11302 6996
rect 12621 6987 12679 6993
rect 12621 6984 12633 6987
rect 11296 6956 12633 6984
rect 11296 6944 11302 6956
rect 12621 6953 12633 6956
rect 12667 6953 12679 6987
rect 12621 6947 12679 6953
rect 10042 6916 10048 6928
rect 8772 6888 10048 6916
rect 10042 6876 10048 6888
rect 10100 6876 10106 6928
rect 11508 6919 11566 6925
rect 11508 6885 11520 6919
rect 11554 6916 11566 6919
rect 11606 6916 11612 6928
rect 11554 6888 11612 6916
rect 11554 6885 11566 6888
rect 11508 6879 11566 6885
rect 11606 6876 11612 6888
rect 11664 6876 11670 6928
rect 11698 6876 11704 6928
rect 11756 6916 11762 6928
rect 12986 6916 12992 6928
rect 11756 6888 12992 6916
rect 11756 6876 11762 6888
rect 12986 6876 12992 6888
rect 13044 6876 13050 6928
rect 7791 6820 7972 6848
rect 8012 6851 8070 6857
rect 7791 6817 7803 6820
rect 7745 6811 7803 6817
rect 8012 6817 8024 6851
rect 8058 6848 8070 6851
rect 8680 6848 8708 6876
rect 8058 6820 8708 6848
rect 8058 6817 8070 6820
rect 8012 6811 8070 6817
rect 9030 6808 9036 6860
rect 9088 6848 9094 6860
rect 10137 6851 10195 6857
rect 10137 6848 10149 6851
rect 9088 6820 10149 6848
rect 9088 6808 9094 6820
rect 10137 6817 10149 6820
rect 10183 6848 10195 6851
rect 10318 6848 10324 6860
rect 10183 6820 10324 6848
rect 10183 6817 10195 6820
rect 10137 6811 10195 6817
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 10505 6851 10563 6857
rect 10505 6817 10517 6851
rect 10551 6848 10563 6851
rect 10873 6851 10931 6857
rect 10873 6848 10885 6851
rect 10551 6820 10885 6848
rect 10551 6817 10563 6820
rect 10505 6811 10563 6817
rect 10873 6817 10885 6820
rect 10919 6817 10931 6851
rect 10873 6811 10931 6817
rect 11241 6851 11299 6857
rect 11241 6817 11253 6851
rect 11287 6848 11299 6851
rect 11330 6848 11336 6860
rect 11287 6820 11336 6848
rect 11287 6817 11299 6820
rect 11241 6811 11299 6817
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 12526 6808 12532 6860
rect 12584 6848 12590 6860
rect 13265 6851 13323 6857
rect 13265 6848 13277 6851
rect 12584 6820 13277 6848
rect 12584 6808 12590 6820
rect 13265 6817 13277 6820
rect 13311 6817 13323 6851
rect 13265 6811 13323 6817
rect 13357 6851 13415 6857
rect 13357 6817 13369 6851
rect 13403 6848 13415 6851
rect 13630 6848 13636 6860
rect 13403 6820 13636 6848
rect 13403 6817 13415 6820
rect 13357 6811 13415 6817
rect 13630 6808 13636 6820
rect 13688 6848 13694 6860
rect 14366 6848 14372 6860
rect 13688 6820 14372 6848
rect 13688 6808 13694 6820
rect 14366 6808 14372 6820
rect 14424 6808 14430 6860
rect 7190 6780 7196 6792
rect 5408 6752 5453 6780
rect 5920 6752 7196 6780
rect 5408 6740 5414 6752
rect 7190 6740 7196 6752
rect 7248 6740 7254 6792
rect 7374 6780 7380 6792
rect 7335 6752 7380 6780
rect 7374 6740 7380 6752
rect 7432 6740 7438 6792
rect 10226 6740 10232 6792
rect 10284 6780 10290 6792
rect 13446 6780 13452 6792
rect 10284 6752 10329 6780
rect 13407 6752 13452 6780
rect 10284 6740 10290 6752
rect 13446 6740 13452 6752
rect 13504 6740 13510 6792
rect 7650 6712 7656 6724
rect 4724 6684 7656 6712
rect 7650 6672 7656 6684
rect 7708 6672 7714 6724
rect 9490 6672 9496 6724
rect 9548 6712 9554 6724
rect 10594 6712 10600 6724
rect 9548 6684 10600 6712
rect 9548 6672 9554 6684
rect 10594 6672 10600 6684
rect 10652 6672 10658 6724
rect 2774 6644 2780 6656
rect 1688 6616 2780 6644
rect 2774 6604 2780 6616
rect 2832 6604 2838 6656
rect 4522 6644 4528 6656
rect 4435 6616 4528 6644
rect 4522 6604 4528 6616
rect 4580 6644 4586 6656
rect 4706 6644 4712 6656
rect 4580 6616 4712 6644
rect 4580 6604 4586 6616
rect 4706 6604 4712 6616
rect 4764 6604 4770 6656
rect 5626 6604 5632 6656
rect 5684 6644 5690 6656
rect 6181 6647 6239 6653
rect 6181 6644 6193 6647
rect 5684 6616 6193 6644
rect 5684 6604 5690 6616
rect 6181 6613 6193 6616
rect 6227 6613 6239 6647
rect 6730 6644 6736 6656
rect 6691 6616 6736 6644
rect 6181 6607 6239 6613
rect 6730 6604 6736 6616
rect 6788 6604 6794 6656
rect 7668 6644 7696 6672
rect 10505 6647 10563 6653
rect 10505 6644 10517 6647
rect 7668 6616 10517 6644
rect 10505 6613 10517 6616
rect 10551 6613 10563 6647
rect 10686 6644 10692 6656
rect 10647 6616 10692 6644
rect 10505 6607 10563 6613
rect 10686 6604 10692 6616
rect 10744 6604 10750 6656
rect 12894 6644 12900 6656
rect 12855 6616 12900 6644
rect 12894 6604 12900 6616
rect 12952 6604 12958 6656
rect 1104 6554 15824 6576
rect 1104 6502 3447 6554
rect 3499 6502 3511 6554
rect 3563 6502 3575 6554
rect 3627 6502 3639 6554
rect 3691 6502 8378 6554
rect 8430 6502 8442 6554
rect 8494 6502 8506 6554
rect 8558 6502 8570 6554
rect 8622 6502 13308 6554
rect 13360 6502 13372 6554
rect 13424 6502 13436 6554
rect 13488 6502 13500 6554
rect 13552 6502 15824 6554
rect 1104 6480 15824 6502
rect 3053 6443 3111 6449
rect 3053 6409 3065 6443
rect 3099 6440 3111 6443
rect 4154 6440 4160 6452
rect 3099 6412 4160 6440
rect 3099 6409 3111 6412
rect 3053 6403 3111 6409
rect 4154 6400 4160 6412
rect 4212 6400 4218 6452
rect 4525 6443 4583 6449
rect 4525 6409 4537 6443
rect 4571 6440 4583 6443
rect 4982 6440 4988 6452
rect 4571 6412 4988 6440
rect 4571 6409 4583 6412
rect 4525 6403 4583 6409
rect 4982 6400 4988 6412
rect 5040 6400 5046 6452
rect 8481 6443 8539 6449
rect 8481 6440 8493 6443
rect 6104 6412 8493 6440
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6304 3939 6307
rect 5077 6307 5135 6313
rect 5077 6304 5089 6307
rect 3927 6276 5089 6304
rect 3927 6273 3939 6276
rect 3881 6267 3939 6273
rect 5077 6273 5089 6276
rect 5123 6304 5135 6307
rect 5350 6304 5356 6316
rect 5123 6276 5356 6304
rect 5123 6273 5135 6276
rect 5077 6267 5135 6273
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 1762 6236 1768 6248
rect 1719 6208 1768 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 1762 6196 1768 6208
rect 1820 6196 1826 6248
rect 3896 6236 3924 6267
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 6104 6304 6132 6412
rect 8481 6409 8493 6412
rect 8527 6409 8539 6443
rect 10134 6440 10140 6452
rect 8481 6403 8539 6409
rect 9508 6412 10140 6440
rect 8205 6375 8263 6381
rect 8205 6341 8217 6375
rect 8251 6341 8263 6375
rect 8205 6335 8263 6341
rect 6181 6307 6239 6313
rect 6181 6304 6193 6307
rect 6104 6276 6193 6304
rect 6181 6273 6193 6276
rect 6227 6273 6239 6307
rect 6362 6304 6368 6316
rect 6275 6276 6368 6304
rect 6181 6267 6239 6273
rect 6362 6264 6368 6276
rect 6420 6304 6426 6316
rect 6420 6276 6960 6304
rect 6420 6264 6426 6276
rect 2424 6208 3924 6236
rect 2424 6180 2452 6208
rect 4062 6196 4068 6248
rect 4120 6196 4126 6248
rect 6089 6239 6147 6245
rect 6089 6205 6101 6239
rect 6135 6236 6147 6239
rect 6730 6236 6736 6248
rect 6135 6208 6736 6236
rect 6135 6205 6147 6208
rect 6089 6199 6147 6205
rect 6730 6196 6736 6208
rect 6788 6196 6794 6248
rect 6825 6239 6883 6245
rect 6825 6205 6837 6239
rect 6871 6205 6883 6239
rect 6932 6236 6960 6276
rect 8220 6236 8248 6335
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6304 9183 6307
rect 9214 6304 9220 6316
rect 9171 6276 9220 6304
rect 9171 6273 9183 6276
rect 9125 6267 9183 6273
rect 9214 6264 9220 6276
rect 9272 6264 9278 6316
rect 9508 6313 9536 6412
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 11333 6443 11391 6449
rect 11333 6409 11345 6443
rect 11379 6440 11391 6443
rect 12066 6440 12072 6452
rect 11379 6412 12072 6440
rect 11379 6409 11391 6412
rect 11333 6403 11391 6409
rect 12066 6400 12072 6412
rect 12124 6400 12130 6452
rect 12434 6400 12440 6452
rect 12492 6400 12498 6452
rect 10873 6375 10931 6381
rect 10873 6341 10885 6375
rect 10919 6372 10931 6375
rect 11606 6372 11612 6384
rect 10919 6344 11612 6372
rect 10919 6341 10931 6344
rect 10873 6335 10931 6341
rect 11606 6332 11612 6344
rect 11664 6332 11670 6384
rect 12452 6372 12480 6400
rect 12452 6344 12664 6372
rect 9493 6307 9551 6313
rect 9493 6273 9505 6307
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 11238 6264 11244 6316
rect 11296 6304 11302 6316
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 11296 6276 11897 6304
rect 11296 6264 11302 6276
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 11885 6267 11943 6273
rect 12437 6307 12495 6313
rect 12437 6273 12449 6307
rect 12483 6304 12495 6307
rect 12526 6304 12532 6316
rect 12483 6276 12532 6304
rect 12483 6273 12495 6276
rect 12437 6267 12495 6273
rect 12526 6264 12532 6276
rect 12584 6264 12590 6316
rect 6932 6208 8248 6236
rect 6825 6199 6883 6205
rect 1940 6171 1998 6177
rect 1940 6137 1952 6171
rect 1986 6168 1998 6171
rect 2406 6168 2412 6180
rect 1986 6140 2412 6168
rect 1986 6137 1998 6140
rect 1940 6131 1998 6137
rect 2406 6128 2412 6140
rect 2464 6128 2470 6180
rect 3697 6171 3755 6177
rect 3697 6137 3709 6171
rect 3743 6168 3755 6171
rect 4080 6168 4108 6196
rect 3743 6140 4108 6168
rect 4985 6171 5043 6177
rect 3743 6137 3755 6140
rect 3697 6131 3755 6137
rect 4985 6137 4997 6171
rect 5031 6168 5043 6171
rect 6178 6168 6184 6180
rect 5031 6140 6184 6168
rect 5031 6137 5043 6140
rect 4985 6131 5043 6137
rect 6178 6128 6184 6140
rect 6236 6128 6242 6180
rect 6270 6128 6276 6180
rect 6328 6168 6334 6180
rect 6840 6168 6868 6199
rect 8386 6196 8392 6248
rect 8444 6236 8450 6248
rect 9760 6239 9818 6245
rect 8444 6208 9076 6236
rect 8444 6196 8450 6208
rect 6328 6140 6868 6168
rect 7092 6171 7150 6177
rect 6328 6128 6334 6140
rect 7092 6137 7104 6171
rect 7138 6168 7150 6171
rect 7374 6168 7380 6180
rect 7138 6140 7380 6168
rect 7138 6137 7150 6140
rect 7092 6131 7150 6137
rect 7374 6128 7380 6140
rect 7432 6168 7438 6180
rect 8294 6168 8300 6180
rect 7432 6140 8300 6168
rect 7432 6128 7438 6140
rect 8294 6128 8300 6140
rect 8352 6128 8358 6180
rect 8941 6171 8999 6177
rect 8941 6168 8953 6171
rect 8404 6140 8953 6168
rect 3326 6100 3332 6112
rect 3287 6072 3332 6100
rect 3326 6060 3332 6072
rect 3384 6060 3390 6112
rect 3789 6103 3847 6109
rect 3789 6069 3801 6103
rect 3835 6100 3847 6103
rect 4062 6100 4068 6112
rect 3835 6072 4068 6100
rect 3835 6069 3847 6072
rect 3789 6063 3847 6069
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 4890 6100 4896 6112
rect 4851 6072 4896 6100
rect 4890 6060 4896 6072
rect 4948 6060 4954 6112
rect 5721 6103 5779 6109
rect 5721 6069 5733 6103
rect 5767 6100 5779 6103
rect 5810 6100 5816 6112
rect 5767 6072 5816 6100
rect 5767 6069 5779 6072
rect 5721 6063 5779 6069
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 6546 6060 6552 6112
rect 6604 6100 6610 6112
rect 8404 6100 8432 6140
rect 8941 6137 8953 6140
rect 8987 6137 8999 6171
rect 9048 6168 9076 6208
rect 9760 6205 9772 6239
rect 9806 6236 9818 6239
rect 10226 6236 10232 6248
rect 9806 6208 10232 6236
rect 9806 6205 9818 6208
rect 9760 6199 9818 6205
rect 10226 6196 10232 6208
rect 10284 6196 10290 6248
rect 11793 6239 11851 6245
rect 11793 6205 11805 6239
rect 11839 6236 11851 6239
rect 12636 6236 12664 6344
rect 13906 6264 13912 6316
rect 13964 6304 13970 6316
rect 14734 6304 14740 6316
rect 13964 6276 14740 6304
rect 13964 6264 13970 6276
rect 14734 6264 14740 6276
rect 14792 6264 14798 6316
rect 11839 6208 12664 6236
rect 11839 6205 11851 6208
rect 11793 6199 11851 6205
rect 11422 6168 11428 6180
rect 9048 6140 11428 6168
rect 8941 6131 8999 6137
rect 11422 6128 11428 6140
rect 11480 6128 11486 6180
rect 11701 6171 11759 6177
rect 11701 6137 11713 6171
rect 11747 6168 11759 6171
rect 12894 6168 12900 6180
rect 11747 6140 12900 6168
rect 11747 6137 11759 6140
rect 11701 6131 11759 6137
rect 12894 6128 12900 6140
rect 12952 6128 12958 6180
rect 6604 6072 8432 6100
rect 6604 6060 6610 6072
rect 8478 6060 8484 6112
rect 8536 6100 8542 6112
rect 8849 6103 8907 6109
rect 8849 6100 8861 6103
rect 8536 6072 8861 6100
rect 8536 6060 8542 6072
rect 8849 6069 8861 6072
rect 8895 6100 8907 6103
rect 9490 6100 9496 6112
rect 8895 6072 9496 6100
rect 8895 6069 8907 6072
rect 8849 6063 8907 6069
rect 9490 6060 9496 6072
rect 9548 6060 9554 6112
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 10226 6100 10232 6112
rect 9732 6072 10232 6100
rect 9732 6060 9738 6072
rect 10226 6060 10232 6072
rect 10284 6060 10290 6112
rect 1104 6010 15824 6032
rect 1104 5958 5912 6010
rect 5964 5958 5976 6010
rect 6028 5958 6040 6010
rect 6092 5958 6104 6010
rect 6156 5958 10843 6010
rect 10895 5958 10907 6010
rect 10959 5958 10971 6010
rect 11023 5958 11035 6010
rect 11087 5958 15824 6010
rect 1104 5936 15824 5958
rect 4062 5896 4068 5908
rect 4023 5868 4068 5896
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 4338 5856 4344 5908
rect 4396 5896 4402 5908
rect 4433 5899 4491 5905
rect 4433 5896 4445 5899
rect 4396 5868 4445 5896
rect 4396 5856 4402 5868
rect 4433 5865 4445 5868
rect 4479 5865 4491 5899
rect 4433 5859 4491 5865
rect 4525 5899 4583 5905
rect 4525 5865 4537 5899
rect 4571 5896 4583 5899
rect 4798 5896 4804 5908
rect 4571 5868 4804 5896
rect 4571 5865 4583 5868
rect 4525 5859 4583 5865
rect 4798 5856 4804 5868
rect 4856 5856 4862 5908
rect 4890 5856 4896 5908
rect 4948 5896 4954 5908
rect 6917 5899 6975 5905
rect 4948 5868 6500 5896
rect 4948 5856 4954 5868
rect 1670 5828 1676 5840
rect 1631 5800 1676 5828
rect 1670 5788 1676 5800
rect 1728 5788 1734 5840
rect 1762 5788 1768 5840
rect 1820 5828 1826 5840
rect 2501 5831 2559 5837
rect 2501 5828 2513 5831
rect 1820 5800 2513 5828
rect 1820 5788 1826 5800
rect 2501 5797 2513 5800
rect 2547 5828 2559 5831
rect 3234 5828 3240 5840
rect 2547 5800 3240 5828
rect 2547 5797 2559 5800
rect 2501 5791 2559 5797
rect 3234 5788 3240 5800
rect 3292 5788 3298 5840
rect 4614 5828 4620 5840
rect 3436 5800 4620 5828
rect 1394 5760 1400 5772
rect 1355 5732 1400 5760
rect 1394 5720 1400 5732
rect 1452 5720 1458 5772
rect 3436 5769 3464 5800
rect 4614 5788 4620 5800
rect 4672 5788 4678 5840
rect 5528 5831 5586 5837
rect 5528 5797 5540 5831
rect 5574 5828 5586 5831
rect 6362 5828 6368 5840
rect 5574 5800 6368 5828
rect 5574 5797 5586 5800
rect 5528 5791 5586 5797
rect 6362 5788 6368 5800
rect 6420 5788 6426 5840
rect 6472 5828 6500 5868
rect 6917 5865 6929 5899
rect 6963 5896 6975 5899
rect 7098 5896 7104 5908
rect 6963 5868 7104 5896
rect 6963 5865 6975 5868
rect 6917 5859 6975 5865
rect 7098 5856 7104 5868
rect 7156 5856 7162 5908
rect 7190 5856 7196 5908
rect 7248 5896 7254 5908
rect 9398 5896 9404 5908
rect 7248 5868 9404 5896
rect 7248 5856 7254 5868
rect 9398 5856 9404 5868
rect 9456 5856 9462 5908
rect 9490 5856 9496 5908
rect 9548 5896 9554 5908
rect 14274 5896 14280 5908
rect 9548 5868 14280 5896
rect 9548 5856 9554 5868
rect 14274 5856 14280 5868
rect 14332 5856 14338 5908
rect 8478 5828 8484 5840
rect 6472 5800 8484 5828
rect 8478 5788 8484 5800
rect 8536 5788 8542 5840
rect 13906 5828 13912 5840
rect 8956 5800 13912 5828
rect 3421 5763 3479 5769
rect 3421 5729 3433 5763
rect 3467 5729 3479 5763
rect 3421 5723 3479 5729
rect 5261 5763 5319 5769
rect 5261 5729 5273 5763
rect 5307 5760 5319 5763
rect 6270 5760 6276 5772
rect 5307 5732 6276 5760
rect 5307 5729 5319 5732
rect 5261 5723 5319 5729
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 7466 5720 7472 5772
rect 7524 5760 7530 5772
rect 7745 5763 7803 5769
rect 7745 5760 7757 5763
rect 7524 5732 7757 5760
rect 7524 5720 7530 5732
rect 7745 5729 7757 5732
rect 7791 5729 7803 5763
rect 7745 5723 7803 5729
rect 2590 5692 2596 5704
rect 2551 5664 2596 5692
rect 2590 5652 2596 5664
rect 2648 5652 2654 5704
rect 2682 5652 2688 5704
rect 2740 5692 2746 5704
rect 2740 5664 2785 5692
rect 2740 5652 2746 5664
rect 4614 5652 4620 5704
rect 4672 5692 4678 5704
rect 7558 5692 7564 5704
rect 4672 5664 4717 5692
rect 6288 5664 7564 5692
rect 4672 5652 4678 5664
rect 2133 5559 2191 5565
rect 2133 5525 2145 5559
rect 2179 5556 2191 5559
rect 2222 5556 2228 5568
rect 2179 5528 2228 5556
rect 2179 5525 2191 5528
rect 2133 5519 2191 5525
rect 2222 5516 2228 5528
rect 2280 5516 2286 5568
rect 3605 5559 3663 5565
rect 3605 5525 3617 5559
rect 3651 5556 3663 5559
rect 3878 5556 3884 5568
rect 3651 5528 3884 5556
rect 3651 5525 3663 5528
rect 3605 5519 3663 5525
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 4338 5516 4344 5568
rect 4396 5556 4402 5568
rect 6288 5556 6316 5664
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 7760 5692 7788 5723
rect 7834 5720 7840 5772
rect 7892 5760 7898 5772
rect 8389 5763 8447 5769
rect 7892 5732 7937 5760
rect 7892 5720 7898 5732
rect 8389 5729 8401 5763
rect 8435 5760 8447 5763
rect 8846 5760 8852 5772
rect 8435 5732 8852 5760
rect 8435 5729 8447 5732
rect 8389 5723 8447 5729
rect 8846 5720 8852 5732
rect 8904 5720 8910 5772
rect 8956 5769 8984 5800
rect 13906 5788 13912 5800
rect 13964 5788 13970 5840
rect 14734 5828 14740 5840
rect 14695 5800 14740 5828
rect 14734 5788 14740 5800
rect 14792 5788 14798 5840
rect 8941 5763 8999 5769
rect 8941 5729 8953 5763
rect 8987 5729 8999 5763
rect 9950 5760 9956 5772
rect 8941 5723 8999 5729
rect 9324 5732 9956 5760
rect 7926 5692 7932 5704
rect 7760 5664 7932 5692
rect 7926 5652 7932 5664
rect 7984 5652 7990 5704
rect 8021 5695 8079 5701
rect 8021 5661 8033 5695
rect 8067 5692 8079 5695
rect 8294 5692 8300 5704
rect 8067 5664 8300 5692
rect 8067 5661 8079 5664
rect 8021 5655 8079 5661
rect 8294 5652 8300 5664
rect 8352 5692 8358 5704
rect 9214 5692 9220 5704
rect 8352 5664 9220 5692
rect 8352 5652 8358 5664
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 7006 5584 7012 5636
rect 7064 5624 7070 5636
rect 8573 5627 8631 5633
rect 8573 5624 8585 5627
rect 7064 5596 8585 5624
rect 7064 5584 7070 5596
rect 8573 5593 8585 5596
rect 8619 5593 8631 5627
rect 9324 5624 9352 5732
rect 9950 5720 9956 5732
rect 10008 5720 10014 5772
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5760 10379 5763
rect 10778 5760 10784 5772
rect 10367 5732 10784 5760
rect 10367 5729 10379 5732
rect 10321 5723 10379 5729
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 13170 5720 13176 5772
rect 13228 5760 13234 5772
rect 13357 5763 13415 5769
rect 13357 5760 13369 5763
rect 13228 5732 13369 5760
rect 13228 5720 13234 5732
rect 13357 5729 13369 5732
rect 13403 5729 13415 5763
rect 13357 5723 13415 5729
rect 14461 5763 14519 5769
rect 14461 5729 14473 5763
rect 14507 5729 14519 5763
rect 14461 5723 14519 5729
rect 10226 5652 10232 5704
rect 10284 5692 10290 5704
rect 10413 5695 10471 5701
rect 10413 5692 10425 5695
rect 10284 5664 10425 5692
rect 10284 5652 10290 5664
rect 10413 5661 10425 5664
rect 10459 5661 10471 5695
rect 10594 5692 10600 5704
rect 10555 5664 10600 5692
rect 10413 5655 10471 5661
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 11330 5652 11336 5704
rect 11388 5692 11394 5704
rect 13449 5695 13507 5701
rect 13449 5692 13461 5695
rect 11388 5664 13461 5692
rect 11388 5652 11394 5664
rect 13449 5661 13461 5664
rect 13495 5661 13507 5695
rect 13630 5692 13636 5704
rect 13591 5664 13636 5692
rect 13449 5655 13507 5661
rect 13630 5652 13636 5664
rect 13688 5652 13694 5704
rect 8573 5587 8631 5593
rect 8680 5596 9352 5624
rect 6638 5556 6644 5568
rect 4396 5528 6316 5556
rect 6599 5528 6644 5556
rect 4396 5516 4402 5528
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 7374 5556 7380 5568
rect 7335 5528 7380 5556
rect 7374 5516 7380 5528
rect 7432 5516 7438 5568
rect 7558 5516 7564 5568
rect 7616 5556 7622 5568
rect 8680 5556 8708 5596
rect 9398 5584 9404 5636
rect 9456 5624 9462 5636
rect 12989 5627 13047 5633
rect 9456 5596 11928 5624
rect 9456 5584 9462 5596
rect 9122 5556 9128 5568
rect 7616 5528 8708 5556
rect 9083 5528 9128 5556
rect 7616 5516 7622 5528
rect 9122 5516 9128 5528
rect 9180 5516 9186 5568
rect 9950 5556 9956 5568
rect 9911 5528 9956 5556
rect 9950 5516 9956 5528
rect 10008 5516 10014 5568
rect 11900 5556 11928 5596
rect 12989 5593 13001 5627
rect 13035 5624 13047 5627
rect 14476 5624 14504 5723
rect 13035 5596 14504 5624
rect 13035 5593 13047 5596
rect 12989 5587 13047 5593
rect 14182 5556 14188 5568
rect 11900 5528 14188 5556
rect 14182 5516 14188 5528
rect 14240 5516 14246 5568
rect 1104 5466 15824 5488
rect 1104 5414 3447 5466
rect 3499 5414 3511 5466
rect 3563 5414 3575 5466
rect 3627 5414 3639 5466
rect 3691 5414 8378 5466
rect 8430 5414 8442 5466
rect 8494 5414 8506 5466
rect 8558 5414 8570 5466
rect 8622 5414 13308 5466
rect 13360 5414 13372 5466
rect 13424 5414 13436 5466
rect 13488 5414 13500 5466
rect 13552 5414 15824 5466
rect 1104 5392 15824 5414
rect 5261 5355 5319 5361
rect 2608 5324 5212 5352
rect 2608 5225 2636 5324
rect 5184 5284 5212 5324
rect 5261 5321 5273 5355
rect 5307 5352 5319 5355
rect 5350 5352 5356 5364
rect 5307 5324 5356 5352
rect 5307 5321 5319 5324
rect 5261 5315 5319 5321
rect 5350 5312 5356 5324
rect 5408 5312 5414 5364
rect 7650 5352 7656 5364
rect 5460 5324 7656 5352
rect 5460 5284 5488 5324
rect 7650 5312 7656 5324
rect 7708 5312 7714 5364
rect 9214 5352 9220 5364
rect 7944 5324 9220 5352
rect 5184 5256 5488 5284
rect 5552 5256 7788 5284
rect 2593 5219 2651 5225
rect 2593 5185 2605 5219
rect 2639 5185 2651 5219
rect 2593 5179 2651 5185
rect 2682 5176 2688 5228
rect 2740 5216 2746 5228
rect 2740 5188 4016 5216
rect 2740 5176 2746 5188
rect 1581 5151 1639 5157
rect 1581 5117 1593 5151
rect 1627 5148 1639 5151
rect 1762 5148 1768 5160
rect 1627 5120 1768 5148
rect 1627 5117 1639 5120
rect 1581 5111 1639 5117
rect 1762 5108 1768 5120
rect 1820 5108 1826 5160
rect 3145 5151 3203 5157
rect 3145 5117 3157 5151
rect 3191 5117 3203 5151
rect 3145 5111 3203 5117
rect 3160 5080 3188 5111
rect 3786 5108 3792 5160
rect 3844 5148 3850 5160
rect 3881 5151 3939 5157
rect 3881 5148 3893 5151
rect 3844 5120 3893 5148
rect 3844 5108 3850 5120
rect 3881 5117 3893 5120
rect 3927 5117 3939 5151
rect 3988 5148 4016 5188
rect 5166 5176 5172 5228
rect 5224 5216 5230 5228
rect 5552 5216 5580 5256
rect 6362 5216 6368 5228
rect 5224 5188 5580 5216
rect 6323 5188 6368 5216
rect 5224 5176 5230 5188
rect 6362 5176 6368 5188
rect 6420 5176 6426 5228
rect 6822 5216 6828 5228
rect 6783 5188 6828 5216
rect 6822 5176 6828 5188
rect 6880 5176 6886 5228
rect 6914 5176 6920 5228
rect 6972 5216 6978 5228
rect 6972 5188 7696 5216
rect 6972 5176 6978 5188
rect 4137 5151 4195 5157
rect 4137 5148 4149 5151
rect 3988 5120 4149 5148
rect 3881 5111 3939 5117
rect 4137 5117 4149 5120
rect 4183 5148 4195 5151
rect 4614 5148 4620 5160
rect 4183 5120 4620 5148
rect 4183 5117 4195 5120
rect 4137 5111 4195 5117
rect 4614 5108 4620 5120
rect 4672 5108 4678 5160
rect 6089 5151 6147 5157
rect 6089 5117 6101 5151
rect 6135 5148 6147 5151
rect 7374 5148 7380 5160
rect 6135 5120 7380 5148
rect 6135 5117 6147 5120
rect 6089 5111 6147 5117
rect 7374 5108 7380 5120
rect 7432 5108 7438 5160
rect 7668 5157 7696 5188
rect 7653 5151 7711 5157
rect 7653 5117 7665 5151
rect 7699 5117 7711 5151
rect 7760 5148 7788 5256
rect 7944 5225 7972 5324
rect 9214 5312 9220 5324
rect 9272 5352 9278 5364
rect 9677 5355 9735 5361
rect 9677 5352 9689 5355
rect 9272 5324 9689 5352
rect 9272 5312 9278 5324
rect 9677 5321 9689 5324
rect 9723 5321 9735 5355
rect 9677 5315 9735 5321
rect 10594 5312 10600 5364
rect 10652 5352 10658 5364
rect 12069 5355 12127 5361
rect 12069 5352 12081 5355
rect 10652 5324 12081 5352
rect 10652 5312 10658 5324
rect 12069 5321 12081 5324
rect 12115 5321 12127 5355
rect 12069 5315 12127 5321
rect 12253 5355 12311 5361
rect 12253 5321 12265 5355
rect 12299 5352 12311 5355
rect 13630 5352 13636 5364
rect 12299 5324 13636 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 13630 5312 13636 5324
rect 13688 5352 13694 5364
rect 13817 5355 13875 5361
rect 13817 5352 13829 5355
rect 13688 5324 13829 5352
rect 13688 5312 13694 5324
rect 13817 5321 13829 5324
rect 13863 5321 13875 5355
rect 13817 5315 13875 5321
rect 14090 5244 14096 5296
rect 14148 5284 14154 5296
rect 15930 5284 15936 5296
rect 14148 5256 15936 5284
rect 14148 5244 14154 5256
rect 15930 5244 15936 5256
rect 15988 5244 15994 5296
rect 7929 5219 7987 5225
rect 7929 5185 7941 5219
rect 7975 5185 7987 5219
rect 14734 5216 14740 5228
rect 14695 5188 14740 5216
rect 7929 5179 7987 5185
rect 14734 5176 14740 5188
rect 14792 5176 14798 5228
rect 8113 5151 8171 5157
rect 8113 5148 8125 5151
rect 7760 5120 8125 5148
rect 7653 5111 7711 5117
rect 8113 5117 8125 5120
rect 8159 5117 8171 5151
rect 8113 5111 8171 5117
rect 8297 5151 8355 5157
rect 8297 5117 8309 5151
rect 8343 5148 8355 5151
rect 9490 5148 9496 5160
rect 8343 5120 9496 5148
rect 8343 5117 8355 5120
rect 8297 5111 8355 5117
rect 6181 5083 6239 5089
rect 3160 5052 6132 5080
rect 1394 4972 1400 5024
rect 1452 5012 1458 5024
rect 1765 5015 1823 5021
rect 1765 5012 1777 5015
rect 1452 4984 1777 5012
rect 1452 4972 1458 4984
rect 1765 4981 1777 4984
rect 1811 4981 1823 5015
rect 1765 4975 1823 4981
rect 2133 5015 2191 5021
rect 2133 4981 2145 5015
rect 2179 5012 2191 5015
rect 2314 5012 2320 5024
rect 2179 4984 2320 5012
rect 2179 4981 2191 4984
rect 2133 4975 2191 4981
rect 2314 4972 2320 4984
rect 2372 4972 2378 5024
rect 2498 5012 2504 5024
rect 2459 4984 2504 5012
rect 2498 4972 2504 4984
rect 2556 4972 2562 5024
rect 2958 4972 2964 5024
rect 3016 5012 3022 5024
rect 3329 5015 3387 5021
rect 3329 5012 3341 5015
rect 3016 4984 3341 5012
rect 3016 4972 3022 4984
rect 3329 4981 3341 4984
rect 3375 4981 3387 5015
rect 5718 5012 5724 5024
rect 5679 4984 5724 5012
rect 3329 4975 3387 4981
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 6104 5012 6132 5052
rect 6181 5049 6193 5083
rect 6227 5080 6239 5083
rect 7668 5080 7696 5111
rect 9490 5108 9496 5120
rect 9548 5108 9554 5160
rect 9858 5108 9864 5160
rect 9916 5148 9922 5160
rect 9953 5151 10011 5157
rect 9953 5148 9965 5151
rect 9916 5120 9965 5148
rect 9916 5108 9922 5120
rect 9953 5117 9965 5120
rect 9999 5117 10011 5151
rect 9953 5111 10011 5117
rect 10134 5108 10140 5160
rect 10192 5148 10198 5160
rect 10689 5151 10747 5157
rect 10689 5148 10701 5151
rect 10192 5120 10701 5148
rect 10192 5108 10198 5120
rect 10689 5117 10701 5120
rect 10735 5148 10747 5151
rect 12437 5151 12495 5157
rect 12437 5148 12449 5151
rect 10735 5120 12449 5148
rect 10735 5117 10747 5120
rect 10689 5111 10747 5117
rect 12437 5117 12449 5120
rect 12483 5148 12495 5151
rect 12526 5148 12532 5160
rect 12483 5120 12532 5148
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 12526 5108 12532 5120
rect 12584 5108 12590 5160
rect 14553 5151 14611 5157
rect 14553 5117 14565 5151
rect 14599 5148 14611 5151
rect 14918 5148 14924 5160
rect 14599 5120 14924 5148
rect 14599 5117 14611 5120
rect 14553 5111 14611 5117
rect 14918 5108 14924 5120
rect 14976 5108 14982 5160
rect 8386 5080 8392 5092
rect 6227 5052 7328 5080
rect 7668 5052 8392 5080
rect 6227 5049 6239 5052
rect 6181 5043 6239 5049
rect 6914 5012 6920 5024
rect 6104 4984 6920 5012
rect 6914 4972 6920 4984
rect 6972 5012 6978 5024
rect 7190 5012 7196 5024
rect 6972 4984 7196 5012
rect 6972 4972 6978 4984
rect 7190 4972 7196 4984
rect 7248 4972 7254 5024
rect 7300 5021 7328 5052
rect 8386 5040 8392 5052
rect 8444 5040 8450 5092
rect 8564 5083 8622 5089
rect 8564 5049 8576 5083
rect 8610 5080 8622 5083
rect 8754 5080 8760 5092
rect 8610 5052 8760 5080
rect 8610 5049 8622 5052
rect 8564 5043 8622 5049
rect 8754 5040 8760 5052
rect 8812 5040 8818 5092
rect 10502 5080 10508 5092
rect 8864 5052 10508 5080
rect 7285 5015 7343 5021
rect 7285 4981 7297 5015
rect 7331 4981 7343 5015
rect 7742 5012 7748 5024
rect 7703 4984 7748 5012
rect 7285 4975 7343 4981
rect 7742 4972 7748 4984
rect 7800 4972 7806 5024
rect 8113 5015 8171 5021
rect 8113 4981 8125 5015
rect 8159 5012 8171 5015
rect 8864 5012 8892 5052
rect 10502 5040 10508 5052
rect 10560 5040 10566 5092
rect 10934 5083 10992 5089
rect 10934 5080 10946 5083
rect 10796 5052 10946 5080
rect 8159 4984 8892 5012
rect 8159 4981 8171 4984
rect 8113 4975 8171 4981
rect 8938 4972 8944 5024
rect 8996 5012 9002 5024
rect 10137 5015 10195 5021
rect 10137 5012 10149 5015
rect 8996 4984 10149 5012
rect 8996 4972 9002 4984
rect 10137 4981 10149 4984
rect 10183 4981 10195 5015
rect 10796 5012 10824 5052
rect 10934 5049 10946 5052
rect 10980 5049 10992 5083
rect 10934 5043 10992 5049
rect 12618 5040 12624 5092
rect 12676 5089 12682 5092
rect 12676 5083 12740 5089
rect 12676 5049 12694 5083
rect 12728 5049 12740 5083
rect 12676 5043 12740 5049
rect 12676 5040 12682 5043
rect 12253 5015 12311 5021
rect 12253 5012 12265 5015
rect 10796 4984 12265 5012
rect 10137 4975 10195 4981
rect 12253 4981 12265 4984
rect 12299 4981 12311 5015
rect 14090 5012 14096 5024
rect 14051 4984 14096 5012
rect 12253 4975 12311 4981
rect 14090 4972 14096 4984
rect 14148 4972 14154 5024
rect 14458 5012 14464 5024
rect 14419 4984 14464 5012
rect 14458 4972 14464 4984
rect 14516 4972 14522 5024
rect 1104 4922 15824 4944
rect 1104 4870 5912 4922
rect 5964 4870 5976 4922
rect 6028 4870 6040 4922
rect 6092 4870 6104 4922
rect 6156 4870 10843 4922
rect 10895 4870 10907 4922
rect 10959 4870 10971 4922
rect 11023 4870 11035 4922
rect 11087 4870 15824 4922
rect 1104 4848 15824 4870
rect 1857 4811 1915 4817
rect 1857 4777 1869 4811
rect 1903 4777 1915 4811
rect 2314 4808 2320 4820
rect 2275 4780 2320 4808
rect 1857 4771 1915 4777
rect 1872 4672 1900 4771
rect 2314 4768 2320 4780
rect 2372 4768 2378 4820
rect 2866 4808 2872 4820
rect 2827 4780 2872 4808
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 3237 4811 3295 4817
rect 3237 4777 3249 4811
rect 3283 4808 3295 4811
rect 3326 4808 3332 4820
rect 3283 4780 3332 4808
rect 3283 4777 3295 4780
rect 3237 4771 3295 4777
rect 3326 4768 3332 4780
rect 3384 4768 3390 4820
rect 5166 4768 5172 4820
rect 5224 4768 5230 4820
rect 6270 4808 6276 4820
rect 5828 4780 6276 4808
rect 2222 4740 2228 4752
rect 2183 4712 2228 4740
rect 2222 4700 2228 4712
rect 2280 4700 2286 4752
rect 5184 4740 5212 4768
rect 4080 4712 5212 4740
rect 4080 4681 4108 4712
rect 3329 4675 3387 4681
rect 3329 4672 3341 4675
rect 1872 4644 3341 4672
rect 3329 4641 3341 4644
rect 3375 4641 3387 4675
rect 3329 4635 3387 4641
rect 4065 4675 4123 4681
rect 4065 4641 4077 4675
rect 4111 4641 4123 4675
rect 4065 4635 4123 4641
rect 4617 4675 4675 4681
rect 4617 4641 4629 4675
rect 4663 4641 4675 4675
rect 4617 4635 4675 4641
rect 2406 4604 2412 4616
rect 2367 4576 2412 4604
rect 2406 4564 2412 4576
rect 2464 4564 2470 4616
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4604 3571 4607
rect 4154 4604 4160 4616
rect 3559 4576 4160 4604
rect 3559 4573 3571 4576
rect 3513 4567 3571 4573
rect 4154 4564 4160 4576
rect 4212 4564 4218 4616
rect 4632 4604 4660 4635
rect 5074 4632 5080 4684
rect 5132 4672 5138 4684
rect 5828 4681 5856 4780
rect 6270 4768 6276 4780
rect 6328 4768 6334 4820
rect 7561 4811 7619 4817
rect 7561 4777 7573 4811
rect 7607 4808 7619 4811
rect 7742 4808 7748 4820
rect 7607 4780 7748 4808
rect 7607 4777 7619 4780
rect 7561 4771 7619 4777
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 8941 4811 8999 4817
rect 8941 4777 8953 4811
rect 8987 4808 8999 4811
rect 9950 4808 9956 4820
rect 8987 4780 9956 4808
rect 8987 4777 8999 4780
rect 8941 4771 8999 4777
rect 9950 4768 9956 4780
rect 10008 4768 10014 4820
rect 12618 4768 12624 4820
rect 12676 4808 12682 4820
rect 13909 4811 13967 4817
rect 13909 4808 13921 4811
rect 12676 4780 13921 4808
rect 12676 4768 12682 4780
rect 13909 4777 13921 4780
rect 13955 4777 13967 4811
rect 14550 4808 14556 4820
rect 14511 4780 14556 4808
rect 13909 4771 13967 4777
rect 14550 4768 14556 4780
rect 14608 4808 14614 4820
rect 15102 4808 15108 4820
rect 14608 4780 15108 4808
rect 14608 4768 14614 4780
rect 15102 4768 15108 4780
rect 15160 4768 15166 4820
rect 6080 4743 6138 4749
rect 6080 4709 6092 4743
rect 6126 4740 6138 4743
rect 6638 4740 6644 4752
rect 6126 4712 6644 4740
rect 6126 4709 6138 4712
rect 6080 4703 6138 4709
rect 6638 4700 6644 4712
rect 6696 4700 6702 4752
rect 7650 4700 7656 4752
rect 7708 4740 7714 4752
rect 8018 4740 8024 4752
rect 7708 4712 8024 4740
rect 7708 4700 7714 4712
rect 8018 4700 8024 4712
rect 8076 4700 8082 4752
rect 9033 4743 9091 4749
rect 9033 4709 9045 4743
rect 9079 4740 9091 4743
rect 9766 4740 9772 4752
rect 9079 4712 9772 4740
rect 9079 4709 9091 4712
rect 9033 4703 9091 4709
rect 9766 4700 9772 4712
rect 9824 4700 9830 4752
rect 10496 4743 10554 4749
rect 10496 4709 10508 4743
rect 10542 4740 10554 4743
rect 10594 4740 10600 4752
rect 10542 4712 10600 4740
rect 10542 4709 10554 4712
rect 10496 4703 10554 4709
rect 10594 4700 10600 4712
rect 10652 4700 10658 4752
rect 12066 4700 12072 4752
rect 12124 4740 12130 4752
rect 14645 4743 14703 4749
rect 14645 4740 14657 4743
rect 12124 4712 14657 4740
rect 12124 4700 12130 4712
rect 14645 4709 14657 4712
rect 14691 4740 14703 4743
rect 15010 4740 15016 4752
rect 14691 4712 15016 4740
rect 14691 4709 14703 4712
rect 14645 4703 14703 4709
rect 15010 4700 15016 4712
rect 15068 4700 15074 4752
rect 5169 4675 5227 4681
rect 5169 4672 5181 4675
rect 5132 4644 5181 4672
rect 5132 4632 5138 4644
rect 5169 4641 5181 4644
rect 5215 4641 5227 4675
rect 5169 4635 5227 4641
rect 5813 4675 5871 4681
rect 5813 4641 5825 4675
rect 5859 4641 5871 4675
rect 6546 4672 6552 4684
rect 5813 4635 5871 4641
rect 5920 4644 6552 4672
rect 5920 4604 5948 4644
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 7834 4632 7840 4684
rect 7892 4672 7898 4684
rect 7929 4675 7987 4681
rect 7929 4672 7941 4675
rect 7892 4644 7941 4672
rect 7892 4632 7898 4644
rect 7929 4641 7941 4644
rect 7975 4641 7987 4675
rect 7929 4635 7987 4641
rect 9398 4632 9404 4684
rect 9456 4672 9462 4684
rect 9677 4675 9735 4681
rect 9677 4672 9689 4675
rect 9456 4644 9689 4672
rect 9456 4632 9462 4644
rect 9677 4641 9689 4644
rect 9723 4641 9735 4675
rect 12796 4675 12854 4681
rect 9677 4635 9735 4641
rect 10152 4644 11652 4672
rect 4632 4576 5948 4604
rect 8205 4607 8263 4613
rect 8205 4573 8217 4607
rect 8251 4604 8263 4607
rect 8754 4604 8760 4616
rect 8251 4576 8760 4604
rect 8251 4573 8263 4576
rect 8205 4567 8263 4573
rect 8754 4564 8760 4576
rect 8812 4604 8818 4616
rect 8938 4604 8944 4616
rect 8812 4576 8944 4604
rect 8812 4564 8818 4576
rect 8938 4564 8944 4576
rect 8996 4564 9002 4616
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4604 9275 4607
rect 10152 4604 10180 4644
rect 9263 4576 10180 4604
rect 10229 4607 10287 4613
rect 9263 4573 9275 4576
rect 9217 4567 9275 4573
rect 10229 4573 10241 4607
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 3050 4496 3056 4548
rect 3108 4536 3114 4548
rect 5353 4539 5411 4545
rect 5353 4536 5365 4539
rect 3108 4508 5365 4536
rect 3108 4496 3114 4508
rect 5353 4505 5365 4508
rect 5399 4505 5411 4539
rect 5353 4499 5411 4505
rect 8110 4496 8116 4548
rect 8168 4536 8174 4548
rect 9861 4539 9919 4545
rect 9861 4536 9873 4539
rect 8168 4508 9873 4536
rect 8168 4496 8174 4508
rect 9861 4505 9873 4508
rect 9907 4505 9919 4539
rect 9861 4499 9919 4505
rect 10134 4496 10140 4548
rect 10192 4536 10198 4548
rect 10244 4536 10272 4567
rect 11624 4548 11652 4644
rect 12796 4641 12808 4675
rect 12842 4672 12854 4675
rect 13722 4672 13728 4684
rect 12842 4644 13728 4672
rect 12842 4641 12854 4644
rect 12796 4635 12854 4641
rect 13722 4632 13728 4644
rect 13780 4632 13786 4684
rect 12526 4604 12532 4616
rect 12487 4576 12532 4604
rect 12526 4564 12532 4576
rect 12584 4564 12590 4616
rect 13740 4604 13768 4632
rect 14734 4604 14740 4616
rect 13740 4576 14740 4604
rect 14734 4564 14740 4576
rect 14792 4564 14798 4616
rect 11606 4536 11612 4548
rect 10192 4508 10272 4536
rect 11567 4508 11612 4536
rect 10192 4496 10198 4508
rect 11606 4496 11612 4508
rect 11664 4496 11670 4548
rect 4246 4468 4252 4480
rect 4207 4440 4252 4468
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 4798 4468 4804 4480
rect 4759 4440 4804 4468
rect 4798 4428 4804 4440
rect 4856 4428 4862 4480
rect 7190 4468 7196 4480
rect 7151 4440 7196 4468
rect 7190 4428 7196 4440
rect 7248 4428 7254 4480
rect 8573 4471 8631 4477
rect 8573 4437 8585 4471
rect 8619 4468 8631 4471
rect 9030 4468 9036 4480
rect 8619 4440 9036 4468
rect 8619 4437 8631 4440
rect 8573 4431 8631 4437
rect 9030 4428 9036 4440
rect 9088 4428 9094 4480
rect 9490 4428 9496 4480
rect 9548 4468 9554 4480
rect 10152 4468 10180 4496
rect 14182 4468 14188 4480
rect 9548 4440 10180 4468
rect 14143 4440 14188 4468
rect 9548 4428 9554 4440
rect 14182 4428 14188 4440
rect 14240 4428 14246 4480
rect 1104 4378 15824 4400
rect 1104 4326 3447 4378
rect 3499 4326 3511 4378
rect 3563 4326 3575 4378
rect 3627 4326 3639 4378
rect 3691 4326 8378 4378
rect 8430 4326 8442 4378
rect 8494 4326 8506 4378
rect 8558 4326 8570 4378
rect 8622 4326 13308 4378
rect 13360 4326 13372 4378
rect 13424 4326 13436 4378
rect 13488 4326 13500 4378
rect 13552 4326 15824 4378
rect 1104 4304 15824 4326
rect 2498 4224 2504 4276
rect 2556 4264 2562 4276
rect 4341 4267 4399 4273
rect 2556 4236 4292 4264
rect 2556 4224 2562 4236
rect 4264 4196 4292 4236
rect 4341 4233 4353 4267
rect 4387 4264 4399 4267
rect 4614 4264 4620 4276
rect 4387 4236 4620 4264
rect 4387 4233 4399 4236
rect 4341 4227 4399 4233
rect 4614 4224 4620 4236
rect 4672 4224 4678 4276
rect 7834 4264 7840 4276
rect 6288 4236 7840 4264
rect 6288 4196 6316 4236
rect 7834 4224 7840 4236
rect 7892 4224 7898 4276
rect 8018 4224 8024 4276
rect 8076 4264 8082 4276
rect 8076 4236 8800 4264
rect 8076 4224 8082 4236
rect 6638 4196 6644 4208
rect 4264 4168 6316 4196
rect 6380 4168 6644 4196
rect 1670 4128 1676 4140
rect 1631 4100 1676 4128
rect 1670 4088 1676 4100
rect 1728 4088 1734 4140
rect 1964 4100 3096 4128
rect 1489 4063 1547 4069
rect 1489 4029 1501 4063
rect 1535 4060 1547 4063
rect 1964 4060 1992 4100
rect 2222 4060 2228 4072
rect 1535 4032 1992 4060
rect 2183 4032 2228 4060
rect 1535 4029 1547 4032
rect 1489 4023 1547 4029
rect 2222 4020 2228 4032
rect 2280 4020 2286 4072
rect 2501 4063 2559 4069
rect 2501 4029 2513 4063
rect 2547 4060 2559 4063
rect 2774 4060 2780 4072
rect 2547 4032 2780 4060
rect 2547 4029 2559 4032
rect 2501 4023 2559 4029
rect 2774 4020 2780 4032
rect 2832 4020 2838 4072
rect 2961 4063 3019 4069
rect 2961 4029 2973 4063
rect 3007 4029 3019 4063
rect 3068 4060 3096 4100
rect 4430 4088 4436 4140
rect 4488 4128 4494 4140
rect 4614 4128 4620 4140
rect 4488 4100 4620 4128
rect 4488 4088 4494 4100
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 5258 4128 5264 4140
rect 5219 4100 5264 4128
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 5718 4088 5724 4140
rect 5776 4128 5782 4140
rect 6380 4137 6408 4168
rect 6638 4156 6644 4168
rect 6696 4156 6702 4208
rect 8772 4196 8800 4236
rect 8938 4224 8944 4276
rect 8996 4264 9002 4276
rect 9217 4267 9275 4273
rect 9217 4264 9229 4267
rect 8996 4236 9229 4264
rect 8996 4224 9002 4236
rect 9217 4233 9229 4236
rect 9263 4233 9275 4267
rect 9490 4264 9496 4276
rect 9451 4236 9496 4264
rect 9217 4227 9275 4233
rect 9490 4224 9496 4236
rect 9548 4224 9554 4276
rect 9766 4264 9772 4276
rect 9727 4236 9772 4264
rect 9766 4224 9772 4236
rect 9824 4224 9830 4276
rect 12618 4196 12624 4208
rect 8772 4168 10732 4196
rect 6181 4131 6239 4137
rect 6181 4128 6193 4131
rect 5776 4100 6193 4128
rect 5776 4088 5782 4100
rect 6181 4097 6193 4100
rect 6227 4097 6239 4131
rect 6181 4091 6239 4097
rect 6365 4131 6423 4137
rect 6365 4097 6377 4131
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 10413 4131 10471 4137
rect 10413 4097 10425 4131
rect 10459 4128 10471 4131
rect 10594 4128 10600 4140
rect 10459 4100 10600 4128
rect 10459 4097 10471 4100
rect 10413 4091 10471 4097
rect 10594 4088 10600 4100
rect 10652 4088 10658 4140
rect 10704 4128 10732 4168
rect 11992 4168 12624 4196
rect 11882 4128 11888 4140
rect 10704 4100 11888 4128
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 11992 4137 12020 4168
rect 12618 4156 12624 4168
rect 12676 4196 12682 4208
rect 12676 4168 14044 4196
rect 12676 4156 12682 4168
rect 11977 4131 12035 4137
rect 11977 4097 11989 4131
rect 12023 4097 12035 4131
rect 11977 4091 12035 4097
rect 13081 4131 13139 4137
rect 13081 4097 13093 4131
rect 13127 4128 13139 4131
rect 13722 4128 13728 4140
rect 13127 4100 13728 4128
rect 13127 4097 13139 4100
rect 13081 4091 13139 4097
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 14016 4137 14044 4168
rect 14001 4131 14059 4137
rect 14001 4097 14013 4131
rect 14047 4097 14059 4131
rect 14458 4128 14464 4140
rect 14419 4100 14464 4128
rect 14001 4091 14059 4097
rect 14458 4088 14464 4100
rect 14516 4088 14522 4140
rect 3068 4032 5764 4060
rect 2961 4023 3019 4029
rect 1946 3884 1952 3936
rect 2004 3924 2010 3936
rect 2976 3924 3004 4023
rect 3228 3995 3286 4001
rect 3228 3961 3240 3995
rect 3274 3992 3286 3995
rect 3326 3992 3332 4004
rect 3274 3964 3332 3992
rect 3274 3961 3286 3964
rect 3228 3955 3286 3961
rect 3326 3952 3332 3964
rect 3384 3952 3390 4004
rect 3694 3952 3700 4004
rect 3752 3992 3758 4004
rect 4982 3992 4988 4004
rect 3752 3964 4988 3992
rect 3752 3952 3758 3964
rect 4982 3952 4988 3964
rect 5040 3952 5046 4004
rect 5077 3995 5135 4001
rect 5077 3961 5089 3995
rect 5123 3992 5135 3995
rect 5442 3992 5448 4004
rect 5123 3964 5448 3992
rect 5123 3961 5135 3964
rect 5077 3955 5135 3961
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 3786 3924 3792 3936
rect 2004 3896 3792 3924
rect 2004 3884 2010 3896
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 4706 3924 4712 3936
rect 4667 3896 4712 3924
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 5166 3884 5172 3936
rect 5224 3924 5230 3936
rect 5736 3933 5764 4032
rect 5810 4020 5816 4072
rect 5868 4060 5874 4072
rect 6089 4063 6147 4069
rect 6089 4060 6101 4063
rect 5868 4032 6101 4060
rect 5868 4020 5874 4032
rect 6089 4029 6101 4032
rect 6135 4029 6147 4063
rect 6089 4023 6147 4029
rect 6730 4020 6736 4072
rect 6788 4060 6794 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6788 4032 6837 4060
rect 6788 4020 6794 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 7834 4060 7840 4072
rect 7795 4032 7840 4060
rect 6825 4023 6883 4029
rect 7834 4020 7840 4032
rect 7892 4020 7898 4072
rect 7944 4032 8331 4060
rect 6546 3952 6552 4004
rect 6604 3992 6610 4004
rect 7944 3992 7972 4032
rect 6604 3964 7972 3992
rect 8104 3995 8162 4001
rect 6604 3952 6610 3964
rect 8104 3961 8116 3995
rect 8150 3992 8162 3995
rect 8202 3992 8208 4004
rect 8150 3964 8208 3992
rect 8150 3961 8162 3964
rect 8104 3955 8162 3961
rect 8202 3952 8208 3964
rect 8260 3952 8266 4004
rect 8303 3992 8331 4032
rect 8662 4020 8668 4072
rect 8720 4060 8726 4072
rect 9214 4060 9220 4072
rect 8720 4032 9220 4060
rect 8720 4020 8726 4032
rect 9214 4020 9220 4032
rect 9272 4020 9278 4072
rect 9677 4063 9735 4069
rect 9677 4029 9689 4063
rect 9723 4060 9735 4063
rect 10686 4060 10692 4072
rect 9723 4032 10692 4060
rect 9723 4029 9735 4032
rect 9677 4023 9735 4029
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 10778 4020 10784 4072
rect 10836 4060 10842 4072
rect 10836 4032 10881 4060
rect 10836 4020 10842 4032
rect 11146 4020 11152 4072
rect 11204 4060 11210 4072
rect 13909 4063 13967 4069
rect 11204 4032 13584 4060
rect 11204 4020 11210 4032
rect 8303 3964 11008 3992
rect 5721 3927 5779 3933
rect 5224 3896 5269 3924
rect 5224 3884 5230 3896
rect 5721 3893 5733 3927
rect 5767 3893 5779 3927
rect 5721 3887 5779 3893
rect 5810 3884 5816 3936
rect 5868 3924 5874 3936
rect 7009 3927 7067 3933
rect 7009 3924 7021 3927
rect 5868 3896 7021 3924
rect 5868 3884 5874 3896
rect 7009 3893 7021 3896
rect 7055 3893 7067 3927
rect 7009 3887 7067 3893
rect 7374 3884 7380 3936
rect 7432 3924 7438 3936
rect 9122 3924 9128 3936
rect 7432 3896 9128 3924
rect 7432 3884 7438 3896
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 9766 3884 9772 3936
rect 9824 3924 9830 3936
rect 10042 3924 10048 3936
rect 9824 3896 10048 3924
rect 9824 3884 9830 3896
rect 10042 3884 10048 3896
rect 10100 3924 10106 3936
rect 10137 3927 10195 3933
rect 10137 3924 10149 3927
rect 10100 3896 10149 3924
rect 10100 3884 10106 3896
rect 10137 3893 10149 3896
rect 10183 3893 10195 3927
rect 10137 3887 10195 3893
rect 10229 3927 10287 3933
rect 10229 3893 10241 3927
rect 10275 3924 10287 3927
rect 10318 3924 10324 3936
rect 10275 3896 10324 3924
rect 10275 3893 10287 3896
rect 10229 3887 10287 3893
rect 10318 3884 10324 3896
rect 10376 3884 10382 3936
rect 10410 3884 10416 3936
rect 10468 3924 10474 3936
rect 10686 3924 10692 3936
rect 10468 3896 10692 3924
rect 10468 3884 10474 3896
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 10980 3933 11008 3964
rect 11882 3952 11888 4004
rect 11940 3992 11946 4004
rect 12342 3992 12348 4004
rect 11940 3964 12348 3992
rect 11940 3952 11946 3964
rect 12342 3952 12348 3964
rect 12400 3952 12406 4004
rect 10965 3927 11023 3933
rect 10965 3893 10977 3927
rect 11011 3893 11023 3927
rect 11330 3924 11336 3936
rect 11291 3896 11336 3924
rect 10965 3887 11023 3893
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 11422 3884 11428 3936
rect 11480 3924 11486 3936
rect 11701 3927 11759 3933
rect 11701 3924 11713 3927
rect 11480 3896 11713 3924
rect 11480 3884 11486 3896
rect 11701 3893 11713 3896
rect 11747 3893 11759 3927
rect 11701 3887 11759 3893
rect 11793 3927 11851 3933
rect 11793 3893 11805 3927
rect 11839 3924 11851 3927
rect 12437 3927 12495 3933
rect 12437 3924 12449 3927
rect 11839 3896 12449 3924
rect 11839 3893 11851 3896
rect 11793 3887 11851 3893
rect 12437 3893 12449 3896
rect 12483 3893 12495 3927
rect 12437 3887 12495 3893
rect 12618 3884 12624 3936
rect 12676 3924 12682 3936
rect 12805 3927 12863 3933
rect 12805 3924 12817 3927
rect 12676 3896 12817 3924
rect 12676 3884 12682 3896
rect 12805 3893 12817 3896
rect 12851 3893 12863 3927
rect 12805 3887 12863 3893
rect 12894 3884 12900 3936
rect 12952 3924 12958 3936
rect 12952 3896 12997 3924
rect 12952 3884 12958 3896
rect 13170 3884 13176 3936
rect 13228 3924 13234 3936
rect 13449 3927 13507 3933
rect 13449 3924 13461 3927
rect 13228 3896 13461 3924
rect 13228 3884 13234 3896
rect 13449 3893 13461 3896
rect 13495 3893 13507 3927
rect 13556 3924 13584 4032
rect 13909 4029 13921 4063
rect 13955 4060 13967 4063
rect 14182 4060 14188 4072
rect 13955 4032 14188 4060
rect 13955 4029 13967 4032
rect 13909 4023 13967 4029
rect 14182 4020 14188 4032
rect 14240 4020 14246 4072
rect 13817 3995 13875 4001
rect 13817 3961 13829 3995
rect 13863 3992 13875 3995
rect 14090 3992 14096 4004
rect 13863 3964 14096 3992
rect 13863 3961 13875 3964
rect 13817 3955 13875 3961
rect 14090 3952 14096 3964
rect 14148 3952 14154 4004
rect 14366 3924 14372 3936
rect 13556 3896 14372 3924
rect 13449 3887 13507 3893
rect 14366 3884 14372 3896
rect 14424 3884 14430 3936
rect 1104 3834 15824 3856
rect 1104 3782 5912 3834
rect 5964 3782 5976 3834
rect 6028 3782 6040 3834
rect 6092 3782 6104 3834
rect 6156 3782 10843 3834
rect 10895 3782 10907 3834
rect 10959 3782 10971 3834
rect 11023 3782 11035 3834
rect 11087 3782 15824 3834
rect 1104 3760 15824 3782
rect 4522 3720 4528 3732
rect 3896 3692 4528 3720
rect 2216 3655 2274 3661
rect 1412 3624 2176 3652
rect 1412 3593 1440 3624
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3553 1455 3587
rect 1946 3584 1952 3596
rect 1907 3556 1952 3584
rect 1397 3547 1455 3553
rect 1946 3544 1952 3556
rect 2004 3544 2010 3596
rect 2148 3584 2176 3624
rect 2216 3621 2228 3655
rect 2262 3652 2274 3655
rect 3234 3652 3240 3664
rect 2262 3624 3240 3652
rect 2262 3621 2274 3624
rect 2216 3615 2274 3621
rect 3234 3612 3240 3624
rect 3292 3612 3298 3664
rect 3694 3584 3700 3596
rect 2148 3556 3700 3584
rect 3694 3544 3700 3556
rect 3752 3544 3758 3596
rect 3896 3593 3924 3692
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 4982 3680 4988 3732
rect 5040 3720 5046 3732
rect 6638 3720 6644 3732
rect 5040 3692 6644 3720
rect 5040 3680 5046 3692
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 6822 3680 6828 3732
rect 6880 3720 6886 3732
rect 6880 3692 7328 3720
rect 6880 3680 6886 3692
rect 4338 3612 4344 3664
rect 4396 3652 4402 3664
rect 5258 3652 5264 3664
rect 4396 3624 5264 3652
rect 4396 3612 4402 3624
rect 5258 3612 5264 3624
rect 5316 3652 5322 3664
rect 6724 3655 6782 3661
rect 5316 3624 5672 3652
rect 5316 3612 5322 3624
rect 3881 3587 3939 3593
rect 3881 3553 3893 3587
rect 3927 3553 3939 3587
rect 3881 3547 3939 3553
rect 4430 3544 4436 3596
rect 4488 3544 4494 3596
rect 4608 3587 4666 3593
rect 4608 3553 4620 3587
rect 4654 3584 4666 3587
rect 4982 3584 4988 3596
rect 4654 3556 4988 3584
rect 4654 3553 4666 3556
rect 4608 3547 4666 3553
rect 4982 3544 4988 3556
rect 5040 3544 5046 3596
rect 3786 3476 3792 3528
rect 3844 3476 3850 3528
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3516 4399 3519
rect 4448 3516 4476 3544
rect 4387 3488 4476 3516
rect 4387 3485 4399 3488
rect 4341 3479 4399 3485
rect 3697 3451 3755 3457
rect 3697 3417 3709 3451
rect 3743 3448 3755 3451
rect 3804 3448 3832 3476
rect 4356 3448 4384 3479
rect 3743 3420 4384 3448
rect 5644 3448 5672 3624
rect 6724 3621 6736 3655
rect 6770 3652 6782 3655
rect 7190 3652 7196 3664
rect 6770 3624 7196 3652
rect 6770 3621 6782 3624
rect 6724 3615 6782 3621
rect 7190 3612 7196 3624
rect 7248 3612 7254 3664
rect 7300 3652 7328 3692
rect 7650 3680 7656 3732
rect 7708 3720 7714 3732
rect 8846 3720 8852 3732
rect 7708 3692 8852 3720
rect 7708 3680 7714 3692
rect 8846 3680 8852 3692
rect 8904 3680 8910 3732
rect 9030 3720 9036 3732
rect 8991 3692 9036 3720
rect 9030 3680 9036 3692
rect 9088 3680 9094 3732
rect 10321 3723 10379 3729
rect 10321 3689 10333 3723
rect 10367 3720 10379 3723
rect 10502 3720 10508 3732
rect 10367 3692 10508 3720
rect 10367 3689 10379 3692
rect 10321 3683 10379 3689
rect 10502 3680 10508 3692
rect 10560 3680 10566 3732
rect 11422 3720 11428 3732
rect 11383 3692 11428 3720
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 11790 3720 11796 3732
rect 11751 3692 11796 3720
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 11882 3680 11888 3732
rect 11940 3720 11946 3732
rect 12897 3723 12955 3729
rect 12897 3720 12909 3723
rect 11940 3692 12909 3720
rect 11940 3680 11946 3692
rect 12897 3689 12909 3692
rect 12943 3689 12955 3723
rect 13906 3720 13912 3732
rect 13867 3692 13912 3720
rect 12897 3683 12955 3689
rect 13906 3680 13912 3692
rect 13964 3680 13970 3732
rect 11146 3652 11152 3664
rect 7300 3624 11152 3652
rect 11146 3612 11152 3624
rect 11204 3612 11210 3664
rect 11808 3652 11836 3680
rect 12342 3652 12348 3664
rect 11808 3624 12348 3652
rect 12342 3612 12348 3624
rect 12400 3612 12406 3664
rect 12434 3612 12440 3664
rect 12492 3652 12498 3664
rect 13817 3655 13875 3661
rect 13817 3652 13829 3655
rect 12492 3624 13829 3652
rect 12492 3612 12498 3624
rect 13817 3621 13829 3624
rect 13863 3621 13875 3655
rect 13817 3615 13875 3621
rect 6270 3544 6276 3596
rect 6328 3584 6334 3596
rect 8110 3584 8116 3596
rect 6328 3556 8116 3584
rect 6328 3544 6334 3556
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 8941 3587 8999 3593
rect 8941 3553 8953 3587
rect 8987 3584 8999 3587
rect 9766 3584 9772 3596
rect 8987 3556 9772 3584
rect 8987 3553 8999 3556
rect 8941 3547 8999 3553
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 12710 3544 12716 3596
rect 12768 3584 12774 3596
rect 12805 3587 12863 3593
rect 12805 3584 12817 3587
rect 12768 3556 12817 3584
rect 12768 3544 12774 3556
rect 12805 3553 12817 3556
rect 12851 3553 12863 3587
rect 13722 3584 13728 3596
rect 12805 3547 12863 3553
rect 13004 3556 13728 3584
rect 6362 3476 6368 3528
rect 6420 3516 6426 3528
rect 6457 3519 6515 3525
rect 6457 3516 6469 3519
rect 6420 3488 6469 3516
rect 6420 3476 6426 3488
rect 6457 3485 6469 3488
rect 6503 3485 6515 3519
rect 6457 3479 6515 3485
rect 7834 3476 7840 3528
rect 7892 3516 7898 3528
rect 9217 3519 9275 3525
rect 7892 3488 9168 3516
rect 7892 3476 7898 3488
rect 5721 3451 5779 3457
rect 5721 3448 5733 3451
rect 5644 3420 5733 3448
rect 3743 3417 3755 3420
rect 3697 3411 3755 3417
rect 5721 3417 5733 3420
rect 5767 3417 5779 3451
rect 5721 3411 5779 3417
rect 7926 3408 7932 3460
rect 7984 3448 7990 3460
rect 9140 3448 9168 3488
rect 9217 3485 9229 3519
rect 9263 3516 9275 3519
rect 9398 3516 9404 3528
rect 9263 3488 9404 3516
rect 9263 3485 9275 3488
rect 9217 3479 9275 3485
rect 9398 3476 9404 3488
rect 9456 3476 9462 3528
rect 9582 3476 9588 3528
rect 9640 3516 9646 3528
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 9640 3488 10425 3516
rect 9640 3476 9646 3488
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 10594 3516 10600 3528
rect 10555 3488 10600 3516
rect 10413 3479 10471 3485
rect 9674 3448 9680 3460
rect 7984 3420 8800 3448
rect 9140 3420 9680 3448
rect 7984 3408 7990 3420
rect 566 3340 572 3392
rect 624 3380 630 3392
rect 1581 3383 1639 3389
rect 1581 3380 1593 3383
rect 624 3352 1593 3380
rect 624 3340 630 3352
rect 1581 3349 1593 3352
rect 1627 3349 1639 3383
rect 3326 3380 3332 3392
rect 3287 3352 3332 3380
rect 1581 3343 1639 3349
rect 3326 3340 3332 3352
rect 3384 3340 3390 3392
rect 3786 3340 3792 3392
rect 3844 3380 3850 3392
rect 5810 3380 5816 3392
rect 3844 3352 5816 3380
rect 3844 3340 3850 3352
rect 5810 3340 5816 3352
rect 5868 3340 5874 3392
rect 6362 3340 6368 3392
rect 6420 3380 6426 3392
rect 6730 3380 6736 3392
rect 6420 3352 6736 3380
rect 6420 3340 6426 3352
rect 6730 3340 6736 3352
rect 6788 3380 6794 3392
rect 7837 3383 7895 3389
rect 7837 3380 7849 3383
rect 6788 3352 7849 3380
rect 6788 3340 6794 3352
rect 7837 3349 7849 3352
rect 7883 3349 7895 3383
rect 7837 3343 7895 3349
rect 8573 3383 8631 3389
rect 8573 3349 8585 3383
rect 8619 3380 8631 3383
rect 8662 3380 8668 3392
rect 8619 3352 8668 3380
rect 8619 3349 8631 3352
rect 8573 3343 8631 3349
rect 8662 3340 8668 3352
rect 8720 3340 8726 3392
rect 8772 3380 8800 3420
rect 9674 3408 9680 3420
rect 9732 3408 9738 3460
rect 10428 3448 10456 3479
rect 10594 3476 10600 3488
rect 10652 3476 10658 3528
rect 11330 3476 11336 3528
rect 11388 3516 11394 3528
rect 11885 3519 11943 3525
rect 11885 3516 11897 3519
rect 11388 3488 11897 3516
rect 11388 3476 11394 3488
rect 11885 3485 11897 3488
rect 11931 3485 11943 3519
rect 11885 3479 11943 3485
rect 12069 3519 12127 3525
rect 12069 3485 12081 3519
rect 12115 3516 12127 3519
rect 13004 3516 13032 3556
rect 13722 3544 13728 3556
rect 13780 3584 13786 3596
rect 14182 3584 14188 3596
rect 13780 3556 14188 3584
rect 13780 3544 13786 3556
rect 14182 3544 14188 3556
rect 14240 3544 14246 3596
rect 12115 3488 13032 3516
rect 13081 3519 13139 3525
rect 12115 3485 12127 3488
rect 12069 3479 12127 3485
rect 13081 3485 13093 3519
rect 13127 3516 13139 3519
rect 13170 3516 13176 3528
rect 13127 3488 13176 3516
rect 13127 3485 13139 3488
rect 13081 3479 13139 3485
rect 13170 3476 13176 3488
rect 13228 3476 13234 3528
rect 13262 3476 13268 3528
rect 13320 3516 13326 3528
rect 14001 3519 14059 3525
rect 14001 3516 14013 3519
rect 13320 3488 14013 3516
rect 13320 3476 13326 3488
rect 14001 3485 14013 3488
rect 14047 3485 14059 3519
rect 14001 3479 14059 3485
rect 10502 3448 10508 3460
rect 10428 3420 10508 3448
rect 10502 3408 10508 3420
rect 10560 3408 10566 3460
rect 12437 3451 12495 3457
rect 12437 3417 12449 3451
rect 12483 3448 12495 3451
rect 12894 3448 12900 3460
rect 12483 3420 12900 3448
rect 12483 3417 12495 3420
rect 12437 3411 12495 3417
rect 12894 3408 12900 3420
rect 12952 3408 12958 3460
rect 9490 3380 9496 3392
rect 8772 3352 9496 3380
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 9950 3380 9956 3392
rect 9911 3352 9956 3380
rect 9950 3340 9956 3352
rect 10008 3340 10014 3392
rect 10042 3340 10048 3392
rect 10100 3380 10106 3392
rect 13449 3383 13507 3389
rect 13449 3380 13461 3383
rect 10100 3352 13461 3380
rect 10100 3340 10106 3352
rect 13449 3349 13461 3352
rect 13495 3349 13507 3383
rect 13449 3343 13507 3349
rect 1104 3290 15824 3312
rect 1104 3238 3447 3290
rect 3499 3238 3511 3290
rect 3563 3238 3575 3290
rect 3627 3238 3639 3290
rect 3691 3238 8378 3290
rect 8430 3238 8442 3290
rect 8494 3238 8506 3290
rect 8558 3238 8570 3290
rect 8622 3238 13308 3290
rect 13360 3238 13372 3290
rect 13424 3238 13436 3290
rect 13488 3238 13500 3290
rect 13552 3238 15824 3290
rect 1104 3216 15824 3238
rect 2222 3176 2228 3188
rect 2183 3148 2228 3176
rect 2222 3136 2228 3148
rect 2280 3136 2286 3188
rect 2682 3136 2688 3188
rect 2740 3176 2746 3188
rect 4798 3176 4804 3188
rect 2740 3148 4804 3176
rect 2740 3136 2746 3148
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 5166 3136 5172 3188
rect 5224 3176 5230 3188
rect 5721 3179 5779 3185
rect 5721 3176 5733 3179
rect 5224 3148 5733 3176
rect 5224 3136 5230 3148
rect 5721 3145 5733 3148
rect 5767 3145 5779 3179
rect 5721 3139 5779 3145
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 7834 3176 7840 3188
rect 5868 3148 7840 3176
rect 5868 3136 5874 3148
rect 7834 3136 7840 3148
rect 7892 3136 7898 3188
rect 8202 3136 8208 3188
rect 8260 3176 8266 3188
rect 9309 3179 9367 3185
rect 9309 3176 9321 3179
rect 8260 3148 9321 3176
rect 8260 3136 8266 3148
rect 9309 3145 9321 3148
rect 9355 3145 9367 3179
rect 9309 3139 9367 3145
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 10965 3179 11023 3185
rect 10965 3176 10977 3179
rect 9456 3148 10977 3176
rect 9456 3136 9462 3148
rect 10965 3145 10977 3148
rect 11011 3145 11023 3179
rect 11330 3176 11336 3188
rect 11291 3148 11336 3176
rect 10965 3139 11023 3145
rect 11330 3136 11336 3148
rect 11388 3136 11394 3188
rect 11790 3136 11796 3188
rect 11848 3176 11854 3188
rect 12250 3176 12256 3188
rect 11848 3148 12256 3176
rect 11848 3136 11854 3148
rect 12250 3136 12256 3148
rect 12308 3136 12314 3188
rect 14182 3136 14188 3188
rect 14240 3176 14246 3188
rect 14277 3179 14335 3185
rect 14277 3176 14289 3179
rect 14240 3148 14289 3176
rect 14240 3136 14246 3148
rect 14277 3145 14289 3148
rect 14323 3145 14335 3179
rect 14277 3139 14335 3145
rect 4706 3108 4712 3120
rect 2700 3080 4712 3108
rect 1670 3040 1676 3052
rect 1631 3012 1676 3040
rect 1670 3000 1676 3012
rect 1728 3000 1734 3052
rect 2700 3049 2728 3080
rect 4706 3068 4712 3080
rect 4764 3068 4770 3120
rect 12526 3068 12532 3120
rect 12584 3108 12590 3120
rect 12584 3080 12940 3108
rect 12584 3068 12590 3080
rect 2685 3043 2743 3049
rect 2685 3009 2697 3043
rect 2731 3009 2743 3043
rect 2685 3003 2743 3009
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3040 2927 3043
rect 3326 3040 3332 3052
rect 2915 3012 3332 3040
rect 2915 3009 2927 3012
rect 2869 3003 2927 3009
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 3418 3000 3424 3052
rect 3476 3040 3482 3052
rect 3789 3043 3847 3049
rect 3789 3040 3801 3043
rect 3476 3012 3801 3040
rect 3476 3000 3482 3012
rect 3789 3009 3801 3012
rect 3835 3040 3847 3043
rect 4338 3040 4344 3052
rect 3835 3012 4344 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 4338 3000 4344 3012
rect 4396 3000 4402 3052
rect 4893 3043 4951 3049
rect 4893 3009 4905 3043
rect 4939 3040 4951 3043
rect 4982 3040 4988 3052
rect 4939 3012 4988 3040
rect 4939 3009 4951 3012
rect 4893 3003 4951 3009
rect 4982 3000 4988 3012
rect 5040 3000 5046 3052
rect 5166 3000 5172 3052
rect 5224 3040 5230 3052
rect 5626 3040 5632 3052
rect 5224 3012 5632 3040
rect 5224 3000 5230 3012
rect 5626 3000 5632 3012
rect 5684 3000 5690 3052
rect 6362 3040 6368 3052
rect 6323 3012 6368 3040
rect 6362 3000 6368 3012
rect 6420 3000 6426 3052
rect 7190 3000 7196 3052
rect 7248 3040 7254 3052
rect 7377 3043 7435 3049
rect 7377 3040 7389 3043
rect 7248 3012 7389 3040
rect 7248 3000 7254 3012
rect 7377 3009 7389 3012
rect 7423 3009 7435 3043
rect 7926 3040 7932 3052
rect 7887 3012 7932 3040
rect 7377 3003 7435 3009
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 9490 3000 9496 3052
rect 9548 3040 9554 3052
rect 9585 3043 9643 3049
rect 9585 3040 9597 3043
rect 9548 3012 9597 3040
rect 9548 3000 9554 3012
rect 9585 3009 9597 3012
rect 9631 3009 9643 3043
rect 9585 3003 9643 3009
rect 11698 3000 11704 3052
rect 11756 3040 11762 3052
rect 11885 3043 11943 3049
rect 11885 3040 11897 3043
rect 11756 3012 11897 3040
rect 11756 3000 11762 3012
rect 11885 3009 11897 3012
rect 11931 3009 11943 3043
rect 11885 3003 11943 3009
rect 12434 3000 12440 3052
rect 12492 3040 12498 3052
rect 12912 3049 12940 3080
rect 12897 3043 12955 3049
rect 12492 3012 12537 3040
rect 12492 3000 12498 3012
rect 12897 3009 12909 3043
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 14642 3000 14648 3052
rect 14700 3040 14706 3052
rect 14700 3012 14872 3040
rect 14700 3000 14706 3012
rect 1489 2975 1547 2981
rect 1489 2941 1501 2975
rect 1535 2972 1547 2975
rect 2038 2972 2044 2984
rect 1535 2944 2044 2972
rect 1535 2941 1547 2944
rect 1489 2935 1547 2941
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 2222 2932 2228 2984
rect 2280 2972 2286 2984
rect 4246 2972 4252 2984
rect 2280 2944 4252 2972
rect 2280 2932 2286 2944
rect 4246 2932 4252 2944
rect 4304 2932 4310 2984
rect 4617 2975 4675 2981
rect 4617 2941 4629 2975
rect 4663 2972 4675 2975
rect 4706 2972 4712 2984
rect 4663 2944 4712 2972
rect 4663 2941 4675 2944
rect 4617 2935 4675 2941
rect 4706 2932 4712 2944
rect 4764 2932 4770 2984
rect 6638 2932 6644 2984
rect 6696 2972 6702 2984
rect 8196 2975 8254 2981
rect 6696 2944 7236 2972
rect 6696 2932 6702 2944
rect 2593 2907 2651 2913
rect 2593 2873 2605 2907
rect 2639 2904 2651 2907
rect 3605 2907 3663 2913
rect 2639 2876 3280 2904
rect 2639 2873 2651 2876
rect 2593 2867 2651 2873
rect 1486 2796 1492 2848
rect 1544 2836 1550 2848
rect 2958 2836 2964 2848
rect 1544 2808 2964 2836
rect 1544 2796 1550 2808
rect 2958 2796 2964 2808
rect 3016 2796 3022 2848
rect 3252 2845 3280 2876
rect 3605 2873 3617 2907
rect 3651 2904 3663 2907
rect 4338 2904 4344 2916
rect 3651 2876 4344 2904
rect 3651 2873 3663 2876
rect 3605 2867 3663 2873
rect 4338 2864 4344 2876
rect 4396 2864 4402 2916
rect 4430 2864 4436 2916
rect 4488 2904 4494 2916
rect 7208 2913 7236 2944
rect 8196 2941 8208 2975
rect 8242 2972 8254 2975
rect 9306 2972 9312 2984
rect 8242 2944 9312 2972
rect 8242 2941 8254 2944
rect 8196 2935 8254 2941
rect 9306 2932 9312 2944
rect 9364 2932 9370 2984
rect 12526 2972 12532 2984
rect 9692 2944 12532 2972
rect 7193 2907 7251 2913
rect 4488 2876 6960 2904
rect 4488 2864 4494 2876
rect 3237 2839 3295 2845
rect 3237 2805 3249 2839
rect 3283 2805 3295 2839
rect 3237 2799 3295 2805
rect 3697 2839 3755 2845
rect 3697 2805 3709 2839
rect 3743 2836 3755 2839
rect 4249 2839 4307 2845
rect 4249 2836 4261 2839
rect 3743 2808 4261 2836
rect 3743 2805 3755 2808
rect 3697 2799 3755 2805
rect 4249 2805 4261 2808
rect 4295 2805 4307 2839
rect 4249 2799 4307 2805
rect 4709 2839 4767 2845
rect 4709 2805 4721 2839
rect 4755 2836 4767 2839
rect 5074 2836 5080 2848
rect 4755 2808 5080 2836
rect 4755 2805 4767 2808
rect 4709 2799 4767 2805
rect 5074 2796 5080 2808
rect 5132 2796 5138 2848
rect 5258 2836 5264 2848
rect 5219 2808 5264 2836
rect 5258 2796 5264 2808
rect 5316 2796 5322 2848
rect 5810 2796 5816 2848
rect 5868 2836 5874 2848
rect 6089 2839 6147 2845
rect 6089 2836 6101 2839
rect 5868 2808 6101 2836
rect 5868 2796 5874 2808
rect 6089 2805 6101 2808
rect 6135 2805 6147 2839
rect 6089 2799 6147 2805
rect 6181 2839 6239 2845
rect 6181 2805 6193 2839
rect 6227 2836 6239 2839
rect 6825 2839 6883 2845
rect 6825 2836 6837 2839
rect 6227 2808 6837 2836
rect 6227 2805 6239 2808
rect 6181 2799 6239 2805
rect 6825 2805 6837 2808
rect 6871 2805 6883 2839
rect 6932 2836 6960 2876
rect 7193 2873 7205 2907
rect 7239 2873 7251 2907
rect 7193 2867 7251 2873
rect 7285 2907 7343 2913
rect 7285 2873 7297 2907
rect 7331 2904 7343 2907
rect 7926 2904 7932 2916
rect 7331 2876 7932 2904
rect 7331 2873 7343 2876
rect 7285 2867 7343 2873
rect 7926 2864 7932 2876
rect 7984 2864 7990 2916
rect 8018 2864 8024 2916
rect 8076 2904 8082 2916
rect 9692 2904 9720 2944
rect 12526 2932 12532 2944
rect 12584 2932 12590 2984
rect 14844 2981 14872 3012
rect 14829 2975 14887 2981
rect 14829 2941 14841 2975
rect 14875 2941 14887 2975
rect 14829 2935 14887 2941
rect 8076 2876 9720 2904
rect 9852 2907 9910 2913
rect 8076 2864 8082 2876
rect 9852 2873 9864 2907
rect 9898 2904 9910 2907
rect 10410 2904 10416 2916
rect 9898 2876 10416 2904
rect 9898 2873 9910 2876
rect 9852 2867 9910 2873
rect 10410 2864 10416 2876
rect 10468 2864 10474 2916
rect 10594 2864 10600 2916
rect 10652 2904 10658 2916
rect 13170 2913 13176 2916
rect 11701 2907 11759 2913
rect 11701 2904 11713 2907
rect 10652 2876 11713 2904
rect 10652 2864 10658 2876
rect 11701 2873 11713 2876
rect 11747 2873 11759 2907
rect 13164 2904 13176 2913
rect 13131 2876 13176 2904
rect 11701 2867 11759 2873
rect 13164 2867 13176 2876
rect 13170 2864 13176 2867
rect 13228 2864 13234 2916
rect 11146 2836 11152 2848
rect 6932 2808 11152 2836
rect 6825 2799 6883 2805
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 11422 2796 11428 2848
rect 11480 2836 11486 2848
rect 11793 2839 11851 2845
rect 11793 2836 11805 2839
rect 11480 2808 11805 2836
rect 11480 2796 11486 2808
rect 11793 2805 11805 2808
rect 11839 2805 11851 2839
rect 11793 2799 11851 2805
rect 14734 2796 14740 2848
rect 14792 2836 14798 2848
rect 14844 2836 14872 2935
rect 15105 2907 15163 2913
rect 15105 2873 15117 2907
rect 15151 2904 15163 2907
rect 16758 2904 16764 2916
rect 15151 2876 16764 2904
rect 15151 2873 15163 2876
rect 15105 2867 15163 2873
rect 16758 2864 16764 2876
rect 16816 2864 16822 2916
rect 14792 2808 14872 2836
rect 14792 2796 14798 2808
rect 1104 2746 15824 2768
rect 1104 2694 5912 2746
rect 5964 2694 5976 2746
rect 6028 2694 6040 2746
rect 6092 2694 6104 2746
rect 6156 2694 10843 2746
rect 10895 2694 10907 2746
rect 10959 2694 10971 2746
rect 11023 2694 11035 2746
rect 11087 2694 15824 2746
rect 1104 2672 15824 2694
rect 4338 2632 4344 2644
rect 4299 2604 4344 2632
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 4801 2635 4859 2641
rect 4801 2601 4813 2635
rect 4847 2632 4859 2635
rect 4890 2632 4896 2644
rect 4847 2604 4896 2632
rect 4847 2601 4859 2604
rect 4801 2595 4859 2601
rect 4890 2592 4896 2604
rect 4948 2592 4954 2644
rect 5442 2632 5448 2644
rect 5403 2604 5448 2632
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 5905 2635 5963 2641
rect 5905 2601 5917 2635
rect 5951 2632 5963 2635
rect 6914 2632 6920 2644
rect 5951 2604 6920 2632
rect 5951 2601 5963 2604
rect 5905 2595 5963 2601
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 7098 2632 7104 2644
rect 7059 2604 7104 2632
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 8665 2635 8723 2641
rect 8665 2632 8677 2635
rect 8067 2604 8677 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 8665 2601 8677 2604
rect 8711 2601 8723 2635
rect 9766 2632 9772 2644
rect 9727 2604 9772 2632
rect 8665 2595 8723 2601
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 9950 2592 9956 2644
rect 10008 2632 10014 2644
rect 10229 2635 10287 2641
rect 10229 2632 10241 2635
rect 10008 2604 10241 2632
rect 10008 2592 10014 2604
rect 10229 2601 10241 2604
rect 10275 2601 10287 2635
rect 10229 2595 10287 2601
rect 11146 2592 11152 2644
rect 11204 2632 11210 2644
rect 12069 2635 12127 2641
rect 12069 2632 12081 2635
rect 11204 2604 12081 2632
rect 11204 2592 11210 2604
rect 12069 2601 12081 2604
rect 12115 2601 12127 2635
rect 12618 2632 12624 2644
rect 12579 2604 12624 2632
rect 12069 2595 12127 2601
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 12986 2592 12992 2644
rect 13044 2632 13050 2644
rect 13081 2635 13139 2641
rect 13081 2632 13093 2635
rect 13044 2604 13093 2632
rect 13044 2592 13050 2604
rect 13081 2601 13093 2604
rect 13127 2601 13139 2635
rect 13081 2595 13139 2601
rect 13817 2635 13875 2641
rect 13817 2601 13829 2635
rect 13863 2632 13875 2635
rect 13906 2632 13912 2644
rect 13863 2604 13912 2632
rect 13863 2601 13875 2604
rect 13817 2595 13875 2601
rect 13906 2592 13912 2604
rect 13964 2592 13970 2644
rect 14366 2632 14372 2644
rect 14327 2604 14372 2632
rect 14366 2592 14372 2604
rect 14424 2592 14430 2644
rect 2498 2564 2504 2576
rect 1504 2536 2504 2564
rect 1504 2505 1532 2536
rect 2498 2524 2504 2536
rect 2556 2524 2562 2576
rect 4709 2567 4767 2573
rect 4709 2533 4721 2567
rect 4755 2564 4767 2567
rect 5258 2564 5264 2576
rect 4755 2536 5264 2564
rect 4755 2533 4767 2536
rect 4709 2527 4767 2533
rect 5258 2524 5264 2536
rect 5316 2524 5322 2576
rect 7558 2564 7564 2576
rect 6932 2536 7564 2564
rect 1489 2499 1547 2505
rect 1489 2465 1501 2499
rect 1535 2465 1547 2499
rect 1489 2459 1547 2465
rect 1946 2456 1952 2508
rect 2004 2496 2010 2508
rect 2041 2499 2099 2505
rect 2041 2496 2053 2499
rect 2004 2468 2053 2496
rect 2004 2456 2010 2468
rect 2041 2465 2053 2468
rect 2087 2465 2099 2499
rect 2041 2459 2099 2465
rect 2308 2499 2366 2505
rect 2308 2465 2320 2499
rect 2354 2496 2366 2499
rect 2774 2496 2780 2508
rect 2354 2468 2780 2496
rect 2354 2465 2366 2468
rect 2308 2459 2366 2465
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 6932 2505 6960 2536
rect 7558 2524 7564 2536
rect 7616 2564 7622 2576
rect 9033 2567 9091 2573
rect 7616 2536 8800 2564
rect 7616 2524 7622 2536
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2496 5871 2499
rect 6917 2499 6975 2505
rect 5859 2468 6868 2496
rect 5859 2465 5871 2468
rect 5813 2459 5871 2465
rect 4982 2428 4988 2440
rect 4895 2400 4988 2428
rect 4982 2388 4988 2400
rect 5040 2428 5046 2440
rect 6089 2431 6147 2437
rect 6089 2428 6101 2431
rect 5040 2400 6101 2428
rect 5040 2388 5046 2400
rect 6089 2397 6101 2400
rect 6135 2428 6147 2431
rect 6638 2428 6644 2440
rect 6135 2400 6644 2428
rect 6135 2397 6147 2400
rect 6089 2391 6147 2397
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 6840 2428 6868 2468
rect 6917 2465 6929 2499
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 8113 2499 8171 2505
rect 8113 2465 8125 2499
rect 8159 2496 8171 2499
rect 8662 2496 8668 2508
rect 8159 2468 8668 2496
rect 8159 2465 8171 2468
rect 8113 2459 8171 2465
rect 8662 2456 8668 2468
rect 8720 2456 8726 2508
rect 8772 2496 8800 2536
rect 9033 2533 9045 2567
rect 9079 2564 9091 2567
rect 10042 2564 10048 2576
rect 9079 2536 10048 2564
rect 9079 2533 9091 2536
rect 9033 2527 9091 2533
rect 10042 2524 10048 2536
rect 10100 2524 10106 2576
rect 10137 2567 10195 2573
rect 10137 2533 10149 2567
rect 10183 2564 10195 2567
rect 11054 2564 11060 2576
rect 10183 2536 11060 2564
rect 10183 2533 10195 2536
rect 10137 2527 10195 2533
rect 11054 2524 11060 2536
rect 11112 2524 11118 2576
rect 11333 2567 11391 2573
rect 11333 2533 11345 2567
rect 11379 2564 11391 2567
rect 14918 2564 14924 2576
rect 11379 2536 13676 2564
rect 11379 2533 11391 2536
rect 11333 2527 11391 2533
rect 13648 2508 13676 2536
rect 14200 2536 14924 2564
rect 10594 2496 10600 2508
rect 8772 2468 9444 2496
rect 6840 2400 7788 2428
rect 7653 2363 7711 2369
rect 7653 2360 7665 2363
rect 3160 2332 7665 2360
rect 198 2252 204 2304
rect 256 2292 262 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 256 2264 1685 2292
rect 256 2252 262 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 2038 2252 2044 2304
rect 2096 2292 2102 2304
rect 3160 2292 3188 2332
rect 7653 2329 7665 2332
rect 7699 2329 7711 2363
rect 7653 2323 7711 2329
rect 2096 2264 3188 2292
rect 3421 2295 3479 2301
rect 2096 2252 2102 2264
rect 3421 2261 3433 2295
rect 3467 2292 3479 2295
rect 7558 2292 7564 2304
rect 3467 2264 7564 2292
rect 3467 2261 3479 2264
rect 3421 2255 3479 2261
rect 7558 2252 7564 2264
rect 7616 2252 7622 2304
rect 7760 2292 7788 2400
rect 8202 2388 8208 2440
rect 8260 2428 8266 2440
rect 9125 2431 9183 2437
rect 8260 2400 8305 2428
rect 8260 2388 8266 2400
rect 9125 2397 9137 2431
rect 9171 2397 9183 2431
rect 9306 2428 9312 2440
rect 9267 2400 9312 2428
rect 9125 2391 9183 2397
rect 9140 2360 9168 2391
rect 9306 2388 9312 2400
rect 9364 2388 9370 2440
rect 9416 2428 9444 2468
rect 10244 2468 10600 2496
rect 10244 2428 10272 2468
rect 10594 2456 10600 2468
rect 10652 2456 10658 2508
rect 11241 2499 11299 2505
rect 11241 2465 11253 2499
rect 11287 2496 11299 2499
rect 11885 2499 11943 2505
rect 11287 2468 11836 2496
rect 11287 2465 11299 2468
rect 11241 2459 11299 2465
rect 10410 2428 10416 2440
rect 9416 2400 10272 2428
rect 10323 2400 10416 2428
rect 10410 2388 10416 2400
rect 10468 2428 10474 2440
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 10468 2400 11529 2428
rect 10468 2388 10474 2400
rect 11517 2397 11529 2400
rect 11563 2428 11575 2431
rect 11606 2428 11612 2440
rect 11563 2400 11612 2428
rect 11563 2397 11575 2400
rect 11517 2391 11575 2397
rect 11606 2388 11612 2400
rect 11664 2388 11670 2440
rect 11808 2428 11836 2468
rect 11885 2465 11897 2499
rect 11931 2496 11943 2499
rect 12066 2496 12072 2508
rect 11931 2468 12072 2496
rect 11931 2465 11943 2468
rect 11885 2459 11943 2465
rect 12066 2456 12072 2468
rect 12124 2456 12130 2508
rect 12802 2456 12808 2508
rect 12860 2496 12866 2508
rect 12989 2499 13047 2505
rect 12989 2496 13001 2499
rect 12860 2468 13001 2496
rect 12860 2456 12866 2468
rect 12989 2465 13001 2468
rect 13035 2465 13047 2499
rect 13630 2496 13636 2508
rect 13591 2468 13636 2496
rect 12989 2459 13047 2465
rect 13630 2456 13636 2468
rect 13688 2456 13694 2508
rect 14200 2505 14228 2536
rect 14918 2524 14924 2536
rect 14976 2524 14982 2576
rect 14185 2499 14243 2505
rect 14185 2465 14197 2499
rect 14231 2465 14243 2499
rect 14185 2459 14243 2465
rect 14550 2456 14556 2508
rect 14608 2496 14614 2508
rect 14737 2499 14795 2505
rect 14737 2496 14749 2499
rect 14608 2468 14749 2496
rect 14608 2456 14614 2468
rect 14737 2465 14749 2468
rect 14783 2465 14795 2499
rect 14737 2459 14795 2465
rect 11974 2428 11980 2440
rect 11808 2400 11980 2428
rect 11974 2388 11980 2400
rect 12032 2388 12038 2440
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 13170 2428 13176 2440
rect 12308 2400 13176 2428
rect 12308 2388 12314 2400
rect 13170 2388 13176 2400
rect 13228 2388 13234 2440
rect 10873 2363 10931 2369
rect 10873 2360 10885 2363
rect 9140 2332 10885 2360
rect 10873 2329 10885 2332
rect 10919 2329 10931 2363
rect 10873 2323 10931 2329
rect 9490 2292 9496 2304
rect 7760 2264 9496 2292
rect 9490 2252 9496 2264
rect 9548 2292 9554 2304
rect 11330 2292 11336 2304
rect 9548 2264 11336 2292
rect 9548 2252 9554 2264
rect 11330 2252 11336 2264
rect 11388 2252 11394 2304
rect 11992 2292 12020 2388
rect 15470 2360 15476 2372
rect 12452 2332 15476 2360
rect 12452 2292 12480 2332
rect 15470 2320 15476 2332
rect 15528 2320 15534 2372
rect 11992 2264 12480 2292
rect 12526 2252 12532 2304
rect 12584 2292 12590 2304
rect 14921 2295 14979 2301
rect 14921 2292 14933 2295
rect 12584 2264 14933 2292
rect 12584 2252 12590 2264
rect 14921 2261 14933 2264
rect 14967 2261 14979 2295
rect 14921 2255 14979 2261
rect 1104 2202 15824 2224
rect 1104 2150 3447 2202
rect 3499 2150 3511 2202
rect 3563 2150 3575 2202
rect 3627 2150 3639 2202
rect 3691 2150 8378 2202
rect 8430 2150 8442 2202
rect 8494 2150 8506 2202
rect 8558 2150 8570 2202
rect 8622 2150 13308 2202
rect 13360 2150 13372 2202
rect 13424 2150 13436 2202
rect 13488 2150 13500 2202
rect 13552 2150 15824 2202
rect 1104 2128 15824 2150
rect 11514 2048 11520 2100
rect 11572 2088 11578 2100
rect 12986 2088 12992 2100
rect 11572 2060 12992 2088
rect 11572 2048 11578 2060
rect 12986 2048 12992 2060
rect 13044 2048 13050 2100
rect 7558 1980 7564 2032
rect 7616 2020 7622 2032
rect 11698 2020 11704 2032
rect 7616 1992 11704 2020
rect 7616 1980 7622 1992
rect 11698 1980 11704 1992
rect 11756 2020 11762 2032
rect 12250 2020 12256 2032
rect 11756 1992 12256 2020
rect 11756 1980 11762 1992
rect 12250 1980 12256 1992
rect 12308 1980 12314 2032
rect 4062 1776 4068 1828
rect 4120 1816 4126 1828
rect 14734 1816 14740 1828
rect 4120 1788 14740 1816
rect 4120 1776 4126 1788
rect 14734 1776 14740 1788
rect 14792 1776 14798 1828
rect 1854 1096 1860 1148
rect 1912 1136 1918 1148
rect 7098 1136 7104 1148
rect 1912 1108 7104 1136
rect 1912 1096 1918 1108
rect 7098 1096 7104 1108
rect 7156 1096 7162 1148
<< via1 >>
rect 4068 17960 4120 18012
rect 14096 17960 14148 18012
rect 8944 17620 8996 17672
rect 9496 17620 9548 17672
rect 5356 17552 5408 17604
rect 11520 17552 11572 17604
rect 204 17484 256 17536
rect 14188 17484 14240 17536
rect 3447 17382 3499 17434
rect 3511 17382 3563 17434
rect 3575 17382 3627 17434
rect 3639 17382 3691 17434
rect 8378 17382 8430 17434
rect 8442 17382 8494 17434
rect 8506 17382 8558 17434
rect 8570 17382 8622 17434
rect 13308 17382 13360 17434
rect 13372 17382 13424 17434
rect 13436 17382 13488 17434
rect 13500 17382 13552 17434
rect 2780 17280 2832 17332
rect 4620 17280 4672 17332
rect 5080 17280 5132 17332
rect 5632 17280 5684 17332
rect 7840 17280 7892 17332
rect 2872 17212 2924 17264
rect 2964 17212 3016 17264
rect 5816 17212 5868 17264
rect 12716 17280 12768 17332
rect 1584 17119 1636 17128
rect 1584 17085 1593 17119
rect 1593 17085 1627 17119
rect 1627 17085 1636 17119
rect 1584 17076 1636 17085
rect 3884 17076 3936 17128
rect 5356 17119 5408 17128
rect 4160 17008 4212 17060
rect 5356 17085 5365 17119
rect 5365 17085 5399 17119
rect 5399 17085 5408 17119
rect 5356 17076 5408 17085
rect 6828 17076 6880 17128
rect 13728 17212 13780 17264
rect 8392 17144 8444 17196
rect 11244 17144 11296 17196
rect 11612 17144 11664 17196
rect 13176 17187 13228 17196
rect 13176 17153 13185 17187
rect 13185 17153 13219 17187
rect 13219 17153 13228 17187
rect 13176 17144 13228 17153
rect 14096 17187 14148 17196
rect 14096 17153 14105 17187
rect 14105 17153 14139 17187
rect 14139 17153 14148 17187
rect 14096 17144 14148 17153
rect 15108 17187 15160 17196
rect 15108 17153 15117 17187
rect 15117 17153 15151 17187
rect 15151 17153 15160 17187
rect 15108 17144 15160 17153
rect 6552 17008 6604 17060
rect 10232 17076 10284 17128
rect 12440 17076 12492 17128
rect 2872 16940 2924 16992
rect 8300 16940 8352 16992
rect 8668 16983 8720 16992
rect 8668 16949 8677 16983
rect 8677 16949 8711 16983
rect 8711 16949 8720 16983
rect 8668 16940 8720 16949
rect 9036 16983 9088 16992
rect 9036 16949 9045 16983
rect 9045 16949 9079 16983
rect 9079 16949 9088 16983
rect 9036 16940 9088 16949
rect 9128 16983 9180 16992
rect 9128 16949 9137 16983
rect 9137 16949 9171 16983
rect 9171 16949 9180 16983
rect 9128 16940 9180 16949
rect 11152 16983 11204 16992
rect 11152 16949 11161 16983
rect 11161 16949 11195 16983
rect 11195 16949 11204 16983
rect 15016 17008 15068 17060
rect 11152 16940 11204 16949
rect 12992 16983 13044 16992
rect 12992 16949 13001 16983
rect 13001 16949 13035 16983
rect 13035 16949 13044 16983
rect 12992 16940 13044 16949
rect 13912 16940 13964 16992
rect 5912 16838 5964 16890
rect 5976 16838 6028 16890
rect 6040 16838 6092 16890
rect 6104 16838 6156 16890
rect 10843 16838 10895 16890
rect 10907 16838 10959 16890
rect 10971 16838 11023 16890
rect 11035 16838 11087 16890
rect 940 16736 992 16788
rect 1400 16668 1452 16720
rect 4252 16736 4304 16788
rect 8392 16779 8444 16788
rect 3148 16711 3200 16720
rect 3148 16677 3157 16711
rect 3157 16677 3191 16711
rect 3191 16677 3200 16711
rect 3148 16668 3200 16677
rect 5724 16668 5776 16720
rect 6368 16668 6420 16720
rect 8392 16745 8401 16779
rect 8401 16745 8435 16779
rect 8435 16745 8444 16779
rect 8392 16736 8444 16745
rect 8668 16736 8720 16788
rect 11152 16736 11204 16788
rect 12624 16736 12676 16788
rect 13084 16736 13136 16788
rect 13176 16736 13228 16788
rect 8300 16668 8352 16720
rect 9496 16668 9548 16720
rect 1676 16600 1728 16652
rect 2504 16600 2556 16652
rect 2872 16643 2924 16652
rect 2872 16609 2881 16643
rect 2881 16609 2915 16643
rect 2915 16609 2924 16643
rect 2872 16600 2924 16609
rect 6736 16600 6788 16652
rect 5356 16396 5408 16448
rect 11796 16668 11848 16720
rect 11428 16643 11480 16652
rect 8116 16532 8168 16584
rect 8024 16464 8076 16516
rect 8944 16464 8996 16516
rect 9588 16532 9640 16584
rect 11428 16609 11437 16643
rect 11437 16609 11471 16643
rect 11471 16609 11480 16643
rect 11428 16600 11480 16609
rect 14004 16600 14056 16652
rect 14188 16643 14240 16652
rect 14188 16609 14197 16643
rect 14197 16609 14231 16643
rect 14231 16609 14240 16643
rect 14188 16600 14240 16609
rect 14832 16600 14884 16652
rect 11704 16575 11756 16584
rect 11704 16541 11713 16575
rect 11713 16541 11747 16575
rect 11747 16541 11756 16575
rect 11704 16532 11756 16541
rect 11980 16532 12032 16584
rect 15016 16532 15068 16584
rect 11336 16464 11388 16516
rect 7656 16396 7708 16448
rect 9772 16396 9824 16448
rect 10600 16396 10652 16448
rect 15200 16396 15252 16448
rect 15936 16396 15988 16448
rect 3447 16294 3499 16346
rect 3511 16294 3563 16346
rect 3575 16294 3627 16346
rect 3639 16294 3691 16346
rect 8378 16294 8430 16346
rect 8442 16294 8494 16346
rect 8506 16294 8558 16346
rect 8570 16294 8622 16346
rect 13308 16294 13360 16346
rect 13372 16294 13424 16346
rect 13436 16294 13488 16346
rect 13500 16294 13552 16346
rect 1860 16192 1912 16244
rect 3332 16192 3384 16244
rect 3792 16192 3844 16244
rect 6276 16192 6328 16244
rect 7012 16192 7064 16244
rect 9036 16192 9088 16244
rect 11428 16192 11480 16244
rect 12440 16235 12492 16244
rect 12440 16201 12449 16235
rect 12449 16201 12483 16235
rect 12483 16201 12492 16235
rect 12440 16192 12492 16201
rect 2228 16124 2280 16176
rect 6460 16124 6512 16176
rect 8116 16124 8168 16176
rect 1768 16099 1820 16108
rect 1768 16065 1777 16099
rect 1777 16065 1811 16099
rect 1811 16065 1820 16099
rect 1768 16056 1820 16065
rect 2320 16031 2372 16040
rect 2320 15997 2329 16031
rect 2329 15997 2363 16031
rect 2363 15997 2372 16031
rect 2320 15988 2372 15997
rect 5540 16056 5592 16108
rect 6368 16099 6420 16108
rect 6368 16065 6377 16099
rect 6377 16065 6411 16099
rect 6411 16065 6420 16099
rect 6368 16056 6420 16065
rect 7656 16056 7708 16108
rect 11704 16056 11756 16108
rect 3332 15988 3384 16040
rect 3792 15988 3844 16040
rect 5172 16031 5224 16040
rect 5172 15997 5181 16031
rect 5181 15997 5215 16031
rect 5215 15997 5224 16031
rect 5172 15988 5224 15997
rect 7840 16031 7892 16040
rect 7840 15997 7849 16031
rect 7849 15997 7883 16031
rect 7883 15997 7892 16031
rect 7840 15988 7892 15997
rect 8392 16031 8444 16040
rect 8392 15997 8401 16031
rect 8401 15997 8435 16031
rect 8435 15997 8444 16031
rect 8392 15988 8444 15997
rect 8668 16031 8720 16040
rect 8668 15997 8702 16031
rect 8702 15997 8720 16031
rect 8668 15988 8720 15997
rect 9128 15988 9180 16040
rect 2780 15920 2832 15972
rect 2596 15852 2648 15904
rect 9588 15920 9640 15972
rect 7012 15852 7064 15904
rect 7288 15895 7340 15904
rect 7288 15861 7297 15895
rect 7297 15861 7331 15895
rect 7331 15861 7340 15895
rect 7288 15852 7340 15861
rect 8392 15852 8444 15904
rect 10140 15920 10192 15972
rect 11980 15988 12032 16040
rect 11244 15920 11296 15972
rect 13544 15920 13596 15972
rect 11612 15852 11664 15904
rect 15292 15920 15344 15972
rect 16396 15920 16448 15972
rect 14832 15895 14884 15904
rect 14832 15861 14841 15895
rect 14841 15861 14875 15895
rect 14875 15861 14884 15895
rect 14832 15852 14884 15861
rect 14924 15852 14976 15904
rect 5912 15750 5964 15802
rect 5976 15750 6028 15802
rect 6040 15750 6092 15802
rect 6104 15750 6156 15802
rect 10843 15750 10895 15802
rect 10907 15750 10959 15802
rect 10971 15750 11023 15802
rect 11035 15750 11087 15802
rect 572 15648 624 15700
rect 6644 15648 6696 15700
rect 7012 15691 7064 15700
rect 7012 15657 7021 15691
rect 7021 15657 7055 15691
rect 7055 15657 7064 15691
rect 7012 15648 7064 15657
rect 7472 15691 7524 15700
rect 7472 15657 7481 15691
rect 7481 15657 7515 15691
rect 7515 15657 7524 15691
rect 7472 15648 7524 15657
rect 7932 15648 7984 15700
rect 10232 15648 10284 15700
rect 11244 15648 11296 15700
rect 1768 15623 1820 15632
rect 1768 15589 1777 15623
rect 1777 15589 1811 15623
rect 1811 15589 1820 15623
rect 1768 15580 1820 15589
rect 2596 15580 2648 15632
rect 3976 15580 4028 15632
rect 8392 15623 8444 15632
rect 3240 15512 3292 15564
rect 4344 15512 4396 15564
rect 5356 15512 5408 15564
rect 6368 15555 6420 15564
rect 6368 15521 6377 15555
rect 6377 15521 6411 15555
rect 6411 15521 6420 15555
rect 6368 15512 6420 15521
rect 6552 15512 6604 15564
rect 7196 15512 7248 15564
rect 8392 15589 8401 15623
rect 8401 15589 8435 15623
rect 8435 15589 8444 15623
rect 8392 15580 8444 15589
rect 12808 15648 12860 15700
rect 13176 15648 13228 15700
rect 13544 15648 13596 15700
rect 13912 15691 13964 15700
rect 13912 15657 13921 15691
rect 13921 15657 13955 15691
rect 13955 15657 13964 15691
rect 13912 15648 13964 15657
rect 15108 15648 15160 15700
rect 16764 15648 16816 15700
rect 13084 15580 13136 15632
rect 2780 15444 2832 15496
rect 2964 15444 3016 15496
rect 8116 15512 8168 15564
rect 8852 15512 8904 15564
rect 9036 15555 9088 15564
rect 9036 15521 9045 15555
rect 9045 15521 9079 15555
rect 9079 15521 9088 15555
rect 9036 15512 9088 15521
rect 9312 15512 9364 15564
rect 10048 15555 10100 15564
rect 10048 15521 10057 15555
rect 10057 15521 10091 15555
rect 10091 15521 10100 15555
rect 10048 15512 10100 15521
rect 10140 15512 10192 15564
rect 10968 15512 11020 15564
rect 11520 15512 11572 15564
rect 14280 15555 14332 15564
rect 14280 15521 14289 15555
rect 14289 15521 14323 15555
rect 14323 15521 14332 15555
rect 14280 15512 14332 15521
rect 8024 15444 8076 15496
rect 2780 15308 2832 15360
rect 5724 15376 5776 15428
rect 7656 15376 7708 15428
rect 10416 15444 10468 15496
rect 11704 15444 11756 15496
rect 11980 15444 12032 15496
rect 12164 15444 12216 15496
rect 14004 15444 14056 15496
rect 14556 15444 14608 15496
rect 8760 15376 8812 15428
rect 9588 15376 9640 15428
rect 11520 15308 11572 15360
rect 12256 15308 12308 15360
rect 3447 15206 3499 15258
rect 3511 15206 3563 15258
rect 3575 15206 3627 15258
rect 3639 15206 3691 15258
rect 8378 15206 8430 15258
rect 8442 15206 8494 15258
rect 8506 15206 8558 15258
rect 8570 15206 8622 15258
rect 13308 15206 13360 15258
rect 13372 15206 13424 15258
rect 13436 15206 13488 15258
rect 13500 15206 13552 15258
rect 4068 15147 4120 15156
rect 4068 15113 4077 15147
rect 4077 15113 4111 15147
rect 4111 15113 4120 15147
rect 4068 15104 4120 15113
rect 4344 15147 4396 15156
rect 4344 15113 4353 15147
rect 4353 15113 4387 15147
rect 4387 15113 4396 15147
rect 4344 15104 4396 15113
rect 5356 15104 5408 15156
rect 7288 15104 7340 15156
rect 8024 15104 8076 15156
rect 10048 15104 10100 15156
rect 10232 15104 10284 15156
rect 4528 14968 4580 15020
rect 5632 14968 5684 15020
rect 1492 14900 1544 14952
rect 2780 14832 2832 14884
rect 2964 14943 3016 14952
rect 2964 14909 2998 14943
rect 2998 14909 3016 14943
rect 4804 14943 4856 14952
rect 2964 14900 3016 14909
rect 4804 14909 4813 14943
rect 4813 14909 4847 14943
rect 4847 14909 4856 14943
rect 4804 14900 4856 14909
rect 6552 14943 6604 14952
rect 6552 14909 6561 14943
rect 6561 14909 6595 14943
rect 6595 14909 6604 14943
rect 6552 14900 6604 14909
rect 7748 14968 7800 15020
rect 8024 15011 8076 15020
rect 8024 14977 8033 15011
rect 8033 14977 8067 15011
rect 8067 14977 8076 15011
rect 8024 14968 8076 14977
rect 9680 14968 9732 15020
rect 10140 14968 10192 15020
rect 10600 15011 10652 15020
rect 10600 14977 10609 15011
rect 10609 14977 10643 15011
rect 10643 14977 10652 15011
rect 10600 14968 10652 14977
rect 12256 15104 12308 15156
rect 12992 15104 13044 15156
rect 14556 15104 14608 15156
rect 11612 14968 11664 15020
rect 12992 15011 13044 15020
rect 12992 14977 13001 15011
rect 13001 14977 13035 15011
rect 13035 14977 13044 15011
rect 12992 14968 13044 14977
rect 14096 15011 14148 15020
rect 14096 14977 14105 15011
rect 14105 14977 14139 15011
rect 14139 14977 14148 15011
rect 14096 14968 14148 14977
rect 5448 14832 5500 14884
rect 5540 14832 5592 14884
rect 7380 14900 7432 14952
rect 8576 14900 8628 14952
rect 11520 14943 11572 14952
rect 11520 14909 11529 14943
rect 11529 14909 11563 14943
rect 11563 14909 11572 14943
rect 11520 14900 11572 14909
rect 13728 14900 13780 14952
rect 8944 14832 8996 14884
rect 9772 14832 9824 14884
rect 1400 14764 1452 14816
rect 1952 14764 2004 14816
rect 4712 14807 4764 14816
rect 4712 14773 4721 14807
rect 4721 14773 4755 14807
rect 4755 14773 4764 14807
rect 4712 14764 4764 14773
rect 5356 14807 5408 14816
rect 5356 14773 5365 14807
rect 5365 14773 5399 14807
rect 5399 14773 5408 14807
rect 5356 14764 5408 14773
rect 5724 14807 5776 14816
rect 5724 14773 5733 14807
rect 5733 14773 5767 14807
rect 5767 14773 5776 14807
rect 5724 14764 5776 14773
rect 5816 14807 5868 14816
rect 5816 14773 5825 14807
rect 5825 14773 5859 14807
rect 5859 14773 5868 14807
rect 5816 14764 5868 14773
rect 7932 14807 7984 14816
rect 7932 14773 7941 14807
rect 7941 14773 7975 14807
rect 7975 14773 7984 14807
rect 7932 14764 7984 14773
rect 9588 14764 9640 14816
rect 10048 14764 10100 14816
rect 10324 14764 10376 14816
rect 13268 14764 13320 14816
rect 5912 14662 5964 14714
rect 5976 14662 6028 14714
rect 6040 14662 6092 14714
rect 6104 14662 6156 14714
rect 10843 14662 10895 14714
rect 10907 14662 10959 14714
rect 10971 14662 11023 14714
rect 11035 14662 11087 14714
rect 2964 14560 3016 14612
rect 5724 14560 5776 14612
rect 6276 14603 6328 14612
rect 6276 14569 6285 14603
rect 6285 14569 6319 14603
rect 6319 14569 6328 14603
rect 6276 14560 6328 14569
rect 7380 14560 7432 14612
rect 7932 14560 7984 14612
rect 3424 14535 3476 14544
rect 3424 14501 3433 14535
rect 3433 14501 3467 14535
rect 3467 14501 3476 14535
rect 3424 14492 3476 14501
rect 4068 14492 4120 14544
rect 8760 14560 8812 14612
rect 14648 14560 14700 14612
rect 1492 14467 1544 14476
rect 1492 14433 1501 14467
rect 1501 14433 1535 14467
rect 1535 14433 1544 14467
rect 1492 14424 1544 14433
rect 2688 14424 2740 14476
rect 10600 14492 10652 14544
rect 12992 14492 13044 14544
rect 14004 14535 14056 14544
rect 14004 14501 14013 14535
rect 14013 14501 14047 14535
rect 14047 14501 14056 14535
rect 14004 14492 14056 14501
rect 7012 14424 7064 14476
rect 7472 14424 7524 14476
rect 8116 14424 8168 14476
rect 9956 14424 10008 14476
rect 11612 14424 11664 14476
rect 4160 14399 4212 14408
rect 4160 14365 4169 14399
rect 4169 14365 4203 14399
rect 4203 14365 4212 14399
rect 4160 14356 4212 14365
rect 6184 14288 6236 14340
rect 3240 14220 3292 14272
rect 4344 14220 4396 14272
rect 5724 14220 5776 14272
rect 9128 14399 9180 14408
rect 9128 14365 9137 14399
rect 9137 14365 9171 14399
rect 9171 14365 9180 14399
rect 9128 14356 9180 14365
rect 8944 14288 8996 14340
rect 9036 14288 9088 14340
rect 10508 14220 10560 14272
rect 13728 14356 13780 14408
rect 10968 14220 11020 14272
rect 12992 14220 13044 14272
rect 14096 14220 14148 14272
rect 3447 14118 3499 14170
rect 3511 14118 3563 14170
rect 3575 14118 3627 14170
rect 3639 14118 3691 14170
rect 8378 14118 8430 14170
rect 8442 14118 8494 14170
rect 8506 14118 8558 14170
rect 8570 14118 8622 14170
rect 13308 14118 13360 14170
rect 13372 14118 13424 14170
rect 13436 14118 13488 14170
rect 13500 14118 13552 14170
rect 1952 14059 2004 14068
rect 1952 14025 1961 14059
rect 1961 14025 1995 14059
rect 1995 14025 2004 14059
rect 1952 14016 2004 14025
rect 3976 14059 4028 14068
rect 3976 14025 3985 14059
rect 3985 14025 4019 14059
rect 4019 14025 4028 14059
rect 3976 14016 4028 14025
rect 4160 14016 4212 14068
rect 5080 14016 5132 14068
rect 5816 14016 5868 14068
rect 5908 14016 5960 14068
rect 9680 14016 9732 14068
rect 9956 14016 10008 14068
rect 14004 14016 14056 14068
rect 2964 13880 3016 13932
rect 5264 13948 5316 14000
rect 5448 13948 5500 14000
rect 4528 13923 4580 13932
rect 2688 13812 2740 13864
rect 3240 13812 3292 13864
rect 4528 13889 4537 13923
rect 4537 13889 4571 13923
rect 4571 13889 4580 13923
rect 4528 13880 4580 13889
rect 4712 13880 4764 13932
rect 5724 13880 5776 13932
rect 6184 13923 6236 13932
rect 6184 13889 6193 13923
rect 6193 13889 6227 13923
rect 6227 13889 6236 13923
rect 6184 13880 6236 13889
rect 4896 13812 4948 13864
rect 5816 13812 5868 13864
rect 3332 13787 3384 13796
rect 3332 13753 3341 13787
rect 3341 13753 3375 13787
rect 3375 13753 3384 13787
rect 3332 13744 3384 13753
rect 4712 13744 4764 13796
rect 6368 13744 6420 13796
rect 8668 13812 8720 13864
rect 9036 13855 9088 13864
rect 9036 13821 9045 13855
rect 9045 13821 9079 13855
rect 9079 13821 9088 13855
rect 9036 13812 9088 13821
rect 9128 13812 9180 13864
rect 10508 13948 10560 14000
rect 12164 13948 12216 14000
rect 7196 13744 7248 13796
rect 8116 13744 8168 13796
rect 11612 13880 11664 13932
rect 14556 13948 14608 14000
rect 10232 13812 10284 13864
rect 12440 13812 12492 13864
rect 15016 13812 15068 13864
rect 12992 13744 13044 13796
rect 13544 13744 13596 13796
rect 14648 13744 14700 13796
rect 15568 13744 15620 13796
rect 2412 13719 2464 13728
rect 2412 13685 2421 13719
rect 2421 13685 2455 13719
rect 2455 13685 2464 13719
rect 2412 13676 2464 13685
rect 7472 13676 7524 13728
rect 11980 13676 12032 13728
rect 5912 13574 5964 13626
rect 5976 13574 6028 13626
rect 6040 13574 6092 13626
rect 6104 13574 6156 13626
rect 10843 13574 10895 13626
rect 10907 13574 10959 13626
rect 10971 13574 11023 13626
rect 11035 13574 11087 13626
rect 2412 13472 2464 13524
rect 5356 13472 5408 13524
rect 6460 13472 6512 13524
rect 8944 13515 8996 13524
rect 8944 13481 8953 13515
rect 8953 13481 8987 13515
rect 8987 13481 8996 13515
rect 8944 13472 8996 13481
rect 10232 13472 10284 13524
rect 11612 13472 11664 13524
rect 11980 13515 12032 13524
rect 11980 13481 11989 13515
rect 11989 13481 12023 13515
rect 12023 13481 12032 13515
rect 11980 13472 12032 13481
rect 2320 13404 2372 13456
rect 3884 13404 3936 13456
rect 1768 13336 1820 13388
rect 5356 13336 5408 13388
rect 2136 13311 2188 13320
rect 2136 13277 2145 13311
rect 2145 13277 2179 13311
rect 2179 13277 2188 13311
rect 2136 13268 2188 13277
rect 2228 13311 2280 13320
rect 2228 13277 2237 13311
rect 2237 13277 2271 13311
rect 2271 13277 2280 13311
rect 3148 13311 3200 13320
rect 2228 13268 2280 13277
rect 3148 13277 3157 13311
rect 3157 13277 3191 13311
rect 3191 13277 3200 13311
rect 3148 13268 3200 13277
rect 3240 13311 3292 13320
rect 3240 13277 3249 13311
rect 3249 13277 3283 13311
rect 3283 13277 3292 13311
rect 3240 13268 3292 13277
rect 5724 13268 5776 13320
rect 6276 13311 6328 13320
rect 6276 13277 6285 13311
rect 6285 13277 6319 13311
rect 6319 13277 6328 13311
rect 6276 13268 6328 13277
rect 5540 13200 5592 13252
rect 6644 13200 6696 13252
rect 7656 13336 7708 13388
rect 9128 13336 9180 13388
rect 9588 13404 9640 13456
rect 12532 13404 12584 13456
rect 14280 13472 14332 13524
rect 10416 13336 10468 13388
rect 10876 13336 10928 13388
rect 12256 13336 12308 13388
rect 12992 13336 13044 13388
rect 13728 13336 13780 13388
rect 1584 13132 1636 13184
rect 3976 13132 4028 13184
rect 4620 13175 4672 13184
rect 4620 13141 4629 13175
rect 4629 13141 4663 13175
rect 4663 13141 4672 13175
rect 4620 13132 4672 13141
rect 5816 13132 5868 13184
rect 9036 13132 9088 13184
rect 13084 13200 13136 13252
rect 13544 13311 13596 13320
rect 13544 13277 13553 13311
rect 13553 13277 13587 13311
rect 13587 13277 13596 13311
rect 13544 13268 13596 13277
rect 14004 13200 14056 13252
rect 14648 13132 14700 13184
rect 3447 13030 3499 13082
rect 3511 13030 3563 13082
rect 3575 13030 3627 13082
rect 3639 13030 3691 13082
rect 8378 13030 8430 13082
rect 8442 13030 8494 13082
rect 8506 13030 8558 13082
rect 8570 13030 8622 13082
rect 13308 13030 13360 13082
rect 13372 13030 13424 13082
rect 13436 13030 13488 13082
rect 13500 13030 13552 13082
rect 3148 12928 3200 12980
rect 3792 12928 3844 12980
rect 4068 12928 4120 12980
rect 4528 12971 4580 12980
rect 4528 12937 4537 12971
rect 4537 12937 4571 12971
rect 4571 12937 4580 12971
rect 4528 12928 4580 12937
rect 5356 12971 5408 12980
rect 5356 12937 5365 12971
rect 5365 12937 5399 12971
rect 5399 12937 5408 12971
rect 5356 12928 5408 12937
rect 10600 12928 10652 12980
rect 12440 12971 12492 12980
rect 12440 12937 12449 12971
rect 12449 12937 12483 12971
rect 12483 12937 12492 12971
rect 12440 12928 12492 12937
rect 12716 12928 12768 12980
rect 13176 12928 13228 12980
rect 5908 12860 5960 12912
rect 1584 12835 1636 12844
rect 1584 12801 1593 12835
rect 1593 12801 1627 12835
rect 1627 12801 1636 12835
rect 1584 12792 1636 12801
rect 1676 12792 1728 12844
rect 5816 12835 5868 12844
rect 5816 12801 5825 12835
rect 5825 12801 5859 12835
rect 5859 12801 5868 12835
rect 5816 12792 5868 12801
rect 6736 12860 6788 12912
rect 7932 12860 7984 12912
rect 7472 12792 7524 12844
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 2872 12724 2924 12776
rect 3240 12724 3292 12776
rect 6368 12724 6420 12776
rect 6644 12724 6696 12776
rect 6828 12724 6880 12776
rect 7196 12724 7248 12776
rect 8024 12767 8076 12776
rect 8024 12733 8033 12767
rect 8033 12733 8067 12767
rect 8067 12733 8076 12767
rect 8024 12724 8076 12733
rect 9036 12724 9088 12776
rect 8300 12699 8352 12708
rect 8300 12665 8334 12699
rect 8334 12665 8352 12699
rect 8300 12656 8352 12665
rect 4252 12588 4304 12640
rect 6552 12588 6604 12640
rect 6828 12631 6880 12640
rect 6828 12597 6837 12631
rect 6837 12597 6871 12631
rect 6871 12597 6880 12631
rect 6828 12588 6880 12597
rect 7840 12588 7892 12640
rect 10416 12835 10468 12844
rect 10416 12801 10425 12835
rect 10425 12801 10459 12835
rect 10459 12801 10468 12835
rect 10416 12792 10468 12801
rect 10876 12792 10928 12844
rect 9496 12724 9548 12776
rect 10324 12767 10376 12776
rect 10324 12733 10333 12767
rect 10333 12733 10367 12767
rect 10367 12733 10376 12767
rect 10324 12724 10376 12733
rect 9772 12588 9824 12640
rect 12808 12860 12860 12912
rect 11612 12792 11664 12844
rect 12256 12792 12308 12844
rect 13268 12792 13320 12844
rect 14556 12835 14608 12844
rect 14556 12801 14565 12835
rect 14565 12801 14599 12835
rect 14599 12801 14608 12835
rect 14556 12792 14608 12801
rect 12440 12724 12492 12776
rect 13820 12724 13872 12776
rect 14556 12656 14608 12708
rect 11336 12631 11388 12640
rect 11336 12597 11345 12631
rect 11345 12597 11379 12631
rect 11379 12597 11388 12631
rect 11336 12588 11388 12597
rect 11796 12588 11848 12640
rect 12256 12588 12308 12640
rect 13912 12631 13964 12640
rect 13912 12597 13921 12631
rect 13921 12597 13955 12631
rect 13955 12597 13964 12631
rect 13912 12588 13964 12597
rect 5912 12486 5964 12538
rect 5976 12486 6028 12538
rect 6040 12486 6092 12538
rect 6104 12486 6156 12538
rect 10843 12486 10895 12538
rect 10907 12486 10959 12538
rect 10971 12486 11023 12538
rect 11035 12486 11087 12538
rect 3240 12384 3292 12436
rect 4620 12384 4672 12436
rect 5724 12384 5776 12436
rect 6276 12384 6328 12436
rect 2228 12291 2280 12300
rect 2228 12257 2262 12291
rect 2262 12257 2280 12291
rect 2228 12248 2280 12257
rect 4252 12248 4304 12300
rect 4436 12291 4488 12300
rect 4436 12257 4445 12291
rect 4445 12257 4479 12291
rect 4479 12257 4488 12291
rect 4436 12248 4488 12257
rect 5080 12291 5132 12300
rect 5080 12257 5089 12291
rect 5089 12257 5123 12291
rect 5123 12257 5132 12291
rect 5080 12248 5132 12257
rect 5816 12248 5868 12300
rect 8300 12384 8352 12436
rect 7196 12316 7248 12368
rect 7564 12316 7616 12368
rect 11336 12384 11388 12436
rect 12532 12427 12584 12436
rect 12532 12393 12541 12427
rect 12541 12393 12575 12427
rect 12575 12393 12584 12427
rect 12532 12384 12584 12393
rect 13176 12427 13228 12436
rect 13176 12393 13185 12427
rect 13185 12393 13219 12427
rect 13219 12393 13228 12427
rect 13176 12384 13228 12393
rect 14924 12384 14976 12436
rect 10968 12316 11020 12368
rect 13912 12316 13964 12368
rect 14740 12316 14792 12368
rect 8668 12248 8720 12300
rect 10692 12248 10744 12300
rect 6736 12223 6788 12232
rect 1400 12044 1452 12096
rect 6736 12189 6745 12223
rect 6745 12189 6779 12223
rect 6779 12189 6788 12223
rect 6736 12180 6788 12189
rect 8208 12223 8260 12232
rect 8208 12189 8217 12223
rect 8217 12189 8251 12223
rect 8251 12189 8260 12223
rect 8208 12180 8260 12189
rect 8944 12223 8996 12232
rect 8944 12189 8953 12223
rect 8953 12189 8987 12223
rect 8987 12189 8996 12223
rect 8944 12180 8996 12189
rect 2872 12044 2924 12096
rect 4252 12112 4304 12164
rect 3792 12044 3844 12096
rect 5264 12044 5316 12096
rect 8852 12112 8904 12164
rect 9680 12180 9732 12232
rect 10416 12180 10468 12232
rect 12348 12248 12400 12300
rect 13084 12248 13136 12300
rect 14464 12248 14516 12300
rect 10876 12223 10928 12232
rect 10876 12189 10885 12223
rect 10885 12189 10919 12223
rect 10919 12189 10928 12223
rect 14924 12248 14976 12300
rect 10876 12180 10928 12189
rect 7932 12044 7984 12096
rect 10416 12044 10468 12096
rect 3447 11942 3499 11994
rect 3511 11942 3563 11994
rect 3575 11942 3627 11994
rect 3639 11942 3691 11994
rect 8378 11942 8430 11994
rect 8442 11942 8494 11994
rect 8506 11942 8558 11994
rect 8570 11942 8622 11994
rect 13308 11942 13360 11994
rect 13372 11942 13424 11994
rect 13436 11942 13488 11994
rect 13500 11942 13552 11994
rect 2136 11840 2188 11892
rect 2504 11747 2556 11756
rect 2504 11713 2513 11747
rect 2513 11713 2547 11747
rect 2547 11713 2556 11747
rect 4436 11840 4488 11892
rect 6368 11840 6420 11892
rect 8668 11883 8720 11892
rect 8668 11849 8677 11883
rect 8677 11849 8711 11883
rect 8711 11849 8720 11883
rect 8668 11840 8720 11849
rect 9036 11840 9088 11892
rect 9588 11840 9640 11892
rect 9680 11883 9732 11892
rect 9680 11849 9689 11883
rect 9689 11849 9723 11883
rect 9723 11849 9732 11883
rect 10692 11883 10744 11892
rect 9680 11840 9732 11849
rect 10692 11849 10701 11883
rect 10701 11849 10735 11883
rect 10735 11849 10744 11883
rect 10692 11840 10744 11849
rect 2872 11747 2924 11756
rect 2504 11704 2556 11713
rect 2872 11713 2881 11747
rect 2881 11713 2915 11747
rect 2915 11713 2924 11747
rect 2872 11704 2924 11713
rect 4896 11704 4948 11756
rect 5172 11704 5224 11756
rect 3148 11679 3200 11688
rect 3148 11645 3182 11679
rect 3182 11645 3200 11679
rect 5448 11704 5500 11756
rect 6276 11747 6328 11756
rect 6276 11713 6285 11747
rect 6285 11713 6319 11747
rect 6319 11713 6328 11747
rect 6276 11704 6328 11713
rect 14924 11772 14976 11824
rect 7472 11747 7524 11756
rect 3148 11636 3200 11645
rect 6828 11636 6880 11688
rect 7472 11713 7481 11747
rect 7481 11713 7515 11747
rect 7515 11713 7524 11747
rect 7472 11704 7524 11713
rect 9220 11747 9272 11756
rect 9220 11713 9229 11747
rect 9229 11713 9263 11747
rect 9263 11713 9272 11747
rect 9220 11704 9272 11713
rect 9772 11704 9824 11756
rect 10692 11704 10744 11756
rect 10968 11704 11020 11756
rect 11152 11747 11204 11756
rect 11152 11713 11161 11747
rect 11161 11713 11195 11747
rect 11195 11713 11204 11747
rect 11152 11704 11204 11713
rect 2780 11568 2832 11620
rect 3240 11568 3292 11620
rect 5632 11568 5684 11620
rect 2320 11543 2372 11552
rect 2320 11509 2329 11543
rect 2329 11509 2363 11543
rect 2363 11509 2372 11543
rect 4620 11543 4672 11552
rect 2320 11500 2372 11509
rect 4620 11509 4629 11543
rect 4629 11509 4663 11543
rect 4663 11509 4672 11543
rect 4620 11500 4672 11509
rect 4896 11500 4948 11552
rect 6460 11500 6512 11552
rect 8208 11636 8260 11688
rect 9956 11636 10008 11688
rect 10416 11636 10468 11688
rect 11520 11704 11572 11756
rect 15108 11747 15160 11756
rect 15108 11713 15117 11747
rect 15117 11713 15151 11747
rect 15151 11713 15160 11747
rect 15108 11704 15160 11713
rect 14648 11636 14700 11688
rect 7196 11568 7248 11620
rect 8300 11568 8352 11620
rect 9864 11568 9916 11620
rect 11060 11611 11112 11620
rect 11060 11577 11069 11611
rect 11069 11577 11103 11611
rect 11103 11577 11112 11611
rect 11060 11568 11112 11577
rect 13084 11568 13136 11620
rect 14004 11568 14056 11620
rect 8668 11500 8720 11552
rect 9496 11500 9548 11552
rect 13912 11500 13964 11552
rect 5912 11398 5964 11450
rect 5976 11398 6028 11450
rect 6040 11398 6092 11450
rect 6104 11398 6156 11450
rect 10843 11398 10895 11450
rect 10907 11398 10959 11450
rect 10971 11398 11023 11450
rect 11035 11398 11087 11450
rect 2228 11296 2280 11348
rect 5724 11296 5776 11348
rect 2504 11228 2556 11280
rect 5264 11271 5316 11280
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 2872 11092 2924 11144
rect 3240 10956 3292 11008
rect 5264 11237 5273 11271
rect 5273 11237 5307 11271
rect 5307 11237 5316 11271
rect 5264 11228 5316 11237
rect 6276 11296 6328 11348
rect 6736 11296 6788 11348
rect 6184 11228 6236 11280
rect 8300 11296 8352 11348
rect 8944 11296 8996 11348
rect 9036 11296 9088 11348
rect 9312 11296 9364 11348
rect 10324 11296 10376 11348
rect 11244 11296 11296 11348
rect 6460 11160 6512 11212
rect 8852 11228 8904 11280
rect 10140 11228 10192 11280
rect 7932 11203 7984 11212
rect 7932 11169 7941 11203
rect 7941 11169 7975 11203
rect 7975 11169 7984 11203
rect 8944 11203 8996 11212
rect 7932 11160 7984 11169
rect 8944 11169 8953 11203
rect 8953 11169 8987 11203
rect 8987 11169 8996 11203
rect 8944 11160 8996 11169
rect 6920 11092 6972 11144
rect 8024 11135 8076 11144
rect 8024 11101 8033 11135
rect 8033 11101 8067 11135
rect 8067 11101 8076 11135
rect 8024 11092 8076 11101
rect 9220 11135 9272 11144
rect 9220 11101 9229 11135
rect 9229 11101 9263 11135
rect 9263 11101 9272 11135
rect 9220 11092 9272 11101
rect 10232 11160 10284 11212
rect 10692 11160 10744 11212
rect 11704 11203 11756 11212
rect 10140 11092 10192 11144
rect 10876 11135 10928 11144
rect 10876 11101 10885 11135
rect 10885 11101 10919 11135
rect 10919 11101 10928 11135
rect 10876 11092 10928 11101
rect 4804 10956 4856 11008
rect 5080 10956 5132 11008
rect 7012 10956 7064 11008
rect 7564 10956 7616 11008
rect 9312 11024 9364 11076
rect 11704 11169 11713 11203
rect 11713 11169 11747 11203
rect 11747 11169 11756 11203
rect 11704 11160 11756 11169
rect 12532 11160 12584 11212
rect 9588 10956 9640 11008
rect 10508 10956 10560 11008
rect 3447 10854 3499 10906
rect 3511 10854 3563 10906
rect 3575 10854 3627 10906
rect 3639 10854 3691 10906
rect 8378 10854 8430 10906
rect 8442 10854 8494 10906
rect 8506 10854 8558 10906
rect 8570 10854 8622 10906
rect 13308 10854 13360 10906
rect 13372 10854 13424 10906
rect 13436 10854 13488 10906
rect 13500 10854 13552 10906
rect 2320 10752 2372 10804
rect 3148 10616 3200 10668
rect 3424 10616 3476 10668
rect 2964 10548 3016 10600
rect 5448 10752 5500 10804
rect 6736 10752 6788 10804
rect 8024 10752 8076 10804
rect 8852 10752 8904 10804
rect 10692 10752 10744 10804
rect 7288 10684 7340 10736
rect 7564 10684 7616 10736
rect 9588 10684 9640 10736
rect 3792 10480 3844 10532
rect 5632 10616 5684 10668
rect 7196 10659 7248 10668
rect 7196 10625 7205 10659
rect 7205 10625 7239 10659
rect 7239 10625 7248 10659
rect 7196 10616 7248 10625
rect 10048 10616 10100 10668
rect 10232 10616 10284 10668
rect 4252 10591 4304 10600
rect 4252 10557 4261 10591
rect 4261 10557 4295 10591
rect 4295 10557 4304 10591
rect 4252 10548 4304 10557
rect 5448 10548 5500 10600
rect 5540 10548 5592 10600
rect 4528 10523 4580 10532
rect 4528 10489 4562 10523
rect 4562 10489 4580 10523
rect 4528 10480 4580 10489
rect 2596 10455 2648 10464
rect 2596 10421 2605 10455
rect 2605 10421 2639 10455
rect 2639 10421 2648 10455
rect 2596 10412 2648 10421
rect 4344 10412 4396 10464
rect 7196 10480 7248 10532
rect 7748 10548 7800 10600
rect 9220 10548 9272 10600
rect 9772 10548 9824 10600
rect 10508 10548 10560 10600
rect 11704 10616 11756 10668
rect 14004 10616 14056 10668
rect 11244 10548 11296 10600
rect 15108 10548 15160 10600
rect 11888 10480 11940 10532
rect 4712 10412 4764 10464
rect 5172 10412 5224 10464
rect 11336 10412 11388 10464
rect 12532 10412 12584 10464
rect 14280 10455 14332 10464
rect 14280 10421 14289 10455
rect 14289 10421 14323 10455
rect 14323 10421 14332 10455
rect 14280 10412 14332 10421
rect 14372 10412 14424 10464
rect 5912 10310 5964 10362
rect 5976 10310 6028 10362
rect 6040 10310 6092 10362
rect 6104 10310 6156 10362
rect 10843 10310 10895 10362
rect 10907 10310 10959 10362
rect 10971 10310 11023 10362
rect 11035 10310 11087 10362
rect 2780 10208 2832 10260
rect 4528 10208 4580 10260
rect 8944 10208 8996 10260
rect 9220 10208 9272 10260
rect 11612 10208 11664 10260
rect 13636 10208 13688 10260
rect 14372 10251 14424 10260
rect 14372 10217 14381 10251
rect 14381 10217 14415 10251
rect 14415 10217 14424 10251
rect 14372 10208 14424 10217
rect 2320 10183 2372 10192
rect 2320 10149 2329 10183
rect 2329 10149 2363 10183
rect 2363 10149 2372 10183
rect 2320 10140 2372 10149
rect 5080 10140 5132 10192
rect 5356 10140 5408 10192
rect 5816 10140 5868 10192
rect 7012 10140 7064 10192
rect 3884 10072 3936 10124
rect 4804 10115 4856 10124
rect 3148 10004 3200 10056
rect 3332 10047 3384 10056
rect 3332 10013 3341 10047
rect 3341 10013 3375 10047
rect 3375 10013 3384 10047
rect 3332 10004 3384 10013
rect 3424 10047 3476 10056
rect 3424 10013 3433 10047
rect 3433 10013 3467 10047
rect 3467 10013 3476 10047
rect 3424 10004 3476 10013
rect 4528 9936 4580 9988
rect 1860 9911 1912 9920
rect 1860 9877 1869 9911
rect 1869 9877 1903 9911
rect 1903 9877 1912 9911
rect 1860 9868 1912 9877
rect 4344 9868 4396 9920
rect 4804 10081 4813 10115
rect 4813 10081 4847 10115
rect 4847 10081 4856 10115
rect 4804 10072 4856 10081
rect 5448 10072 5500 10124
rect 6276 10072 6328 10124
rect 8668 10072 8720 10124
rect 5080 10047 5132 10056
rect 5080 10013 5089 10047
rect 5089 10013 5123 10047
rect 5123 10013 5132 10047
rect 5080 10004 5132 10013
rect 8852 10004 8904 10056
rect 8760 9936 8812 9988
rect 9404 10140 9456 10192
rect 9680 10140 9732 10192
rect 9864 10072 9916 10124
rect 10508 10140 10560 10192
rect 15108 10140 15160 10192
rect 12164 10072 12216 10124
rect 14096 10072 14148 10124
rect 9128 10004 9180 10056
rect 9312 10047 9364 10056
rect 9312 10013 9321 10047
rect 9321 10013 9355 10047
rect 9355 10013 9364 10047
rect 9312 10004 9364 10013
rect 9772 10004 9824 10056
rect 7472 9868 7524 9920
rect 9772 9868 9824 9920
rect 11612 9868 11664 9920
rect 11704 9868 11756 9920
rect 12808 10004 12860 10056
rect 12992 10004 13044 10056
rect 14004 10047 14056 10056
rect 14004 10013 14013 10047
rect 14013 10013 14047 10047
rect 14047 10013 14056 10047
rect 14004 10004 14056 10013
rect 12624 9868 12676 9920
rect 12900 9868 12952 9920
rect 13084 9868 13136 9920
rect 14372 9868 14424 9920
rect 3447 9766 3499 9818
rect 3511 9766 3563 9818
rect 3575 9766 3627 9818
rect 3639 9766 3691 9818
rect 8378 9766 8430 9818
rect 8442 9766 8494 9818
rect 8506 9766 8558 9818
rect 8570 9766 8622 9818
rect 13308 9766 13360 9818
rect 13372 9766 13424 9818
rect 13436 9766 13488 9818
rect 13500 9766 13552 9818
rect 3148 9664 3200 9716
rect 7104 9664 7156 9716
rect 7840 9664 7892 9716
rect 1768 9639 1820 9648
rect 1768 9605 1777 9639
rect 1777 9605 1811 9639
rect 1811 9605 1820 9639
rect 1768 9596 1820 9605
rect 3884 9596 3936 9648
rect 7656 9596 7708 9648
rect 8024 9596 8076 9648
rect 8944 9596 8996 9648
rect 10140 9639 10192 9648
rect 2504 9528 2556 9580
rect 5080 9571 5132 9580
rect 5080 9537 5089 9571
rect 5089 9537 5123 9571
rect 5123 9537 5132 9571
rect 5080 9528 5132 9537
rect 7748 9528 7800 9580
rect 10140 9605 10149 9639
rect 10149 9605 10183 9639
rect 10183 9605 10192 9639
rect 10140 9596 10192 9605
rect 12624 9664 12676 9716
rect 11336 9639 11388 9648
rect 1860 9460 1912 9512
rect 2780 9503 2832 9512
rect 2780 9469 2789 9503
rect 2789 9469 2823 9503
rect 2823 9469 2832 9503
rect 2780 9460 2832 9469
rect 4620 9460 4672 9512
rect 4712 9460 4764 9512
rect 8392 9460 8444 9512
rect 8852 9460 8904 9512
rect 3516 9392 3568 9444
rect 6920 9392 6972 9444
rect 9404 9392 9456 9444
rect 9680 9460 9732 9512
rect 10324 9528 10376 9580
rect 10692 9571 10744 9580
rect 10692 9537 10701 9571
rect 10701 9537 10735 9571
rect 10735 9537 10744 9571
rect 10692 9528 10744 9537
rect 11336 9605 11345 9639
rect 11345 9605 11379 9639
rect 11379 9605 11388 9639
rect 11336 9596 11388 9605
rect 11796 9528 11848 9580
rect 12532 9528 12584 9580
rect 13084 9571 13136 9580
rect 13084 9537 13093 9571
rect 13093 9537 13127 9571
rect 13127 9537 13136 9571
rect 13084 9528 13136 9537
rect 10416 9460 10468 9512
rect 11704 9503 11756 9512
rect 11704 9469 11713 9503
rect 11713 9469 11747 9503
rect 11747 9469 11756 9503
rect 11704 9460 11756 9469
rect 11888 9460 11940 9512
rect 14280 9460 14332 9512
rect 13268 9392 13320 9444
rect 14372 9392 14424 9444
rect 2412 9324 2464 9376
rect 3792 9324 3844 9376
rect 4436 9367 4488 9376
rect 4436 9333 4445 9367
rect 4445 9333 4479 9367
rect 4479 9333 4488 9367
rect 4436 9324 4488 9333
rect 4620 9324 4672 9376
rect 5172 9324 5224 9376
rect 5816 9324 5868 9376
rect 8300 9324 8352 9376
rect 8944 9324 8996 9376
rect 9128 9324 9180 9376
rect 9864 9324 9916 9376
rect 10048 9324 10100 9376
rect 12072 9324 12124 9376
rect 12900 9367 12952 9376
rect 12900 9333 12909 9367
rect 12909 9333 12943 9367
rect 12943 9333 12952 9367
rect 12900 9324 12952 9333
rect 5912 9222 5964 9274
rect 5976 9222 6028 9274
rect 6040 9222 6092 9274
rect 6104 9222 6156 9274
rect 10843 9222 10895 9274
rect 10907 9222 10959 9274
rect 10971 9222 11023 9274
rect 11035 9222 11087 9274
rect 3516 9163 3568 9172
rect 3516 9129 3525 9163
rect 3525 9129 3559 9163
rect 3559 9129 3568 9163
rect 3516 9120 3568 9129
rect 3792 9120 3844 9172
rect 1676 9027 1728 9036
rect 1676 8993 1685 9027
rect 1685 8993 1719 9027
rect 1719 8993 1728 9027
rect 1676 8984 1728 8993
rect 2780 9052 2832 9104
rect 3884 9052 3936 9104
rect 4804 9120 4856 9172
rect 4252 8984 4304 9036
rect 4528 9027 4580 9036
rect 4528 8993 4537 9027
rect 4537 8993 4571 9027
rect 4571 8993 4580 9027
rect 4528 8984 4580 8993
rect 8668 9120 8720 9172
rect 9128 9120 9180 9172
rect 9864 9120 9916 9172
rect 8300 9052 8352 9104
rect 8944 9052 8996 9104
rect 12348 9120 12400 9172
rect 11612 9052 11664 9104
rect 12992 9052 13044 9104
rect 13636 9052 13688 9104
rect 15292 9052 15344 9104
rect 3884 8916 3936 8968
rect 7380 8984 7432 9036
rect 8392 8984 8444 9036
rect 9036 8984 9088 9036
rect 10784 8984 10836 9036
rect 11336 8984 11388 9036
rect 11520 8984 11572 9036
rect 11980 8984 12032 9036
rect 12440 8984 12492 9036
rect 12808 9027 12860 9036
rect 12808 8993 12817 9027
rect 12817 8993 12851 9027
rect 12851 8993 12860 9027
rect 12808 8984 12860 8993
rect 13820 9027 13872 9036
rect 13820 8993 13829 9027
rect 13829 8993 13863 9027
rect 13863 8993 13872 9027
rect 13820 8984 13872 8993
rect 6644 8959 6696 8968
rect 6644 8925 6653 8959
rect 6653 8925 6687 8959
rect 6687 8925 6696 8959
rect 6644 8916 6696 8925
rect 7840 8916 7892 8968
rect 9036 8848 9088 8900
rect 9864 8916 9916 8968
rect 10692 8959 10744 8968
rect 10692 8925 10701 8959
rect 10701 8925 10735 8959
rect 10735 8925 10744 8959
rect 10692 8916 10744 8925
rect 13084 8959 13136 8968
rect 13084 8925 13093 8959
rect 13093 8925 13127 8959
rect 13127 8925 13136 8959
rect 13084 8916 13136 8925
rect 14004 8959 14056 8968
rect 14004 8925 14013 8959
rect 14013 8925 14047 8959
rect 14047 8925 14056 8959
rect 14004 8916 14056 8925
rect 13268 8848 13320 8900
rect 11704 8780 11756 8832
rect 12164 8780 12216 8832
rect 13728 8780 13780 8832
rect 3447 8678 3499 8730
rect 3511 8678 3563 8730
rect 3575 8678 3627 8730
rect 3639 8678 3691 8730
rect 8378 8678 8430 8730
rect 8442 8678 8494 8730
rect 8506 8678 8558 8730
rect 8570 8678 8622 8730
rect 13308 8678 13360 8730
rect 13372 8678 13424 8730
rect 13436 8678 13488 8730
rect 13500 8678 13552 8730
rect 2412 8483 2464 8492
rect 2412 8449 2421 8483
rect 2421 8449 2455 8483
rect 2455 8449 2464 8483
rect 2412 8440 2464 8449
rect 3332 8483 3384 8492
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 4436 8576 4488 8628
rect 5724 8619 5776 8628
rect 5724 8585 5733 8619
rect 5733 8585 5767 8619
rect 5767 8585 5776 8619
rect 5724 8576 5776 8585
rect 6736 8576 6788 8628
rect 8760 8576 8812 8628
rect 8668 8508 8720 8560
rect 8852 8508 8904 8560
rect 4252 8440 4304 8492
rect 5080 8440 5132 8492
rect 5448 8483 5500 8492
rect 5448 8449 5457 8483
rect 5457 8449 5491 8483
rect 5491 8449 5500 8483
rect 5448 8440 5500 8449
rect 5816 8440 5868 8492
rect 6460 8440 6512 8492
rect 6644 8440 6696 8492
rect 7932 8440 7984 8492
rect 9036 8440 9088 8492
rect 6828 8372 6880 8424
rect 2964 8304 3016 8356
rect 4344 8304 4396 8356
rect 4436 8304 4488 8356
rect 5080 8304 5132 8356
rect 5540 8304 5592 8356
rect 6368 8304 6420 8356
rect 7288 8304 7340 8356
rect 10692 8576 10744 8628
rect 10876 8576 10928 8628
rect 12624 8576 12676 8628
rect 14004 8576 14056 8628
rect 11244 8508 11296 8560
rect 12164 8508 12216 8560
rect 11612 8483 11664 8492
rect 11612 8449 11621 8483
rect 11621 8449 11655 8483
rect 11655 8449 11664 8483
rect 11612 8440 11664 8449
rect 10600 8372 10652 8424
rect 10692 8372 10744 8424
rect 1492 8236 1544 8288
rect 3792 8279 3844 8288
rect 3792 8245 3801 8279
rect 3801 8245 3835 8279
rect 3835 8245 3844 8279
rect 3792 8236 3844 8245
rect 4252 8279 4304 8288
rect 4252 8245 4261 8279
rect 4261 8245 4295 8279
rect 4295 8245 4304 8279
rect 4252 8236 4304 8245
rect 4804 8279 4856 8288
rect 4804 8245 4813 8279
rect 4813 8245 4847 8279
rect 4847 8245 4856 8279
rect 4804 8236 4856 8245
rect 8760 8236 8812 8288
rect 9404 8236 9456 8288
rect 11060 8304 11112 8356
rect 12532 8304 12584 8356
rect 13084 8347 13136 8356
rect 13084 8313 13118 8347
rect 13118 8313 13136 8347
rect 13084 8304 13136 8313
rect 13268 8304 13320 8356
rect 11336 8279 11388 8288
rect 11336 8245 11345 8279
rect 11345 8245 11379 8279
rect 11379 8245 11388 8279
rect 11336 8236 11388 8245
rect 11612 8236 11664 8288
rect 12256 8236 12308 8288
rect 12900 8236 12952 8288
rect 5912 8134 5964 8186
rect 5976 8134 6028 8186
rect 6040 8134 6092 8186
rect 6104 8134 6156 8186
rect 10843 8134 10895 8186
rect 10907 8134 10959 8186
rect 10971 8134 11023 8186
rect 11035 8134 11087 8186
rect 2964 8075 3016 8084
rect 2964 8041 2973 8075
rect 2973 8041 3007 8075
rect 3007 8041 3016 8075
rect 2964 8032 3016 8041
rect 3792 8032 3844 8084
rect 4252 8032 4304 8084
rect 5172 8032 5224 8084
rect 5448 8032 5500 8084
rect 7288 8032 7340 8084
rect 9680 8032 9732 8084
rect 10324 8032 10376 8084
rect 13820 8032 13872 8084
rect 2504 8007 2556 8016
rect 2504 7973 2513 8007
rect 2513 7973 2547 8007
rect 2547 7973 2556 8007
rect 2504 7964 2556 7973
rect 4344 7964 4396 8016
rect 1492 7939 1544 7948
rect 1492 7905 1501 7939
rect 1501 7905 1535 7939
rect 1535 7905 1544 7939
rect 1492 7896 1544 7905
rect 1676 7871 1728 7880
rect 1676 7837 1685 7871
rect 1685 7837 1719 7871
rect 1719 7837 1728 7871
rect 1676 7828 1728 7837
rect 3332 7896 3384 7948
rect 4160 7896 4212 7948
rect 8484 7964 8536 8016
rect 9956 7964 10008 8016
rect 10784 7964 10836 8016
rect 12992 7964 13044 8016
rect 6184 7896 6236 7948
rect 7564 7896 7616 7948
rect 7748 7896 7800 7948
rect 8852 7896 8904 7948
rect 9312 7896 9364 7948
rect 11060 7939 11112 7948
rect 7288 7871 7340 7880
rect 3884 7760 3936 7812
rect 7288 7837 7297 7871
rect 7297 7837 7331 7871
rect 7331 7837 7340 7871
rect 7288 7828 7340 7837
rect 7380 7871 7432 7880
rect 7380 7837 7389 7871
rect 7389 7837 7423 7871
rect 7423 7837 7432 7871
rect 7380 7828 7432 7837
rect 7564 7760 7616 7812
rect 9128 7871 9180 7880
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 11060 7905 11069 7939
rect 11069 7905 11103 7939
rect 11103 7905 11112 7939
rect 11060 7896 11112 7905
rect 11428 7896 11480 7948
rect 11888 7896 11940 7948
rect 12072 7939 12124 7948
rect 12072 7905 12081 7939
rect 12081 7905 12115 7939
rect 12115 7905 12124 7939
rect 12072 7896 12124 7905
rect 12532 7896 12584 7948
rect 12900 7896 12952 7948
rect 9128 7828 9180 7837
rect 11152 7828 11204 7880
rect 11336 7828 11388 7880
rect 13268 7871 13320 7880
rect 13268 7837 13277 7871
rect 13277 7837 13311 7871
rect 13311 7837 13320 7871
rect 13268 7828 13320 7837
rect 9956 7760 10008 7812
rect 10140 7760 10192 7812
rect 11704 7803 11756 7812
rect 11704 7769 11713 7803
rect 11713 7769 11747 7803
rect 11747 7769 11756 7803
rect 11704 7760 11756 7769
rect 13176 7692 13228 7744
rect 15016 7692 15068 7744
rect 3447 7590 3499 7642
rect 3511 7590 3563 7642
rect 3575 7590 3627 7642
rect 3639 7590 3691 7642
rect 8378 7590 8430 7642
rect 8442 7590 8494 7642
rect 8506 7590 8558 7642
rect 8570 7590 8622 7642
rect 13308 7590 13360 7642
rect 13372 7590 13424 7642
rect 13436 7590 13488 7642
rect 13500 7590 13552 7642
rect 5540 7531 5592 7540
rect 5540 7497 5549 7531
rect 5549 7497 5583 7531
rect 5583 7497 5592 7531
rect 5540 7488 5592 7497
rect 6828 7531 6880 7540
rect 6828 7497 6837 7531
rect 6837 7497 6871 7531
rect 6871 7497 6880 7531
rect 6828 7488 6880 7497
rect 4160 7352 4212 7404
rect 6184 7395 6236 7404
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 2872 7327 2924 7336
rect 2872 7293 2881 7327
rect 2881 7293 2915 7327
rect 2915 7293 2924 7327
rect 2872 7284 2924 7293
rect 9036 7488 9088 7540
rect 10784 7488 10836 7540
rect 11060 7531 11112 7540
rect 11060 7497 11069 7531
rect 11069 7497 11103 7531
rect 11103 7497 11112 7531
rect 11060 7488 11112 7497
rect 10232 7420 10284 7472
rect 11612 7352 11664 7404
rect 13452 7352 13504 7404
rect 8024 7327 8076 7336
rect 8024 7293 8033 7327
rect 8033 7293 8067 7327
rect 8067 7293 8076 7327
rect 8024 7284 8076 7293
rect 8300 7327 8352 7336
rect 8300 7293 8309 7327
rect 8309 7293 8343 7327
rect 8343 7293 8352 7327
rect 8300 7284 8352 7293
rect 10140 7284 10192 7336
rect 10324 7284 10376 7336
rect 11520 7284 11572 7336
rect 11888 7284 11940 7336
rect 12716 7284 12768 7336
rect 3056 7216 3108 7268
rect 4896 7259 4948 7268
rect 4896 7225 4905 7259
rect 4905 7225 4939 7259
rect 4939 7225 4948 7259
rect 4896 7216 4948 7225
rect 1400 7148 1452 7200
rect 2872 7148 2924 7200
rect 4988 7191 5040 7200
rect 4988 7157 4997 7191
rect 4997 7157 5031 7191
rect 5031 7157 5040 7191
rect 4988 7148 5040 7157
rect 6276 7148 6328 7200
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 7656 7148 7708 7200
rect 9312 7216 9364 7268
rect 9404 7216 9456 7268
rect 11704 7216 11756 7268
rect 13084 7216 13136 7268
rect 9220 7148 9272 7200
rect 9680 7148 9732 7200
rect 10600 7148 10652 7200
rect 12440 7191 12492 7200
rect 12440 7157 12449 7191
rect 12449 7157 12483 7191
rect 12483 7157 12492 7191
rect 12440 7148 12492 7157
rect 12624 7148 12676 7200
rect 16304 7148 16356 7200
rect 5912 7046 5964 7098
rect 5976 7046 6028 7098
rect 6040 7046 6092 7098
rect 6104 7046 6156 7098
rect 10843 7046 10895 7098
rect 10907 7046 10959 7098
rect 10971 7046 11023 7098
rect 11035 7046 11087 7098
rect 3056 6987 3108 6996
rect 3056 6953 3065 6987
rect 3065 6953 3099 6987
rect 3099 6953 3108 6987
rect 3056 6944 3108 6953
rect 4896 6944 4948 6996
rect 6276 6944 6328 6996
rect 6828 6876 6880 6928
rect 4160 6808 4212 6860
rect 5264 6851 5316 6860
rect 5264 6817 5273 6851
rect 5273 6817 5307 6851
rect 5307 6817 5316 6851
rect 5264 6808 5316 6817
rect 5356 6783 5408 6792
rect 5356 6749 5365 6783
rect 5365 6749 5399 6783
rect 5399 6749 5408 6783
rect 6920 6808 6972 6860
rect 7104 6851 7156 6860
rect 7104 6817 7113 6851
rect 7113 6817 7147 6851
rect 7147 6817 7156 6851
rect 7104 6808 7156 6817
rect 8300 6876 8352 6928
rect 8668 6876 8720 6928
rect 9312 6944 9364 6996
rect 10324 6944 10376 6996
rect 11244 6944 11296 6996
rect 10048 6919 10100 6928
rect 10048 6885 10057 6919
rect 10057 6885 10091 6919
rect 10091 6885 10100 6919
rect 10048 6876 10100 6885
rect 11612 6876 11664 6928
rect 11704 6876 11756 6928
rect 12992 6876 13044 6928
rect 9036 6808 9088 6860
rect 10324 6808 10376 6860
rect 11336 6808 11388 6860
rect 12532 6808 12584 6860
rect 13636 6808 13688 6860
rect 14372 6808 14424 6860
rect 7196 6783 7248 6792
rect 5356 6740 5408 6749
rect 7196 6749 7205 6783
rect 7205 6749 7239 6783
rect 7239 6749 7248 6783
rect 7196 6740 7248 6749
rect 7380 6783 7432 6792
rect 7380 6749 7389 6783
rect 7389 6749 7423 6783
rect 7423 6749 7432 6783
rect 7380 6740 7432 6749
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 13452 6783 13504 6792
rect 10232 6740 10284 6749
rect 13452 6749 13461 6783
rect 13461 6749 13495 6783
rect 13495 6749 13504 6783
rect 13452 6740 13504 6749
rect 7656 6672 7708 6724
rect 9496 6672 9548 6724
rect 10600 6672 10652 6724
rect 2780 6604 2832 6656
rect 4528 6647 4580 6656
rect 4528 6613 4537 6647
rect 4537 6613 4571 6647
rect 4571 6613 4580 6647
rect 4528 6604 4580 6613
rect 4712 6604 4764 6656
rect 5632 6604 5684 6656
rect 6736 6647 6788 6656
rect 6736 6613 6745 6647
rect 6745 6613 6779 6647
rect 6779 6613 6788 6647
rect 6736 6604 6788 6613
rect 10692 6647 10744 6656
rect 10692 6613 10701 6647
rect 10701 6613 10735 6647
rect 10735 6613 10744 6647
rect 10692 6604 10744 6613
rect 12900 6647 12952 6656
rect 12900 6613 12909 6647
rect 12909 6613 12943 6647
rect 12943 6613 12952 6647
rect 12900 6604 12952 6613
rect 3447 6502 3499 6554
rect 3511 6502 3563 6554
rect 3575 6502 3627 6554
rect 3639 6502 3691 6554
rect 8378 6502 8430 6554
rect 8442 6502 8494 6554
rect 8506 6502 8558 6554
rect 8570 6502 8622 6554
rect 13308 6502 13360 6554
rect 13372 6502 13424 6554
rect 13436 6502 13488 6554
rect 13500 6502 13552 6554
rect 4160 6400 4212 6452
rect 4988 6400 5040 6452
rect 1768 6196 1820 6248
rect 5356 6264 5408 6316
rect 6368 6307 6420 6316
rect 6368 6273 6377 6307
rect 6377 6273 6411 6307
rect 6411 6273 6420 6307
rect 6368 6264 6420 6273
rect 4068 6196 4120 6248
rect 6736 6196 6788 6248
rect 9220 6264 9272 6316
rect 10140 6400 10192 6452
rect 12072 6400 12124 6452
rect 12440 6400 12492 6452
rect 11612 6332 11664 6384
rect 11244 6264 11296 6316
rect 12532 6264 12584 6316
rect 2412 6128 2464 6180
rect 6184 6128 6236 6180
rect 6276 6128 6328 6180
rect 8392 6196 8444 6248
rect 7380 6128 7432 6180
rect 8300 6128 8352 6180
rect 3332 6103 3384 6112
rect 3332 6069 3341 6103
rect 3341 6069 3375 6103
rect 3375 6069 3384 6103
rect 3332 6060 3384 6069
rect 4068 6060 4120 6112
rect 4896 6103 4948 6112
rect 4896 6069 4905 6103
rect 4905 6069 4939 6103
rect 4939 6069 4948 6103
rect 4896 6060 4948 6069
rect 5816 6060 5868 6112
rect 6552 6060 6604 6112
rect 10232 6196 10284 6248
rect 13912 6264 13964 6316
rect 14740 6264 14792 6316
rect 11428 6128 11480 6180
rect 12900 6128 12952 6180
rect 8484 6060 8536 6112
rect 9496 6060 9548 6112
rect 9680 6060 9732 6112
rect 10232 6060 10284 6112
rect 5912 5958 5964 6010
rect 5976 5958 6028 6010
rect 6040 5958 6092 6010
rect 6104 5958 6156 6010
rect 10843 5958 10895 6010
rect 10907 5958 10959 6010
rect 10971 5958 11023 6010
rect 11035 5958 11087 6010
rect 4068 5899 4120 5908
rect 4068 5865 4077 5899
rect 4077 5865 4111 5899
rect 4111 5865 4120 5899
rect 4068 5856 4120 5865
rect 4344 5856 4396 5908
rect 4804 5856 4856 5908
rect 4896 5856 4948 5908
rect 1676 5831 1728 5840
rect 1676 5797 1685 5831
rect 1685 5797 1719 5831
rect 1719 5797 1728 5831
rect 1676 5788 1728 5797
rect 1768 5788 1820 5840
rect 3240 5788 3292 5840
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 4620 5788 4672 5840
rect 6368 5788 6420 5840
rect 7104 5856 7156 5908
rect 7196 5856 7248 5908
rect 9404 5856 9456 5908
rect 9496 5856 9548 5908
rect 14280 5856 14332 5908
rect 8484 5788 8536 5840
rect 6276 5720 6328 5772
rect 7472 5720 7524 5772
rect 2596 5695 2648 5704
rect 2596 5661 2605 5695
rect 2605 5661 2639 5695
rect 2639 5661 2648 5695
rect 2596 5652 2648 5661
rect 2688 5695 2740 5704
rect 2688 5661 2697 5695
rect 2697 5661 2731 5695
rect 2731 5661 2740 5695
rect 2688 5652 2740 5661
rect 4620 5695 4672 5704
rect 4620 5661 4629 5695
rect 4629 5661 4663 5695
rect 4663 5661 4672 5695
rect 4620 5652 4672 5661
rect 2228 5516 2280 5568
rect 3884 5516 3936 5568
rect 4344 5516 4396 5568
rect 7564 5652 7616 5704
rect 7840 5763 7892 5772
rect 7840 5729 7849 5763
rect 7849 5729 7883 5763
rect 7883 5729 7892 5763
rect 7840 5720 7892 5729
rect 8852 5720 8904 5772
rect 13912 5788 13964 5840
rect 14740 5831 14792 5840
rect 14740 5797 14749 5831
rect 14749 5797 14783 5831
rect 14783 5797 14792 5831
rect 14740 5788 14792 5797
rect 7932 5652 7984 5704
rect 8300 5652 8352 5704
rect 9220 5652 9272 5704
rect 7012 5584 7064 5636
rect 9956 5720 10008 5772
rect 10784 5720 10836 5772
rect 13176 5720 13228 5772
rect 10232 5652 10284 5704
rect 10600 5695 10652 5704
rect 10600 5661 10609 5695
rect 10609 5661 10643 5695
rect 10643 5661 10652 5695
rect 10600 5652 10652 5661
rect 11336 5652 11388 5704
rect 13636 5695 13688 5704
rect 13636 5661 13645 5695
rect 13645 5661 13679 5695
rect 13679 5661 13688 5695
rect 13636 5652 13688 5661
rect 6644 5559 6696 5568
rect 6644 5525 6653 5559
rect 6653 5525 6687 5559
rect 6687 5525 6696 5559
rect 6644 5516 6696 5525
rect 7380 5559 7432 5568
rect 7380 5525 7389 5559
rect 7389 5525 7423 5559
rect 7423 5525 7432 5559
rect 7380 5516 7432 5525
rect 7564 5516 7616 5568
rect 9404 5584 9456 5636
rect 9128 5559 9180 5568
rect 9128 5525 9137 5559
rect 9137 5525 9171 5559
rect 9171 5525 9180 5559
rect 9128 5516 9180 5525
rect 9956 5559 10008 5568
rect 9956 5525 9965 5559
rect 9965 5525 9999 5559
rect 9999 5525 10008 5559
rect 9956 5516 10008 5525
rect 14188 5516 14240 5568
rect 3447 5414 3499 5466
rect 3511 5414 3563 5466
rect 3575 5414 3627 5466
rect 3639 5414 3691 5466
rect 8378 5414 8430 5466
rect 8442 5414 8494 5466
rect 8506 5414 8558 5466
rect 8570 5414 8622 5466
rect 13308 5414 13360 5466
rect 13372 5414 13424 5466
rect 13436 5414 13488 5466
rect 13500 5414 13552 5466
rect 5356 5312 5408 5364
rect 7656 5312 7708 5364
rect 2688 5219 2740 5228
rect 2688 5185 2697 5219
rect 2697 5185 2731 5219
rect 2731 5185 2740 5219
rect 2688 5176 2740 5185
rect 1768 5108 1820 5160
rect 3792 5108 3844 5160
rect 5172 5176 5224 5228
rect 6368 5219 6420 5228
rect 6368 5185 6377 5219
rect 6377 5185 6411 5219
rect 6411 5185 6420 5219
rect 6368 5176 6420 5185
rect 6828 5219 6880 5228
rect 6828 5185 6837 5219
rect 6837 5185 6871 5219
rect 6871 5185 6880 5219
rect 6828 5176 6880 5185
rect 6920 5176 6972 5228
rect 4620 5108 4672 5160
rect 7380 5108 7432 5160
rect 9220 5312 9272 5364
rect 10600 5312 10652 5364
rect 13636 5312 13688 5364
rect 14096 5244 14148 5296
rect 15936 5244 15988 5296
rect 14740 5219 14792 5228
rect 14740 5185 14749 5219
rect 14749 5185 14783 5219
rect 14783 5185 14792 5219
rect 14740 5176 14792 5185
rect 1400 4972 1452 5024
rect 2320 4972 2372 5024
rect 2504 5015 2556 5024
rect 2504 4981 2513 5015
rect 2513 4981 2547 5015
rect 2547 4981 2556 5015
rect 2504 4972 2556 4981
rect 2964 4972 3016 5024
rect 5724 5015 5776 5024
rect 5724 4981 5733 5015
rect 5733 4981 5767 5015
rect 5767 4981 5776 5015
rect 5724 4972 5776 4981
rect 9496 5108 9548 5160
rect 9864 5108 9916 5160
rect 10140 5108 10192 5160
rect 12532 5108 12584 5160
rect 14924 5108 14976 5160
rect 6920 4972 6972 5024
rect 7196 4972 7248 5024
rect 8392 5040 8444 5092
rect 8760 5040 8812 5092
rect 7748 5015 7800 5024
rect 7748 4981 7757 5015
rect 7757 4981 7791 5015
rect 7791 4981 7800 5015
rect 7748 4972 7800 4981
rect 10508 5040 10560 5092
rect 8944 4972 8996 5024
rect 12624 5040 12676 5092
rect 14096 5015 14148 5024
rect 14096 4981 14105 5015
rect 14105 4981 14139 5015
rect 14139 4981 14148 5015
rect 14096 4972 14148 4981
rect 14464 5015 14516 5024
rect 14464 4981 14473 5015
rect 14473 4981 14507 5015
rect 14507 4981 14516 5015
rect 14464 4972 14516 4981
rect 5912 4870 5964 4922
rect 5976 4870 6028 4922
rect 6040 4870 6092 4922
rect 6104 4870 6156 4922
rect 10843 4870 10895 4922
rect 10907 4870 10959 4922
rect 10971 4870 11023 4922
rect 11035 4870 11087 4922
rect 2320 4811 2372 4820
rect 2320 4777 2329 4811
rect 2329 4777 2363 4811
rect 2363 4777 2372 4811
rect 2320 4768 2372 4777
rect 2872 4811 2924 4820
rect 2872 4777 2881 4811
rect 2881 4777 2915 4811
rect 2915 4777 2924 4811
rect 2872 4768 2924 4777
rect 3332 4768 3384 4820
rect 5172 4768 5224 4820
rect 2228 4743 2280 4752
rect 2228 4709 2237 4743
rect 2237 4709 2271 4743
rect 2271 4709 2280 4743
rect 2228 4700 2280 4709
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 2412 4564 2464 4573
rect 4160 4564 4212 4616
rect 5080 4632 5132 4684
rect 6276 4768 6328 4820
rect 7748 4768 7800 4820
rect 9956 4768 10008 4820
rect 12624 4768 12676 4820
rect 14556 4811 14608 4820
rect 14556 4777 14565 4811
rect 14565 4777 14599 4811
rect 14599 4777 14608 4811
rect 14556 4768 14608 4777
rect 15108 4768 15160 4820
rect 6644 4700 6696 4752
rect 7656 4700 7708 4752
rect 8024 4743 8076 4752
rect 8024 4709 8033 4743
rect 8033 4709 8067 4743
rect 8067 4709 8076 4743
rect 8024 4700 8076 4709
rect 9772 4700 9824 4752
rect 10600 4700 10652 4752
rect 12072 4700 12124 4752
rect 15016 4700 15068 4752
rect 6552 4632 6604 4684
rect 7840 4632 7892 4684
rect 9404 4632 9456 4684
rect 8760 4564 8812 4616
rect 8944 4564 8996 4616
rect 3056 4496 3108 4548
rect 8116 4496 8168 4548
rect 10140 4496 10192 4548
rect 13728 4632 13780 4684
rect 12532 4607 12584 4616
rect 12532 4573 12541 4607
rect 12541 4573 12575 4607
rect 12575 4573 12584 4607
rect 12532 4564 12584 4573
rect 14740 4607 14792 4616
rect 14740 4573 14749 4607
rect 14749 4573 14783 4607
rect 14783 4573 14792 4607
rect 14740 4564 14792 4573
rect 11612 4539 11664 4548
rect 11612 4505 11621 4539
rect 11621 4505 11655 4539
rect 11655 4505 11664 4539
rect 11612 4496 11664 4505
rect 4252 4471 4304 4480
rect 4252 4437 4261 4471
rect 4261 4437 4295 4471
rect 4295 4437 4304 4471
rect 4252 4428 4304 4437
rect 4804 4471 4856 4480
rect 4804 4437 4813 4471
rect 4813 4437 4847 4471
rect 4847 4437 4856 4471
rect 4804 4428 4856 4437
rect 7196 4471 7248 4480
rect 7196 4437 7205 4471
rect 7205 4437 7239 4471
rect 7239 4437 7248 4471
rect 7196 4428 7248 4437
rect 9036 4428 9088 4480
rect 9496 4428 9548 4480
rect 14188 4471 14240 4480
rect 14188 4437 14197 4471
rect 14197 4437 14231 4471
rect 14231 4437 14240 4471
rect 14188 4428 14240 4437
rect 3447 4326 3499 4378
rect 3511 4326 3563 4378
rect 3575 4326 3627 4378
rect 3639 4326 3691 4378
rect 8378 4326 8430 4378
rect 8442 4326 8494 4378
rect 8506 4326 8558 4378
rect 8570 4326 8622 4378
rect 13308 4326 13360 4378
rect 13372 4326 13424 4378
rect 13436 4326 13488 4378
rect 13500 4326 13552 4378
rect 2504 4224 2556 4276
rect 4620 4224 4672 4276
rect 7840 4224 7892 4276
rect 8024 4224 8076 4276
rect 1676 4131 1728 4140
rect 1676 4097 1685 4131
rect 1685 4097 1719 4131
rect 1719 4097 1728 4131
rect 1676 4088 1728 4097
rect 2228 4063 2280 4072
rect 2228 4029 2237 4063
rect 2237 4029 2271 4063
rect 2271 4029 2280 4063
rect 2228 4020 2280 4029
rect 2780 4020 2832 4072
rect 4436 4088 4488 4140
rect 4620 4088 4672 4140
rect 5264 4131 5316 4140
rect 5264 4097 5273 4131
rect 5273 4097 5307 4131
rect 5307 4097 5316 4131
rect 5264 4088 5316 4097
rect 5724 4088 5776 4140
rect 6644 4156 6696 4208
rect 8944 4224 8996 4276
rect 9496 4267 9548 4276
rect 9496 4233 9505 4267
rect 9505 4233 9539 4267
rect 9539 4233 9548 4267
rect 9496 4224 9548 4233
rect 9772 4267 9824 4276
rect 9772 4233 9781 4267
rect 9781 4233 9815 4267
rect 9815 4233 9824 4267
rect 9772 4224 9824 4233
rect 10600 4088 10652 4140
rect 11888 4088 11940 4140
rect 12624 4156 12676 4208
rect 13728 4088 13780 4140
rect 14464 4131 14516 4140
rect 14464 4097 14473 4131
rect 14473 4097 14507 4131
rect 14507 4097 14516 4131
rect 14464 4088 14516 4097
rect 1952 3884 2004 3936
rect 3332 3952 3384 4004
rect 3700 3952 3752 4004
rect 4988 3952 5040 4004
rect 5448 3952 5500 4004
rect 3792 3884 3844 3936
rect 4712 3927 4764 3936
rect 4712 3893 4721 3927
rect 4721 3893 4755 3927
rect 4755 3893 4764 3927
rect 4712 3884 4764 3893
rect 5172 3927 5224 3936
rect 5172 3893 5181 3927
rect 5181 3893 5215 3927
rect 5215 3893 5224 3927
rect 5816 4020 5868 4072
rect 6736 4020 6788 4072
rect 7840 4063 7892 4072
rect 7840 4029 7849 4063
rect 7849 4029 7883 4063
rect 7883 4029 7892 4063
rect 7840 4020 7892 4029
rect 6552 3952 6604 4004
rect 8208 3952 8260 4004
rect 8668 4020 8720 4072
rect 9220 4020 9272 4072
rect 10692 4020 10744 4072
rect 10784 4063 10836 4072
rect 10784 4029 10793 4063
rect 10793 4029 10827 4063
rect 10827 4029 10836 4063
rect 10784 4020 10836 4029
rect 11152 4020 11204 4072
rect 5172 3884 5224 3893
rect 5816 3884 5868 3936
rect 7380 3884 7432 3936
rect 9128 3884 9180 3936
rect 9772 3884 9824 3936
rect 10048 3884 10100 3936
rect 10324 3884 10376 3936
rect 10416 3884 10468 3936
rect 10692 3884 10744 3936
rect 11888 3952 11940 4004
rect 12348 3952 12400 4004
rect 11336 3927 11388 3936
rect 11336 3893 11345 3927
rect 11345 3893 11379 3927
rect 11379 3893 11388 3927
rect 11336 3884 11388 3893
rect 11428 3884 11480 3936
rect 12624 3884 12676 3936
rect 12900 3927 12952 3936
rect 12900 3893 12909 3927
rect 12909 3893 12943 3927
rect 12943 3893 12952 3927
rect 12900 3884 12952 3893
rect 13176 3884 13228 3936
rect 14188 4020 14240 4072
rect 14096 3952 14148 4004
rect 14372 3884 14424 3936
rect 5912 3782 5964 3834
rect 5976 3782 6028 3834
rect 6040 3782 6092 3834
rect 6104 3782 6156 3834
rect 10843 3782 10895 3834
rect 10907 3782 10959 3834
rect 10971 3782 11023 3834
rect 11035 3782 11087 3834
rect 1952 3587 2004 3596
rect 1952 3553 1961 3587
rect 1961 3553 1995 3587
rect 1995 3553 2004 3587
rect 1952 3544 2004 3553
rect 3240 3612 3292 3664
rect 3700 3544 3752 3596
rect 4528 3680 4580 3732
rect 4988 3680 5040 3732
rect 6644 3680 6696 3732
rect 6828 3680 6880 3732
rect 4344 3612 4396 3664
rect 5264 3612 5316 3664
rect 4436 3544 4488 3596
rect 4988 3544 5040 3596
rect 3792 3476 3844 3528
rect 7196 3612 7248 3664
rect 7656 3680 7708 3732
rect 8852 3680 8904 3732
rect 9036 3723 9088 3732
rect 9036 3689 9045 3723
rect 9045 3689 9079 3723
rect 9079 3689 9088 3723
rect 9036 3680 9088 3689
rect 10508 3680 10560 3732
rect 11428 3723 11480 3732
rect 11428 3689 11437 3723
rect 11437 3689 11471 3723
rect 11471 3689 11480 3723
rect 11428 3680 11480 3689
rect 11796 3723 11848 3732
rect 11796 3689 11805 3723
rect 11805 3689 11839 3723
rect 11839 3689 11848 3723
rect 11796 3680 11848 3689
rect 11888 3680 11940 3732
rect 13912 3723 13964 3732
rect 13912 3689 13921 3723
rect 13921 3689 13955 3723
rect 13955 3689 13964 3723
rect 13912 3680 13964 3689
rect 11152 3612 11204 3664
rect 12348 3612 12400 3664
rect 12440 3612 12492 3664
rect 6276 3544 6328 3596
rect 8116 3544 8168 3596
rect 9772 3544 9824 3596
rect 12716 3544 12768 3596
rect 6368 3476 6420 3528
rect 7840 3476 7892 3528
rect 7932 3408 7984 3460
rect 9404 3476 9456 3528
rect 9588 3476 9640 3528
rect 10600 3519 10652 3528
rect 572 3340 624 3392
rect 3332 3383 3384 3392
rect 3332 3349 3341 3383
rect 3341 3349 3375 3383
rect 3375 3349 3384 3383
rect 3332 3340 3384 3349
rect 3792 3340 3844 3392
rect 5816 3340 5868 3392
rect 6368 3340 6420 3392
rect 6736 3340 6788 3392
rect 8668 3340 8720 3392
rect 9680 3408 9732 3460
rect 10600 3485 10609 3519
rect 10609 3485 10643 3519
rect 10643 3485 10652 3519
rect 10600 3476 10652 3485
rect 11336 3476 11388 3528
rect 13728 3544 13780 3596
rect 14188 3544 14240 3596
rect 13176 3476 13228 3528
rect 13268 3476 13320 3528
rect 10508 3408 10560 3460
rect 12900 3408 12952 3460
rect 9496 3340 9548 3392
rect 9956 3383 10008 3392
rect 9956 3349 9965 3383
rect 9965 3349 9999 3383
rect 9999 3349 10008 3383
rect 9956 3340 10008 3349
rect 10048 3340 10100 3392
rect 3447 3238 3499 3290
rect 3511 3238 3563 3290
rect 3575 3238 3627 3290
rect 3639 3238 3691 3290
rect 8378 3238 8430 3290
rect 8442 3238 8494 3290
rect 8506 3238 8558 3290
rect 8570 3238 8622 3290
rect 13308 3238 13360 3290
rect 13372 3238 13424 3290
rect 13436 3238 13488 3290
rect 13500 3238 13552 3290
rect 2228 3179 2280 3188
rect 2228 3145 2237 3179
rect 2237 3145 2271 3179
rect 2271 3145 2280 3179
rect 2228 3136 2280 3145
rect 2688 3136 2740 3188
rect 4804 3136 4856 3188
rect 5172 3136 5224 3188
rect 5816 3136 5868 3188
rect 7840 3136 7892 3188
rect 8208 3136 8260 3188
rect 9404 3136 9456 3188
rect 11336 3179 11388 3188
rect 11336 3145 11345 3179
rect 11345 3145 11379 3179
rect 11379 3145 11388 3179
rect 11336 3136 11388 3145
rect 11796 3136 11848 3188
rect 12256 3136 12308 3188
rect 14188 3136 14240 3188
rect 1676 3043 1728 3052
rect 1676 3009 1685 3043
rect 1685 3009 1719 3043
rect 1719 3009 1728 3043
rect 1676 3000 1728 3009
rect 4712 3068 4764 3120
rect 12532 3068 12584 3120
rect 3332 3000 3384 3052
rect 3424 3000 3476 3052
rect 4344 3000 4396 3052
rect 4988 3000 5040 3052
rect 5172 3000 5224 3052
rect 5632 3000 5684 3052
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 7196 3000 7248 3052
rect 7932 3043 7984 3052
rect 7932 3009 7941 3043
rect 7941 3009 7975 3043
rect 7975 3009 7984 3043
rect 7932 3000 7984 3009
rect 9496 3000 9548 3052
rect 11704 3000 11756 3052
rect 12440 3043 12492 3052
rect 12440 3009 12449 3043
rect 12449 3009 12483 3043
rect 12483 3009 12492 3043
rect 12440 3000 12492 3009
rect 14648 3000 14700 3052
rect 2044 2932 2096 2984
rect 2228 2932 2280 2984
rect 4252 2932 4304 2984
rect 4712 2932 4764 2984
rect 6644 2932 6696 2984
rect 1492 2796 1544 2848
rect 2964 2796 3016 2848
rect 4344 2864 4396 2916
rect 4436 2864 4488 2916
rect 9312 2932 9364 2984
rect 5080 2796 5132 2848
rect 5264 2839 5316 2848
rect 5264 2805 5273 2839
rect 5273 2805 5307 2839
rect 5307 2805 5316 2839
rect 5264 2796 5316 2805
rect 5816 2796 5868 2848
rect 7932 2864 7984 2916
rect 8024 2864 8076 2916
rect 12532 2932 12584 2984
rect 10416 2864 10468 2916
rect 10600 2864 10652 2916
rect 13176 2907 13228 2916
rect 13176 2873 13210 2907
rect 13210 2873 13228 2907
rect 13176 2864 13228 2873
rect 11152 2796 11204 2848
rect 11428 2796 11480 2848
rect 14740 2796 14792 2848
rect 16764 2864 16816 2916
rect 5912 2694 5964 2746
rect 5976 2694 6028 2746
rect 6040 2694 6092 2746
rect 6104 2694 6156 2746
rect 10843 2694 10895 2746
rect 10907 2694 10959 2746
rect 10971 2694 11023 2746
rect 11035 2694 11087 2746
rect 4344 2635 4396 2644
rect 4344 2601 4353 2635
rect 4353 2601 4387 2635
rect 4387 2601 4396 2635
rect 4344 2592 4396 2601
rect 4896 2592 4948 2644
rect 5448 2635 5500 2644
rect 5448 2601 5457 2635
rect 5457 2601 5491 2635
rect 5491 2601 5500 2635
rect 5448 2592 5500 2601
rect 6920 2592 6972 2644
rect 7104 2635 7156 2644
rect 7104 2601 7113 2635
rect 7113 2601 7147 2635
rect 7147 2601 7156 2635
rect 7104 2592 7156 2601
rect 9772 2635 9824 2644
rect 9772 2601 9781 2635
rect 9781 2601 9815 2635
rect 9815 2601 9824 2635
rect 9772 2592 9824 2601
rect 9956 2592 10008 2644
rect 11152 2592 11204 2644
rect 12624 2635 12676 2644
rect 12624 2601 12633 2635
rect 12633 2601 12667 2635
rect 12667 2601 12676 2635
rect 12624 2592 12676 2601
rect 12992 2592 13044 2644
rect 13912 2592 13964 2644
rect 14372 2635 14424 2644
rect 14372 2601 14381 2635
rect 14381 2601 14415 2635
rect 14415 2601 14424 2635
rect 14372 2592 14424 2601
rect 2504 2524 2556 2576
rect 5264 2524 5316 2576
rect 1952 2456 2004 2508
rect 2780 2456 2832 2508
rect 7564 2524 7616 2576
rect 4988 2431 5040 2440
rect 4988 2397 4997 2431
rect 4997 2397 5031 2431
rect 5031 2397 5040 2431
rect 4988 2388 5040 2397
rect 6644 2388 6696 2440
rect 8668 2456 8720 2508
rect 10048 2524 10100 2576
rect 11060 2524 11112 2576
rect 204 2252 256 2304
rect 2044 2252 2096 2304
rect 7564 2252 7616 2304
rect 8208 2431 8260 2440
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 8208 2388 8260 2397
rect 9312 2431 9364 2440
rect 9312 2397 9321 2431
rect 9321 2397 9355 2431
rect 9355 2397 9364 2431
rect 9312 2388 9364 2397
rect 10600 2456 10652 2508
rect 10416 2431 10468 2440
rect 10416 2397 10425 2431
rect 10425 2397 10459 2431
rect 10459 2397 10468 2431
rect 10416 2388 10468 2397
rect 11612 2388 11664 2440
rect 12072 2456 12124 2508
rect 12808 2456 12860 2508
rect 13636 2499 13688 2508
rect 13636 2465 13645 2499
rect 13645 2465 13679 2499
rect 13679 2465 13688 2499
rect 13636 2456 13688 2465
rect 14924 2524 14976 2576
rect 14556 2456 14608 2508
rect 11980 2388 12032 2440
rect 12256 2388 12308 2440
rect 13176 2431 13228 2440
rect 13176 2397 13185 2431
rect 13185 2397 13219 2431
rect 13219 2397 13228 2431
rect 13176 2388 13228 2397
rect 9496 2252 9548 2304
rect 11336 2252 11388 2304
rect 15476 2320 15528 2372
rect 12532 2252 12584 2304
rect 3447 2150 3499 2202
rect 3511 2150 3563 2202
rect 3575 2150 3627 2202
rect 3639 2150 3691 2202
rect 8378 2150 8430 2202
rect 8442 2150 8494 2202
rect 8506 2150 8558 2202
rect 8570 2150 8622 2202
rect 13308 2150 13360 2202
rect 13372 2150 13424 2202
rect 13436 2150 13488 2202
rect 13500 2150 13552 2202
rect 11520 2048 11572 2100
rect 12992 2048 13044 2100
rect 7564 1980 7616 2032
rect 11704 1980 11756 2032
rect 12256 1980 12308 2032
rect 4068 1776 4120 1828
rect 14740 1776 14792 1828
rect 1860 1096 1912 1148
rect 7104 1096 7156 1148
<< metal2 >>
rect 202 19200 258 20000
rect 570 19200 626 20000
rect 938 19200 994 20000
rect 1398 19200 1454 20000
rect 1766 19200 1822 20000
rect 2226 19200 2282 20000
rect 2594 19200 2650 20000
rect 2870 19544 2926 19553
rect 2870 19479 2926 19488
rect 216 17542 244 19200
rect 204 17536 256 17542
rect 204 17478 256 17484
rect 584 15706 612 19200
rect 952 16794 980 19200
rect 940 16788 992 16794
rect 940 16730 992 16736
rect 1412 16726 1440 19200
rect 1584 17128 1636 17134
rect 1584 17070 1636 17076
rect 1400 16720 1452 16726
rect 1400 16662 1452 16668
rect 572 15700 624 15706
rect 572 15642 624 15648
rect 1492 14952 1544 14958
rect 1492 14894 1544 14900
rect 1400 14816 1452 14822
rect 1400 14758 1452 14764
rect 1412 12782 1440 14758
rect 1504 14482 1532 14894
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1596 13190 1624 17070
rect 1780 16810 1808 19200
rect 1780 16782 1900 16810
rect 1766 16688 1822 16697
rect 1676 16652 1728 16658
rect 1766 16623 1822 16632
rect 1676 16594 1728 16600
rect 1688 16561 1716 16594
rect 1674 16552 1730 16561
rect 1674 16487 1730 16496
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1582 12880 1638 12889
rect 1688 12850 1716 16487
rect 1780 16114 1808 16623
rect 1872 16250 1900 16782
rect 1860 16244 1912 16250
rect 1860 16186 1912 16192
rect 2240 16182 2268 19200
rect 2608 17354 2636 19200
rect 2608 17338 2820 17354
rect 2608 17332 2832 17338
rect 2608 17326 2780 17332
rect 2780 17274 2832 17280
rect 2884 17270 2912 19479
rect 2962 19200 3018 20000
rect 3422 19200 3478 20000
rect 3790 19200 3846 20000
rect 4250 19200 4306 20000
rect 4618 19200 4674 20000
rect 4986 19200 5042 20000
rect 5446 19200 5502 20000
rect 5814 19200 5870 20000
rect 6274 19200 6330 20000
rect 6642 19200 6698 20000
rect 7010 19200 7066 20000
rect 7470 19200 7526 20000
rect 7838 19200 7894 20000
rect 8298 19200 8354 20000
rect 8666 19200 8722 20000
rect 9034 19200 9090 20000
rect 9494 19200 9550 20000
rect 9862 19200 9918 20000
rect 10322 19200 10378 20000
rect 10690 19200 10746 20000
rect 11058 19200 11114 20000
rect 11518 19200 11574 20000
rect 11886 19200 11942 20000
rect 12346 19200 12402 20000
rect 12714 19200 12770 20000
rect 13082 19200 13138 20000
rect 13542 19200 13598 20000
rect 13910 19200 13966 20000
rect 14370 19200 14426 20000
rect 14738 19200 14794 20000
rect 15106 19200 15162 20000
rect 15566 19200 15622 20000
rect 15934 19200 15990 20000
rect 16394 19200 16450 20000
rect 16762 19200 16818 20000
rect 2976 17270 3004 19200
rect 3146 17640 3202 17649
rect 3436 17626 3464 19200
rect 3146 17575 3202 17584
rect 3344 17598 3464 17626
rect 2872 17264 2924 17270
rect 2872 17206 2924 17212
rect 2964 17264 3016 17270
rect 2964 17206 3016 17212
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2884 16658 2912 16934
rect 3160 16726 3188 17575
rect 3148 16720 3200 16726
rect 3148 16662 3200 16668
rect 2504 16652 2556 16658
rect 2504 16594 2556 16600
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2228 16176 2280 16182
rect 2228 16118 2280 16124
rect 2318 16144 2374 16153
rect 1768 16108 1820 16114
rect 2318 16079 2374 16088
rect 1768 16050 1820 16056
rect 2332 16046 2360 16079
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 1766 15736 1822 15745
rect 1766 15671 1822 15680
rect 1780 15638 1808 15671
rect 1768 15632 1820 15638
rect 1768 15574 1820 15580
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1964 14074 1992 14758
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 2332 13462 2360 15982
rect 2516 15484 2544 16594
rect 3344 16250 3372 17598
rect 3421 17436 3717 17456
rect 3477 17434 3501 17436
rect 3557 17434 3581 17436
rect 3637 17434 3661 17436
rect 3499 17382 3501 17434
rect 3563 17382 3575 17434
rect 3637 17382 3639 17434
rect 3477 17380 3501 17382
rect 3557 17380 3581 17382
rect 3637 17380 3661 17382
rect 3421 17360 3717 17380
rect 3421 16348 3717 16368
rect 3477 16346 3501 16348
rect 3557 16346 3581 16348
rect 3637 16346 3661 16348
rect 3499 16294 3501 16346
rect 3563 16294 3575 16346
rect 3637 16294 3639 16346
rect 3477 16292 3501 16294
rect 3557 16292 3581 16294
rect 3637 16292 3661 16294
rect 3421 16272 3717 16292
rect 3804 16250 3832 19200
rect 4066 18592 4122 18601
rect 4066 18527 4122 18536
rect 4080 18018 4108 18527
rect 4068 18012 4120 18018
rect 4068 17954 4120 17960
rect 3884 17128 3936 17134
rect 3884 17070 3936 17076
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 3792 16244 3844 16250
rect 3792 16186 3844 16192
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 2780 15972 2832 15978
rect 2780 15914 2832 15920
rect 2596 15904 2648 15910
rect 2596 15846 2648 15852
rect 2608 15638 2636 15846
rect 2596 15632 2648 15638
rect 2596 15574 2648 15580
rect 2792 15502 2820 15914
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 2780 15496 2832 15502
rect 2516 15456 2636 15484
rect 2608 14521 2636 15456
rect 2780 15438 2832 15444
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2792 14890 2820 15302
rect 2976 14958 3004 15438
rect 2964 14952 3016 14958
rect 2964 14894 3016 14900
rect 2780 14884 2832 14890
rect 2780 14826 2832 14832
rect 2976 14618 3004 14894
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 2594 14512 2650 14521
rect 2594 14447 2650 14456
rect 2688 14476 2740 14482
rect 2412 13728 2464 13734
rect 2412 13670 2464 13676
rect 2424 13530 2452 13670
rect 2412 13524 2464 13530
rect 2412 13466 2464 13472
rect 2320 13456 2372 13462
rect 2320 13398 2372 13404
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 1582 12815 1584 12824
rect 1636 12815 1638 12824
rect 1676 12844 1728 12850
rect 1584 12786 1636 12792
rect 1676 12786 1728 12792
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1400 12096 1452 12102
rect 1400 12038 1452 12044
rect 1412 11218 1440 12038
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1780 9654 1808 13330
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2228 13320 2280 13326
rect 2228 13262 2280 13268
rect 2148 11898 2176 13262
rect 2240 12306 2268 13262
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 2240 11354 2268 12242
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2332 10810 2360 11494
rect 2516 11286 2544 11698
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2320 10192 2372 10198
rect 2318 10160 2320 10169
rect 2372 10160 2374 10169
rect 2318 10095 2374 10104
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 1768 9648 1820 9654
rect 1768 9590 1820 9596
rect 1872 9518 1900 9862
rect 2516 9586 2544 11222
rect 2608 10470 2636 14447
rect 2688 14418 2740 14424
rect 2700 13870 2728 14418
rect 2976 13938 3004 14554
rect 3252 14278 3280 15506
rect 3240 14272 3292 14278
rect 3240 14214 3292 14220
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2688 13864 2740 13870
rect 3240 13864 3292 13870
rect 2688 13806 2740 13812
rect 2962 13832 3018 13841
rect 3240 13806 3292 13812
rect 2962 13767 3018 13776
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2884 12102 2912 12718
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2884 11762 2912 12038
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 1860 9512 1912 9518
rect 1860 9454 1912 9460
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 1674 9072 1730 9081
rect 1674 9007 1676 9016
rect 1728 9007 1730 9016
rect 1676 8978 1728 8984
rect 2424 8498 2452 9318
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 1492 8288 1544 8294
rect 1492 8230 1544 8236
rect 1504 7954 1532 8230
rect 2502 8120 2558 8129
rect 2502 8055 2558 8064
rect 2516 8022 2544 8055
rect 2504 8016 2556 8022
rect 2504 7958 2556 7964
rect 1492 7948 1544 7954
rect 1492 7890 1544 7896
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1400 7200 1452 7206
rect 1688 7177 1716 7822
rect 1400 7142 1452 7148
rect 1674 7168 1730 7177
rect 1412 5778 1440 7142
rect 1674 7103 1730 7112
rect 1768 6248 1820 6254
rect 1674 6216 1730 6225
rect 1820 6208 1900 6236
rect 1768 6190 1820 6196
rect 1674 6151 1730 6160
rect 1688 5846 1716 6151
rect 1676 5840 1728 5846
rect 1676 5782 1728 5788
rect 1768 5840 1820 5846
rect 1768 5782 1820 5788
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1780 5166 1808 5782
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 572 3392 624 3398
rect 572 3334 624 3340
rect 204 2304 256 2310
rect 204 2246 256 2252
rect 216 800 244 2246
rect 584 800 612 3334
rect 1412 2802 1440 4966
rect 1674 4312 1730 4321
rect 1674 4247 1730 4256
rect 1688 4146 1716 4247
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1872 3924 1900 6208
rect 2412 6180 2464 6186
rect 2412 6122 2464 6128
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 2240 4758 2268 5510
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2332 4826 2360 4966
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2228 4752 2280 4758
rect 2228 4694 2280 4700
rect 2424 4622 2452 6122
rect 2608 5710 2636 10406
rect 2792 10266 2820 11562
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2884 10033 2912 11086
rect 2976 10606 3004 13767
rect 3252 13326 3280 13806
rect 3344 13802 3372 15982
rect 3421 15260 3717 15280
rect 3477 15258 3501 15260
rect 3557 15258 3581 15260
rect 3637 15258 3661 15260
rect 3499 15206 3501 15258
rect 3563 15206 3575 15258
rect 3637 15206 3639 15258
rect 3477 15204 3501 15206
rect 3557 15204 3581 15206
rect 3637 15204 3661 15206
rect 3421 15184 3717 15204
rect 3422 14784 3478 14793
rect 3422 14719 3478 14728
rect 3436 14550 3464 14719
rect 3424 14544 3476 14550
rect 3424 14486 3476 14492
rect 3421 14172 3717 14192
rect 3477 14170 3501 14172
rect 3557 14170 3581 14172
rect 3637 14170 3661 14172
rect 3499 14118 3501 14170
rect 3563 14118 3575 14170
rect 3637 14118 3639 14170
rect 3477 14116 3501 14118
rect 3557 14116 3581 14118
rect 3637 14116 3661 14118
rect 3421 14096 3717 14116
rect 3332 13796 3384 13802
rect 3332 13738 3384 13744
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3160 12986 3188 13262
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3252 12442 3280 12718
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3238 11928 3294 11937
rect 3238 11863 3294 11872
rect 3148 11688 3200 11694
rect 3148 11630 3200 11636
rect 3160 10674 3188 11630
rect 3252 11626 3280 11863
rect 3240 11620 3292 11626
rect 3240 11562 3292 11568
rect 3344 11121 3372 13738
rect 3421 13084 3717 13104
rect 3477 13082 3501 13084
rect 3557 13082 3581 13084
rect 3637 13082 3661 13084
rect 3499 13030 3501 13082
rect 3563 13030 3575 13082
rect 3637 13030 3639 13082
rect 3477 13028 3501 13030
rect 3557 13028 3581 13030
rect 3637 13028 3661 13030
rect 3421 13008 3717 13028
rect 3804 12986 3832 15982
rect 3896 13462 3924 17070
rect 4160 17060 4212 17066
rect 4160 17002 4212 17008
rect 3976 15632 4028 15638
rect 3976 15574 4028 15580
rect 3988 14074 4016 15574
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4080 14550 4108 15098
rect 4068 14544 4120 14550
rect 4068 14486 4120 14492
rect 4172 14498 4200 17002
rect 4264 16794 4292 19200
rect 4632 17338 4660 19200
rect 4620 17332 4672 17338
rect 5000 17320 5028 19200
rect 5356 17604 5408 17610
rect 5356 17546 5408 17552
rect 5080 17332 5132 17338
rect 5000 17292 5080 17320
rect 4620 17274 4672 17280
rect 5080 17274 5132 17280
rect 5368 17134 5396 17546
rect 5460 17320 5488 19200
rect 5632 17332 5684 17338
rect 5460 17292 5632 17320
rect 5632 17274 5684 17280
rect 5828 17270 5856 19200
rect 5816 17264 5868 17270
rect 5816 17206 5868 17212
rect 5356 17128 5408 17134
rect 5356 17070 5408 17076
rect 5886 16892 6182 16912
rect 5942 16890 5966 16892
rect 6022 16890 6046 16892
rect 6102 16890 6126 16892
rect 5964 16838 5966 16890
rect 6028 16838 6040 16890
rect 6102 16838 6104 16890
rect 5942 16836 5966 16838
rect 6022 16836 6046 16838
rect 6102 16836 6126 16838
rect 5886 16816 6182 16836
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 5724 16720 5776 16726
rect 5724 16662 5776 16668
rect 5356 16448 5408 16454
rect 5356 16390 5408 16396
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 4344 15564 4396 15570
rect 4344 15506 4396 15512
rect 4356 15162 4384 15506
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4172 14470 4292 14498
rect 4160 14408 4212 14414
rect 4066 14376 4122 14385
rect 4160 14350 4212 14356
rect 4066 14311 4122 14320
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 3884 13456 3936 13462
rect 3884 13398 3936 13404
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3421 11996 3717 12016
rect 3477 11994 3501 11996
rect 3557 11994 3581 11996
rect 3637 11994 3661 11996
rect 3499 11942 3501 11994
rect 3563 11942 3575 11994
rect 3637 11942 3639 11994
rect 3477 11940 3501 11942
rect 3557 11940 3581 11942
rect 3637 11940 3661 11942
rect 3421 11920 3717 11940
rect 3330 11112 3386 11121
rect 3330 11047 3386 11056
rect 3240 11008 3292 11014
rect 3238 10976 3240 10985
rect 3292 10976 3294 10985
rect 3238 10911 3294 10920
rect 3421 10908 3717 10928
rect 3477 10906 3501 10908
rect 3557 10906 3581 10908
rect 3637 10906 3661 10908
rect 3499 10854 3501 10906
rect 3563 10854 3575 10906
rect 3637 10854 3639 10906
rect 3477 10852 3501 10854
rect 3557 10852 3581 10854
rect 3637 10852 3661 10854
rect 3421 10832 3717 10852
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 3160 10062 3188 10610
rect 3436 10062 3464 10610
rect 3804 10538 3832 12038
rect 3792 10532 3844 10538
rect 3792 10474 3844 10480
rect 3896 10130 3924 13398
rect 3976 13184 4028 13190
rect 4080 13172 4108 14311
rect 4172 14074 4200 14350
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4264 13410 4292 14470
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4028 13144 4108 13172
rect 4172 13382 4292 13410
rect 3976 13126 4028 13132
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3148 10056 3200 10062
rect 2870 10024 2926 10033
rect 3332 10056 3384 10062
rect 3148 9998 3200 10004
rect 3252 10004 3332 10010
rect 3252 9998 3384 10004
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 2870 9959 2926 9968
rect 3252 9982 3372 9998
rect 3148 9716 3200 9722
rect 3252 9704 3280 9982
rect 3421 9820 3717 9840
rect 3477 9818 3501 9820
rect 3557 9818 3581 9820
rect 3637 9818 3661 9820
rect 3499 9766 3501 9818
rect 3563 9766 3575 9818
rect 3637 9766 3639 9818
rect 3477 9764 3501 9766
rect 3557 9764 3581 9766
rect 3637 9764 3661 9766
rect 3421 9744 3717 9764
rect 3200 9676 3280 9704
rect 3148 9658 3200 9664
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2792 9110 2820 9454
rect 2780 9104 2832 9110
rect 2780 9046 2832 9052
rect 2792 7324 2820 9046
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 2976 8090 3004 8298
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2872 7336 2924 7342
rect 2792 7296 2872 7324
rect 2792 6662 2820 7296
rect 2872 7278 2924 7284
rect 3056 7268 3108 7274
rect 3056 7210 3108 7216
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2596 5704 2648 5710
rect 2594 5672 2596 5681
rect 2688 5704 2740 5710
rect 2648 5672 2650 5681
rect 2688 5646 2740 5652
rect 2594 5607 2650 5616
rect 2700 5234 2728 5646
rect 2778 5264 2834 5273
rect 2688 5228 2740 5234
rect 2778 5199 2834 5208
rect 2688 5170 2740 5176
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2516 4282 2544 4966
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 2228 4072 2280 4078
rect 2228 4014 2280 4020
rect 1952 3936 2004 3942
rect 1872 3896 1952 3924
rect 1952 3878 2004 3884
rect 1964 3602 1992 3878
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1674 3360 1730 3369
rect 1674 3295 1730 3304
rect 1688 3058 1716 3295
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1044 2774 1440 2802
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 1044 800 1072 2774
rect 1504 2530 1532 2790
rect 1412 2502 1532 2530
rect 1964 2514 1992 3538
rect 2240 3194 2268 4014
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 2228 2984 2280 2990
rect 2228 2926 2280 2932
rect 1952 2508 2004 2514
rect 1412 800 1440 2502
rect 1952 2450 2004 2456
rect 2056 2310 2084 2926
rect 2044 2304 2096 2310
rect 2044 2246 2096 2252
rect 1860 1148 1912 1154
rect 1860 1090 1912 1096
rect 1872 800 1900 1090
rect 2240 800 2268 2926
rect 2516 2582 2544 4218
rect 2792 4078 2820 5199
rect 2884 4826 2912 7142
rect 3068 7002 3096 7210
rect 3056 6996 3108 7002
rect 3056 6938 3108 6944
rect 3252 5846 3280 9676
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 3516 9444 3568 9450
rect 3516 9386 3568 9392
rect 3528 9178 3556 9386
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3804 9178 3832 9318
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3528 8922 3556 9114
rect 3896 9110 3924 9590
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3896 8974 3924 9046
rect 3344 8894 3556 8922
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 3344 8498 3372 8894
rect 3421 8732 3717 8752
rect 3477 8730 3501 8732
rect 3557 8730 3581 8732
rect 3637 8730 3661 8732
rect 3499 8678 3501 8730
rect 3563 8678 3575 8730
rect 3637 8678 3639 8730
rect 3477 8676 3501 8678
rect 3557 8676 3581 8678
rect 3637 8676 3661 8678
rect 3421 8656 3717 8676
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3344 7954 3372 8434
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3804 8090 3832 8230
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3896 7818 3924 8910
rect 3884 7812 3936 7818
rect 3884 7754 3936 7760
rect 3421 7644 3717 7664
rect 3477 7642 3501 7644
rect 3557 7642 3581 7644
rect 3637 7642 3661 7644
rect 3499 7590 3501 7642
rect 3563 7590 3575 7642
rect 3637 7590 3639 7642
rect 3477 7588 3501 7590
rect 3557 7588 3581 7590
rect 3637 7588 3661 7590
rect 3421 7568 3717 7588
rect 3421 6556 3717 6576
rect 3477 6554 3501 6556
rect 3557 6554 3581 6556
rect 3637 6554 3661 6556
rect 3499 6502 3501 6554
rect 3563 6502 3575 6554
rect 3637 6502 3639 6554
rect 3477 6500 3501 6502
rect 3557 6500 3581 6502
rect 3637 6500 3661 6502
rect 3421 6480 3717 6500
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3240 5840 3292 5846
rect 3240 5782 3292 5788
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2504 2576 2556 2582
rect 2504 2518 2556 2524
rect 2700 800 2728 3130
rect 2976 2854 3004 4966
rect 3344 4826 3372 6054
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3421 5468 3717 5488
rect 3477 5466 3501 5468
rect 3557 5466 3581 5468
rect 3637 5466 3661 5468
rect 3499 5414 3501 5466
rect 3563 5414 3575 5466
rect 3637 5414 3639 5466
rect 3477 5412 3501 5414
rect 3557 5412 3581 5414
rect 3637 5412 3661 5414
rect 3421 5392 3717 5412
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 2964 2848 3016 2854
rect 2964 2790 3016 2796
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2792 1465 2820 2450
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 3068 800 3096 4490
rect 3421 4380 3717 4400
rect 3477 4378 3501 4380
rect 3557 4378 3581 4380
rect 3637 4378 3661 4380
rect 3499 4326 3501 4378
rect 3563 4326 3575 4378
rect 3637 4326 3639 4378
rect 3477 4324 3501 4326
rect 3557 4324 3581 4326
rect 3637 4324 3661 4326
rect 3421 4304 3717 4324
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 3700 4004 3752 4010
rect 3700 3946 3752 3952
rect 3240 3664 3292 3670
rect 3240 3606 3292 3612
rect 3252 2938 3280 3606
rect 3344 3398 3372 3946
rect 3712 3602 3740 3946
rect 3804 3942 3832 5102
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 3804 3534 3832 3878
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3344 3058 3372 3334
rect 3421 3292 3717 3312
rect 3477 3290 3501 3292
rect 3557 3290 3581 3292
rect 3637 3290 3661 3292
rect 3499 3238 3501 3290
rect 3563 3238 3575 3290
rect 3637 3238 3639 3290
rect 3477 3236 3501 3238
rect 3557 3236 3581 3238
rect 3637 3236 3661 3238
rect 3421 3216 3717 3236
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 3436 2938 3464 2994
rect 3252 2910 3464 2938
rect 3421 2204 3717 2224
rect 3477 2202 3501 2204
rect 3557 2202 3581 2204
rect 3637 2202 3661 2204
rect 3499 2150 3501 2202
rect 3563 2150 3575 2202
rect 3637 2150 3639 2202
rect 3477 2148 3501 2150
rect 3557 2148 3581 2150
rect 3637 2148 3661 2150
rect 3421 2128 3717 2148
rect 3804 1442 3832 3334
rect 3528 1414 3832 1442
rect 3528 800 3556 1414
rect 3896 800 3924 5510
rect 3988 2836 4016 13126
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 4080 7993 4108 12922
rect 4066 7984 4122 7993
rect 4172 7954 4200 13382
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4264 12306 4292 12582
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 4264 10606 4292 12106
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4356 10470 4384 14214
rect 4540 13938 4568 14962
rect 4804 14952 4856 14958
rect 4802 14920 4804 14929
rect 4856 14920 4858 14929
rect 4802 14855 4858 14864
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4724 13938 4752 14758
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 4540 12986 4568 13874
rect 4712 13796 4764 13802
rect 4712 13738 4764 13744
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4632 12442 4660 13126
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4448 11898 4476 12242
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4528 10532 4580 10538
rect 4528 10474 4580 10480
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4540 10266 4568 10474
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4264 8498 4292 8978
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4356 8362 4384 9862
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4448 8634 4476 9318
rect 4540 9042 4568 9930
rect 4632 9518 4660 11494
rect 4724 10470 4752 13738
rect 4816 11014 4844 14855
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 4896 13864 4948 13870
rect 4948 13824 5028 13852
rect 4896 13806 4948 13812
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 4908 11558 4936 11698
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4264 8090 4292 8230
rect 4342 8120 4398 8129
rect 4252 8084 4304 8090
rect 4342 8055 4398 8064
rect 4252 8026 4304 8032
rect 4356 8022 4384 8055
rect 4344 8016 4396 8022
rect 4344 7958 4396 7964
rect 4066 7919 4122 7928
rect 4160 7948 4212 7954
rect 4080 6254 4108 7919
rect 4160 7890 4212 7896
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4172 6866 4200 7346
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4172 6458 4200 6802
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4080 5914 4108 6054
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 4172 4622 4200 6394
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4356 5574 4384 5850
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4264 2990 4292 4422
rect 4448 4146 4476 8298
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4540 3738 4568 6598
rect 4632 5846 4660 9318
rect 4724 6662 4752 9454
rect 4816 9178 4844 10066
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4816 8129 4844 8230
rect 4802 8120 4858 8129
rect 4802 8055 4858 8064
rect 4908 8004 4936 11494
rect 4816 7976 4936 8004
rect 4816 6882 4844 7976
rect 5000 7290 5028 13824
rect 5092 12306 5120 14010
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 5184 11762 5212 15982
rect 5368 15570 5396 16390
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 5262 15464 5318 15473
rect 5262 15399 5318 15408
rect 5276 14006 5304 15399
rect 5368 15162 5396 15506
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5368 14906 5396 15098
rect 5368 14890 5488 14906
rect 5552 14890 5580 16050
rect 5736 15434 5764 16662
rect 6288 16250 6316 19200
rect 6552 17060 6604 17066
rect 6552 17002 6604 17008
rect 6368 16720 6420 16726
rect 6368 16662 6420 16668
rect 6276 16244 6328 16250
rect 6276 16186 6328 16192
rect 6380 16114 6408 16662
rect 6460 16176 6512 16182
rect 6460 16118 6512 16124
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 5886 15804 6182 15824
rect 5942 15802 5966 15804
rect 6022 15802 6046 15804
rect 6102 15802 6126 15804
rect 5964 15750 5966 15802
rect 6028 15750 6040 15802
rect 6102 15750 6104 15802
rect 5942 15748 5966 15750
rect 6022 15748 6046 15750
rect 6102 15748 6126 15750
rect 5886 15728 6182 15748
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 5724 15428 5776 15434
rect 5724 15370 5776 15376
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 5368 14884 5500 14890
rect 5368 14878 5448 14884
rect 5448 14826 5500 14832
rect 5540 14884 5592 14890
rect 5540 14826 5592 14832
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5264 14000 5316 14006
rect 5264 13942 5316 13948
rect 5368 13530 5396 14758
rect 5460 14006 5488 14826
rect 5448 14000 5500 14006
rect 5448 13942 5500 13948
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5552 13410 5580 14826
rect 5644 13512 5672 14962
rect 5724 14816 5776 14822
rect 5724 14758 5776 14764
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5736 14618 5764 14758
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5736 13938 5764 14214
rect 5828 14074 5856 14758
rect 5886 14716 6182 14736
rect 5942 14714 5966 14716
rect 6022 14714 6046 14716
rect 6102 14714 6126 14716
rect 5964 14662 5966 14714
rect 6028 14662 6040 14714
rect 6102 14662 6104 14714
rect 5942 14660 5966 14662
rect 6022 14660 6046 14662
rect 6102 14660 6126 14662
rect 5886 14640 6182 14660
rect 6276 14612 6328 14618
rect 6276 14554 6328 14560
rect 6288 14521 6316 14554
rect 6274 14512 6330 14521
rect 6274 14447 6330 14456
rect 6184 14340 6236 14346
rect 6184 14282 6236 14288
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5816 13864 5868 13870
rect 5920 13852 5948 14010
rect 6196 13938 6224 14282
rect 6184 13932 6236 13938
rect 6236 13892 6316 13920
rect 6184 13874 6236 13880
rect 5868 13824 5948 13852
rect 5816 13806 5868 13812
rect 5886 13628 6182 13648
rect 5942 13626 5966 13628
rect 6022 13626 6046 13628
rect 6102 13626 6126 13628
rect 5964 13574 5966 13626
rect 6028 13574 6040 13626
rect 6102 13574 6104 13626
rect 5942 13572 5966 13574
rect 6022 13572 6046 13574
rect 6102 13572 6126 13574
rect 5886 13552 6182 13572
rect 5644 13484 5948 13512
rect 5356 13388 5408 13394
rect 5552 13382 5672 13410
rect 5356 13330 5408 13336
rect 5368 12986 5396 13330
rect 5540 13252 5592 13258
rect 5540 13194 5592 13200
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 5276 11286 5304 12038
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5264 11280 5316 11286
rect 5264 11222 5316 11228
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 5092 10198 5120 10950
rect 5460 10810 5488 11698
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5552 10606 5580 13194
rect 5644 12889 5672 13382
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5630 12880 5686 12889
rect 5630 12815 5686 12824
rect 5736 12442 5764 13262
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5828 12850 5856 13126
rect 5920 12918 5948 13484
rect 6288 13326 6316 13892
rect 6380 13802 6408 15506
rect 6368 13796 6420 13802
rect 6368 13738 6420 13744
rect 6472 13530 6500 16118
rect 6564 15570 6592 17002
rect 6656 15706 6684 19200
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6736 16652 6788 16658
rect 6736 16594 6788 16600
rect 6644 15700 6696 15706
rect 6644 15642 6696 15648
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 6460 13524 6512 13530
rect 6460 13466 6512 13472
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 5908 12912 5960 12918
rect 5908 12854 5960 12860
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 5920 12628 5948 12854
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 5828 12600 5948 12628
rect 6380 12617 6408 12718
rect 6366 12608 6422 12617
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5828 12306 5856 12600
rect 5886 12540 6182 12560
rect 6366 12543 6422 12552
rect 5942 12538 5966 12540
rect 6022 12538 6046 12540
rect 6102 12538 6126 12540
rect 5964 12486 5966 12538
rect 6028 12486 6040 12538
rect 6102 12486 6104 12538
rect 5942 12484 5966 12486
rect 6022 12484 6046 12486
rect 6102 12484 6126 12486
rect 5886 12464 6182 12484
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 6288 11762 6316 12378
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6276 11756 6328 11762
rect 6276 11698 6328 11704
rect 5632 11620 5684 11626
rect 5632 11562 5684 11568
rect 5644 10674 5672 11562
rect 5886 11452 6182 11472
rect 5942 11450 5966 11452
rect 6022 11450 6046 11452
rect 6102 11450 6126 11452
rect 5964 11398 5966 11450
rect 6028 11398 6040 11450
rect 6102 11398 6104 11450
rect 5942 11396 5966 11398
rect 6022 11396 6046 11398
rect 6102 11396 6126 11398
rect 5886 11376 6182 11396
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5080 10192 5132 10198
rect 5080 10134 5132 10140
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 5092 9586 5120 9998
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 5092 8498 5120 9522
rect 5184 9382 5212 10406
rect 5356 10192 5408 10198
rect 5262 10160 5318 10169
rect 5356 10134 5408 10140
rect 5262 10095 5318 10104
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 5080 8356 5132 8362
rect 5184 8344 5212 9318
rect 5132 8316 5212 8344
rect 5080 8298 5132 8304
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 4896 7268 4948 7274
rect 5000 7262 5120 7290
rect 4896 7210 4948 7216
rect 4908 7002 4936 7210
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4816 6854 4936 6882
rect 4802 6760 4858 6769
rect 4802 6695 4858 6704
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4816 5914 4844 6695
rect 4908 6118 4936 6854
rect 5000 6458 5028 7142
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4908 5914 4936 6054
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4620 5840 4672 5846
rect 4620 5782 4672 5788
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4632 5166 4660 5646
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4632 4282 4660 5102
rect 5092 4690 5120 7262
rect 5184 5234 5212 8026
rect 5276 6866 5304 10095
rect 5368 7970 5396 10134
rect 5460 10130 5488 10542
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5736 8634 5764 11290
rect 6184 11280 6236 11286
rect 5828 11240 6184 11268
rect 5828 10198 5856 11240
rect 6184 11222 6236 11228
rect 5886 10364 6182 10384
rect 5942 10362 5966 10364
rect 6022 10362 6046 10364
rect 6102 10362 6126 10364
rect 5964 10310 5966 10362
rect 6028 10310 6040 10362
rect 6102 10310 6104 10362
rect 5942 10308 5966 10310
rect 6022 10308 6046 10310
rect 6102 10308 6126 10310
rect 5886 10288 6182 10308
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 6288 10130 6316 11290
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5828 8498 5856 9318
rect 5886 9276 6182 9296
rect 5942 9274 5966 9276
rect 6022 9274 6046 9276
rect 6102 9274 6126 9276
rect 5964 9222 5966 9274
rect 6028 9222 6040 9274
rect 6102 9222 6104 9274
rect 5942 9220 5966 9222
rect 6022 9220 6046 9222
rect 6102 9220 6126 9222
rect 5886 9200 6182 9220
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5460 8090 5488 8434
rect 6380 8362 6408 11834
rect 6472 11558 6500 13466
rect 6564 12646 6592 14894
rect 6644 13252 6696 13258
rect 6644 13194 6696 13200
rect 6656 12782 6684 13194
rect 6748 12918 6776 16594
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6840 12782 6868 17070
rect 7024 16250 7052 19200
rect 7484 16674 7512 19200
rect 7852 17338 7880 19200
rect 8312 17626 8340 19200
rect 8680 17762 8708 19200
rect 8680 17734 8892 17762
rect 8312 17598 8800 17626
rect 8352 17436 8648 17456
rect 8408 17434 8432 17436
rect 8488 17434 8512 17436
rect 8568 17434 8592 17436
rect 8430 17382 8432 17434
rect 8494 17382 8506 17434
rect 8568 17382 8570 17434
rect 8408 17380 8432 17382
rect 8488 17380 8512 17382
rect 8568 17380 8592 17382
rect 8352 17360 8648 17380
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8312 16726 8340 16934
rect 8404 16794 8432 17138
rect 8668 16992 8720 16998
rect 8668 16934 8720 16940
rect 8680 16794 8708 16934
rect 8392 16788 8444 16794
rect 8668 16788 8720 16794
rect 8444 16748 8616 16776
rect 8392 16730 8444 16736
rect 8300 16720 8352 16726
rect 7484 16646 7696 16674
rect 8300 16662 8352 16668
rect 7668 16454 7696 16646
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 8588 16538 8616 16748
rect 8668 16730 8720 16736
rect 8024 16516 8076 16522
rect 8024 16458 8076 16464
rect 7656 16448 7708 16454
rect 7656 16390 7708 16396
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7024 15706 7052 15846
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 7208 14521 7236 15506
rect 7300 15162 7328 15846
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7392 14618 7420 14894
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7194 14512 7250 14521
rect 7012 14476 7064 14482
rect 7484 14482 7512 15642
rect 7668 15434 7696 16050
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7656 15428 7708 15434
rect 7656 15370 7708 15376
rect 7746 15056 7802 15065
rect 7746 14991 7748 15000
rect 7800 14991 7802 15000
rect 7748 14962 7800 14968
rect 7194 14447 7250 14456
rect 7472 14476 7524 14482
rect 7012 14418 7064 14424
rect 7472 14418 7524 14424
rect 6644 12776 6696 12782
rect 6644 12718 6696 12724
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6918 12744 6974 12753
rect 6918 12679 6974 12688
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 6460 11552 6512 11558
rect 6512 11512 6592 11540
rect 6460 11494 6512 11500
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6472 8498 6500 11154
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5368 7942 5488 7970
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5368 6322 5396 6734
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5368 5370 5396 6258
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5460 5250 5488 7942
rect 5552 7546 5580 8298
rect 5886 8188 6182 8208
rect 5942 8186 5966 8188
rect 6022 8186 6046 8188
rect 6102 8186 6126 8188
rect 5964 8134 5966 8186
rect 6028 8134 6040 8186
rect 6102 8134 6104 8186
rect 5942 8132 5966 8134
rect 6022 8132 6046 8134
rect 6102 8132 6126 8134
rect 5886 8112 6182 8132
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 6196 7410 6224 7890
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 5886 7100 6182 7120
rect 5942 7098 5966 7100
rect 6022 7098 6046 7100
rect 6102 7098 6126 7100
rect 5964 7046 5966 7098
rect 6028 7046 6040 7098
rect 6102 7046 6104 7098
rect 5942 7044 5966 7046
rect 6022 7044 6046 7046
rect 6102 7044 6126 7046
rect 5886 7024 6182 7044
rect 6288 7002 6316 7142
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5368 5222 5488 5250
rect 5184 4826 5212 5170
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4344 3664 4396 3670
rect 4344 3606 4396 3612
rect 4434 3632 4490 3641
rect 4356 3058 4384 3606
rect 4434 3567 4436 3576
rect 4488 3567 4490 3576
rect 4436 3538 4488 3544
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 4252 2984 4304 2990
rect 4632 2972 4660 4082
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4724 3126 4752 3878
rect 4816 3194 4844 4422
rect 4894 4040 4950 4049
rect 4894 3975 4950 3984
rect 4988 4004 5040 4010
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 4802 3088 4858 3097
rect 4802 3023 4858 3032
rect 4712 2984 4764 2990
rect 4632 2952 4712 2972
rect 4764 2952 4766 2961
rect 4632 2944 4710 2952
rect 4252 2926 4304 2932
rect 4344 2916 4396 2922
rect 4344 2858 4396 2864
rect 4436 2916 4488 2922
rect 4710 2887 4766 2896
rect 4436 2858 4488 2864
rect 3988 2808 4200 2836
rect 4066 2408 4122 2417
rect 4066 2343 4122 2352
rect 4080 1834 4108 2343
rect 4068 1828 4120 1834
rect 4068 1770 4120 1776
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1398 0 1454 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2686 0 2742 800
rect 3054 0 3110 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4172 513 4200 2808
rect 4356 2650 4384 2858
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4448 1442 4476 2858
rect 4356 1414 4476 1442
rect 4356 800 4384 1414
rect 4816 898 4844 3023
rect 4908 2650 4936 3975
rect 4988 3946 5040 3952
rect 5000 3738 5028 3946
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 5000 3058 5028 3538
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 5000 2446 5028 2994
rect 5092 2854 5120 4626
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 5184 3194 5212 3878
rect 5276 3670 5304 4082
rect 5368 4049 5396 5222
rect 5354 4040 5410 4049
rect 5354 3975 5410 3984
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 4724 870 4844 898
rect 4724 800 4752 870
rect 5184 800 5212 2994
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 5276 2582 5304 2790
rect 5460 2650 5488 3946
rect 5644 3058 5672 6598
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6182 6216 6238 6225
rect 6182 6151 6184 6160
rect 6236 6151 6238 6160
rect 6276 6180 6328 6186
rect 6184 6122 6236 6128
rect 6276 6122 6328 6128
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5736 4146 5764 4966
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5828 4078 5856 6054
rect 5886 6012 6182 6032
rect 5942 6010 5966 6012
rect 6022 6010 6046 6012
rect 6102 6010 6126 6012
rect 5964 5958 5966 6010
rect 6028 5958 6040 6010
rect 6102 5958 6104 6010
rect 5942 5956 5966 5958
rect 6022 5956 6046 5958
rect 6102 5956 6126 5958
rect 5886 5936 6182 5956
rect 6288 5778 6316 6122
rect 6380 5846 6408 6258
rect 6564 6118 6592 11512
rect 6748 11354 6776 12174
rect 6840 11694 6868 12582
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6932 11540 6960 12679
rect 7024 11778 7052 14418
rect 7196 13796 7248 13802
rect 7196 13738 7248 13744
rect 7208 13682 7236 13738
rect 7116 13654 7236 13682
rect 7472 13728 7524 13734
rect 7472 13670 7524 13676
rect 7116 12050 7144 13654
rect 7484 12850 7512 13670
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7208 12374 7236 12718
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7116 12022 7328 12050
rect 7024 11750 7144 11778
rect 6840 11512 6960 11540
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6656 8498 6684 8910
rect 6748 8634 6776 10746
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6840 8514 6868 11512
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6932 9450 6960 11086
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 7024 10198 7052 10950
rect 7012 10192 7064 10198
rect 7012 10134 7064 10140
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6748 8486 6868 8514
rect 6748 6769 6776 8486
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6840 7546 6868 8366
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 6734 6760 6790 6769
rect 6734 6695 6790 6704
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6748 6254 6776 6598
rect 6736 6248 6788 6254
rect 6642 6216 6698 6225
rect 6736 6190 6788 6196
rect 6642 6151 6698 6160
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6368 5840 6420 5846
rect 6368 5782 6420 5788
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 5886 4924 6182 4944
rect 5942 4922 5966 4924
rect 6022 4922 6046 4924
rect 6102 4922 6126 4924
rect 5964 4870 5966 4922
rect 6028 4870 6040 4922
rect 6102 4870 6104 4922
rect 5942 4868 5966 4870
rect 6022 4868 6046 4870
rect 6102 4868 6126 4870
rect 5886 4848 6182 4868
rect 6288 4826 6316 5714
rect 6380 5234 6408 5782
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6276 4820 6328 4826
rect 6328 4780 6408 4808
rect 6276 4762 6328 4768
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5828 3398 5856 3878
rect 5886 3836 6182 3856
rect 5942 3834 5966 3836
rect 6022 3834 6046 3836
rect 6102 3834 6126 3836
rect 5964 3782 5966 3834
rect 6028 3782 6040 3834
rect 6102 3782 6104 3834
rect 5942 3780 5966 3782
rect 6022 3780 6046 3782
rect 6102 3780 6126 3782
rect 5886 3760 6182 3780
rect 6380 3641 6408 4780
rect 6564 4690 6592 6054
rect 6656 5658 6684 6151
rect 6656 5630 6776 5658
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6656 4758 6684 5510
rect 6644 4752 6696 4758
rect 6644 4694 6696 4700
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6656 4214 6684 4694
rect 6644 4208 6696 4214
rect 6644 4150 6696 4156
rect 6748 4078 6776 5630
rect 6840 5234 6868 6870
rect 6920 6860 6972 6866
rect 7024 6848 7052 10134
rect 7116 9722 7144 11750
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 7208 10674 7236 11562
rect 7300 10742 7328 12022
rect 7484 11762 7512 12786
rect 7564 12368 7616 12374
rect 7564 12310 7616 12316
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7576 11014 7604 12310
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7288 10736 7340 10742
rect 7288 10678 7340 10684
rect 7564 10736 7616 10742
rect 7564 10678 7616 10684
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7196 10532 7248 10538
rect 7196 10474 7248 10480
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7208 7970 7236 10474
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 7300 8090 7328 8298
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7208 7942 7328 7970
rect 7300 7886 7328 7942
rect 7392 7886 7420 8978
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7196 7200 7248 7206
rect 7248 7160 7328 7188
rect 7196 7142 7248 7148
rect 6972 6820 7052 6848
rect 7104 6860 7156 6866
rect 6920 6802 6972 6808
rect 7104 6802 7156 6808
rect 7116 5914 7144 6802
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7208 5914 7236 6734
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7300 5817 7328 7160
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7392 6186 7420 6734
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 7286 5808 7342 5817
rect 7484 5778 7512 9862
rect 7576 8537 7604 10678
rect 7668 9654 7696 13330
rect 7852 12646 7880 15982
rect 7932 15700 7984 15706
rect 8036 15688 8064 16458
rect 8128 16182 8156 16526
rect 8588 16510 8708 16538
rect 8352 16348 8648 16368
rect 8408 16346 8432 16348
rect 8488 16346 8512 16348
rect 8568 16346 8592 16348
rect 8430 16294 8432 16346
rect 8494 16294 8506 16346
rect 8568 16294 8570 16346
rect 8408 16292 8432 16294
rect 8488 16292 8512 16294
rect 8568 16292 8592 16294
rect 8352 16272 8648 16292
rect 8116 16176 8168 16182
rect 8116 16118 8168 16124
rect 8680 16046 8708 16510
rect 8392 16040 8444 16046
rect 8668 16040 8720 16046
rect 8444 15988 8524 15994
rect 8392 15982 8524 15988
rect 8668 15982 8720 15988
rect 8404 15966 8524 15982
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8496 15858 8524 15966
rect 7984 15660 8064 15688
rect 7932 15642 7984 15648
rect 8404 15638 8432 15846
rect 8496 15830 8708 15858
rect 8392 15632 8444 15638
rect 8392 15574 8444 15580
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 8036 15162 8064 15438
rect 8024 15156 8076 15162
rect 8024 15098 8076 15104
rect 8036 15026 8064 15098
rect 8024 15020 8076 15026
rect 8024 14962 8076 14968
rect 7932 14816 7984 14822
rect 7932 14758 7984 14764
rect 7944 14618 7972 14758
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 8128 14482 8156 15506
rect 8352 15260 8648 15280
rect 8408 15258 8432 15260
rect 8488 15258 8512 15260
rect 8568 15258 8592 15260
rect 8430 15206 8432 15258
rect 8494 15206 8506 15258
rect 8568 15206 8570 15258
rect 8408 15204 8432 15206
rect 8488 15204 8512 15206
rect 8568 15204 8592 15206
rect 8352 15184 8648 15204
rect 8576 14952 8628 14958
rect 8680 14906 8708 15830
rect 8772 15434 8800 17598
rect 8864 15570 8892 17734
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 8956 16522 8984 17614
rect 9048 16998 9076 19200
rect 9508 17678 9536 19200
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 9876 17082 9904 19200
rect 10232 17128 10284 17134
rect 9876 17054 9996 17082
rect 10232 17070 10284 17076
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 8944 16516 8996 16522
rect 8944 16458 8996 16464
rect 9048 16402 9076 16934
rect 9140 16561 9168 16934
rect 9496 16720 9548 16726
rect 9496 16662 9548 16668
rect 9126 16552 9182 16561
rect 9126 16487 9182 16496
rect 9048 16374 9260 16402
rect 9036 16244 9088 16250
rect 9036 16186 9088 16192
rect 9048 15570 9076 16186
rect 9128 16040 9180 16046
rect 9128 15982 9180 15988
rect 8852 15564 8904 15570
rect 8852 15506 8904 15512
rect 9036 15564 9088 15570
rect 9036 15506 9088 15512
rect 8760 15428 8812 15434
rect 8760 15370 8812 15376
rect 9140 15042 9168 15982
rect 9048 15014 9168 15042
rect 8628 14900 8708 14906
rect 8576 14894 8708 14900
rect 8588 14878 8708 14894
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8128 13802 8156 14418
rect 8352 14172 8648 14192
rect 8408 14170 8432 14172
rect 8488 14170 8512 14172
rect 8568 14170 8592 14172
rect 8430 14118 8432 14170
rect 8494 14118 8506 14170
rect 8568 14118 8570 14170
rect 8408 14116 8432 14118
rect 8488 14116 8512 14118
rect 8568 14116 8592 14118
rect 8352 14096 8648 14116
rect 8680 13870 8708 14878
rect 8758 14920 8814 14929
rect 8758 14855 8814 14864
rect 8944 14884 8996 14890
rect 8772 14618 8800 14855
rect 8944 14826 8996 14832
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 8850 14512 8906 14521
rect 8850 14447 8906 14456
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 8116 13796 8168 13802
rect 8116 13738 8168 13744
rect 8352 13084 8648 13104
rect 8408 13082 8432 13084
rect 8488 13082 8512 13084
rect 8568 13082 8592 13084
rect 8430 13030 8432 13082
rect 8494 13030 8506 13082
rect 8568 13030 8570 13082
rect 8408 13028 8432 13030
rect 8488 13028 8512 13030
rect 8568 13028 8592 13030
rect 8352 13008 8648 13028
rect 7932 12912 7984 12918
rect 7932 12854 7984 12860
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7944 12186 7972 12854
rect 8024 12776 8076 12782
rect 8024 12718 8076 12724
rect 8036 12345 8064 12718
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 8312 12442 8340 12650
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8022 12336 8078 12345
rect 8022 12271 8078 12280
rect 8668 12300 8720 12306
rect 8864 12288 8892 14447
rect 8956 14346 8984 14826
rect 9048 14346 9076 15014
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 8944 14340 8996 14346
rect 8944 14282 8996 14288
rect 9036 14340 9088 14346
rect 9036 14282 9088 14288
rect 8956 13530 8984 14282
rect 9048 13870 9076 14282
rect 9140 13870 9168 14350
rect 9036 13864 9088 13870
rect 9036 13806 9088 13812
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 8944 13524 8996 13530
rect 8944 13466 8996 13472
rect 9048 13190 9076 13806
rect 9140 13394 9168 13806
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 9126 12744 9182 12753
rect 8668 12242 8720 12248
rect 8772 12260 8892 12288
rect 8208 12232 8260 12238
rect 7944 12158 8064 12186
rect 8208 12174 8260 12180
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7944 11218 7972 12038
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 8036 11150 8064 12158
rect 8220 11694 8248 12174
rect 8352 11996 8648 12016
rect 8408 11994 8432 11996
rect 8488 11994 8512 11996
rect 8568 11994 8592 11996
rect 8430 11942 8432 11994
rect 8494 11942 8506 11994
rect 8568 11942 8570 11994
rect 8408 11940 8432 11942
rect 8488 11940 8512 11942
rect 8568 11940 8592 11942
rect 8352 11920 8648 11940
rect 8680 11898 8708 12242
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8666 11792 8722 11801
rect 8666 11727 8722 11736
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8300 11620 8352 11626
rect 8300 11562 8352 11568
rect 8312 11354 8340 11562
rect 8680 11558 8708 11727
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 8036 10810 8064 11086
rect 8352 10908 8648 10928
rect 8408 10906 8432 10908
rect 8488 10906 8512 10908
rect 8568 10906 8592 10908
rect 8430 10854 8432 10906
rect 8494 10854 8506 10906
rect 8568 10854 8570 10906
rect 8408 10852 8432 10854
rect 8488 10852 8512 10854
rect 8568 10852 8592 10854
rect 8352 10832 8648 10852
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 7760 9586 7788 10542
rect 8036 10169 8064 10746
rect 8022 10160 8078 10169
rect 8772 10146 8800 12260
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8852 12164 8904 12170
rect 8852 12106 8904 12112
rect 8864 11286 8892 12106
rect 8956 11354 8984 12174
rect 9048 11898 9076 12718
rect 9126 12679 9182 12688
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 8864 10810 8892 11222
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 8956 10266 8984 11154
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 8022 10095 8078 10104
rect 8668 10124 8720 10130
rect 8772 10118 8984 10146
rect 8668 10066 8720 10072
rect 8352 9820 8648 9840
rect 8408 9818 8432 9820
rect 8488 9818 8512 9820
rect 8568 9818 8592 9820
rect 8430 9766 8432 9818
rect 8494 9766 8506 9818
rect 8568 9766 8570 9818
rect 8408 9764 8432 9766
rect 8488 9764 8512 9766
rect 8568 9764 8592 9766
rect 8352 9744 8648 9764
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7852 8974 7880 9658
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7562 8528 7618 8537
rect 7562 8463 7618 8472
rect 7852 8480 7880 8910
rect 7932 8492 7984 8498
rect 7576 7954 7604 8463
rect 7852 8452 7932 8480
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7564 7812 7616 7818
rect 7564 7754 7616 7760
rect 7576 5794 7604 7754
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7668 6730 7696 7142
rect 7656 6724 7708 6730
rect 7656 6666 7708 6672
rect 7286 5743 7342 5752
rect 7472 5772 7524 5778
rect 6918 5672 6974 5681
rect 6918 5607 6974 5616
rect 7012 5636 7064 5642
rect 6932 5234 6960 5607
rect 7012 5578 7064 5584
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6366 3632 6422 3641
rect 6276 3596 6328 3602
rect 6366 3567 6422 3576
rect 6276 3538 6328 3544
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5828 2854 5856 3130
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 5886 2748 6182 2768
rect 5942 2746 5966 2748
rect 6022 2746 6046 2748
rect 6102 2746 6126 2748
rect 5964 2694 5966 2746
rect 6028 2694 6040 2746
rect 6102 2694 6104 2746
rect 5942 2692 5966 2694
rect 6022 2692 6046 2694
rect 6102 2692 6126 2694
rect 5886 2672 6182 2692
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5264 2576 5316 2582
rect 5264 2518 5316 2524
rect 6288 1442 6316 3538
rect 6380 3534 6408 3567
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 6380 3058 6408 3334
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 6564 2938 6592 3946
rect 6642 3768 6698 3777
rect 6642 3703 6644 3712
rect 6696 3703 6698 3712
rect 6828 3732 6880 3738
rect 6644 3674 6696 3680
rect 6828 3674 6880 3680
rect 6656 2990 6684 3674
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6012 1414 6316 1442
rect 6380 2910 6592 2938
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 5538 912 5594 921
rect 5538 847 5594 856
rect 5552 800 5580 847
rect 6012 800 6040 1414
rect 6380 800 6408 2910
rect 6748 2836 6776 3334
rect 6656 2808 6776 2836
rect 6656 2446 6684 2808
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6840 800 6868 3674
rect 6932 2650 6960 4966
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 7024 921 7052 5578
rect 7196 5024 7248 5030
rect 7300 5012 7328 5743
rect 7576 5766 7696 5794
rect 7472 5714 7524 5720
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7576 5574 7604 5646
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7392 5166 7420 5510
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7248 4984 7328 5012
rect 7196 4966 7248 4972
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 7208 3670 7236 4422
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7196 3664 7248 3670
rect 7196 3606 7248 3612
rect 7208 3058 7236 3606
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7116 1154 7144 2586
rect 7392 1986 7420 3878
rect 7576 2582 7604 5510
rect 7668 5370 7696 5766
rect 7760 5658 7788 7890
rect 7852 5778 7880 8452
rect 7932 8434 7984 8440
rect 8036 7342 8064 9590
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8312 9110 8340 9318
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 8404 9042 8432 9454
rect 8680 9178 8708 10066
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8760 9988 8812 9994
rect 8760 9930 8812 9936
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8352 8732 8648 8752
rect 8408 8730 8432 8732
rect 8488 8730 8512 8732
rect 8568 8730 8592 8732
rect 8430 8678 8432 8730
rect 8494 8678 8506 8730
rect 8568 8678 8570 8730
rect 8408 8676 8432 8678
rect 8488 8676 8512 8678
rect 8568 8676 8592 8678
rect 8352 8656 8648 8676
rect 8772 8634 8800 9930
rect 8864 9518 8892 9998
rect 8956 9654 8984 10118
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8864 8566 8892 9454
rect 8956 9382 8984 9590
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8944 9104 8996 9110
rect 8944 9046 8996 9052
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8852 8560 8904 8566
rect 8852 8502 8904 8508
rect 8484 8016 8536 8022
rect 8484 7958 8536 7964
rect 8496 7857 8524 7958
rect 8482 7848 8538 7857
rect 8482 7783 8538 7792
rect 8352 7644 8648 7664
rect 8408 7642 8432 7644
rect 8488 7642 8512 7644
rect 8568 7642 8592 7644
rect 8430 7590 8432 7642
rect 8494 7590 8506 7642
rect 8568 7590 8570 7642
rect 8408 7588 8432 7590
rect 8488 7588 8512 7590
rect 8568 7588 8592 7590
rect 8352 7568 8648 7588
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8312 6934 8340 7278
rect 8680 6934 8708 8502
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 8668 6928 8720 6934
rect 8668 6870 8720 6876
rect 8772 6746 8800 8230
rect 8850 8120 8906 8129
rect 8850 8055 8906 8064
rect 8864 7954 8892 8055
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8680 6718 8800 6746
rect 8352 6556 8648 6576
rect 8408 6554 8432 6556
rect 8488 6554 8512 6556
rect 8568 6554 8592 6556
rect 8430 6502 8432 6554
rect 8494 6502 8506 6554
rect 8568 6502 8570 6554
rect 8408 6500 8432 6502
rect 8488 6500 8512 6502
rect 8568 6500 8592 6502
rect 8352 6480 8648 6500
rect 8392 6248 8444 6254
rect 8390 6216 8392 6225
rect 8444 6216 8446 6225
rect 8300 6180 8352 6186
rect 8390 6151 8446 6160
rect 8300 6122 8352 6128
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 8312 5710 8340 6122
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8496 5846 8524 6054
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 7932 5704 7984 5710
rect 7930 5672 7932 5681
rect 8300 5704 8352 5710
rect 7984 5672 7986 5681
rect 7760 5630 7880 5658
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7668 4758 7696 5306
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7760 4826 7788 4966
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7656 4752 7708 4758
rect 7656 4694 7708 4700
rect 7852 4690 7880 5630
rect 8300 5646 8352 5652
rect 7930 5607 7986 5616
rect 8352 5468 8648 5488
rect 8408 5466 8432 5468
rect 8488 5466 8512 5468
rect 8568 5466 8592 5468
rect 8430 5414 8432 5466
rect 8494 5414 8506 5466
rect 8568 5414 8570 5466
rect 8408 5412 8432 5414
rect 8488 5412 8512 5414
rect 8568 5412 8592 5414
rect 8352 5392 8648 5412
rect 8392 5092 8444 5098
rect 8680 5080 8708 6718
rect 8956 5794 8984 9046
rect 9048 9042 9076 11290
rect 9140 10062 9168 12679
rect 9232 12617 9260 16374
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9218 12608 9274 12617
rect 9218 12543 9274 12552
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 9232 11150 9260 11698
rect 9324 11354 9352 15506
rect 9402 15464 9458 15473
rect 9402 15399 9458 15408
rect 9416 11665 9444 15399
rect 9508 12782 9536 16662
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9862 16552 9918 16561
rect 9600 16153 9628 16526
rect 9862 16487 9918 16496
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9586 16144 9642 16153
rect 9586 16079 9642 16088
rect 9588 15972 9640 15978
rect 9588 15914 9640 15920
rect 9600 15434 9628 15914
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9600 13462 9628 14758
rect 9692 14074 9720 14962
rect 9784 14890 9812 16390
rect 9772 14884 9824 14890
rect 9772 14826 9824 14832
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9402 11656 9458 11665
rect 9402 11591 9458 11600
rect 9508 11558 9536 12718
rect 9876 12696 9904 16487
rect 9968 15473 9996 17054
rect 10244 15994 10272 17070
rect 10152 15978 10272 15994
rect 10140 15972 10272 15978
rect 10192 15966 10272 15972
rect 10140 15914 10192 15920
rect 10244 15706 10272 15966
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 10140 15564 10192 15570
rect 10140 15506 10192 15512
rect 9954 15464 10010 15473
rect 9954 15399 10010 15408
rect 10060 15162 10088 15506
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 10152 15026 10180 15506
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10244 15065 10272 15098
rect 10230 15056 10286 15065
rect 10140 15020 10192 15026
rect 10230 14991 10286 15000
rect 10140 14962 10192 14968
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9968 14074 9996 14418
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9876 12668 9996 12696
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9862 12608 9918 12617
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9692 11898 9720 12174
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9494 11112 9550 11121
rect 9232 10606 9260 11086
rect 9312 11076 9364 11082
rect 9600 11098 9628 11834
rect 9784 11762 9812 12582
rect 9862 12543 9918 12552
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9876 11626 9904 12543
rect 9968 11694 9996 12668
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9600 11070 9720 11098
rect 9494 11047 9550 11056
rect 9312 11018 9364 11024
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9232 10266 9260 10542
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9324 10062 9352 11018
rect 9402 10296 9458 10305
rect 9402 10231 9458 10240
rect 9508 10248 9536 11047
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9600 10742 9628 10950
rect 9588 10736 9640 10742
rect 9588 10678 9640 10684
rect 9416 10198 9444 10231
rect 9508 10220 9628 10248
rect 9404 10192 9456 10198
rect 9456 10152 9536 10180
rect 9404 10134 9456 10140
rect 9128 10056 9180 10062
rect 9312 10056 9364 10062
rect 9180 10016 9260 10044
rect 9128 9998 9180 10004
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 9140 9178 9168 9318
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 9036 8900 9088 8906
rect 9036 8842 9088 8848
rect 9048 8498 9076 8842
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 9048 8072 9076 8434
rect 9048 8044 9168 8072
rect 9140 7886 9168 8044
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 9048 6866 9076 7482
rect 9232 7206 9260 10016
rect 9312 9998 9364 10004
rect 9402 10024 9458 10033
rect 9402 9959 9458 9968
rect 9416 9450 9444 9959
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9324 7274 9352 7890
rect 9416 7274 9444 8230
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 9404 7268 9456 7274
rect 9404 7210 9456 7216
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9324 7002 9352 7210
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 9508 6730 9536 10152
rect 9600 8265 9628 10220
rect 9692 10198 9720 11070
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9876 10554 9904 11562
rect 10060 10674 10088 14758
rect 10152 11286 10180 14962
rect 10336 14822 10364 19200
rect 10600 16448 10652 16454
rect 10600 16390 10652 16396
rect 10416 15496 10468 15502
rect 10414 15464 10416 15473
rect 10468 15464 10470 15473
rect 10414 15399 10470 15408
rect 10612 15026 10640 16390
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10600 14544 10652 14550
rect 10600 14486 10652 14492
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10520 14006 10548 14214
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 10244 13530 10272 13806
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10140 11280 10192 11286
rect 10140 11222 10192 11228
rect 10244 11218 10272 13466
rect 10416 13388 10468 13394
rect 10468 13348 10548 13376
rect 10416 13330 10468 13336
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 10336 11354 10364 12718
rect 10428 12238 10456 12786
rect 10520 12345 10548 13348
rect 10612 12986 10640 14486
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10704 12866 10732 19200
rect 11072 17320 11100 19200
rect 11532 17762 11560 19200
rect 11440 17734 11560 17762
rect 11072 17292 11376 17320
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 10817 16892 11113 16912
rect 10873 16890 10897 16892
rect 10953 16890 10977 16892
rect 11033 16890 11057 16892
rect 10895 16838 10897 16890
rect 10959 16838 10971 16890
rect 11033 16838 11035 16890
rect 10873 16836 10897 16838
rect 10953 16836 10977 16838
rect 11033 16836 11057 16838
rect 10817 16816 11113 16836
rect 11164 16794 11192 16934
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11150 16688 11206 16697
rect 11150 16623 11206 16632
rect 10817 15804 11113 15824
rect 10873 15802 10897 15804
rect 10953 15802 10977 15804
rect 11033 15802 11057 15804
rect 10895 15750 10897 15802
rect 10959 15750 10971 15802
rect 11033 15750 11035 15802
rect 10873 15748 10897 15750
rect 10953 15748 10977 15750
rect 11033 15748 11057 15750
rect 10817 15728 11113 15748
rect 11164 15586 11192 16623
rect 11256 15978 11284 17138
rect 11348 16522 11376 17292
rect 11440 16833 11468 17734
rect 11520 17604 11572 17610
rect 11520 17546 11572 17552
rect 11426 16824 11482 16833
rect 11426 16759 11482 16768
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11336 16516 11388 16522
rect 11336 16458 11388 16464
rect 11440 16250 11468 16594
rect 11428 16244 11480 16250
rect 11428 16186 11480 16192
rect 11244 15972 11296 15978
rect 11244 15914 11296 15920
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 10980 15570 11192 15586
rect 10968 15564 11192 15570
rect 11020 15558 11192 15564
rect 10968 15506 11020 15512
rect 10817 14716 11113 14736
rect 10873 14714 10897 14716
rect 10953 14714 10977 14716
rect 11033 14714 11057 14716
rect 10895 14662 10897 14714
rect 10959 14662 10971 14714
rect 11033 14662 11035 14714
rect 10873 14660 10897 14662
rect 10953 14660 10977 14662
rect 11033 14660 11057 14662
rect 10817 14640 11113 14660
rect 10966 14376 11022 14385
rect 10966 14311 11022 14320
rect 10980 14278 11008 14311
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10817 13628 11113 13648
rect 10873 13626 10897 13628
rect 10953 13626 10977 13628
rect 11033 13626 11057 13628
rect 10895 13574 10897 13626
rect 10959 13574 10971 13626
rect 11033 13574 11035 13626
rect 10873 13572 10897 13574
rect 10953 13572 10977 13574
rect 11033 13572 11057 13574
rect 10817 13552 11113 13572
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10612 12838 10732 12866
rect 10888 12850 10916 13330
rect 10876 12844 10928 12850
rect 10612 12458 10640 12838
rect 10876 12786 10928 12792
rect 11150 12744 11206 12753
rect 11150 12679 11206 12688
rect 10817 12540 11113 12560
rect 10873 12538 10897 12540
rect 10953 12538 10977 12540
rect 11033 12538 11057 12540
rect 10895 12486 10897 12538
rect 10959 12486 10971 12538
rect 11033 12486 11035 12538
rect 10873 12484 10897 12486
rect 10953 12484 10977 12486
rect 11033 12484 11057 12486
rect 10817 12464 11113 12484
rect 10603 12430 10640 12458
rect 10603 12356 10631 12430
rect 10968 12368 11020 12374
rect 10506 12336 10562 12345
rect 10603 12328 10640 12356
rect 10506 12271 10562 12280
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10428 12102 10456 12174
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10416 11688 10468 11694
rect 10416 11630 10468 11636
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 9784 10062 9812 10542
rect 9876 10526 10088 10554
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9784 9466 9812 9862
rect 9876 9761 9904 10066
rect 9862 9752 9918 9761
rect 9862 9687 9918 9696
rect 9586 8256 9642 8265
rect 9586 8191 9642 8200
rect 9692 8090 9720 9454
rect 9784 9438 9996 9466
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9876 9178 9904 9318
rect 9864 9172 9916 9178
rect 9864 9114 9916 9120
rect 9862 9072 9918 9081
rect 9862 9007 9918 9016
rect 9876 8974 9904 9007
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9586 7848 9642 7857
rect 9586 7783 9642 7792
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 8864 5778 8984 5794
rect 8852 5772 8984 5778
rect 8904 5766 8984 5772
rect 8852 5714 8904 5720
rect 9232 5710 9260 6258
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9508 5914 9536 6054
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 8444 5052 8708 5080
rect 8392 5034 8444 5040
rect 8024 4752 8076 4758
rect 8024 4694 8076 4700
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 7852 4282 7880 4626
rect 8036 4282 8064 4694
rect 8116 4548 8168 4554
rect 8116 4490 8168 4496
rect 7840 4276 7892 4282
rect 7840 4218 7892 4224
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 7840 4072 7892 4078
rect 7892 4020 7972 4026
rect 7840 4014 7972 4020
rect 7852 3998 7972 4014
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7564 2576 7616 2582
rect 7564 2518 7616 2524
rect 7564 2304 7616 2310
rect 7564 2246 7616 2252
rect 7576 2038 7604 2246
rect 7208 1958 7420 1986
rect 7564 2032 7616 2038
rect 7564 1974 7616 1980
rect 7104 1148 7156 1154
rect 7104 1090 7156 1096
rect 7010 912 7066 921
rect 7010 847 7066 856
rect 7208 800 7236 1958
rect 7668 800 7696 3674
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7852 3194 7880 3470
rect 7944 3466 7972 3998
rect 7932 3460 7984 3466
rect 7932 3402 7984 3408
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7944 3058 7972 3402
rect 8036 3346 8064 4218
rect 8128 3602 8156 4490
rect 8352 4380 8648 4400
rect 8408 4378 8432 4380
rect 8488 4378 8512 4380
rect 8568 4378 8592 4380
rect 8430 4326 8432 4378
rect 8494 4326 8506 4378
rect 8568 4326 8570 4378
rect 8408 4324 8432 4326
rect 8488 4324 8512 4326
rect 8568 4324 8592 4326
rect 8352 4304 8648 4324
rect 8680 4078 8708 5052
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8772 4622 8800 5034
rect 8944 5024 8996 5030
rect 8864 4984 8944 5012
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 8036 3318 8156 3346
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7932 2916 7984 2922
rect 7932 2858 7984 2864
rect 8024 2916 8076 2922
rect 8024 2858 8076 2864
rect 7944 2825 7972 2858
rect 7930 2816 7986 2825
rect 7930 2751 7986 2760
rect 8036 800 8064 2858
rect 8128 1986 8156 3318
rect 8220 3194 8248 3946
rect 8864 3738 8892 4984
rect 8944 4966 8996 4972
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 8956 4282 8984 4558
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 9048 3738 9076 4422
rect 9140 3942 9168 5510
rect 9232 5370 9260 5646
rect 9416 5642 9444 5850
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9416 4690 9444 5578
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 9404 4684 9456 4690
rect 9404 4626 9456 4632
rect 9508 4486 9536 5102
rect 9496 4480 9548 4486
rect 9496 4422 9548 4428
rect 9508 4282 9536 4422
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8352 3292 8648 3312
rect 8408 3290 8432 3292
rect 8488 3290 8512 3292
rect 8568 3290 8592 3292
rect 8430 3238 8432 3290
rect 8494 3238 8506 3290
rect 8568 3238 8570 3290
rect 8408 3236 8432 3238
rect 8488 3236 8512 3238
rect 8568 3236 8592 3238
rect 8352 3216 8648 3236
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8220 2446 8248 3130
rect 8680 2514 8708 3334
rect 8850 2816 8906 2825
rect 8850 2751 8906 2760
rect 8668 2508 8720 2514
rect 8668 2450 8720 2456
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 8352 2204 8648 2224
rect 8408 2202 8432 2204
rect 8488 2202 8512 2204
rect 8568 2202 8592 2204
rect 8430 2150 8432 2202
rect 8494 2150 8506 2202
rect 8568 2150 8570 2202
rect 8408 2148 8432 2150
rect 8488 2148 8512 2150
rect 8568 2148 8592 2150
rect 8352 2128 8648 2148
rect 8128 1958 8524 1986
rect 8496 800 8524 1958
rect 8864 800 8892 2751
rect 9232 1034 9260 4014
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9416 3194 9444 3470
rect 9508 3398 9536 4218
rect 9600 3534 9628 7783
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 6118 9720 7142
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9692 3466 9720 6054
rect 9876 5166 9904 8910
rect 9968 8022 9996 9438
rect 10060 9382 10088 10526
rect 10152 9654 10180 11086
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 9956 7812 10008 7818
rect 9956 7754 10008 7760
rect 9968 5778 9996 7754
rect 10060 6934 10088 9318
rect 10140 7812 10192 7818
rect 10244 7800 10272 10610
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10336 8090 10364 9522
rect 10428 9518 10456 11630
rect 10520 11014 10548 12271
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10520 10606 10548 10950
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10508 10192 10560 10198
rect 10508 10134 10560 10140
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10192 7772 10272 7800
rect 10140 7754 10192 7760
rect 10232 7472 10284 7478
rect 10138 7440 10194 7449
rect 10232 7414 10284 7420
rect 10138 7375 10194 7384
rect 10152 7342 10180 7375
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 10048 6928 10100 6934
rect 10048 6870 10100 6876
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9968 4826 9996 5510
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9784 4282 9812 4694
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 10060 3942 10088 6870
rect 10152 6458 10180 7278
rect 10244 6798 10272 7414
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10336 7002 10364 7278
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10324 6860 10376 6866
rect 10428 6848 10456 9454
rect 10520 9081 10548 10134
rect 10506 9072 10562 9081
rect 10506 9007 10562 9016
rect 10612 8514 10640 12328
rect 10874 12336 10930 12345
rect 10692 12300 10744 12306
rect 10968 12310 11020 12316
rect 10874 12271 10930 12280
rect 10692 12242 10744 12248
rect 10704 11898 10732 12242
rect 10888 12238 10916 12271
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10980 11762 11008 12310
rect 11164 11762 11192 12679
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 10704 11218 10732 11698
rect 11058 11656 11114 11665
rect 11058 11591 11060 11600
rect 11112 11591 11114 11600
rect 11060 11562 11112 11568
rect 11256 11506 11284 15642
rect 11532 15570 11560 17546
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11624 15910 11652 17138
rect 11796 16720 11848 16726
rect 11796 16662 11848 16668
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11716 16114 11744 16526
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 11532 15450 11560 15506
rect 11440 15422 11560 15450
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 11348 12442 11376 12582
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11164 11478 11284 11506
rect 10817 11452 11113 11472
rect 10873 11450 10897 11452
rect 10953 11450 10977 11452
rect 11033 11450 11057 11452
rect 10895 11398 10897 11450
rect 10959 11398 10971 11450
rect 11033 11398 11035 11450
rect 10873 11396 10897 11398
rect 10953 11396 10977 11398
rect 11033 11396 11057 11398
rect 10817 11376 11113 11396
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10876 11144 10928 11150
rect 10874 11112 10876 11121
rect 10928 11112 10930 11121
rect 10874 11047 10930 11056
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10704 9761 10732 10746
rect 10817 10364 11113 10384
rect 10873 10362 10897 10364
rect 10953 10362 10977 10364
rect 11033 10362 11057 10364
rect 10895 10310 10897 10362
rect 10959 10310 10971 10362
rect 11033 10310 11035 10362
rect 10873 10308 10897 10310
rect 10953 10308 10977 10310
rect 11033 10308 11057 10310
rect 10817 10288 11113 10308
rect 10690 9752 10746 9761
rect 10690 9687 10746 9696
rect 10704 9586 10732 9687
rect 11164 9625 11192 11478
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11256 10606 11284 11290
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11242 10160 11298 10169
rect 11242 10095 11298 10104
rect 11150 9616 11206 9625
rect 10692 9580 10744 9586
rect 11150 9551 11206 9560
rect 10692 9522 10744 9528
rect 10817 9276 11113 9296
rect 10873 9274 10897 9276
rect 10953 9274 10977 9276
rect 11033 9274 11057 9276
rect 10895 9222 10897 9274
rect 10959 9222 10971 9274
rect 11033 9222 11035 9274
rect 10873 9220 10897 9222
rect 10953 9220 10977 9222
rect 11033 9220 11057 9222
rect 10817 9200 11113 9220
rect 10784 9036 10836 9042
rect 10836 8996 10916 9024
rect 10784 8978 10836 8984
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10704 8634 10732 8910
rect 10888 8634 10916 8996
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10376 6820 10456 6848
rect 10520 8486 10640 8514
rect 10324 6802 10376 6808
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10138 6352 10194 6361
rect 10138 6287 10194 6296
rect 10152 5250 10180 6287
rect 10244 6254 10272 6734
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10244 5710 10272 6054
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10152 5222 10272 5250
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 10152 4554 10180 5102
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9784 3777 9812 3878
rect 9770 3768 9826 3777
rect 9770 3703 9826 3712
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9404 3188 9456 3194
rect 9324 3148 9404 3176
rect 9324 2990 9352 3148
rect 9404 3130 9456 3136
rect 9508 3058 9536 3334
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9324 2446 9352 2926
rect 9494 2680 9550 2689
rect 9494 2615 9550 2624
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9508 2310 9536 2615
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 9232 1006 9352 1034
rect 9324 800 9352 1006
rect 9692 800 9720 3402
rect 9784 2650 9812 3538
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 9968 2650 9996 3334
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 10060 2582 10088 3334
rect 10244 3233 10272 5222
rect 10336 3942 10364 6802
rect 10414 5672 10470 5681
rect 10414 5607 10470 5616
rect 10428 3942 10456 5607
rect 10520 5098 10548 8486
rect 10704 8430 10732 8570
rect 11256 8566 11284 10095
rect 11348 9654 11376 10406
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11244 8560 11296 8566
rect 11244 8502 11296 8508
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10612 7324 10640 8366
rect 10704 7449 10732 8366
rect 11060 8356 11112 8362
rect 11112 8316 11192 8344
rect 11060 8298 11112 8304
rect 10817 8188 11113 8208
rect 10873 8186 10897 8188
rect 10953 8186 10977 8188
rect 11033 8186 11057 8188
rect 10895 8134 10897 8186
rect 10959 8134 10971 8186
rect 11033 8134 11035 8186
rect 10873 8132 10897 8134
rect 10953 8132 10977 8134
rect 11033 8132 11057 8134
rect 10817 8112 11113 8132
rect 10784 8016 10836 8022
rect 10784 7958 10836 7964
rect 10796 7546 10824 7958
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 11072 7546 11100 7890
rect 11164 7886 11192 8316
rect 11348 8294 11376 8978
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11348 7886 11376 8230
rect 11440 7954 11468 15422
rect 11520 15360 11572 15366
rect 11520 15302 11572 15308
rect 11532 14958 11560 15302
rect 11624 15026 11652 15846
rect 11716 15502 11744 16050
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11520 14952 11572 14958
rect 11520 14894 11572 14900
rect 11624 14482 11652 14962
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11624 13530 11652 13874
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11624 12850 11652 13466
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11808 12646 11836 16662
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11900 12458 11928 19200
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 11992 16046 12020 16526
rect 11980 16040 12032 16046
rect 11980 15982 12032 15988
rect 11992 15502 12020 15982
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12176 14006 12204 15438
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12268 15162 12296 15302
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12164 14000 12216 14006
rect 12164 13942 12216 13948
rect 11980 13728 12032 13734
rect 11980 13670 12032 13676
rect 11992 13530 12020 13670
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12268 12850 12296 13330
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 11900 12430 12011 12458
rect 11983 12424 12011 12430
rect 11983 12396 12020 12424
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11532 10033 11560 11698
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11716 10674 11744 11154
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11888 10532 11940 10538
rect 11888 10474 11940 10480
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11518 10024 11574 10033
rect 11518 9959 11574 9968
rect 11624 9926 11652 10202
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11716 9518 11744 9862
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 11152 7880 11204 7886
rect 11336 7880 11388 7886
rect 11204 7840 11284 7868
rect 11152 7822 11204 7828
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 10690 7440 10746 7449
rect 10690 7375 10746 7384
rect 10612 7296 10732 7324
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10612 6730 10640 7142
rect 10600 6724 10652 6730
rect 10600 6666 10652 6672
rect 10612 5817 10640 6666
rect 10704 6662 10732 7296
rect 10817 7100 11113 7120
rect 10873 7098 10897 7100
rect 10953 7098 10977 7100
rect 11033 7098 11057 7100
rect 10895 7046 10897 7098
rect 10959 7046 10971 7098
rect 11033 7046 11035 7098
rect 10873 7044 10897 7046
rect 10953 7044 10977 7046
rect 11033 7044 11057 7046
rect 10817 7024 11113 7044
rect 11256 7002 11284 7840
rect 11532 7834 11560 8978
rect 11624 8498 11652 9046
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11624 7993 11652 8230
rect 11610 7984 11666 7993
rect 11610 7919 11666 7928
rect 11336 7822 11388 7828
rect 11440 7806 11560 7834
rect 11716 7818 11744 8774
rect 11704 7812 11756 7818
rect 11334 7440 11390 7449
rect 11334 7375 11390 7384
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10598 5808 10654 5817
rect 10598 5743 10654 5752
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10612 5370 10640 5646
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10508 5092 10560 5098
rect 10508 5034 10560 5040
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10230 3224 10286 3233
rect 10230 3159 10286 3168
rect 10244 3074 10272 3159
rect 10152 3046 10272 3074
rect 10048 2576 10100 2582
rect 10048 2518 10100 2524
rect 10152 800 10180 3046
rect 10336 2825 10364 3878
rect 10520 3738 10548 5034
rect 10612 4758 10640 5306
rect 10600 4752 10652 4758
rect 10600 4694 10652 4700
rect 10612 4146 10640 4694
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10508 3732 10560 3738
rect 10508 3674 10560 3680
rect 10612 3534 10640 4082
rect 10704 4078 10732 6598
rect 11256 6322 11284 6938
rect 11348 6866 11376 7375
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11440 6186 11468 7806
rect 11704 7754 11756 7760
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11428 6180 11480 6186
rect 11428 6122 11480 6128
rect 10817 6012 11113 6032
rect 10873 6010 10897 6012
rect 10953 6010 10977 6012
rect 11033 6010 11057 6012
rect 10895 5958 10897 6010
rect 10959 5958 10971 6010
rect 11033 5958 11035 6010
rect 10873 5956 10897 5958
rect 10953 5956 10977 5958
rect 11033 5956 11057 5958
rect 10817 5936 11113 5956
rect 10782 5808 10838 5817
rect 10782 5743 10784 5752
rect 10836 5743 10838 5752
rect 10784 5714 10836 5720
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 10817 4924 11113 4944
rect 10873 4922 10897 4924
rect 10953 4922 10977 4924
rect 11033 4922 11057 4924
rect 10895 4870 10897 4922
rect 10959 4870 10971 4922
rect 11033 4870 11035 4922
rect 10873 4868 10897 4870
rect 10953 4868 10977 4870
rect 11033 4868 11057 4870
rect 10817 4848 11113 4868
rect 10692 4072 10744 4078
rect 10784 4072 10836 4078
rect 10692 4014 10744 4020
rect 10782 4040 10784 4049
rect 11152 4072 11204 4078
rect 10836 4040 10838 4049
rect 11152 4014 11204 4020
rect 10782 3975 10838 3984
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10508 3460 10560 3466
rect 10508 3402 10560 3408
rect 10416 2916 10468 2922
rect 10416 2858 10468 2864
rect 10322 2816 10378 2825
rect 10322 2751 10378 2760
rect 10428 2446 10456 2858
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 10520 800 10548 3402
rect 10600 2916 10652 2922
rect 10600 2858 10652 2864
rect 10612 2514 10640 2858
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 10704 1034 10732 3878
rect 10817 3836 11113 3856
rect 10873 3834 10897 3836
rect 10953 3834 10977 3836
rect 11033 3834 11057 3836
rect 10895 3782 10897 3834
rect 10959 3782 10971 3834
rect 11033 3782 11035 3834
rect 10873 3780 10897 3782
rect 10953 3780 10977 3782
rect 11033 3780 11057 3782
rect 10817 3760 11113 3780
rect 11164 3670 11192 4014
rect 11348 3942 11376 5646
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11440 3738 11468 3878
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11348 3194 11376 3470
rect 11426 3224 11482 3233
rect 11336 3188 11388 3194
rect 11426 3159 11482 3168
rect 11336 3130 11388 3136
rect 11440 2854 11468 3159
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 11428 2848 11480 2854
rect 11428 2790 11480 2796
rect 10817 2748 11113 2768
rect 10873 2746 10897 2748
rect 10953 2746 10977 2748
rect 11033 2746 11057 2748
rect 10895 2694 10897 2746
rect 10959 2694 10971 2746
rect 11033 2694 11035 2746
rect 10873 2692 10897 2694
rect 10953 2692 10977 2694
rect 11033 2692 11057 2694
rect 10817 2672 11113 2692
rect 11164 2650 11192 2790
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11060 2576 11112 2582
rect 11532 2530 11560 7278
rect 11624 6934 11652 7346
rect 11704 7268 11756 7274
rect 11704 7210 11756 7216
rect 11716 6934 11744 7210
rect 11612 6928 11664 6934
rect 11612 6870 11664 6876
rect 11704 6928 11756 6934
rect 11704 6870 11756 6876
rect 11624 6390 11652 6870
rect 11612 6384 11664 6390
rect 11612 6326 11664 6332
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 11624 3641 11652 4490
rect 11808 3738 11836 9522
rect 11900 9518 11928 10474
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11992 9364 12020 12396
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12072 9376 12124 9382
rect 11992 9336 12072 9364
rect 11992 9042 12020 9336
rect 12072 9318 12124 9324
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 12176 8838 12204 10066
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12268 8650 12296 12582
rect 12360 12306 12388 19200
rect 12728 17490 12756 19200
rect 12728 17462 12848 17490
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12452 16250 12480 17070
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12452 12986 12480 13806
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12452 12186 12480 12718
rect 12544 12442 12572 13398
rect 12636 12458 12664 16730
rect 12728 12986 12756 17274
rect 12820 15706 12848 17462
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12820 12918 12848 15642
rect 13004 15162 13032 16934
rect 13096 16794 13124 19200
rect 13556 17524 13584 19200
rect 13556 17496 13676 17524
rect 13282 17436 13578 17456
rect 13338 17434 13362 17436
rect 13418 17434 13442 17436
rect 13498 17434 13522 17436
rect 13360 17382 13362 17434
rect 13424 17382 13436 17434
rect 13498 17382 13500 17434
rect 13338 17380 13362 17382
rect 13418 17380 13442 17382
rect 13498 17380 13522 17382
rect 13282 17360 13578 17380
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13188 16794 13216 17138
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 13176 16788 13228 16794
rect 13176 16730 13228 16736
rect 13188 15706 13216 16730
rect 13282 16348 13578 16368
rect 13338 16346 13362 16348
rect 13418 16346 13442 16348
rect 13498 16346 13522 16348
rect 13360 16294 13362 16346
rect 13424 16294 13436 16346
rect 13498 16294 13500 16346
rect 13338 16292 13362 16294
rect 13418 16292 13442 16294
rect 13498 16292 13522 16294
rect 13282 16272 13578 16292
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 13556 15706 13584 15914
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 13004 14550 13032 14962
rect 12992 14544 13044 14550
rect 12992 14486 13044 14492
rect 12992 14272 13044 14278
rect 12992 14214 13044 14220
rect 13004 13802 13032 14214
rect 12992 13796 13044 13802
rect 12992 13738 13044 13744
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 12808 12912 12860 12918
rect 12808 12854 12860 12860
rect 12532 12436 12584 12442
rect 12636 12430 12756 12458
rect 12532 12378 12584 12384
rect 12360 12158 12480 12186
rect 12360 9178 12388 12158
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12544 10470 12572 11154
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12544 9586 12572 10406
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12636 9722 12664 9862
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 11992 8622 12296 8650
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11900 7342 11928 7890
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11900 4010 11928 4082
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 11900 3738 11928 3946
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11610 3632 11666 3641
rect 11610 3567 11666 3576
rect 11112 2524 11560 2530
rect 11060 2518 11560 2524
rect 11072 2502 11560 2518
rect 11336 2304 11388 2310
rect 11336 2246 11388 2252
rect 10704 1006 11008 1034
rect 10980 800 11008 1006
rect 11348 800 11376 2246
rect 11532 2106 11560 2502
rect 11624 2446 11652 3567
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11520 2100 11572 2106
rect 11520 2042 11572 2048
rect 11716 2038 11744 2994
rect 11704 2032 11756 2038
rect 11704 1974 11756 1980
rect 11808 800 11836 3130
rect 11992 2446 12020 8622
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 12084 6458 12112 7890
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 12084 2514 12112 4694
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 12176 800 12204 8502
rect 12452 8344 12480 8978
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12360 8316 12480 8344
rect 12532 8356 12584 8362
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12268 3194 12296 8230
rect 12360 4010 12388 8316
rect 12532 8298 12584 8304
rect 12544 7954 12572 8298
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12636 7206 12664 8570
rect 12728 7342 12756 12430
rect 13004 10062 13032 13330
rect 13096 13258 13124 15574
rect 13084 13252 13136 13258
rect 13084 13194 13136 13200
rect 13188 13138 13216 15642
rect 13282 15260 13578 15280
rect 13338 15258 13362 15260
rect 13418 15258 13442 15260
rect 13498 15258 13522 15260
rect 13360 15206 13362 15258
rect 13424 15206 13436 15258
rect 13498 15206 13500 15258
rect 13338 15204 13362 15206
rect 13418 15204 13442 15206
rect 13498 15204 13522 15206
rect 13282 15184 13578 15204
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13280 14521 13308 14758
rect 13266 14512 13322 14521
rect 13266 14447 13322 14456
rect 13282 14172 13578 14192
rect 13338 14170 13362 14172
rect 13418 14170 13442 14172
rect 13498 14170 13522 14172
rect 13360 14118 13362 14170
rect 13424 14118 13436 14170
rect 13498 14118 13500 14170
rect 13338 14116 13362 14118
rect 13418 14116 13442 14118
rect 13498 14116 13522 14118
rect 13282 14096 13578 14116
rect 13544 13796 13596 13802
rect 13544 13738 13596 13744
rect 13556 13326 13584 13738
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13096 13110 13216 13138
rect 13096 12306 13124 13110
rect 13282 13084 13578 13104
rect 13338 13082 13362 13084
rect 13418 13082 13442 13084
rect 13498 13082 13522 13084
rect 13360 13030 13362 13082
rect 13424 13030 13436 13082
rect 13498 13030 13500 13082
rect 13338 13028 13362 13030
rect 13418 13028 13442 13030
rect 13498 13028 13522 13030
rect 13282 13008 13578 13028
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13188 12442 13216 12922
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 13280 12322 13308 12786
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 13188 12294 13308 12322
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 12820 9042 12848 9998
rect 13096 9926 13124 11562
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 12903 9704 12931 9862
rect 12903 9676 13032 9704
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12820 8537 12848 8978
rect 12806 8528 12862 8537
rect 12806 8463 12862 8472
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12624 7200 12676 7206
rect 12820 7188 12848 8463
rect 12912 8294 12940 9318
rect 13004 9110 13032 9676
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 13096 8974 13124 9522
rect 13084 8968 13136 8974
rect 12990 8936 13046 8945
rect 13084 8910 13136 8916
rect 12990 8871 13046 8880
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 13004 8106 13032 8871
rect 13096 8362 13124 8910
rect 13084 8356 13136 8362
rect 13084 8298 13136 8304
rect 12912 8078 13032 8106
rect 12912 7954 12940 8078
rect 12992 8016 13044 8022
rect 12992 7958 13044 7964
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12624 7142 12676 7148
rect 12728 7160 12848 7188
rect 12452 6458 12480 7142
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12544 6322 12572 6802
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12544 4622 12572 5102
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12636 4826 12664 5034
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12348 4004 12400 4010
rect 12348 3946 12400 3952
rect 12348 3664 12400 3670
rect 12348 3606 12400 3612
rect 12440 3664 12492 3670
rect 12440 3606 12492 3612
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12360 2938 12388 3606
rect 12452 3058 12480 3606
rect 12544 3126 12572 4558
rect 12636 4214 12664 4762
rect 12624 4208 12676 4214
rect 12624 4150 12676 4156
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12532 2984 12584 2990
rect 12360 2910 12480 2938
rect 12532 2926 12584 2932
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 12268 2038 12296 2382
rect 12256 2032 12308 2038
rect 12256 1974 12308 1980
rect 12452 1442 12480 2910
rect 12544 2310 12572 2926
rect 12636 2650 12664 3878
rect 12728 3602 12756 7160
rect 12912 7018 12940 7890
rect 12820 6990 12940 7018
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 12820 2514 12848 6990
rect 13004 6934 13032 7958
rect 13188 7750 13216 12294
rect 13282 11996 13578 12016
rect 13338 11994 13362 11996
rect 13418 11994 13442 11996
rect 13498 11994 13522 11996
rect 13360 11942 13362 11994
rect 13424 11942 13436 11994
rect 13498 11942 13500 11994
rect 13338 11940 13362 11942
rect 13418 11940 13442 11942
rect 13498 11940 13522 11942
rect 13282 11920 13578 11940
rect 13282 10908 13578 10928
rect 13338 10906 13362 10908
rect 13418 10906 13442 10908
rect 13498 10906 13522 10908
rect 13360 10854 13362 10906
rect 13424 10854 13436 10906
rect 13498 10854 13500 10906
rect 13338 10852 13362 10854
rect 13418 10852 13442 10854
rect 13498 10852 13522 10854
rect 13282 10832 13578 10852
rect 13648 10266 13676 17496
rect 13728 17264 13780 17270
rect 13728 17206 13780 17212
rect 13740 14958 13768 17206
rect 13924 17082 13952 19200
rect 14096 18012 14148 18018
rect 14096 17954 14148 17960
rect 14108 17202 14136 17954
rect 14188 17536 14240 17542
rect 14188 17478 14240 17484
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 13832 17054 13952 17082
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13740 13977 13768 14350
rect 13726 13968 13782 13977
rect 13726 13903 13782 13912
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13282 9820 13578 9840
rect 13338 9818 13362 9820
rect 13418 9818 13442 9820
rect 13498 9818 13522 9820
rect 13360 9766 13362 9818
rect 13424 9766 13436 9818
rect 13498 9766 13500 9818
rect 13338 9764 13362 9766
rect 13418 9764 13442 9766
rect 13498 9764 13522 9766
rect 13282 9744 13578 9764
rect 13268 9444 13320 9450
rect 13268 9386 13320 9392
rect 13280 8906 13308 9386
rect 13636 9104 13688 9110
rect 13636 9046 13688 9052
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13282 8732 13578 8752
rect 13338 8730 13362 8732
rect 13418 8730 13442 8732
rect 13498 8730 13522 8732
rect 13360 8678 13362 8730
rect 13424 8678 13436 8730
rect 13498 8678 13500 8730
rect 13338 8676 13362 8678
rect 13418 8676 13442 8678
rect 13498 8676 13522 8678
rect 13282 8656 13578 8676
rect 13268 8356 13320 8362
rect 13268 8298 13320 8304
rect 13280 7886 13308 8298
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 13282 7644 13578 7664
rect 13338 7642 13362 7644
rect 13418 7642 13442 7644
rect 13498 7642 13522 7644
rect 13360 7590 13362 7642
rect 13424 7590 13436 7642
rect 13498 7590 13500 7642
rect 13338 7588 13362 7590
rect 13418 7588 13442 7590
rect 13498 7588 13522 7590
rect 13282 7568 13578 7588
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13084 7268 13136 7274
rect 13084 7210 13136 7216
rect 12992 6928 13044 6934
rect 12992 6870 13044 6876
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 12912 6186 12940 6598
rect 12900 6180 12952 6186
rect 12900 6122 12952 6128
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12912 3466 12940 3878
rect 12900 3460 12952 3466
rect 12900 3402 12952 3408
rect 13004 2650 13032 6870
rect 13096 3754 13124 7210
rect 13464 6798 13492 7346
rect 13648 6866 13676 9046
rect 13740 8945 13768 13330
rect 13832 12782 13860 17054
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13924 15706 13952 16934
rect 14200 16658 14228 17478
rect 14004 16652 14056 16658
rect 14004 16594 14056 16600
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 14016 15502 14044 16594
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 14004 15496 14056 15502
rect 14004 15438 14056 15444
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 14016 14074 14044 14486
rect 14108 14278 14136 14962
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 14292 13530 14320 15506
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14004 13252 14056 13258
rect 14004 13194 14056 13200
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13924 12374 13952 12582
rect 13912 12368 13964 12374
rect 13912 12310 13964 12316
rect 14016 11626 14044 13194
rect 14384 12458 14412 19200
rect 14752 18170 14780 19200
rect 14660 18142 14780 18170
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14568 15162 14596 15438
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14568 14006 14596 15098
rect 14660 14618 14688 18142
rect 15120 18000 15148 19200
rect 14752 17972 15148 18000
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14556 14000 14608 14006
rect 14556 13942 14608 13948
rect 14568 12850 14596 13942
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14660 13190 14688 13738
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14556 12844 14608 12850
rect 14292 12430 14412 12458
rect 14476 12804 14556 12832
rect 14292 12424 14320 12430
rect 14200 12396 14320 12424
rect 14004 11620 14056 11626
rect 14004 11562 14056 11568
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13726 8936 13782 8945
rect 13726 8871 13782 8880
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13282 6556 13578 6576
rect 13338 6554 13362 6556
rect 13418 6554 13442 6556
rect 13498 6554 13522 6556
rect 13360 6502 13362 6554
rect 13424 6502 13436 6554
rect 13498 6502 13500 6554
rect 13338 6500 13362 6502
rect 13418 6500 13442 6502
rect 13498 6500 13522 6502
rect 13282 6480 13578 6500
rect 13176 5772 13228 5778
rect 13176 5714 13228 5720
rect 13188 3942 13216 5714
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 13282 5468 13578 5488
rect 13338 5466 13362 5468
rect 13418 5466 13442 5468
rect 13498 5466 13522 5468
rect 13360 5414 13362 5466
rect 13424 5414 13436 5466
rect 13498 5414 13500 5466
rect 13338 5412 13362 5414
rect 13418 5412 13442 5414
rect 13498 5412 13522 5414
rect 13282 5392 13578 5412
rect 13648 5370 13676 5646
rect 13740 5386 13768 8774
rect 13832 8090 13860 8978
rect 13924 8514 13952 11494
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14016 10062 14044 10610
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 14016 8974 14044 9998
rect 14108 9625 14136 10066
rect 14094 9616 14150 9625
rect 14094 9551 14150 9560
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 14016 8634 14044 8910
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 13924 8486 14044 8514
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 13924 5846 13952 6258
rect 13912 5840 13964 5846
rect 13912 5782 13964 5788
rect 13636 5364 13688 5370
rect 13740 5358 13860 5386
rect 13636 5306 13688 5312
rect 13728 4684 13780 4690
rect 13728 4626 13780 4632
rect 13282 4380 13578 4400
rect 13338 4378 13362 4380
rect 13418 4378 13442 4380
rect 13498 4378 13522 4380
rect 13360 4326 13362 4378
rect 13424 4326 13436 4378
rect 13498 4326 13500 4378
rect 13338 4324 13362 4326
rect 13418 4324 13442 4326
rect 13498 4324 13522 4326
rect 13282 4304 13578 4324
rect 13740 4146 13768 4626
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 13096 3726 13676 3754
rect 13266 3632 13322 3641
rect 13266 3567 13322 3576
rect 13280 3534 13308 3567
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13188 2922 13216 3470
rect 13282 3292 13578 3312
rect 13338 3290 13362 3292
rect 13418 3290 13442 3292
rect 13498 3290 13522 3292
rect 13360 3238 13362 3290
rect 13424 3238 13436 3290
rect 13498 3238 13500 3290
rect 13338 3236 13362 3238
rect 13418 3236 13442 3238
rect 13498 3236 13522 3238
rect 13282 3216 13578 3236
rect 13176 2916 13228 2922
rect 13176 2858 13228 2864
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 13188 2446 13216 2858
rect 13648 2514 13676 3726
rect 13740 3602 13768 4082
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13832 2802 13860 5358
rect 13924 3738 13952 5782
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13910 3088 13966 3097
rect 13910 3023 13966 3032
rect 13740 2774 13860 2802
rect 13636 2508 13688 2514
rect 13636 2450 13688 2456
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 12532 2304 12584 2310
rect 12532 2246 12584 2252
rect 13282 2204 13578 2224
rect 13338 2202 13362 2204
rect 13418 2202 13442 2204
rect 13498 2202 13522 2204
rect 13360 2150 13362 2202
rect 13424 2150 13436 2202
rect 13498 2150 13500 2202
rect 13338 2148 13362 2150
rect 13418 2148 13442 2150
rect 13498 2148 13522 2150
rect 13282 2128 13578 2148
rect 12992 2100 13044 2106
rect 12992 2042 13044 2048
rect 12452 1414 12664 1442
rect 12636 800 12664 1414
rect 13004 800 13032 2042
rect 13740 1306 13768 2774
rect 13924 2650 13952 3023
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 13464 1278 13768 1306
rect 13464 800 13492 1278
rect 14016 898 14044 8486
rect 14108 5302 14136 9551
rect 14200 5574 14228 12396
rect 14476 12306 14504 12804
rect 14556 12786 14608 12792
rect 14556 12708 14608 12714
rect 14556 12650 14608 12656
rect 14464 12300 14516 12306
rect 14464 12242 14516 12248
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14292 9518 14320 10406
rect 14384 10266 14412 10406
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14384 9450 14412 9862
rect 14372 9444 14424 9450
rect 14372 9386 14424 9392
rect 14372 6860 14424 6866
rect 14372 6802 14424 6808
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 14096 5296 14148 5302
rect 14096 5238 14148 5244
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 14108 4010 14136 4966
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 14200 4078 14228 4422
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14096 4004 14148 4010
rect 14096 3946 14148 3952
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 14200 3194 14228 3538
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 13832 870 14044 898
rect 13832 800 13860 870
rect 14292 800 14320 5850
rect 14384 4026 14412 6802
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14476 4146 14504 4966
rect 14568 4826 14596 12650
rect 14660 11778 14688 13126
rect 14752 12374 14780 17972
rect 15106 17912 15162 17921
rect 15106 17847 15162 17856
rect 15120 17202 15148 17847
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 15016 17060 15068 17066
rect 15016 17002 15068 17008
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 14844 15910 14872 16594
rect 15028 16590 15056 17002
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 14832 15904 14884 15910
rect 14832 15846 14884 15852
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 14740 12368 14792 12374
rect 14740 12310 14792 12316
rect 14660 11750 14780 11778
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14556 4820 14608 4826
rect 14556 4762 14608 4768
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14384 3998 14596 4026
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14384 2650 14412 3878
rect 14462 2952 14518 2961
rect 14462 2887 14518 2896
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14476 2394 14504 2887
rect 14568 2514 14596 3998
rect 14660 3058 14688 11630
rect 14752 6322 14780 11750
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14738 5944 14794 5953
rect 14738 5879 14794 5888
rect 14752 5846 14780 5879
rect 14740 5840 14792 5846
rect 14740 5782 14792 5788
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14752 4622 14780 5170
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 14476 2366 14688 2394
rect 14660 800 14688 2366
rect 14752 1834 14780 2790
rect 14844 2009 14872 15846
rect 14936 12442 14964 15846
rect 15028 13870 15056 16526
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15108 15700 15160 15706
rect 15108 15642 15160 15648
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 14924 12436 14976 12442
rect 14924 12378 14976 12384
rect 14924 12300 14976 12306
rect 14924 12242 14976 12248
rect 14936 11830 14964 12242
rect 14924 11824 14976 11830
rect 14924 11766 14976 11772
rect 14936 5166 14964 11766
rect 15028 9897 15056 13806
rect 15120 11762 15148 15642
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15212 10690 15240 16390
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 15304 11801 15332 15914
rect 15580 13802 15608 19200
rect 15948 16454 15976 19200
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 16408 15978 16436 19200
rect 16396 15972 16448 15978
rect 16396 15914 16448 15920
rect 16776 15706 16804 19200
rect 16764 15700 16816 15706
rect 16764 15642 16816 15648
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15290 11792 15346 11801
rect 15290 11727 15346 11736
rect 15120 10662 15240 10690
rect 15120 10606 15148 10662
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15120 10198 15148 10542
rect 15108 10192 15160 10198
rect 15108 10134 15160 10140
rect 15014 9888 15070 9897
rect 15014 9823 15070 9832
rect 15304 9110 15332 11727
rect 15292 9104 15344 9110
rect 15292 9046 15344 9052
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 14936 2582 14964 5102
rect 15028 4758 15056 7686
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 15936 5296 15988 5302
rect 15936 5238 15988 5244
rect 15108 4820 15160 4826
rect 15108 4762 15160 4768
rect 15016 4752 15068 4758
rect 15016 4694 15068 4700
rect 14924 2576 14976 2582
rect 14924 2518 14976 2524
rect 14830 2000 14886 2009
rect 14830 1935 14886 1944
rect 14740 1828 14792 1834
rect 14740 1770 14792 1776
rect 15120 800 15148 4762
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 15488 800 15516 2314
rect 15948 800 15976 5238
rect 16316 800 16344 7142
rect 16764 2916 16816 2922
rect 16764 2858 16816 2864
rect 16776 800 16804 2858
rect 4158 504 4214 513
rect 4158 439 4214 448
rect 4342 0 4398 800
rect 4710 0 4766 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6366 0 6422 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9310 0 9366 800
rect 9678 0 9734 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12622 0 12678 800
rect 12990 0 13046 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 14646 0 14702 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15934 0 15990 800
rect 16302 0 16358 800
rect 16762 0 16818 800
<< via2 >>
rect 2870 19488 2926 19544
rect 1766 16632 1822 16688
rect 1674 16496 1730 16552
rect 1582 12844 1638 12880
rect 3146 17584 3202 17640
rect 2318 16088 2374 16144
rect 1766 15680 1822 15736
rect 3421 17434 3477 17436
rect 3501 17434 3557 17436
rect 3581 17434 3637 17436
rect 3661 17434 3717 17436
rect 3421 17382 3447 17434
rect 3447 17382 3477 17434
rect 3501 17382 3511 17434
rect 3511 17382 3557 17434
rect 3581 17382 3627 17434
rect 3627 17382 3637 17434
rect 3661 17382 3691 17434
rect 3691 17382 3717 17434
rect 3421 17380 3477 17382
rect 3501 17380 3557 17382
rect 3581 17380 3637 17382
rect 3661 17380 3717 17382
rect 3421 16346 3477 16348
rect 3501 16346 3557 16348
rect 3581 16346 3637 16348
rect 3661 16346 3717 16348
rect 3421 16294 3447 16346
rect 3447 16294 3477 16346
rect 3501 16294 3511 16346
rect 3511 16294 3557 16346
rect 3581 16294 3627 16346
rect 3627 16294 3637 16346
rect 3661 16294 3691 16346
rect 3691 16294 3717 16346
rect 3421 16292 3477 16294
rect 3501 16292 3557 16294
rect 3581 16292 3637 16294
rect 3661 16292 3717 16294
rect 4066 18536 4122 18592
rect 2594 14456 2650 14512
rect 1582 12824 1584 12844
rect 1584 12824 1636 12844
rect 1636 12824 1638 12844
rect 2318 10140 2320 10160
rect 2320 10140 2372 10160
rect 2372 10140 2374 10160
rect 2318 10104 2374 10140
rect 2962 13776 3018 13832
rect 1674 9036 1730 9072
rect 1674 9016 1676 9036
rect 1676 9016 1728 9036
rect 1728 9016 1730 9036
rect 2502 8064 2558 8120
rect 1674 7112 1730 7168
rect 1674 6160 1730 6216
rect 1674 4256 1730 4312
rect 3421 15258 3477 15260
rect 3501 15258 3557 15260
rect 3581 15258 3637 15260
rect 3661 15258 3717 15260
rect 3421 15206 3447 15258
rect 3447 15206 3477 15258
rect 3501 15206 3511 15258
rect 3511 15206 3557 15258
rect 3581 15206 3627 15258
rect 3627 15206 3637 15258
rect 3661 15206 3691 15258
rect 3691 15206 3717 15258
rect 3421 15204 3477 15206
rect 3501 15204 3557 15206
rect 3581 15204 3637 15206
rect 3661 15204 3717 15206
rect 3422 14728 3478 14784
rect 3421 14170 3477 14172
rect 3501 14170 3557 14172
rect 3581 14170 3637 14172
rect 3661 14170 3717 14172
rect 3421 14118 3447 14170
rect 3447 14118 3477 14170
rect 3501 14118 3511 14170
rect 3511 14118 3557 14170
rect 3581 14118 3627 14170
rect 3627 14118 3637 14170
rect 3661 14118 3691 14170
rect 3691 14118 3717 14170
rect 3421 14116 3477 14118
rect 3501 14116 3557 14118
rect 3581 14116 3637 14118
rect 3661 14116 3717 14118
rect 3238 11872 3294 11928
rect 3421 13082 3477 13084
rect 3501 13082 3557 13084
rect 3581 13082 3637 13084
rect 3661 13082 3717 13084
rect 3421 13030 3447 13082
rect 3447 13030 3477 13082
rect 3501 13030 3511 13082
rect 3511 13030 3557 13082
rect 3581 13030 3627 13082
rect 3627 13030 3637 13082
rect 3661 13030 3691 13082
rect 3691 13030 3717 13082
rect 3421 13028 3477 13030
rect 3501 13028 3557 13030
rect 3581 13028 3637 13030
rect 3661 13028 3717 13030
rect 5886 16890 5942 16892
rect 5966 16890 6022 16892
rect 6046 16890 6102 16892
rect 6126 16890 6182 16892
rect 5886 16838 5912 16890
rect 5912 16838 5942 16890
rect 5966 16838 5976 16890
rect 5976 16838 6022 16890
rect 6046 16838 6092 16890
rect 6092 16838 6102 16890
rect 6126 16838 6156 16890
rect 6156 16838 6182 16890
rect 5886 16836 5942 16838
rect 5966 16836 6022 16838
rect 6046 16836 6102 16838
rect 6126 16836 6182 16838
rect 4066 14320 4122 14376
rect 3421 11994 3477 11996
rect 3501 11994 3557 11996
rect 3581 11994 3637 11996
rect 3661 11994 3717 11996
rect 3421 11942 3447 11994
rect 3447 11942 3477 11994
rect 3501 11942 3511 11994
rect 3511 11942 3557 11994
rect 3581 11942 3627 11994
rect 3627 11942 3637 11994
rect 3661 11942 3691 11994
rect 3691 11942 3717 11994
rect 3421 11940 3477 11942
rect 3501 11940 3557 11942
rect 3581 11940 3637 11942
rect 3661 11940 3717 11942
rect 3330 11056 3386 11112
rect 3238 10956 3240 10976
rect 3240 10956 3292 10976
rect 3292 10956 3294 10976
rect 3238 10920 3294 10956
rect 3421 10906 3477 10908
rect 3501 10906 3557 10908
rect 3581 10906 3637 10908
rect 3661 10906 3717 10908
rect 3421 10854 3447 10906
rect 3447 10854 3477 10906
rect 3501 10854 3511 10906
rect 3511 10854 3557 10906
rect 3581 10854 3627 10906
rect 3627 10854 3637 10906
rect 3661 10854 3691 10906
rect 3691 10854 3717 10906
rect 3421 10852 3477 10854
rect 3501 10852 3557 10854
rect 3581 10852 3637 10854
rect 3661 10852 3717 10854
rect 2870 9968 2926 10024
rect 3421 9818 3477 9820
rect 3501 9818 3557 9820
rect 3581 9818 3637 9820
rect 3661 9818 3717 9820
rect 3421 9766 3447 9818
rect 3447 9766 3477 9818
rect 3501 9766 3511 9818
rect 3511 9766 3557 9818
rect 3581 9766 3627 9818
rect 3627 9766 3637 9818
rect 3661 9766 3691 9818
rect 3691 9766 3717 9818
rect 3421 9764 3477 9766
rect 3501 9764 3557 9766
rect 3581 9764 3637 9766
rect 3661 9764 3717 9766
rect 2594 5652 2596 5672
rect 2596 5652 2648 5672
rect 2648 5652 2650 5672
rect 2594 5616 2650 5652
rect 2778 5208 2834 5264
rect 1674 3304 1730 3360
rect 3421 8730 3477 8732
rect 3501 8730 3557 8732
rect 3581 8730 3637 8732
rect 3661 8730 3717 8732
rect 3421 8678 3447 8730
rect 3447 8678 3477 8730
rect 3501 8678 3511 8730
rect 3511 8678 3557 8730
rect 3581 8678 3627 8730
rect 3627 8678 3637 8730
rect 3661 8678 3691 8730
rect 3691 8678 3717 8730
rect 3421 8676 3477 8678
rect 3501 8676 3557 8678
rect 3581 8676 3637 8678
rect 3661 8676 3717 8678
rect 3421 7642 3477 7644
rect 3501 7642 3557 7644
rect 3581 7642 3637 7644
rect 3661 7642 3717 7644
rect 3421 7590 3447 7642
rect 3447 7590 3477 7642
rect 3501 7590 3511 7642
rect 3511 7590 3557 7642
rect 3581 7590 3627 7642
rect 3627 7590 3637 7642
rect 3661 7590 3691 7642
rect 3691 7590 3717 7642
rect 3421 7588 3477 7590
rect 3501 7588 3557 7590
rect 3581 7588 3637 7590
rect 3661 7588 3717 7590
rect 3421 6554 3477 6556
rect 3501 6554 3557 6556
rect 3581 6554 3637 6556
rect 3661 6554 3717 6556
rect 3421 6502 3447 6554
rect 3447 6502 3477 6554
rect 3501 6502 3511 6554
rect 3511 6502 3557 6554
rect 3581 6502 3627 6554
rect 3627 6502 3637 6554
rect 3661 6502 3691 6554
rect 3691 6502 3717 6554
rect 3421 6500 3477 6502
rect 3501 6500 3557 6502
rect 3581 6500 3637 6502
rect 3661 6500 3717 6502
rect 3421 5466 3477 5468
rect 3501 5466 3557 5468
rect 3581 5466 3637 5468
rect 3661 5466 3717 5468
rect 3421 5414 3447 5466
rect 3447 5414 3477 5466
rect 3501 5414 3511 5466
rect 3511 5414 3557 5466
rect 3581 5414 3627 5466
rect 3627 5414 3637 5466
rect 3661 5414 3691 5466
rect 3691 5414 3717 5466
rect 3421 5412 3477 5414
rect 3501 5412 3557 5414
rect 3581 5412 3637 5414
rect 3661 5412 3717 5414
rect 2778 1400 2834 1456
rect 3421 4378 3477 4380
rect 3501 4378 3557 4380
rect 3581 4378 3637 4380
rect 3661 4378 3717 4380
rect 3421 4326 3447 4378
rect 3447 4326 3477 4378
rect 3501 4326 3511 4378
rect 3511 4326 3557 4378
rect 3581 4326 3627 4378
rect 3627 4326 3637 4378
rect 3661 4326 3691 4378
rect 3691 4326 3717 4378
rect 3421 4324 3477 4326
rect 3501 4324 3557 4326
rect 3581 4324 3637 4326
rect 3661 4324 3717 4326
rect 3421 3290 3477 3292
rect 3501 3290 3557 3292
rect 3581 3290 3637 3292
rect 3661 3290 3717 3292
rect 3421 3238 3447 3290
rect 3447 3238 3477 3290
rect 3501 3238 3511 3290
rect 3511 3238 3557 3290
rect 3581 3238 3627 3290
rect 3627 3238 3637 3290
rect 3661 3238 3691 3290
rect 3691 3238 3717 3290
rect 3421 3236 3477 3238
rect 3501 3236 3557 3238
rect 3581 3236 3637 3238
rect 3661 3236 3717 3238
rect 3421 2202 3477 2204
rect 3501 2202 3557 2204
rect 3581 2202 3637 2204
rect 3661 2202 3717 2204
rect 3421 2150 3447 2202
rect 3447 2150 3477 2202
rect 3501 2150 3511 2202
rect 3511 2150 3557 2202
rect 3581 2150 3627 2202
rect 3627 2150 3637 2202
rect 3661 2150 3691 2202
rect 3691 2150 3717 2202
rect 3421 2148 3477 2150
rect 3501 2148 3557 2150
rect 3581 2148 3637 2150
rect 3661 2148 3717 2150
rect 4066 7928 4122 7984
rect 4802 14900 4804 14920
rect 4804 14900 4856 14920
rect 4856 14900 4858 14920
rect 4802 14864 4858 14900
rect 4342 8064 4398 8120
rect 4802 8064 4858 8120
rect 5262 15408 5318 15464
rect 5886 15802 5942 15804
rect 5966 15802 6022 15804
rect 6046 15802 6102 15804
rect 6126 15802 6182 15804
rect 5886 15750 5912 15802
rect 5912 15750 5942 15802
rect 5966 15750 5976 15802
rect 5976 15750 6022 15802
rect 6046 15750 6092 15802
rect 6092 15750 6102 15802
rect 6126 15750 6156 15802
rect 6156 15750 6182 15802
rect 5886 15748 5942 15750
rect 5966 15748 6022 15750
rect 6046 15748 6102 15750
rect 6126 15748 6182 15750
rect 5886 14714 5942 14716
rect 5966 14714 6022 14716
rect 6046 14714 6102 14716
rect 6126 14714 6182 14716
rect 5886 14662 5912 14714
rect 5912 14662 5942 14714
rect 5966 14662 5976 14714
rect 5976 14662 6022 14714
rect 6046 14662 6092 14714
rect 6092 14662 6102 14714
rect 6126 14662 6156 14714
rect 6156 14662 6182 14714
rect 5886 14660 5942 14662
rect 5966 14660 6022 14662
rect 6046 14660 6102 14662
rect 6126 14660 6182 14662
rect 6274 14456 6330 14512
rect 5886 13626 5942 13628
rect 5966 13626 6022 13628
rect 6046 13626 6102 13628
rect 6126 13626 6182 13628
rect 5886 13574 5912 13626
rect 5912 13574 5942 13626
rect 5966 13574 5976 13626
rect 5976 13574 6022 13626
rect 6046 13574 6092 13626
rect 6092 13574 6102 13626
rect 6126 13574 6156 13626
rect 6156 13574 6182 13626
rect 5886 13572 5942 13574
rect 5966 13572 6022 13574
rect 6046 13572 6102 13574
rect 6126 13572 6182 13574
rect 5630 12824 5686 12880
rect 6366 12552 6422 12608
rect 5886 12538 5942 12540
rect 5966 12538 6022 12540
rect 6046 12538 6102 12540
rect 6126 12538 6182 12540
rect 5886 12486 5912 12538
rect 5912 12486 5942 12538
rect 5966 12486 5976 12538
rect 5976 12486 6022 12538
rect 6046 12486 6092 12538
rect 6092 12486 6102 12538
rect 6126 12486 6156 12538
rect 6156 12486 6182 12538
rect 5886 12484 5942 12486
rect 5966 12484 6022 12486
rect 6046 12484 6102 12486
rect 6126 12484 6182 12486
rect 5886 11450 5942 11452
rect 5966 11450 6022 11452
rect 6046 11450 6102 11452
rect 6126 11450 6182 11452
rect 5886 11398 5912 11450
rect 5912 11398 5942 11450
rect 5966 11398 5976 11450
rect 5976 11398 6022 11450
rect 6046 11398 6092 11450
rect 6092 11398 6102 11450
rect 6126 11398 6156 11450
rect 6156 11398 6182 11450
rect 5886 11396 5942 11398
rect 5966 11396 6022 11398
rect 6046 11396 6102 11398
rect 6126 11396 6182 11398
rect 5262 10104 5318 10160
rect 4802 6704 4858 6760
rect 5886 10362 5942 10364
rect 5966 10362 6022 10364
rect 6046 10362 6102 10364
rect 6126 10362 6182 10364
rect 5886 10310 5912 10362
rect 5912 10310 5942 10362
rect 5966 10310 5976 10362
rect 5976 10310 6022 10362
rect 6046 10310 6092 10362
rect 6092 10310 6102 10362
rect 6126 10310 6156 10362
rect 6156 10310 6182 10362
rect 5886 10308 5942 10310
rect 5966 10308 6022 10310
rect 6046 10308 6102 10310
rect 6126 10308 6182 10310
rect 5886 9274 5942 9276
rect 5966 9274 6022 9276
rect 6046 9274 6102 9276
rect 6126 9274 6182 9276
rect 5886 9222 5912 9274
rect 5912 9222 5942 9274
rect 5966 9222 5976 9274
rect 5976 9222 6022 9274
rect 6046 9222 6092 9274
rect 6092 9222 6102 9274
rect 6126 9222 6156 9274
rect 6156 9222 6182 9274
rect 5886 9220 5942 9222
rect 5966 9220 6022 9222
rect 6046 9220 6102 9222
rect 6126 9220 6182 9222
rect 8352 17434 8408 17436
rect 8432 17434 8488 17436
rect 8512 17434 8568 17436
rect 8592 17434 8648 17436
rect 8352 17382 8378 17434
rect 8378 17382 8408 17434
rect 8432 17382 8442 17434
rect 8442 17382 8488 17434
rect 8512 17382 8558 17434
rect 8558 17382 8568 17434
rect 8592 17382 8622 17434
rect 8622 17382 8648 17434
rect 8352 17380 8408 17382
rect 8432 17380 8488 17382
rect 8512 17380 8568 17382
rect 8592 17380 8648 17382
rect 7194 14456 7250 14512
rect 7746 15020 7802 15056
rect 7746 15000 7748 15020
rect 7748 15000 7800 15020
rect 7800 15000 7802 15020
rect 6918 12688 6974 12744
rect 5886 8186 5942 8188
rect 5966 8186 6022 8188
rect 6046 8186 6102 8188
rect 6126 8186 6182 8188
rect 5886 8134 5912 8186
rect 5912 8134 5942 8186
rect 5966 8134 5976 8186
rect 5976 8134 6022 8186
rect 6046 8134 6092 8186
rect 6092 8134 6102 8186
rect 6126 8134 6156 8186
rect 6156 8134 6182 8186
rect 5886 8132 5942 8134
rect 5966 8132 6022 8134
rect 6046 8132 6102 8134
rect 6126 8132 6182 8134
rect 5886 7098 5942 7100
rect 5966 7098 6022 7100
rect 6046 7098 6102 7100
rect 6126 7098 6182 7100
rect 5886 7046 5912 7098
rect 5912 7046 5942 7098
rect 5966 7046 5976 7098
rect 5976 7046 6022 7098
rect 6046 7046 6092 7098
rect 6092 7046 6102 7098
rect 6126 7046 6156 7098
rect 6156 7046 6182 7098
rect 5886 7044 5942 7046
rect 5966 7044 6022 7046
rect 6046 7044 6102 7046
rect 6126 7044 6182 7046
rect 4434 3596 4490 3632
rect 4434 3576 4436 3596
rect 4436 3576 4488 3596
rect 4488 3576 4490 3596
rect 4894 3984 4950 4040
rect 4802 3032 4858 3088
rect 4710 2932 4712 2952
rect 4712 2932 4764 2952
rect 4764 2932 4766 2952
rect 4710 2896 4766 2932
rect 4066 2352 4122 2408
rect 5354 3984 5410 4040
rect 6182 6180 6238 6216
rect 6182 6160 6184 6180
rect 6184 6160 6236 6180
rect 6236 6160 6238 6180
rect 5886 6010 5942 6012
rect 5966 6010 6022 6012
rect 6046 6010 6102 6012
rect 6126 6010 6182 6012
rect 5886 5958 5912 6010
rect 5912 5958 5942 6010
rect 5966 5958 5976 6010
rect 5976 5958 6022 6010
rect 6046 5958 6092 6010
rect 6092 5958 6102 6010
rect 6126 5958 6156 6010
rect 6156 5958 6182 6010
rect 5886 5956 5942 5958
rect 5966 5956 6022 5958
rect 6046 5956 6102 5958
rect 6126 5956 6182 5958
rect 6734 6704 6790 6760
rect 6642 6160 6698 6216
rect 5886 4922 5942 4924
rect 5966 4922 6022 4924
rect 6046 4922 6102 4924
rect 6126 4922 6182 4924
rect 5886 4870 5912 4922
rect 5912 4870 5942 4922
rect 5966 4870 5976 4922
rect 5976 4870 6022 4922
rect 6046 4870 6092 4922
rect 6092 4870 6102 4922
rect 6126 4870 6156 4922
rect 6156 4870 6182 4922
rect 5886 4868 5942 4870
rect 5966 4868 6022 4870
rect 6046 4868 6102 4870
rect 6126 4868 6182 4870
rect 5886 3834 5942 3836
rect 5966 3834 6022 3836
rect 6046 3834 6102 3836
rect 6126 3834 6182 3836
rect 5886 3782 5912 3834
rect 5912 3782 5942 3834
rect 5966 3782 5976 3834
rect 5976 3782 6022 3834
rect 6046 3782 6092 3834
rect 6092 3782 6102 3834
rect 6126 3782 6156 3834
rect 6156 3782 6182 3834
rect 5886 3780 5942 3782
rect 5966 3780 6022 3782
rect 6046 3780 6102 3782
rect 6126 3780 6182 3782
rect 7286 5752 7342 5808
rect 8352 16346 8408 16348
rect 8432 16346 8488 16348
rect 8512 16346 8568 16348
rect 8592 16346 8648 16348
rect 8352 16294 8378 16346
rect 8378 16294 8408 16346
rect 8432 16294 8442 16346
rect 8442 16294 8488 16346
rect 8512 16294 8558 16346
rect 8558 16294 8568 16346
rect 8592 16294 8622 16346
rect 8622 16294 8648 16346
rect 8352 16292 8408 16294
rect 8432 16292 8488 16294
rect 8512 16292 8568 16294
rect 8592 16292 8648 16294
rect 8352 15258 8408 15260
rect 8432 15258 8488 15260
rect 8512 15258 8568 15260
rect 8592 15258 8648 15260
rect 8352 15206 8378 15258
rect 8378 15206 8408 15258
rect 8432 15206 8442 15258
rect 8442 15206 8488 15258
rect 8512 15206 8558 15258
rect 8558 15206 8568 15258
rect 8592 15206 8622 15258
rect 8622 15206 8648 15258
rect 8352 15204 8408 15206
rect 8432 15204 8488 15206
rect 8512 15204 8568 15206
rect 8592 15204 8648 15206
rect 9126 16496 9182 16552
rect 8352 14170 8408 14172
rect 8432 14170 8488 14172
rect 8512 14170 8568 14172
rect 8592 14170 8648 14172
rect 8352 14118 8378 14170
rect 8378 14118 8408 14170
rect 8432 14118 8442 14170
rect 8442 14118 8488 14170
rect 8512 14118 8558 14170
rect 8558 14118 8568 14170
rect 8592 14118 8622 14170
rect 8622 14118 8648 14170
rect 8352 14116 8408 14118
rect 8432 14116 8488 14118
rect 8512 14116 8568 14118
rect 8592 14116 8648 14118
rect 8758 14864 8814 14920
rect 8850 14456 8906 14512
rect 8352 13082 8408 13084
rect 8432 13082 8488 13084
rect 8512 13082 8568 13084
rect 8592 13082 8648 13084
rect 8352 13030 8378 13082
rect 8378 13030 8408 13082
rect 8432 13030 8442 13082
rect 8442 13030 8488 13082
rect 8512 13030 8558 13082
rect 8558 13030 8568 13082
rect 8592 13030 8622 13082
rect 8622 13030 8648 13082
rect 8352 13028 8408 13030
rect 8432 13028 8488 13030
rect 8512 13028 8568 13030
rect 8592 13028 8648 13030
rect 8022 12280 8078 12336
rect 8352 11994 8408 11996
rect 8432 11994 8488 11996
rect 8512 11994 8568 11996
rect 8592 11994 8648 11996
rect 8352 11942 8378 11994
rect 8378 11942 8408 11994
rect 8432 11942 8442 11994
rect 8442 11942 8488 11994
rect 8512 11942 8558 11994
rect 8558 11942 8568 11994
rect 8592 11942 8622 11994
rect 8622 11942 8648 11994
rect 8352 11940 8408 11942
rect 8432 11940 8488 11942
rect 8512 11940 8568 11942
rect 8592 11940 8648 11942
rect 8666 11736 8722 11792
rect 8352 10906 8408 10908
rect 8432 10906 8488 10908
rect 8512 10906 8568 10908
rect 8592 10906 8648 10908
rect 8352 10854 8378 10906
rect 8378 10854 8408 10906
rect 8432 10854 8442 10906
rect 8442 10854 8488 10906
rect 8512 10854 8558 10906
rect 8558 10854 8568 10906
rect 8592 10854 8622 10906
rect 8622 10854 8648 10906
rect 8352 10852 8408 10854
rect 8432 10852 8488 10854
rect 8512 10852 8568 10854
rect 8592 10852 8648 10854
rect 8022 10104 8078 10160
rect 9126 12688 9182 12744
rect 8352 9818 8408 9820
rect 8432 9818 8488 9820
rect 8512 9818 8568 9820
rect 8592 9818 8648 9820
rect 8352 9766 8378 9818
rect 8378 9766 8408 9818
rect 8432 9766 8442 9818
rect 8442 9766 8488 9818
rect 8512 9766 8558 9818
rect 8558 9766 8568 9818
rect 8592 9766 8622 9818
rect 8622 9766 8648 9818
rect 8352 9764 8408 9766
rect 8432 9764 8488 9766
rect 8512 9764 8568 9766
rect 8592 9764 8648 9766
rect 7562 8472 7618 8528
rect 6918 5616 6974 5672
rect 6366 3576 6422 3632
rect 5886 2746 5942 2748
rect 5966 2746 6022 2748
rect 6046 2746 6102 2748
rect 6126 2746 6182 2748
rect 5886 2694 5912 2746
rect 5912 2694 5942 2746
rect 5966 2694 5976 2746
rect 5976 2694 6022 2746
rect 6046 2694 6092 2746
rect 6092 2694 6102 2746
rect 6126 2694 6156 2746
rect 6156 2694 6182 2746
rect 5886 2692 5942 2694
rect 5966 2692 6022 2694
rect 6046 2692 6102 2694
rect 6126 2692 6182 2694
rect 6642 3732 6698 3768
rect 6642 3712 6644 3732
rect 6644 3712 6696 3732
rect 6696 3712 6698 3732
rect 5538 856 5594 912
rect 8352 8730 8408 8732
rect 8432 8730 8488 8732
rect 8512 8730 8568 8732
rect 8592 8730 8648 8732
rect 8352 8678 8378 8730
rect 8378 8678 8408 8730
rect 8432 8678 8442 8730
rect 8442 8678 8488 8730
rect 8512 8678 8558 8730
rect 8558 8678 8568 8730
rect 8592 8678 8622 8730
rect 8622 8678 8648 8730
rect 8352 8676 8408 8678
rect 8432 8676 8488 8678
rect 8512 8676 8568 8678
rect 8592 8676 8648 8678
rect 8482 7792 8538 7848
rect 8352 7642 8408 7644
rect 8432 7642 8488 7644
rect 8512 7642 8568 7644
rect 8592 7642 8648 7644
rect 8352 7590 8378 7642
rect 8378 7590 8408 7642
rect 8432 7590 8442 7642
rect 8442 7590 8488 7642
rect 8512 7590 8558 7642
rect 8558 7590 8568 7642
rect 8592 7590 8622 7642
rect 8622 7590 8648 7642
rect 8352 7588 8408 7590
rect 8432 7588 8488 7590
rect 8512 7588 8568 7590
rect 8592 7588 8648 7590
rect 8850 8064 8906 8120
rect 8352 6554 8408 6556
rect 8432 6554 8488 6556
rect 8512 6554 8568 6556
rect 8592 6554 8648 6556
rect 8352 6502 8378 6554
rect 8378 6502 8408 6554
rect 8432 6502 8442 6554
rect 8442 6502 8488 6554
rect 8512 6502 8558 6554
rect 8558 6502 8568 6554
rect 8592 6502 8622 6554
rect 8622 6502 8648 6554
rect 8352 6500 8408 6502
rect 8432 6500 8488 6502
rect 8512 6500 8568 6502
rect 8592 6500 8648 6502
rect 8390 6196 8392 6216
rect 8392 6196 8444 6216
rect 8444 6196 8446 6216
rect 8390 6160 8446 6196
rect 7930 5652 7932 5672
rect 7932 5652 7984 5672
rect 7984 5652 7986 5672
rect 7930 5616 7986 5652
rect 8352 5466 8408 5468
rect 8432 5466 8488 5468
rect 8512 5466 8568 5468
rect 8592 5466 8648 5468
rect 8352 5414 8378 5466
rect 8378 5414 8408 5466
rect 8432 5414 8442 5466
rect 8442 5414 8488 5466
rect 8512 5414 8558 5466
rect 8558 5414 8568 5466
rect 8592 5414 8622 5466
rect 8622 5414 8648 5466
rect 8352 5412 8408 5414
rect 8432 5412 8488 5414
rect 8512 5412 8568 5414
rect 8592 5412 8648 5414
rect 9218 12552 9274 12608
rect 9402 15408 9458 15464
rect 9862 16496 9918 16552
rect 9586 16088 9642 16144
rect 9402 11600 9458 11656
rect 9954 15408 10010 15464
rect 10230 15000 10286 15056
rect 9494 11056 9550 11112
rect 9862 12552 9918 12608
rect 9402 10240 9458 10296
rect 9402 9968 9458 10024
rect 10414 15444 10416 15464
rect 10416 15444 10468 15464
rect 10468 15444 10470 15464
rect 10414 15408 10470 15444
rect 10817 16890 10873 16892
rect 10897 16890 10953 16892
rect 10977 16890 11033 16892
rect 11057 16890 11113 16892
rect 10817 16838 10843 16890
rect 10843 16838 10873 16890
rect 10897 16838 10907 16890
rect 10907 16838 10953 16890
rect 10977 16838 11023 16890
rect 11023 16838 11033 16890
rect 11057 16838 11087 16890
rect 11087 16838 11113 16890
rect 10817 16836 10873 16838
rect 10897 16836 10953 16838
rect 10977 16836 11033 16838
rect 11057 16836 11113 16838
rect 11150 16632 11206 16688
rect 10817 15802 10873 15804
rect 10897 15802 10953 15804
rect 10977 15802 11033 15804
rect 11057 15802 11113 15804
rect 10817 15750 10843 15802
rect 10843 15750 10873 15802
rect 10897 15750 10907 15802
rect 10907 15750 10953 15802
rect 10977 15750 11023 15802
rect 11023 15750 11033 15802
rect 11057 15750 11087 15802
rect 11087 15750 11113 15802
rect 10817 15748 10873 15750
rect 10897 15748 10953 15750
rect 10977 15748 11033 15750
rect 11057 15748 11113 15750
rect 11426 16768 11482 16824
rect 10817 14714 10873 14716
rect 10897 14714 10953 14716
rect 10977 14714 11033 14716
rect 11057 14714 11113 14716
rect 10817 14662 10843 14714
rect 10843 14662 10873 14714
rect 10897 14662 10907 14714
rect 10907 14662 10953 14714
rect 10977 14662 11023 14714
rect 11023 14662 11033 14714
rect 11057 14662 11087 14714
rect 11087 14662 11113 14714
rect 10817 14660 10873 14662
rect 10897 14660 10953 14662
rect 10977 14660 11033 14662
rect 11057 14660 11113 14662
rect 10966 14320 11022 14376
rect 10817 13626 10873 13628
rect 10897 13626 10953 13628
rect 10977 13626 11033 13628
rect 11057 13626 11113 13628
rect 10817 13574 10843 13626
rect 10843 13574 10873 13626
rect 10897 13574 10907 13626
rect 10907 13574 10953 13626
rect 10977 13574 11023 13626
rect 11023 13574 11033 13626
rect 11057 13574 11087 13626
rect 11087 13574 11113 13626
rect 10817 13572 10873 13574
rect 10897 13572 10953 13574
rect 10977 13572 11033 13574
rect 11057 13572 11113 13574
rect 11150 12688 11206 12744
rect 10817 12538 10873 12540
rect 10897 12538 10953 12540
rect 10977 12538 11033 12540
rect 11057 12538 11113 12540
rect 10817 12486 10843 12538
rect 10843 12486 10873 12538
rect 10897 12486 10907 12538
rect 10907 12486 10953 12538
rect 10977 12486 11023 12538
rect 11023 12486 11033 12538
rect 11057 12486 11087 12538
rect 11087 12486 11113 12538
rect 10817 12484 10873 12486
rect 10897 12484 10953 12486
rect 10977 12484 11033 12486
rect 11057 12484 11113 12486
rect 10506 12280 10562 12336
rect 9862 9696 9918 9752
rect 9586 8200 9642 8256
rect 9862 9016 9918 9072
rect 9586 7792 9642 7848
rect 7010 856 7066 912
rect 8352 4378 8408 4380
rect 8432 4378 8488 4380
rect 8512 4378 8568 4380
rect 8592 4378 8648 4380
rect 8352 4326 8378 4378
rect 8378 4326 8408 4378
rect 8432 4326 8442 4378
rect 8442 4326 8488 4378
rect 8512 4326 8558 4378
rect 8558 4326 8568 4378
rect 8592 4326 8622 4378
rect 8622 4326 8648 4378
rect 8352 4324 8408 4326
rect 8432 4324 8488 4326
rect 8512 4324 8568 4326
rect 8592 4324 8648 4326
rect 7930 2760 7986 2816
rect 8352 3290 8408 3292
rect 8432 3290 8488 3292
rect 8512 3290 8568 3292
rect 8592 3290 8648 3292
rect 8352 3238 8378 3290
rect 8378 3238 8408 3290
rect 8432 3238 8442 3290
rect 8442 3238 8488 3290
rect 8512 3238 8558 3290
rect 8558 3238 8568 3290
rect 8592 3238 8622 3290
rect 8622 3238 8648 3290
rect 8352 3236 8408 3238
rect 8432 3236 8488 3238
rect 8512 3236 8568 3238
rect 8592 3236 8648 3238
rect 8850 2760 8906 2816
rect 8352 2202 8408 2204
rect 8432 2202 8488 2204
rect 8512 2202 8568 2204
rect 8592 2202 8648 2204
rect 8352 2150 8378 2202
rect 8378 2150 8408 2202
rect 8432 2150 8442 2202
rect 8442 2150 8488 2202
rect 8512 2150 8558 2202
rect 8558 2150 8568 2202
rect 8592 2150 8622 2202
rect 8622 2150 8648 2202
rect 8352 2148 8408 2150
rect 8432 2148 8488 2150
rect 8512 2148 8568 2150
rect 8592 2148 8648 2150
rect 10138 7384 10194 7440
rect 10506 9016 10562 9072
rect 10874 12280 10930 12336
rect 11058 11620 11114 11656
rect 11058 11600 11060 11620
rect 11060 11600 11112 11620
rect 11112 11600 11114 11620
rect 10817 11450 10873 11452
rect 10897 11450 10953 11452
rect 10977 11450 11033 11452
rect 11057 11450 11113 11452
rect 10817 11398 10843 11450
rect 10843 11398 10873 11450
rect 10897 11398 10907 11450
rect 10907 11398 10953 11450
rect 10977 11398 11023 11450
rect 11023 11398 11033 11450
rect 11057 11398 11087 11450
rect 11087 11398 11113 11450
rect 10817 11396 10873 11398
rect 10897 11396 10953 11398
rect 10977 11396 11033 11398
rect 11057 11396 11113 11398
rect 10874 11092 10876 11112
rect 10876 11092 10928 11112
rect 10928 11092 10930 11112
rect 10874 11056 10930 11092
rect 10817 10362 10873 10364
rect 10897 10362 10953 10364
rect 10977 10362 11033 10364
rect 11057 10362 11113 10364
rect 10817 10310 10843 10362
rect 10843 10310 10873 10362
rect 10897 10310 10907 10362
rect 10907 10310 10953 10362
rect 10977 10310 11023 10362
rect 11023 10310 11033 10362
rect 11057 10310 11087 10362
rect 11087 10310 11113 10362
rect 10817 10308 10873 10310
rect 10897 10308 10953 10310
rect 10977 10308 11033 10310
rect 11057 10308 11113 10310
rect 10690 9696 10746 9752
rect 11242 10104 11298 10160
rect 11150 9560 11206 9616
rect 10817 9274 10873 9276
rect 10897 9274 10953 9276
rect 10977 9274 11033 9276
rect 11057 9274 11113 9276
rect 10817 9222 10843 9274
rect 10843 9222 10873 9274
rect 10897 9222 10907 9274
rect 10907 9222 10953 9274
rect 10977 9222 11023 9274
rect 11023 9222 11033 9274
rect 11057 9222 11087 9274
rect 11087 9222 11113 9274
rect 10817 9220 10873 9222
rect 10897 9220 10953 9222
rect 10977 9220 11033 9222
rect 11057 9220 11113 9222
rect 10138 6296 10194 6352
rect 9770 3712 9826 3768
rect 9494 2624 9550 2680
rect 10414 5616 10470 5672
rect 10817 8186 10873 8188
rect 10897 8186 10953 8188
rect 10977 8186 11033 8188
rect 11057 8186 11113 8188
rect 10817 8134 10843 8186
rect 10843 8134 10873 8186
rect 10897 8134 10907 8186
rect 10907 8134 10953 8186
rect 10977 8134 11023 8186
rect 11023 8134 11033 8186
rect 11057 8134 11087 8186
rect 11087 8134 11113 8186
rect 10817 8132 10873 8134
rect 10897 8132 10953 8134
rect 10977 8132 11033 8134
rect 11057 8132 11113 8134
rect 11518 9968 11574 10024
rect 10690 7384 10746 7440
rect 10817 7098 10873 7100
rect 10897 7098 10953 7100
rect 10977 7098 11033 7100
rect 11057 7098 11113 7100
rect 10817 7046 10843 7098
rect 10843 7046 10873 7098
rect 10897 7046 10907 7098
rect 10907 7046 10953 7098
rect 10977 7046 11023 7098
rect 11023 7046 11033 7098
rect 11057 7046 11087 7098
rect 11087 7046 11113 7098
rect 10817 7044 10873 7046
rect 10897 7044 10953 7046
rect 10977 7044 11033 7046
rect 11057 7044 11113 7046
rect 11610 7928 11666 7984
rect 11334 7384 11390 7440
rect 10598 5752 10654 5808
rect 10230 3168 10286 3224
rect 10817 6010 10873 6012
rect 10897 6010 10953 6012
rect 10977 6010 11033 6012
rect 11057 6010 11113 6012
rect 10817 5958 10843 6010
rect 10843 5958 10873 6010
rect 10897 5958 10907 6010
rect 10907 5958 10953 6010
rect 10977 5958 11023 6010
rect 11023 5958 11033 6010
rect 11057 5958 11087 6010
rect 11087 5958 11113 6010
rect 10817 5956 10873 5958
rect 10897 5956 10953 5958
rect 10977 5956 11033 5958
rect 11057 5956 11113 5958
rect 10782 5772 10838 5808
rect 10782 5752 10784 5772
rect 10784 5752 10836 5772
rect 10836 5752 10838 5772
rect 10817 4922 10873 4924
rect 10897 4922 10953 4924
rect 10977 4922 11033 4924
rect 11057 4922 11113 4924
rect 10817 4870 10843 4922
rect 10843 4870 10873 4922
rect 10897 4870 10907 4922
rect 10907 4870 10953 4922
rect 10977 4870 11023 4922
rect 11023 4870 11033 4922
rect 11057 4870 11087 4922
rect 11087 4870 11113 4922
rect 10817 4868 10873 4870
rect 10897 4868 10953 4870
rect 10977 4868 11033 4870
rect 11057 4868 11113 4870
rect 10782 4020 10784 4040
rect 10784 4020 10836 4040
rect 10836 4020 10838 4040
rect 10782 3984 10838 4020
rect 10322 2760 10378 2816
rect 10817 3834 10873 3836
rect 10897 3834 10953 3836
rect 10977 3834 11033 3836
rect 11057 3834 11113 3836
rect 10817 3782 10843 3834
rect 10843 3782 10873 3834
rect 10897 3782 10907 3834
rect 10907 3782 10953 3834
rect 10977 3782 11023 3834
rect 11023 3782 11033 3834
rect 11057 3782 11087 3834
rect 11087 3782 11113 3834
rect 10817 3780 10873 3782
rect 10897 3780 10953 3782
rect 10977 3780 11033 3782
rect 11057 3780 11113 3782
rect 11426 3168 11482 3224
rect 10817 2746 10873 2748
rect 10897 2746 10953 2748
rect 10977 2746 11033 2748
rect 11057 2746 11113 2748
rect 10817 2694 10843 2746
rect 10843 2694 10873 2746
rect 10897 2694 10907 2746
rect 10907 2694 10953 2746
rect 10977 2694 11023 2746
rect 11023 2694 11033 2746
rect 11057 2694 11087 2746
rect 11087 2694 11113 2746
rect 10817 2692 10873 2694
rect 10897 2692 10953 2694
rect 10977 2692 11033 2694
rect 11057 2692 11113 2694
rect 13282 17434 13338 17436
rect 13362 17434 13418 17436
rect 13442 17434 13498 17436
rect 13522 17434 13578 17436
rect 13282 17382 13308 17434
rect 13308 17382 13338 17434
rect 13362 17382 13372 17434
rect 13372 17382 13418 17434
rect 13442 17382 13488 17434
rect 13488 17382 13498 17434
rect 13522 17382 13552 17434
rect 13552 17382 13578 17434
rect 13282 17380 13338 17382
rect 13362 17380 13418 17382
rect 13442 17380 13498 17382
rect 13522 17380 13578 17382
rect 13282 16346 13338 16348
rect 13362 16346 13418 16348
rect 13442 16346 13498 16348
rect 13522 16346 13578 16348
rect 13282 16294 13308 16346
rect 13308 16294 13338 16346
rect 13362 16294 13372 16346
rect 13372 16294 13418 16346
rect 13442 16294 13488 16346
rect 13488 16294 13498 16346
rect 13522 16294 13552 16346
rect 13552 16294 13578 16346
rect 13282 16292 13338 16294
rect 13362 16292 13418 16294
rect 13442 16292 13498 16294
rect 13522 16292 13578 16294
rect 11610 3576 11666 3632
rect 13282 15258 13338 15260
rect 13362 15258 13418 15260
rect 13442 15258 13498 15260
rect 13522 15258 13578 15260
rect 13282 15206 13308 15258
rect 13308 15206 13338 15258
rect 13362 15206 13372 15258
rect 13372 15206 13418 15258
rect 13442 15206 13488 15258
rect 13488 15206 13498 15258
rect 13522 15206 13552 15258
rect 13552 15206 13578 15258
rect 13282 15204 13338 15206
rect 13362 15204 13418 15206
rect 13442 15204 13498 15206
rect 13522 15204 13578 15206
rect 13266 14456 13322 14512
rect 13282 14170 13338 14172
rect 13362 14170 13418 14172
rect 13442 14170 13498 14172
rect 13522 14170 13578 14172
rect 13282 14118 13308 14170
rect 13308 14118 13338 14170
rect 13362 14118 13372 14170
rect 13372 14118 13418 14170
rect 13442 14118 13488 14170
rect 13488 14118 13498 14170
rect 13522 14118 13552 14170
rect 13552 14118 13578 14170
rect 13282 14116 13338 14118
rect 13362 14116 13418 14118
rect 13442 14116 13498 14118
rect 13522 14116 13578 14118
rect 13282 13082 13338 13084
rect 13362 13082 13418 13084
rect 13442 13082 13498 13084
rect 13522 13082 13578 13084
rect 13282 13030 13308 13082
rect 13308 13030 13338 13082
rect 13362 13030 13372 13082
rect 13372 13030 13418 13082
rect 13442 13030 13488 13082
rect 13488 13030 13498 13082
rect 13522 13030 13552 13082
rect 13552 13030 13578 13082
rect 13282 13028 13338 13030
rect 13362 13028 13418 13030
rect 13442 13028 13498 13030
rect 13522 13028 13578 13030
rect 12806 8472 12862 8528
rect 12990 8880 13046 8936
rect 13282 11994 13338 11996
rect 13362 11994 13418 11996
rect 13442 11994 13498 11996
rect 13522 11994 13578 11996
rect 13282 11942 13308 11994
rect 13308 11942 13338 11994
rect 13362 11942 13372 11994
rect 13372 11942 13418 11994
rect 13442 11942 13488 11994
rect 13488 11942 13498 11994
rect 13522 11942 13552 11994
rect 13552 11942 13578 11994
rect 13282 11940 13338 11942
rect 13362 11940 13418 11942
rect 13442 11940 13498 11942
rect 13522 11940 13578 11942
rect 13282 10906 13338 10908
rect 13362 10906 13418 10908
rect 13442 10906 13498 10908
rect 13522 10906 13578 10908
rect 13282 10854 13308 10906
rect 13308 10854 13338 10906
rect 13362 10854 13372 10906
rect 13372 10854 13418 10906
rect 13442 10854 13488 10906
rect 13488 10854 13498 10906
rect 13522 10854 13552 10906
rect 13552 10854 13578 10906
rect 13282 10852 13338 10854
rect 13362 10852 13418 10854
rect 13442 10852 13498 10854
rect 13522 10852 13578 10854
rect 13726 13912 13782 13968
rect 13282 9818 13338 9820
rect 13362 9818 13418 9820
rect 13442 9818 13498 9820
rect 13522 9818 13578 9820
rect 13282 9766 13308 9818
rect 13308 9766 13338 9818
rect 13362 9766 13372 9818
rect 13372 9766 13418 9818
rect 13442 9766 13488 9818
rect 13488 9766 13498 9818
rect 13522 9766 13552 9818
rect 13552 9766 13578 9818
rect 13282 9764 13338 9766
rect 13362 9764 13418 9766
rect 13442 9764 13498 9766
rect 13522 9764 13578 9766
rect 13282 8730 13338 8732
rect 13362 8730 13418 8732
rect 13442 8730 13498 8732
rect 13522 8730 13578 8732
rect 13282 8678 13308 8730
rect 13308 8678 13338 8730
rect 13362 8678 13372 8730
rect 13372 8678 13418 8730
rect 13442 8678 13488 8730
rect 13488 8678 13498 8730
rect 13522 8678 13552 8730
rect 13552 8678 13578 8730
rect 13282 8676 13338 8678
rect 13362 8676 13418 8678
rect 13442 8676 13498 8678
rect 13522 8676 13578 8678
rect 13282 7642 13338 7644
rect 13362 7642 13418 7644
rect 13442 7642 13498 7644
rect 13522 7642 13578 7644
rect 13282 7590 13308 7642
rect 13308 7590 13338 7642
rect 13362 7590 13372 7642
rect 13372 7590 13418 7642
rect 13442 7590 13488 7642
rect 13488 7590 13498 7642
rect 13522 7590 13552 7642
rect 13552 7590 13578 7642
rect 13282 7588 13338 7590
rect 13362 7588 13418 7590
rect 13442 7588 13498 7590
rect 13522 7588 13578 7590
rect 13726 8880 13782 8936
rect 13282 6554 13338 6556
rect 13362 6554 13418 6556
rect 13442 6554 13498 6556
rect 13522 6554 13578 6556
rect 13282 6502 13308 6554
rect 13308 6502 13338 6554
rect 13362 6502 13372 6554
rect 13372 6502 13418 6554
rect 13442 6502 13488 6554
rect 13488 6502 13498 6554
rect 13522 6502 13552 6554
rect 13552 6502 13578 6554
rect 13282 6500 13338 6502
rect 13362 6500 13418 6502
rect 13442 6500 13498 6502
rect 13522 6500 13578 6502
rect 13282 5466 13338 5468
rect 13362 5466 13418 5468
rect 13442 5466 13498 5468
rect 13522 5466 13578 5468
rect 13282 5414 13308 5466
rect 13308 5414 13338 5466
rect 13362 5414 13372 5466
rect 13372 5414 13418 5466
rect 13442 5414 13488 5466
rect 13488 5414 13498 5466
rect 13522 5414 13552 5466
rect 13552 5414 13578 5466
rect 13282 5412 13338 5414
rect 13362 5412 13418 5414
rect 13442 5412 13498 5414
rect 13522 5412 13578 5414
rect 14094 9560 14150 9616
rect 13282 4378 13338 4380
rect 13362 4378 13418 4380
rect 13442 4378 13498 4380
rect 13522 4378 13578 4380
rect 13282 4326 13308 4378
rect 13308 4326 13338 4378
rect 13362 4326 13372 4378
rect 13372 4326 13418 4378
rect 13442 4326 13488 4378
rect 13488 4326 13498 4378
rect 13522 4326 13552 4378
rect 13552 4326 13578 4378
rect 13282 4324 13338 4326
rect 13362 4324 13418 4326
rect 13442 4324 13498 4326
rect 13522 4324 13578 4326
rect 13266 3576 13322 3632
rect 13282 3290 13338 3292
rect 13362 3290 13418 3292
rect 13442 3290 13498 3292
rect 13522 3290 13578 3292
rect 13282 3238 13308 3290
rect 13308 3238 13338 3290
rect 13362 3238 13372 3290
rect 13372 3238 13418 3290
rect 13442 3238 13488 3290
rect 13488 3238 13498 3290
rect 13522 3238 13552 3290
rect 13552 3238 13578 3290
rect 13282 3236 13338 3238
rect 13362 3236 13418 3238
rect 13442 3236 13498 3238
rect 13522 3236 13578 3238
rect 13910 3032 13966 3088
rect 13282 2202 13338 2204
rect 13362 2202 13418 2204
rect 13442 2202 13498 2204
rect 13522 2202 13578 2204
rect 13282 2150 13308 2202
rect 13308 2150 13338 2202
rect 13362 2150 13372 2202
rect 13372 2150 13418 2202
rect 13442 2150 13488 2202
rect 13488 2150 13498 2202
rect 13522 2150 13552 2202
rect 13552 2150 13578 2202
rect 13282 2148 13338 2150
rect 13362 2148 13418 2150
rect 13442 2148 13498 2150
rect 13522 2148 13578 2150
rect 15106 17856 15162 17912
rect 14462 2896 14518 2952
rect 14738 5888 14794 5944
rect 15290 11736 15346 11792
rect 15014 9832 15070 9888
rect 14830 1944 14886 2000
rect 4158 448 4214 504
<< metal3 >>
rect 0 19546 800 19576
rect 2865 19546 2931 19549
rect 0 19544 2931 19546
rect 0 19488 2870 19544
rect 2926 19488 2931 19544
rect 0 19486 2931 19488
rect 0 19456 800 19486
rect 2865 19483 2931 19486
rect 0 18594 800 18624
rect 4061 18594 4127 18597
rect 0 18592 4127 18594
rect 0 18536 4066 18592
rect 4122 18536 4127 18592
rect 0 18534 4127 18536
rect 0 18504 800 18534
rect 4061 18531 4127 18534
rect 15101 17914 15167 17917
rect 16200 17914 17000 17944
rect 15101 17912 17000 17914
rect 15101 17856 15106 17912
rect 15162 17856 17000 17912
rect 15101 17854 17000 17856
rect 15101 17851 15167 17854
rect 16200 17824 17000 17854
rect 0 17642 800 17672
rect 3141 17642 3207 17645
rect 0 17640 3207 17642
rect 0 17584 3146 17640
rect 3202 17584 3207 17640
rect 0 17582 3207 17584
rect 0 17552 800 17582
rect 3141 17579 3207 17582
rect 3409 17440 3729 17441
rect 3409 17376 3417 17440
rect 3481 17376 3497 17440
rect 3561 17376 3577 17440
rect 3641 17376 3657 17440
rect 3721 17376 3729 17440
rect 3409 17375 3729 17376
rect 8340 17440 8660 17441
rect 8340 17376 8348 17440
rect 8412 17376 8428 17440
rect 8492 17376 8508 17440
rect 8572 17376 8588 17440
rect 8652 17376 8660 17440
rect 8340 17375 8660 17376
rect 13270 17440 13590 17441
rect 13270 17376 13278 17440
rect 13342 17376 13358 17440
rect 13422 17376 13438 17440
rect 13502 17376 13518 17440
rect 13582 17376 13590 17440
rect 13270 17375 13590 17376
rect 5874 16896 6194 16897
rect 5874 16832 5882 16896
rect 5946 16832 5962 16896
rect 6026 16832 6042 16896
rect 6106 16832 6122 16896
rect 6186 16832 6194 16896
rect 5874 16831 6194 16832
rect 10805 16896 11125 16897
rect 10805 16832 10813 16896
rect 10877 16832 10893 16896
rect 10957 16832 10973 16896
rect 11037 16832 11053 16896
rect 11117 16832 11125 16896
rect 10805 16831 11125 16832
rect 11421 16826 11487 16829
rect 11286 16824 11487 16826
rect 11286 16768 11426 16824
rect 11482 16768 11487 16824
rect 11286 16766 11487 16768
rect 0 16690 800 16720
rect 1761 16690 1827 16693
rect 0 16688 1827 16690
rect 0 16632 1766 16688
rect 1822 16632 1827 16688
rect 0 16630 1827 16632
rect 0 16600 800 16630
rect 1761 16627 1827 16630
rect 11145 16690 11211 16693
rect 11286 16690 11346 16766
rect 11421 16763 11487 16766
rect 11145 16688 11346 16690
rect 11145 16632 11150 16688
rect 11206 16632 11346 16688
rect 11145 16630 11346 16632
rect 11145 16627 11211 16630
rect 1669 16554 1735 16557
rect 9121 16554 9187 16557
rect 9857 16554 9923 16557
rect 1669 16552 9923 16554
rect 1669 16496 1674 16552
rect 1730 16496 9126 16552
rect 9182 16496 9862 16552
rect 9918 16496 9923 16552
rect 1669 16494 9923 16496
rect 1669 16491 1735 16494
rect 9121 16491 9187 16494
rect 9857 16491 9923 16494
rect 3409 16352 3729 16353
rect 3409 16288 3417 16352
rect 3481 16288 3497 16352
rect 3561 16288 3577 16352
rect 3641 16288 3657 16352
rect 3721 16288 3729 16352
rect 3409 16287 3729 16288
rect 8340 16352 8660 16353
rect 8340 16288 8348 16352
rect 8412 16288 8428 16352
rect 8492 16288 8508 16352
rect 8572 16288 8588 16352
rect 8652 16288 8660 16352
rect 8340 16287 8660 16288
rect 13270 16352 13590 16353
rect 13270 16288 13278 16352
rect 13342 16288 13358 16352
rect 13422 16288 13438 16352
rect 13502 16288 13518 16352
rect 13582 16288 13590 16352
rect 13270 16287 13590 16288
rect 2313 16146 2379 16149
rect 9438 16146 9444 16148
rect 2313 16144 9444 16146
rect 2313 16088 2318 16144
rect 2374 16088 9444 16144
rect 2313 16086 9444 16088
rect 2313 16083 2379 16086
rect 9438 16084 9444 16086
rect 9508 16146 9514 16148
rect 9581 16146 9647 16149
rect 9508 16144 9647 16146
rect 9508 16088 9586 16144
rect 9642 16088 9647 16144
rect 9508 16086 9647 16088
rect 9508 16084 9514 16086
rect 9581 16083 9647 16086
rect 5874 15808 6194 15809
rect 0 15738 800 15768
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6194 15808
rect 5874 15743 6194 15744
rect 10805 15808 11125 15809
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 15743 11125 15744
rect 1761 15738 1827 15741
rect 0 15736 1827 15738
rect 0 15680 1766 15736
rect 1822 15680 1827 15736
rect 0 15678 1827 15680
rect 0 15648 800 15678
rect 1761 15675 1827 15678
rect 5257 15466 5323 15469
rect 9397 15466 9463 15469
rect 9949 15466 10015 15469
rect 10409 15466 10475 15469
rect 5257 15464 10475 15466
rect 5257 15408 5262 15464
rect 5318 15408 9402 15464
rect 9458 15408 9954 15464
rect 10010 15408 10414 15464
rect 10470 15408 10475 15464
rect 5257 15406 10475 15408
rect 5257 15403 5323 15406
rect 9397 15403 9463 15406
rect 9949 15403 10015 15406
rect 10409 15403 10475 15406
rect 3409 15264 3729 15265
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 15199 3729 15200
rect 8340 15264 8660 15265
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 15199 8660 15200
rect 13270 15264 13590 15265
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 15199 13590 15200
rect 7741 15058 7807 15061
rect 10225 15058 10291 15061
rect 7741 15056 10291 15058
rect 7741 15000 7746 15056
rect 7802 15000 10230 15056
rect 10286 15000 10291 15056
rect 7741 14998 10291 15000
rect 7741 14995 7807 14998
rect 10225 14995 10291 14998
rect 4797 14922 4863 14925
rect 8753 14922 8819 14925
rect 4797 14920 8819 14922
rect 4797 14864 4802 14920
rect 4858 14864 8758 14920
rect 8814 14864 8819 14920
rect 4797 14862 8819 14864
rect 4797 14859 4863 14862
rect 8753 14859 8819 14862
rect 0 14786 800 14816
rect 3417 14786 3483 14789
rect 0 14784 3483 14786
rect 0 14728 3422 14784
rect 3478 14728 3483 14784
rect 0 14726 3483 14728
rect 0 14696 800 14726
rect 3417 14723 3483 14726
rect 5874 14720 6194 14721
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6194 14720
rect 5874 14655 6194 14656
rect 10805 14720 11125 14721
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 14655 11125 14656
rect 2589 14514 2655 14517
rect 6269 14514 6335 14517
rect 2589 14512 6335 14514
rect 2589 14456 2594 14512
rect 2650 14456 6274 14512
rect 6330 14456 6335 14512
rect 2589 14454 6335 14456
rect 2589 14451 2655 14454
rect 6269 14451 6335 14454
rect 7189 14514 7255 14517
rect 8845 14514 8911 14517
rect 13261 14514 13327 14517
rect 7189 14512 13327 14514
rect 7189 14456 7194 14512
rect 7250 14456 8850 14512
rect 8906 14456 13266 14512
rect 13322 14456 13327 14512
rect 7189 14454 13327 14456
rect 7189 14451 7255 14454
rect 8845 14451 8911 14454
rect 13261 14451 13327 14454
rect 4061 14378 4127 14381
rect 10961 14378 11027 14381
rect 4061 14376 11027 14378
rect 4061 14320 4066 14376
rect 4122 14320 10966 14376
rect 11022 14320 11027 14376
rect 4061 14318 11027 14320
rect 4061 14315 4127 14318
rect 10961 14315 11027 14318
rect 3409 14176 3729 14177
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 14111 3729 14112
rect 8340 14176 8660 14177
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 14111 8660 14112
rect 13270 14176 13590 14177
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 14111 13590 14112
rect 13721 13970 13787 13973
rect 16200 13970 17000 14000
rect 13721 13968 17000 13970
rect 13721 13912 13726 13968
rect 13782 13912 17000 13968
rect 13721 13910 17000 13912
rect 13721 13907 13787 13910
rect 16200 13880 17000 13910
rect 0 13834 800 13864
rect 2957 13834 3023 13837
rect 0 13832 3023 13834
rect 0 13776 2962 13832
rect 3018 13776 3023 13832
rect 0 13774 3023 13776
rect 0 13744 800 13774
rect 2957 13771 3023 13774
rect 5874 13632 6194 13633
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6194 13632
rect 5874 13567 6194 13568
rect 10805 13632 11125 13633
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 13567 11125 13568
rect 3409 13088 3729 13089
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 13023 3729 13024
rect 8340 13088 8660 13089
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 13023 8660 13024
rect 13270 13088 13590 13089
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 13023 13590 13024
rect 0 12882 800 12912
rect 1577 12882 1643 12885
rect 0 12880 1643 12882
rect 0 12824 1582 12880
rect 1638 12824 1643 12880
rect 0 12822 1643 12824
rect 0 12792 800 12822
rect 1577 12819 1643 12822
rect 5625 12882 5691 12885
rect 5625 12880 6378 12882
rect 5625 12824 5630 12880
rect 5686 12824 6378 12880
rect 5625 12822 6378 12824
rect 5625 12819 5691 12822
rect 6318 12746 6378 12822
rect 6913 12746 6979 12749
rect 6318 12744 6979 12746
rect 6318 12688 6918 12744
rect 6974 12688 6979 12744
rect 6318 12686 6979 12688
rect 6913 12683 6979 12686
rect 9121 12746 9187 12749
rect 9438 12746 9444 12748
rect 9121 12744 9444 12746
rect 9121 12688 9126 12744
rect 9182 12688 9444 12744
rect 9121 12686 9444 12688
rect 9121 12683 9187 12686
rect 9438 12684 9444 12686
rect 9508 12746 9514 12748
rect 11145 12746 11211 12749
rect 9508 12744 11211 12746
rect 9508 12688 11150 12744
rect 11206 12688 11211 12744
rect 9508 12686 11211 12688
rect 9508 12684 9514 12686
rect 11145 12683 11211 12686
rect 6361 12610 6427 12613
rect 9213 12610 9279 12613
rect 9857 12610 9923 12613
rect 6361 12608 9923 12610
rect 6361 12552 6366 12608
rect 6422 12552 9218 12608
rect 9274 12552 9862 12608
rect 9918 12552 9923 12608
rect 6361 12550 9923 12552
rect 6361 12547 6427 12550
rect 9213 12547 9279 12550
rect 9857 12547 9923 12550
rect 5874 12544 6194 12545
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6194 12544
rect 5874 12479 6194 12480
rect 10805 12544 11125 12545
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10805 12479 11125 12480
rect 8017 12338 8083 12341
rect 10501 12338 10567 12341
rect 10869 12338 10935 12341
rect 8017 12336 10935 12338
rect 8017 12280 8022 12336
rect 8078 12280 10506 12336
rect 10562 12280 10874 12336
rect 10930 12280 10935 12336
rect 8017 12278 10935 12280
rect 8017 12275 8083 12278
rect 10501 12275 10567 12278
rect 10869 12275 10935 12278
rect 3409 12000 3729 12001
rect 0 11930 800 11960
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 11935 3729 11936
rect 8340 12000 8660 12001
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 11935 8660 11936
rect 13270 12000 13590 12001
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 11935 13590 11936
rect 3233 11930 3299 11933
rect 0 11928 3299 11930
rect 0 11872 3238 11928
rect 3294 11872 3299 11928
rect 0 11870 3299 11872
rect 0 11840 800 11870
rect 3233 11867 3299 11870
rect 8661 11794 8727 11797
rect 15285 11794 15351 11797
rect 8661 11792 15351 11794
rect 8661 11736 8666 11792
rect 8722 11736 15290 11792
rect 15346 11736 15351 11792
rect 8661 11734 15351 11736
rect 8661 11731 8727 11734
rect 15285 11731 15351 11734
rect 9397 11660 9463 11661
rect 9397 11658 9444 11660
rect 9316 11656 9444 11658
rect 9508 11658 9514 11660
rect 11053 11658 11119 11661
rect 9508 11656 11119 11658
rect 9316 11600 9402 11656
rect 9508 11600 11058 11656
rect 11114 11600 11119 11656
rect 9316 11598 9444 11600
rect 9397 11596 9444 11598
rect 9508 11598 11119 11600
rect 9508 11596 9514 11598
rect 9397 11595 9463 11596
rect 11053 11595 11119 11598
rect 5874 11456 6194 11457
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6194 11456
rect 5874 11391 6194 11392
rect 10805 11456 11125 11457
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 11391 11125 11392
rect 3325 11114 3391 11117
rect 9489 11114 9555 11117
rect 10869 11114 10935 11117
rect 3325 11112 10935 11114
rect 3325 11056 3330 11112
rect 3386 11056 9494 11112
rect 9550 11056 10874 11112
rect 10930 11056 10935 11112
rect 3325 11054 10935 11056
rect 3325 11051 3391 11054
rect 9489 11051 9555 11054
rect 10869 11051 10935 11054
rect 0 10978 800 11008
rect 3233 10978 3299 10981
rect 0 10976 3299 10978
rect 0 10920 3238 10976
rect 3294 10920 3299 10976
rect 0 10918 3299 10920
rect 0 10888 800 10918
rect 3233 10915 3299 10918
rect 3409 10912 3729 10913
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 10847 3729 10848
rect 8340 10912 8660 10913
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 10847 8660 10848
rect 13270 10912 13590 10913
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 10847 13590 10848
rect 5874 10368 6194 10369
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6194 10368
rect 5874 10303 6194 10304
rect 10805 10368 11125 10369
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10805 10303 11125 10304
rect 9397 10300 9463 10301
rect 9397 10298 9444 10300
rect 9352 10296 9444 10298
rect 9352 10240 9402 10296
rect 9352 10238 9444 10240
rect 9397 10236 9444 10238
rect 9508 10236 9514 10300
rect 9397 10235 9463 10236
rect 2313 10162 2379 10165
rect 5257 10162 5323 10165
rect 2313 10160 5323 10162
rect 2313 10104 2318 10160
rect 2374 10104 5262 10160
rect 5318 10104 5323 10160
rect 2313 10102 5323 10104
rect 2313 10099 2379 10102
rect 5257 10099 5323 10102
rect 8017 10162 8083 10165
rect 11237 10162 11303 10165
rect 8017 10160 11303 10162
rect 8017 10104 8022 10160
rect 8078 10104 11242 10160
rect 11298 10104 11303 10160
rect 8017 10102 11303 10104
rect 8017 10099 8083 10102
rect 11237 10099 11303 10102
rect 0 10026 800 10056
rect 2865 10026 2931 10029
rect 0 10024 2931 10026
rect 0 9968 2870 10024
rect 2926 9968 2931 10024
rect 0 9966 2931 9968
rect 0 9936 800 9966
rect 2865 9963 2931 9966
rect 9397 10026 9463 10029
rect 11513 10026 11579 10029
rect 9397 10024 11579 10026
rect 9397 9968 9402 10024
rect 9458 9968 11518 10024
rect 11574 9968 11579 10024
rect 9397 9966 11579 9968
rect 9397 9963 9463 9966
rect 11513 9963 11579 9966
rect 15009 9890 15075 9893
rect 16200 9890 17000 9920
rect 15009 9888 17000 9890
rect 15009 9832 15014 9888
rect 15070 9832 17000 9888
rect 15009 9830 17000 9832
rect 15009 9827 15075 9830
rect 3409 9824 3729 9825
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 9759 3729 9760
rect 8340 9824 8660 9825
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 9759 8660 9760
rect 13270 9824 13590 9825
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 16200 9800 17000 9830
rect 13270 9759 13590 9760
rect 9857 9754 9923 9757
rect 10685 9754 10751 9757
rect 9857 9752 10751 9754
rect 9857 9696 9862 9752
rect 9918 9696 10690 9752
rect 10746 9696 10751 9752
rect 9857 9694 10751 9696
rect 9857 9691 9923 9694
rect 10685 9691 10751 9694
rect 9806 9556 9812 9620
rect 9876 9618 9882 9620
rect 11145 9618 11211 9621
rect 14089 9618 14155 9621
rect 9876 9616 14155 9618
rect 9876 9560 11150 9616
rect 11206 9560 14094 9616
rect 14150 9560 14155 9616
rect 9876 9558 14155 9560
rect 9876 9556 9882 9558
rect 11145 9555 11211 9558
rect 14089 9555 14155 9558
rect 5874 9280 6194 9281
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6194 9280
rect 5874 9215 6194 9216
rect 10805 9280 11125 9281
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 9215 11125 9216
rect 0 9074 800 9104
rect 1669 9074 1735 9077
rect 0 9072 1735 9074
rect 0 9016 1674 9072
rect 1730 9016 1735 9072
rect 0 9014 1735 9016
rect 0 8984 800 9014
rect 1669 9011 1735 9014
rect 9857 9074 9923 9077
rect 10501 9074 10567 9077
rect 9857 9072 10567 9074
rect 9857 9016 9862 9072
rect 9918 9016 10506 9072
rect 10562 9016 10567 9072
rect 9857 9014 10567 9016
rect 9857 9011 9923 9014
rect 10501 9011 10567 9014
rect 12985 8938 13051 8941
rect 13721 8938 13787 8941
rect 12985 8936 13787 8938
rect 12985 8880 12990 8936
rect 13046 8880 13726 8936
rect 13782 8880 13787 8936
rect 12985 8878 13787 8880
rect 12985 8875 13051 8878
rect 13721 8875 13787 8878
rect 3409 8736 3729 8737
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 8671 3729 8672
rect 8340 8736 8660 8737
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 8671 8660 8672
rect 13270 8736 13590 8737
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 8671 13590 8672
rect 7557 8530 7623 8533
rect 12801 8530 12867 8533
rect 7557 8528 12867 8530
rect 7557 8472 7562 8528
rect 7618 8472 12806 8528
rect 12862 8472 12867 8528
rect 7557 8470 12867 8472
rect 7557 8467 7623 8470
rect 12801 8467 12867 8470
rect 9581 8260 9647 8261
rect 9581 8258 9628 8260
rect 9536 8256 9628 8258
rect 9536 8200 9586 8256
rect 9536 8198 9628 8200
rect 9581 8196 9628 8198
rect 9692 8196 9698 8260
rect 9581 8195 9647 8196
rect 5874 8192 6194 8193
rect 0 8122 800 8152
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6194 8192
rect 5874 8127 6194 8128
rect 10805 8192 11125 8193
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 8127 11125 8128
rect 2497 8122 2563 8125
rect 0 8120 2563 8122
rect 0 8064 2502 8120
rect 2558 8064 2563 8120
rect 0 8062 2563 8064
rect 0 8032 800 8062
rect 2497 8059 2563 8062
rect 4337 8122 4403 8125
rect 4797 8122 4863 8125
rect 4337 8120 4863 8122
rect 4337 8064 4342 8120
rect 4398 8064 4802 8120
rect 4858 8064 4863 8120
rect 4337 8062 4863 8064
rect 4337 8059 4403 8062
rect 4797 8059 4863 8062
rect 8845 8122 8911 8125
rect 9806 8122 9812 8124
rect 8845 8120 9812 8122
rect 8845 8064 8850 8120
rect 8906 8064 9812 8120
rect 8845 8062 9812 8064
rect 8845 8059 8911 8062
rect 9806 8060 9812 8062
rect 9876 8060 9882 8124
rect 4061 7986 4127 7989
rect 11605 7986 11671 7989
rect 4061 7984 11671 7986
rect 4061 7928 4066 7984
rect 4122 7928 11610 7984
rect 11666 7928 11671 7984
rect 4061 7926 11671 7928
rect 4061 7923 4127 7926
rect 11605 7923 11671 7926
rect 8477 7850 8543 7853
rect 9581 7850 9647 7853
rect 8477 7848 9647 7850
rect 8477 7792 8482 7848
rect 8538 7792 9586 7848
rect 9642 7792 9647 7848
rect 8477 7790 9647 7792
rect 8477 7787 8543 7790
rect 9581 7787 9647 7790
rect 3409 7648 3729 7649
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 7583 3729 7584
rect 8340 7648 8660 7649
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 7583 8660 7584
rect 13270 7648 13590 7649
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 7583 13590 7584
rect 10133 7442 10199 7445
rect 10685 7442 10751 7445
rect 11329 7442 11395 7445
rect 10133 7440 11395 7442
rect 10133 7384 10138 7440
rect 10194 7384 10690 7440
rect 10746 7384 11334 7440
rect 11390 7384 11395 7440
rect 10133 7382 11395 7384
rect 10133 7379 10199 7382
rect 10685 7379 10751 7382
rect 11329 7379 11395 7382
rect 0 7170 800 7200
rect 1669 7170 1735 7173
rect 0 7168 1735 7170
rect 0 7112 1674 7168
rect 1730 7112 1735 7168
rect 0 7110 1735 7112
rect 0 7080 800 7110
rect 1669 7107 1735 7110
rect 5874 7104 6194 7105
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6194 7104
rect 5874 7039 6194 7040
rect 10805 7104 11125 7105
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 7039 11125 7040
rect 4797 6762 4863 6765
rect 6729 6762 6795 6765
rect 4797 6760 6930 6762
rect 4797 6704 4802 6760
rect 4858 6704 6734 6760
rect 6790 6704 6930 6760
rect 4797 6702 6930 6704
rect 4797 6699 4863 6702
rect 6729 6699 6795 6702
rect 3409 6560 3729 6561
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 6495 3729 6496
rect 6870 6354 6930 6702
rect 8340 6560 8660 6561
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 6495 8660 6496
rect 13270 6560 13590 6561
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 6495 13590 6496
rect 10133 6354 10199 6357
rect 6870 6352 10199 6354
rect 6870 6296 10138 6352
rect 10194 6296 10199 6352
rect 6870 6294 10199 6296
rect 10133 6291 10199 6294
rect 0 6218 800 6248
rect 1669 6218 1735 6221
rect 0 6216 1735 6218
rect 0 6160 1674 6216
rect 1730 6160 1735 6216
rect 0 6158 1735 6160
rect 0 6128 800 6158
rect 1669 6155 1735 6158
rect 6177 6218 6243 6221
rect 6637 6218 6703 6221
rect 8385 6218 8451 6221
rect 6177 6216 8451 6218
rect 6177 6160 6182 6216
rect 6238 6160 6642 6216
rect 6698 6160 8390 6216
rect 8446 6160 8451 6216
rect 6177 6158 8451 6160
rect 6177 6155 6243 6158
rect 6637 6155 6703 6158
rect 8385 6155 8451 6158
rect 5874 6016 6194 6017
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6194 6016
rect 5874 5951 6194 5952
rect 10805 6016 11125 6017
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 5951 11125 5952
rect 14733 5946 14799 5949
rect 16200 5946 17000 5976
rect 14733 5944 17000 5946
rect 14733 5888 14738 5944
rect 14794 5888 17000 5944
rect 14733 5886 17000 5888
rect 14733 5883 14799 5886
rect 16200 5856 17000 5886
rect 7281 5810 7347 5813
rect 10593 5810 10659 5813
rect 10777 5810 10843 5813
rect 7281 5808 10843 5810
rect 7281 5752 7286 5808
rect 7342 5752 10598 5808
rect 10654 5752 10782 5808
rect 10838 5752 10843 5808
rect 7281 5750 10843 5752
rect 7281 5747 7347 5750
rect 10593 5747 10659 5750
rect 10777 5747 10843 5750
rect 2589 5674 2655 5677
rect 6913 5674 6979 5677
rect 2589 5672 6979 5674
rect 2589 5616 2594 5672
rect 2650 5616 6918 5672
rect 6974 5616 6979 5672
rect 2589 5614 6979 5616
rect 2589 5611 2655 5614
rect 6913 5611 6979 5614
rect 7925 5674 7991 5677
rect 10409 5674 10475 5677
rect 7925 5672 10475 5674
rect 7925 5616 7930 5672
rect 7986 5616 10414 5672
rect 10470 5616 10475 5672
rect 7925 5614 10475 5616
rect 7925 5611 7991 5614
rect 10409 5611 10475 5614
rect 3409 5472 3729 5473
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 5407 3729 5408
rect 8340 5472 8660 5473
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 5407 8660 5408
rect 13270 5472 13590 5473
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 5407 13590 5408
rect 0 5266 800 5296
rect 2773 5266 2839 5269
rect 0 5264 2839 5266
rect 0 5208 2778 5264
rect 2834 5208 2839 5264
rect 0 5206 2839 5208
rect 0 5176 800 5206
rect 2773 5203 2839 5206
rect 5874 4928 6194 4929
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6194 4928
rect 5874 4863 6194 4864
rect 10805 4928 11125 4929
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 4863 11125 4864
rect 3409 4384 3729 4385
rect 0 4314 800 4344
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 4319 3729 4320
rect 8340 4384 8660 4385
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 4319 8660 4320
rect 13270 4384 13590 4385
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 4319 13590 4320
rect 1669 4314 1735 4317
rect 0 4312 1735 4314
rect 0 4256 1674 4312
rect 1730 4256 1735 4312
rect 0 4254 1735 4256
rect 0 4224 800 4254
rect 1669 4251 1735 4254
rect 4889 4042 4955 4045
rect 5349 4042 5415 4045
rect 10777 4042 10843 4045
rect 4889 4040 10843 4042
rect 4889 3984 4894 4040
rect 4950 3984 5354 4040
rect 5410 3984 10782 4040
rect 10838 3984 10843 4040
rect 4889 3982 10843 3984
rect 4889 3979 4955 3982
rect 5349 3979 5415 3982
rect 10777 3979 10843 3982
rect 5874 3840 6194 3841
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6194 3840
rect 5874 3775 6194 3776
rect 10805 3840 11125 3841
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 3775 11125 3776
rect 6637 3770 6703 3773
rect 9765 3770 9831 3773
rect 6637 3768 9831 3770
rect 6637 3712 6642 3768
rect 6698 3712 9770 3768
rect 9826 3712 9831 3768
rect 6637 3710 9831 3712
rect 6637 3707 6703 3710
rect 9765 3707 9831 3710
rect 4429 3634 4495 3637
rect 6361 3634 6427 3637
rect 4429 3632 6427 3634
rect 4429 3576 4434 3632
rect 4490 3576 6366 3632
rect 6422 3576 6427 3632
rect 4429 3574 6427 3576
rect 4429 3571 4495 3574
rect 6361 3571 6427 3574
rect 11605 3634 11671 3637
rect 13261 3634 13327 3637
rect 11605 3632 13327 3634
rect 11605 3576 11610 3632
rect 11666 3576 13266 3632
rect 13322 3576 13327 3632
rect 11605 3574 13327 3576
rect 11605 3571 11671 3574
rect 13261 3571 13327 3574
rect 0 3362 800 3392
rect 1669 3362 1735 3365
rect 0 3360 1735 3362
rect 0 3304 1674 3360
rect 1730 3304 1735 3360
rect 0 3302 1735 3304
rect 0 3272 800 3302
rect 1669 3299 1735 3302
rect 3409 3296 3729 3297
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 3231 3729 3232
rect 8340 3296 8660 3297
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 3231 8660 3232
rect 13270 3296 13590 3297
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13270 3231 13590 3232
rect 10225 3226 10291 3229
rect 11421 3226 11487 3229
rect 10225 3224 11487 3226
rect 10225 3168 10230 3224
rect 10286 3168 11426 3224
rect 11482 3168 11487 3224
rect 10225 3166 11487 3168
rect 10225 3163 10291 3166
rect 11421 3163 11487 3166
rect 4797 3090 4863 3093
rect 13905 3090 13971 3093
rect 4797 3088 13971 3090
rect 4797 3032 4802 3088
rect 4858 3032 13910 3088
rect 13966 3032 13971 3088
rect 4797 3030 13971 3032
rect 4797 3027 4863 3030
rect 13905 3027 13971 3030
rect 4705 2954 4771 2957
rect 14457 2954 14523 2957
rect 4705 2952 14523 2954
rect 4705 2896 4710 2952
rect 4766 2896 14462 2952
rect 14518 2896 14523 2952
rect 4705 2894 14523 2896
rect 4705 2891 4771 2894
rect 14457 2891 14523 2894
rect 7925 2818 7991 2821
rect 8845 2818 8911 2821
rect 10317 2818 10383 2821
rect 7925 2816 10383 2818
rect 7925 2760 7930 2816
rect 7986 2760 8850 2816
rect 8906 2760 10322 2816
rect 10378 2760 10383 2816
rect 7925 2758 10383 2760
rect 7925 2755 7991 2758
rect 8845 2755 8911 2758
rect 10317 2755 10383 2758
rect 5874 2752 6194 2753
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6194 2752
rect 5874 2687 6194 2688
rect 10805 2752 11125 2753
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2687 11125 2688
rect 9489 2682 9555 2685
rect 9622 2682 9628 2684
rect 9489 2680 9628 2682
rect 9489 2624 9494 2680
rect 9550 2624 9628 2680
rect 9489 2622 9628 2624
rect 9489 2619 9555 2622
rect 9622 2620 9628 2622
rect 9692 2620 9698 2684
rect 0 2410 800 2440
rect 4061 2410 4127 2413
rect 0 2408 4127 2410
rect 0 2352 4066 2408
rect 4122 2352 4127 2408
rect 0 2350 4127 2352
rect 0 2320 800 2350
rect 4061 2347 4127 2350
rect 3409 2208 3729 2209
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2143 3729 2144
rect 8340 2208 8660 2209
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2143 8660 2144
rect 13270 2208 13590 2209
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2143 13590 2144
rect 14825 2002 14891 2005
rect 16200 2002 17000 2032
rect 14825 2000 17000 2002
rect 14825 1944 14830 2000
rect 14886 1944 17000 2000
rect 14825 1942 17000 1944
rect 14825 1939 14891 1942
rect 16200 1912 17000 1942
rect 0 1458 800 1488
rect 2773 1458 2839 1461
rect 0 1456 2839 1458
rect 0 1400 2778 1456
rect 2834 1400 2839 1456
rect 0 1398 2839 1400
rect 0 1368 800 1398
rect 2773 1395 2839 1398
rect 5533 914 5599 917
rect 7005 914 7071 917
rect 5533 912 7071 914
rect 5533 856 5538 912
rect 5594 856 7010 912
rect 7066 856 7071 912
rect 5533 854 7071 856
rect 5533 851 5599 854
rect 7005 851 7071 854
rect 0 506 800 536
rect 4153 506 4219 509
rect 0 504 4219 506
rect 0 448 4158 504
rect 4214 448 4219 504
rect 0 446 4219 448
rect 0 416 800 446
rect 4153 443 4219 446
<< via3 >>
rect 3417 17436 3481 17440
rect 3417 17380 3421 17436
rect 3421 17380 3477 17436
rect 3477 17380 3481 17436
rect 3417 17376 3481 17380
rect 3497 17436 3561 17440
rect 3497 17380 3501 17436
rect 3501 17380 3557 17436
rect 3557 17380 3561 17436
rect 3497 17376 3561 17380
rect 3577 17436 3641 17440
rect 3577 17380 3581 17436
rect 3581 17380 3637 17436
rect 3637 17380 3641 17436
rect 3577 17376 3641 17380
rect 3657 17436 3721 17440
rect 3657 17380 3661 17436
rect 3661 17380 3717 17436
rect 3717 17380 3721 17436
rect 3657 17376 3721 17380
rect 8348 17436 8412 17440
rect 8348 17380 8352 17436
rect 8352 17380 8408 17436
rect 8408 17380 8412 17436
rect 8348 17376 8412 17380
rect 8428 17436 8492 17440
rect 8428 17380 8432 17436
rect 8432 17380 8488 17436
rect 8488 17380 8492 17436
rect 8428 17376 8492 17380
rect 8508 17436 8572 17440
rect 8508 17380 8512 17436
rect 8512 17380 8568 17436
rect 8568 17380 8572 17436
rect 8508 17376 8572 17380
rect 8588 17436 8652 17440
rect 8588 17380 8592 17436
rect 8592 17380 8648 17436
rect 8648 17380 8652 17436
rect 8588 17376 8652 17380
rect 13278 17436 13342 17440
rect 13278 17380 13282 17436
rect 13282 17380 13338 17436
rect 13338 17380 13342 17436
rect 13278 17376 13342 17380
rect 13358 17436 13422 17440
rect 13358 17380 13362 17436
rect 13362 17380 13418 17436
rect 13418 17380 13422 17436
rect 13358 17376 13422 17380
rect 13438 17436 13502 17440
rect 13438 17380 13442 17436
rect 13442 17380 13498 17436
rect 13498 17380 13502 17436
rect 13438 17376 13502 17380
rect 13518 17436 13582 17440
rect 13518 17380 13522 17436
rect 13522 17380 13578 17436
rect 13578 17380 13582 17436
rect 13518 17376 13582 17380
rect 5882 16892 5946 16896
rect 5882 16836 5886 16892
rect 5886 16836 5942 16892
rect 5942 16836 5946 16892
rect 5882 16832 5946 16836
rect 5962 16892 6026 16896
rect 5962 16836 5966 16892
rect 5966 16836 6022 16892
rect 6022 16836 6026 16892
rect 5962 16832 6026 16836
rect 6042 16892 6106 16896
rect 6042 16836 6046 16892
rect 6046 16836 6102 16892
rect 6102 16836 6106 16892
rect 6042 16832 6106 16836
rect 6122 16892 6186 16896
rect 6122 16836 6126 16892
rect 6126 16836 6182 16892
rect 6182 16836 6186 16892
rect 6122 16832 6186 16836
rect 10813 16892 10877 16896
rect 10813 16836 10817 16892
rect 10817 16836 10873 16892
rect 10873 16836 10877 16892
rect 10813 16832 10877 16836
rect 10893 16892 10957 16896
rect 10893 16836 10897 16892
rect 10897 16836 10953 16892
rect 10953 16836 10957 16892
rect 10893 16832 10957 16836
rect 10973 16892 11037 16896
rect 10973 16836 10977 16892
rect 10977 16836 11033 16892
rect 11033 16836 11037 16892
rect 10973 16832 11037 16836
rect 11053 16892 11117 16896
rect 11053 16836 11057 16892
rect 11057 16836 11113 16892
rect 11113 16836 11117 16892
rect 11053 16832 11117 16836
rect 3417 16348 3481 16352
rect 3417 16292 3421 16348
rect 3421 16292 3477 16348
rect 3477 16292 3481 16348
rect 3417 16288 3481 16292
rect 3497 16348 3561 16352
rect 3497 16292 3501 16348
rect 3501 16292 3557 16348
rect 3557 16292 3561 16348
rect 3497 16288 3561 16292
rect 3577 16348 3641 16352
rect 3577 16292 3581 16348
rect 3581 16292 3637 16348
rect 3637 16292 3641 16348
rect 3577 16288 3641 16292
rect 3657 16348 3721 16352
rect 3657 16292 3661 16348
rect 3661 16292 3717 16348
rect 3717 16292 3721 16348
rect 3657 16288 3721 16292
rect 8348 16348 8412 16352
rect 8348 16292 8352 16348
rect 8352 16292 8408 16348
rect 8408 16292 8412 16348
rect 8348 16288 8412 16292
rect 8428 16348 8492 16352
rect 8428 16292 8432 16348
rect 8432 16292 8488 16348
rect 8488 16292 8492 16348
rect 8428 16288 8492 16292
rect 8508 16348 8572 16352
rect 8508 16292 8512 16348
rect 8512 16292 8568 16348
rect 8568 16292 8572 16348
rect 8508 16288 8572 16292
rect 8588 16348 8652 16352
rect 8588 16292 8592 16348
rect 8592 16292 8648 16348
rect 8648 16292 8652 16348
rect 8588 16288 8652 16292
rect 13278 16348 13342 16352
rect 13278 16292 13282 16348
rect 13282 16292 13338 16348
rect 13338 16292 13342 16348
rect 13278 16288 13342 16292
rect 13358 16348 13422 16352
rect 13358 16292 13362 16348
rect 13362 16292 13418 16348
rect 13418 16292 13422 16348
rect 13358 16288 13422 16292
rect 13438 16348 13502 16352
rect 13438 16292 13442 16348
rect 13442 16292 13498 16348
rect 13498 16292 13502 16348
rect 13438 16288 13502 16292
rect 13518 16348 13582 16352
rect 13518 16292 13522 16348
rect 13522 16292 13578 16348
rect 13578 16292 13582 16348
rect 13518 16288 13582 16292
rect 9444 16084 9508 16148
rect 5882 15804 5946 15808
rect 5882 15748 5886 15804
rect 5886 15748 5942 15804
rect 5942 15748 5946 15804
rect 5882 15744 5946 15748
rect 5962 15804 6026 15808
rect 5962 15748 5966 15804
rect 5966 15748 6022 15804
rect 6022 15748 6026 15804
rect 5962 15744 6026 15748
rect 6042 15804 6106 15808
rect 6042 15748 6046 15804
rect 6046 15748 6102 15804
rect 6102 15748 6106 15804
rect 6042 15744 6106 15748
rect 6122 15804 6186 15808
rect 6122 15748 6126 15804
rect 6126 15748 6182 15804
rect 6182 15748 6186 15804
rect 6122 15744 6186 15748
rect 10813 15804 10877 15808
rect 10813 15748 10817 15804
rect 10817 15748 10873 15804
rect 10873 15748 10877 15804
rect 10813 15744 10877 15748
rect 10893 15804 10957 15808
rect 10893 15748 10897 15804
rect 10897 15748 10953 15804
rect 10953 15748 10957 15804
rect 10893 15744 10957 15748
rect 10973 15804 11037 15808
rect 10973 15748 10977 15804
rect 10977 15748 11033 15804
rect 11033 15748 11037 15804
rect 10973 15744 11037 15748
rect 11053 15804 11117 15808
rect 11053 15748 11057 15804
rect 11057 15748 11113 15804
rect 11113 15748 11117 15804
rect 11053 15744 11117 15748
rect 3417 15260 3481 15264
rect 3417 15204 3421 15260
rect 3421 15204 3477 15260
rect 3477 15204 3481 15260
rect 3417 15200 3481 15204
rect 3497 15260 3561 15264
rect 3497 15204 3501 15260
rect 3501 15204 3557 15260
rect 3557 15204 3561 15260
rect 3497 15200 3561 15204
rect 3577 15260 3641 15264
rect 3577 15204 3581 15260
rect 3581 15204 3637 15260
rect 3637 15204 3641 15260
rect 3577 15200 3641 15204
rect 3657 15260 3721 15264
rect 3657 15204 3661 15260
rect 3661 15204 3717 15260
rect 3717 15204 3721 15260
rect 3657 15200 3721 15204
rect 8348 15260 8412 15264
rect 8348 15204 8352 15260
rect 8352 15204 8408 15260
rect 8408 15204 8412 15260
rect 8348 15200 8412 15204
rect 8428 15260 8492 15264
rect 8428 15204 8432 15260
rect 8432 15204 8488 15260
rect 8488 15204 8492 15260
rect 8428 15200 8492 15204
rect 8508 15260 8572 15264
rect 8508 15204 8512 15260
rect 8512 15204 8568 15260
rect 8568 15204 8572 15260
rect 8508 15200 8572 15204
rect 8588 15260 8652 15264
rect 8588 15204 8592 15260
rect 8592 15204 8648 15260
rect 8648 15204 8652 15260
rect 8588 15200 8652 15204
rect 13278 15260 13342 15264
rect 13278 15204 13282 15260
rect 13282 15204 13338 15260
rect 13338 15204 13342 15260
rect 13278 15200 13342 15204
rect 13358 15260 13422 15264
rect 13358 15204 13362 15260
rect 13362 15204 13418 15260
rect 13418 15204 13422 15260
rect 13358 15200 13422 15204
rect 13438 15260 13502 15264
rect 13438 15204 13442 15260
rect 13442 15204 13498 15260
rect 13498 15204 13502 15260
rect 13438 15200 13502 15204
rect 13518 15260 13582 15264
rect 13518 15204 13522 15260
rect 13522 15204 13578 15260
rect 13578 15204 13582 15260
rect 13518 15200 13582 15204
rect 5882 14716 5946 14720
rect 5882 14660 5886 14716
rect 5886 14660 5942 14716
rect 5942 14660 5946 14716
rect 5882 14656 5946 14660
rect 5962 14716 6026 14720
rect 5962 14660 5966 14716
rect 5966 14660 6022 14716
rect 6022 14660 6026 14716
rect 5962 14656 6026 14660
rect 6042 14716 6106 14720
rect 6042 14660 6046 14716
rect 6046 14660 6102 14716
rect 6102 14660 6106 14716
rect 6042 14656 6106 14660
rect 6122 14716 6186 14720
rect 6122 14660 6126 14716
rect 6126 14660 6182 14716
rect 6182 14660 6186 14716
rect 6122 14656 6186 14660
rect 10813 14716 10877 14720
rect 10813 14660 10817 14716
rect 10817 14660 10873 14716
rect 10873 14660 10877 14716
rect 10813 14656 10877 14660
rect 10893 14716 10957 14720
rect 10893 14660 10897 14716
rect 10897 14660 10953 14716
rect 10953 14660 10957 14716
rect 10893 14656 10957 14660
rect 10973 14716 11037 14720
rect 10973 14660 10977 14716
rect 10977 14660 11033 14716
rect 11033 14660 11037 14716
rect 10973 14656 11037 14660
rect 11053 14716 11117 14720
rect 11053 14660 11057 14716
rect 11057 14660 11113 14716
rect 11113 14660 11117 14716
rect 11053 14656 11117 14660
rect 3417 14172 3481 14176
rect 3417 14116 3421 14172
rect 3421 14116 3477 14172
rect 3477 14116 3481 14172
rect 3417 14112 3481 14116
rect 3497 14172 3561 14176
rect 3497 14116 3501 14172
rect 3501 14116 3557 14172
rect 3557 14116 3561 14172
rect 3497 14112 3561 14116
rect 3577 14172 3641 14176
rect 3577 14116 3581 14172
rect 3581 14116 3637 14172
rect 3637 14116 3641 14172
rect 3577 14112 3641 14116
rect 3657 14172 3721 14176
rect 3657 14116 3661 14172
rect 3661 14116 3717 14172
rect 3717 14116 3721 14172
rect 3657 14112 3721 14116
rect 8348 14172 8412 14176
rect 8348 14116 8352 14172
rect 8352 14116 8408 14172
rect 8408 14116 8412 14172
rect 8348 14112 8412 14116
rect 8428 14172 8492 14176
rect 8428 14116 8432 14172
rect 8432 14116 8488 14172
rect 8488 14116 8492 14172
rect 8428 14112 8492 14116
rect 8508 14172 8572 14176
rect 8508 14116 8512 14172
rect 8512 14116 8568 14172
rect 8568 14116 8572 14172
rect 8508 14112 8572 14116
rect 8588 14172 8652 14176
rect 8588 14116 8592 14172
rect 8592 14116 8648 14172
rect 8648 14116 8652 14172
rect 8588 14112 8652 14116
rect 13278 14172 13342 14176
rect 13278 14116 13282 14172
rect 13282 14116 13338 14172
rect 13338 14116 13342 14172
rect 13278 14112 13342 14116
rect 13358 14172 13422 14176
rect 13358 14116 13362 14172
rect 13362 14116 13418 14172
rect 13418 14116 13422 14172
rect 13358 14112 13422 14116
rect 13438 14172 13502 14176
rect 13438 14116 13442 14172
rect 13442 14116 13498 14172
rect 13498 14116 13502 14172
rect 13438 14112 13502 14116
rect 13518 14172 13582 14176
rect 13518 14116 13522 14172
rect 13522 14116 13578 14172
rect 13578 14116 13582 14172
rect 13518 14112 13582 14116
rect 5882 13628 5946 13632
rect 5882 13572 5886 13628
rect 5886 13572 5942 13628
rect 5942 13572 5946 13628
rect 5882 13568 5946 13572
rect 5962 13628 6026 13632
rect 5962 13572 5966 13628
rect 5966 13572 6022 13628
rect 6022 13572 6026 13628
rect 5962 13568 6026 13572
rect 6042 13628 6106 13632
rect 6042 13572 6046 13628
rect 6046 13572 6102 13628
rect 6102 13572 6106 13628
rect 6042 13568 6106 13572
rect 6122 13628 6186 13632
rect 6122 13572 6126 13628
rect 6126 13572 6182 13628
rect 6182 13572 6186 13628
rect 6122 13568 6186 13572
rect 10813 13628 10877 13632
rect 10813 13572 10817 13628
rect 10817 13572 10873 13628
rect 10873 13572 10877 13628
rect 10813 13568 10877 13572
rect 10893 13628 10957 13632
rect 10893 13572 10897 13628
rect 10897 13572 10953 13628
rect 10953 13572 10957 13628
rect 10893 13568 10957 13572
rect 10973 13628 11037 13632
rect 10973 13572 10977 13628
rect 10977 13572 11033 13628
rect 11033 13572 11037 13628
rect 10973 13568 11037 13572
rect 11053 13628 11117 13632
rect 11053 13572 11057 13628
rect 11057 13572 11113 13628
rect 11113 13572 11117 13628
rect 11053 13568 11117 13572
rect 3417 13084 3481 13088
rect 3417 13028 3421 13084
rect 3421 13028 3477 13084
rect 3477 13028 3481 13084
rect 3417 13024 3481 13028
rect 3497 13084 3561 13088
rect 3497 13028 3501 13084
rect 3501 13028 3557 13084
rect 3557 13028 3561 13084
rect 3497 13024 3561 13028
rect 3577 13084 3641 13088
rect 3577 13028 3581 13084
rect 3581 13028 3637 13084
rect 3637 13028 3641 13084
rect 3577 13024 3641 13028
rect 3657 13084 3721 13088
rect 3657 13028 3661 13084
rect 3661 13028 3717 13084
rect 3717 13028 3721 13084
rect 3657 13024 3721 13028
rect 8348 13084 8412 13088
rect 8348 13028 8352 13084
rect 8352 13028 8408 13084
rect 8408 13028 8412 13084
rect 8348 13024 8412 13028
rect 8428 13084 8492 13088
rect 8428 13028 8432 13084
rect 8432 13028 8488 13084
rect 8488 13028 8492 13084
rect 8428 13024 8492 13028
rect 8508 13084 8572 13088
rect 8508 13028 8512 13084
rect 8512 13028 8568 13084
rect 8568 13028 8572 13084
rect 8508 13024 8572 13028
rect 8588 13084 8652 13088
rect 8588 13028 8592 13084
rect 8592 13028 8648 13084
rect 8648 13028 8652 13084
rect 8588 13024 8652 13028
rect 13278 13084 13342 13088
rect 13278 13028 13282 13084
rect 13282 13028 13338 13084
rect 13338 13028 13342 13084
rect 13278 13024 13342 13028
rect 13358 13084 13422 13088
rect 13358 13028 13362 13084
rect 13362 13028 13418 13084
rect 13418 13028 13422 13084
rect 13358 13024 13422 13028
rect 13438 13084 13502 13088
rect 13438 13028 13442 13084
rect 13442 13028 13498 13084
rect 13498 13028 13502 13084
rect 13438 13024 13502 13028
rect 13518 13084 13582 13088
rect 13518 13028 13522 13084
rect 13522 13028 13578 13084
rect 13578 13028 13582 13084
rect 13518 13024 13582 13028
rect 9444 12684 9508 12748
rect 5882 12540 5946 12544
rect 5882 12484 5886 12540
rect 5886 12484 5942 12540
rect 5942 12484 5946 12540
rect 5882 12480 5946 12484
rect 5962 12540 6026 12544
rect 5962 12484 5966 12540
rect 5966 12484 6022 12540
rect 6022 12484 6026 12540
rect 5962 12480 6026 12484
rect 6042 12540 6106 12544
rect 6042 12484 6046 12540
rect 6046 12484 6102 12540
rect 6102 12484 6106 12540
rect 6042 12480 6106 12484
rect 6122 12540 6186 12544
rect 6122 12484 6126 12540
rect 6126 12484 6182 12540
rect 6182 12484 6186 12540
rect 6122 12480 6186 12484
rect 10813 12540 10877 12544
rect 10813 12484 10817 12540
rect 10817 12484 10873 12540
rect 10873 12484 10877 12540
rect 10813 12480 10877 12484
rect 10893 12540 10957 12544
rect 10893 12484 10897 12540
rect 10897 12484 10953 12540
rect 10953 12484 10957 12540
rect 10893 12480 10957 12484
rect 10973 12540 11037 12544
rect 10973 12484 10977 12540
rect 10977 12484 11033 12540
rect 11033 12484 11037 12540
rect 10973 12480 11037 12484
rect 11053 12540 11117 12544
rect 11053 12484 11057 12540
rect 11057 12484 11113 12540
rect 11113 12484 11117 12540
rect 11053 12480 11117 12484
rect 3417 11996 3481 12000
rect 3417 11940 3421 11996
rect 3421 11940 3477 11996
rect 3477 11940 3481 11996
rect 3417 11936 3481 11940
rect 3497 11996 3561 12000
rect 3497 11940 3501 11996
rect 3501 11940 3557 11996
rect 3557 11940 3561 11996
rect 3497 11936 3561 11940
rect 3577 11996 3641 12000
rect 3577 11940 3581 11996
rect 3581 11940 3637 11996
rect 3637 11940 3641 11996
rect 3577 11936 3641 11940
rect 3657 11996 3721 12000
rect 3657 11940 3661 11996
rect 3661 11940 3717 11996
rect 3717 11940 3721 11996
rect 3657 11936 3721 11940
rect 8348 11996 8412 12000
rect 8348 11940 8352 11996
rect 8352 11940 8408 11996
rect 8408 11940 8412 11996
rect 8348 11936 8412 11940
rect 8428 11996 8492 12000
rect 8428 11940 8432 11996
rect 8432 11940 8488 11996
rect 8488 11940 8492 11996
rect 8428 11936 8492 11940
rect 8508 11996 8572 12000
rect 8508 11940 8512 11996
rect 8512 11940 8568 11996
rect 8568 11940 8572 11996
rect 8508 11936 8572 11940
rect 8588 11996 8652 12000
rect 8588 11940 8592 11996
rect 8592 11940 8648 11996
rect 8648 11940 8652 11996
rect 8588 11936 8652 11940
rect 13278 11996 13342 12000
rect 13278 11940 13282 11996
rect 13282 11940 13338 11996
rect 13338 11940 13342 11996
rect 13278 11936 13342 11940
rect 13358 11996 13422 12000
rect 13358 11940 13362 11996
rect 13362 11940 13418 11996
rect 13418 11940 13422 11996
rect 13358 11936 13422 11940
rect 13438 11996 13502 12000
rect 13438 11940 13442 11996
rect 13442 11940 13498 11996
rect 13498 11940 13502 11996
rect 13438 11936 13502 11940
rect 13518 11996 13582 12000
rect 13518 11940 13522 11996
rect 13522 11940 13578 11996
rect 13578 11940 13582 11996
rect 13518 11936 13582 11940
rect 9444 11656 9508 11660
rect 9444 11600 9458 11656
rect 9458 11600 9508 11656
rect 9444 11596 9508 11600
rect 5882 11452 5946 11456
rect 5882 11396 5886 11452
rect 5886 11396 5942 11452
rect 5942 11396 5946 11452
rect 5882 11392 5946 11396
rect 5962 11452 6026 11456
rect 5962 11396 5966 11452
rect 5966 11396 6022 11452
rect 6022 11396 6026 11452
rect 5962 11392 6026 11396
rect 6042 11452 6106 11456
rect 6042 11396 6046 11452
rect 6046 11396 6102 11452
rect 6102 11396 6106 11452
rect 6042 11392 6106 11396
rect 6122 11452 6186 11456
rect 6122 11396 6126 11452
rect 6126 11396 6182 11452
rect 6182 11396 6186 11452
rect 6122 11392 6186 11396
rect 10813 11452 10877 11456
rect 10813 11396 10817 11452
rect 10817 11396 10873 11452
rect 10873 11396 10877 11452
rect 10813 11392 10877 11396
rect 10893 11452 10957 11456
rect 10893 11396 10897 11452
rect 10897 11396 10953 11452
rect 10953 11396 10957 11452
rect 10893 11392 10957 11396
rect 10973 11452 11037 11456
rect 10973 11396 10977 11452
rect 10977 11396 11033 11452
rect 11033 11396 11037 11452
rect 10973 11392 11037 11396
rect 11053 11452 11117 11456
rect 11053 11396 11057 11452
rect 11057 11396 11113 11452
rect 11113 11396 11117 11452
rect 11053 11392 11117 11396
rect 3417 10908 3481 10912
rect 3417 10852 3421 10908
rect 3421 10852 3477 10908
rect 3477 10852 3481 10908
rect 3417 10848 3481 10852
rect 3497 10908 3561 10912
rect 3497 10852 3501 10908
rect 3501 10852 3557 10908
rect 3557 10852 3561 10908
rect 3497 10848 3561 10852
rect 3577 10908 3641 10912
rect 3577 10852 3581 10908
rect 3581 10852 3637 10908
rect 3637 10852 3641 10908
rect 3577 10848 3641 10852
rect 3657 10908 3721 10912
rect 3657 10852 3661 10908
rect 3661 10852 3717 10908
rect 3717 10852 3721 10908
rect 3657 10848 3721 10852
rect 8348 10908 8412 10912
rect 8348 10852 8352 10908
rect 8352 10852 8408 10908
rect 8408 10852 8412 10908
rect 8348 10848 8412 10852
rect 8428 10908 8492 10912
rect 8428 10852 8432 10908
rect 8432 10852 8488 10908
rect 8488 10852 8492 10908
rect 8428 10848 8492 10852
rect 8508 10908 8572 10912
rect 8508 10852 8512 10908
rect 8512 10852 8568 10908
rect 8568 10852 8572 10908
rect 8508 10848 8572 10852
rect 8588 10908 8652 10912
rect 8588 10852 8592 10908
rect 8592 10852 8648 10908
rect 8648 10852 8652 10908
rect 8588 10848 8652 10852
rect 13278 10908 13342 10912
rect 13278 10852 13282 10908
rect 13282 10852 13338 10908
rect 13338 10852 13342 10908
rect 13278 10848 13342 10852
rect 13358 10908 13422 10912
rect 13358 10852 13362 10908
rect 13362 10852 13418 10908
rect 13418 10852 13422 10908
rect 13358 10848 13422 10852
rect 13438 10908 13502 10912
rect 13438 10852 13442 10908
rect 13442 10852 13498 10908
rect 13498 10852 13502 10908
rect 13438 10848 13502 10852
rect 13518 10908 13582 10912
rect 13518 10852 13522 10908
rect 13522 10852 13578 10908
rect 13578 10852 13582 10908
rect 13518 10848 13582 10852
rect 5882 10364 5946 10368
rect 5882 10308 5886 10364
rect 5886 10308 5942 10364
rect 5942 10308 5946 10364
rect 5882 10304 5946 10308
rect 5962 10364 6026 10368
rect 5962 10308 5966 10364
rect 5966 10308 6022 10364
rect 6022 10308 6026 10364
rect 5962 10304 6026 10308
rect 6042 10364 6106 10368
rect 6042 10308 6046 10364
rect 6046 10308 6102 10364
rect 6102 10308 6106 10364
rect 6042 10304 6106 10308
rect 6122 10364 6186 10368
rect 6122 10308 6126 10364
rect 6126 10308 6182 10364
rect 6182 10308 6186 10364
rect 6122 10304 6186 10308
rect 10813 10364 10877 10368
rect 10813 10308 10817 10364
rect 10817 10308 10873 10364
rect 10873 10308 10877 10364
rect 10813 10304 10877 10308
rect 10893 10364 10957 10368
rect 10893 10308 10897 10364
rect 10897 10308 10953 10364
rect 10953 10308 10957 10364
rect 10893 10304 10957 10308
rect 10973 10364 11037 10368
rect 10973 10308 10977 10364
rect 10977 10308 11033 10364
rect 11033 10308 11037 10364
rect 10973 10304 11037 10308
rect 11053 10364 11117 10368
rect 11053 10308 11057 10364
rect 11057 10308 11113 10364
rect 11113 10308 11117 10364
rect 11053 10304 11117 10308
rect 9444 10296 9508 10300
rect 9444 10240 9458 10296
rect 9458 10240 9508 10296
rect 9444 10236 9508 10240
rect 3417 9820 3481 9824
rect 3417 9764 3421 9820
rect 3421 9764 3477 9820
rect 3477 9764 3481 9820
rect 3417 9760 3481 9764
rect 3497 9820 3561 9824
rect 3497 9764 3501 9820
rect 3501 9764 3557 9820
rect 3557 9764 3561 9820
rect 3497 9760 3561 9764
rect 3577 9820 3641 9824
rect 3577 9764 3581 9820
rect 3581 9764 3637 9820
rect 3637 9764 3641 9820
rect 3577 9760 3641 9764
rect 3657 9820 3721 9824
rect 3657 9764 3661 9820
rect 3661 9764 3717 9820
rect 3717 9764 3721 9820
rect 3657 9760 3721 9764
rect 8348 9820 8412 9824
rect 8348 9764 8352 9820
rect 8352 9764 8408 9820
rect 8408 9764 8412 9820
rect 8348 9760 8412 9764
rect 8428 9820 8492 9824
rect 8428 9764 8432 9820
rect 8432 9764 8488 9820
rect 8488 9764 8492 9820
rect 8428 9760 8492 9764
rect 8508 9820 8572 9824
rect 8508 9764 8512 9820
rect 8512 9764 8568 9820
rect 8568 9764 8572 9820
rect 8508 9760 8572 9764
rect 8588 9820 8652 9824
rect 8588 9764 8592 9820
rect 8592 9764 8648 9820
rect 8648 9764 8652 9820
rect 8588 9760 8652 9764
rect 13278 9820 13342 9824
rect 13278 9764 13282 9820
rect 13282 9764 13338 9820
rect 13338 9764 13342 9820
rect 13278 9760 13342 9764
rect 13358 9820 13422 9824
rect 13358 9764 13362 9820
rect 13362 9764 13418 9820
rect 13418 9764 13422 9820
rect 13358 9760 13422 9764
rect 13438 9820 13502 9824
rect 13438 9764 13442 9820
rect 13442 9764 13498 9820
rect 13498 9764 13502 9820
rect 13438 9760 13502 9764
rect 13518 9820 13582 9824
rect 13518 9764 13522 9820
rect 13522 9764 13578 9820
rect 13578 9764 13582 9820
rect 13518 9760 13582 9764
rect 9812 9556 9876 9620
rect 5882 9276 5946 9280
rect 5882 9220 5886 9276
rect 5886 9220 5942 9276
rect 5942 9220 5946 9276
rect 5882 9216 5946 9220
rect 5962 9276 6026 9280
rect 5962 9220 5966 9276
rect 5966 9220 6022 9276
rect 6022 9220 6026 9276
rect 5962 9216 6026 9220
rect 6042 9276 6106 9280
rect 6042 9220 6046 9276
rect 6046 9220 6102 9276
rect 6102 9220 6106 9276
rect 6042 9216 6106 9220
rect 6122 9276 6186 9280
rect 6122 9220 6126 9276
rect 6126 9220 6182 9276
rect 6182 9220 6186 9276
rect 6122 9216 6186 9220
rect 10813 9276 10877 9280
rect 10813 9220 10817 9276
rect 10817 9220 10873 9276
rect 10873 9220 10877 9276
rect 10813 9216 10877 9220
rect 10893 9276 10957 9280
rect 10893 9220 10897 9276
rect 10897 9220 10953 9276
rect 10953 9220 10957 9276
rect 10893 9216 10957 9220
rect 10973 9276 11037 9280
rect 10973 9220 10977 9276
rect 10977 9220 11033 9276
rect 11033 9220 11037 9276
rect 10973 9216 11037 9220
rect 11053 9276 11117 9280
rect 11053 9220 11057 9276
rect 11057 9220 11113 9276
rect 11113 9220 11117 9276
rect 11053 9216 11117 9220
rect 3417 8732 3481 8736
rect 3417 8676 3421 8732
rect 3421 8676 3477 8732
rect 3477 8676 3481 8732
rect 3417 8672 3481 8676
rect 3497 8732 3561 8736
rect 3497 8676 3501 8732
rect 3501 8676 3557 8732
rect 3557 8676 3561 8732
rect 3497 8672 3561 8676
rect 3577 8732 3641 8736
rect 3577 8676 3581 8732
rect 3581 8676 3637 8732
rect 3637 8676 3641 8732
rect 3577 8672 3641 8676
rect 3657 8732 3721 8736
rect 3657 8676 3661 8732
rect 3661 8676 3717 8732
rect 3717 8676 3721 8732
rect 3657 8672 3721 8676
rect 8348 8732 8412 8736
rect 8348 8676 8352 8732
rect 8352 8676 8408 8732
rect 8408 8676 8412 8732
rect 8348 8672 8412 8676
rect 8428 8732 8492 8736
rect 8428 8676 8432 8732
rect 8432 8676 8488 8732
rect 8488 8676 8492 8732
rect 8428 8672 8492 8676
rect 8508 8732 8572 8736
rect 8508 8676 8512 8732
rect 8512 8676 8568 8732
rect 8568 8676 8572 8732
rect 8508 8672 8572 8676
rect 8588 8732 8652 8736
rect 8588 8676 8592 8732
rect 8592 8676 8648 8732
rect 8648 8676 8652 8732
rect 8588 8672 8652 8676
rect 13278 8732 13342 8736
rect 13278 8676 13282 8732
rect 13282 8676 13338 8732
rect 13338 8676 13342 8732
rect 13278 8672 13342 8676
rect 13358 8732 13422 8736
rect 13358 8676 13362 8732
rect 13362 8676 13418 8732
rect 13418 8676 13422 8732
rect 13358 8672 13422 8676
rect 13438 8732 13502 8736
rect 13438 8676 13442 8732
rect 13442 8676 13498 8732
rect 13498 8676 13502 8732
rect 13438 8672 13502 8676
rect 13518 8732 13582 8736
rect 13518 8676 13522 8732
rect 13522 8676 13578 8732
rect 13578 8676 13582 8732
rect 13518 8672 13582 8676
rect 9628 8256 9692 8260
rect 9628 8200 9642 8256
rect 9642 8200 9692 8256
rect 9628 8196 9692 8200
rect 5882 8188 5946 8192
rect 5882 8132 5886 8188
rect 5886 8132 5942 8188
rect 5942 8132 5946 8188
rect 5882 8128 5946 8132
rect 5962 8188 6026 8192
rect 5962 8132 5966 8188
rect 5966 8132 6022 8188
rect 6022 8132 6026 8188
rect 5962 8128 6026 8132
rect 6042 8188 6106 8192
rect 6042 8132 6046 8188
rect 6046 8132 6102 8188
rect 6102 8132 6106 8188
rect 6042 8128 6106 8132
rect 6122 8188 6186 8192
rect 6122 8132 6126 8188
rect 6126 8132 6182 8188
rect 6182 8132 6186 8188
rect 6122 8128 6186 8132
rect 10813 8188 10877 8192
rect 10813 8132 10817 8188
rect 10817 8132 10873 8188
rect 10873 8132 10877 8188
rect 10813 8128 10877 8132
rect 10893 8188 10957 8192
rect 10893 8132 10897 8188
rect 10897 8132 10953 8188
rect 10953 8132 10957 8188
rect 10893 8128 10957 8132
rect 10973 8188 11037 8192
rect 10973 8132 10977 8188
rect 10977 8132 11033 8188
rect 11033 8132 11037 8188
rect 10973 8128 11037 8132
rect 11053 8188 11117 8192
rect 11053 8132 11057 8188
rect 11057 8132 11113 8188
rect 11113 8132 11117 8188
rect 11053 8128 11117 8132
rect 9812 8060 9876 8124
rect 3417 7644 3481 7648
rect 3417 7588 3421 7644
rect 3421 7588 3477 7644
rect 3477 7588 3481 7644
rect 3417 7584 3481 7588
rect 3497 7644 3561 7648
rect 3497 7588 3501 7644
rect 3501 7588 3557 7644
rect 3557 7588 3561 7644
rect 3497 7584 3561 7588
rect 3577 7644 3641 7648
rect 3577 7588 3581 7644
rect 3581 7588 3637 7644
rect 3637 7588 3641 7644
rect 3577 7584 3641 7588
rect 3657 7644 3721 7648
rect 3657 7588 3661 7644
rect 3661 7588 3717 7644
rect 3717 7588 3721 7644
rect 3657 7584 3721 7588
rect 8348 7644 8412 7648
rect 8348 7588 8352 7644
rect 8352 7588 8408 7644
rect 8408 7588 8412 7644
rect 8348 7584 8412 7588
rect 8428 7644 8492 7648
rect 8428 7588 8432 7644
rect 8432 7588 8488 7644
rect 8488 7588 8492 7644
rect 8428 7584 8492 7588
rect 8508 7644 8572 7648
rect 8508 7588 8512 7644
rect 8512 7588 8568 7644
rect 8568 7588 8572 7644
rect 8508 7584 8572 7588
rect 8588 7644 8652 7648
rect 8588 7588 8592 7644
rect 8592 7588 8648 7644
rect 8648 7588 8652 7644
rect 8588 7584 8652 7588
rect 13278 7644 13342 7648
rect 13278 7588 13282 7644
rect 13282 7588 13338 7644
rect 13338 7588 13342 7644
rect 13278 7584 13342 7588
rect 13358 7644 13422 7648
rect 13358 7588 13362 7644
rect 13362 7588 13418 7644
rect 13418 7588 13422 7644
rect 13358 7584 13422 7588
rect 13438 7644 13502 7648
rect 13438 7588 13442 7644
rect 13442 7588 13498 7644
rect 13498 7588 13502 7644
rect 13438 7584 13502 7588
rect 13518 7644 13582 7648
rect 13518 7588 13522 7644
rect 13522 7588 13578 7644
rect 13578 7588 13582 7644
rect 13518 7584 13582 7588
rect 5882 7100 5946 7104
rect 5882 7044 5886 7100
rect 5886 7044 5942 7100
rect 5942 7044 5946 7100
rect 5882 7040 5946 7044
rect 5962 7100 6026 7104
rect 5962 7044 5966 7100
rect 5966 7044 6022 7100
rect 6022 7044 6026 7100
rect 5962 7040 6026 7044
rect 6042 7100 6106 7104
rect 6042 7044 6046 7100
rect 6046 7044 6102 7100
rect 6102 7044 6106 7100
rect 6042 7040 6106 7044
rect 6122 7100 6186 7104
rect 6122 7044 6126 7100
rect 6126 7044 6182 7100
rect 6182 7044 6186 7100
rect 6122 7040 6186 7044
rect 10813 7100 10877 7104
rect 10813 7044 10817 7100
rect 10817 7044 10873 7100
rect 10873 7044 10877 7100
rect 10813 7040 10877 7044
rect 10893 7100 10957 7104
rect 10893 7044 10897 7100
rect 10897 7044 10953 7100
rect 10953 7044 10957 7100
rect 10893 7040 10957 7044
rect 10973 7100 11037 7104
rect 10973 7044 10977 7100
rect 10977 7044 11033 7100
rect 11033 7044 11037 7100
rect 10973 7040 11037 7044
rect 11053 7100 11117 7104
rect 11053 7044 11057 7100
rect 11057 7044 11113 7100
rect 11113 7044 11117 7100
rect 11053 7040 11117 7044
rect 3417 6556 3481 6560
rect 3417 6500 3421 6556
rect 3421 6500 3477 6556
rect 3477 6500 3481 6556
rect 3417 6496 3481 6500
rect 3497 6556 3561 6560
rect 3497 6500 3501 6556
rect 3501 6500 3557 6556
rect 3557 6500 3561 6556
rect 3497 6496 3561 6500
rect 3577 6556 3641 6560
rect 3577 6500 3581 6556
rect 3581 6500 3637 6556
rect 3637 6500 3641 6556
rect 3577 6496 3641 6500
rect 3657 6556 3721 6560
rect 3657 6500 3661 6556
rect 3661 6500 3717 6556
rect 3717 6500 3721 6556
rect 3657 6496 3721 6500
rect 8348 6556 8412 6560
rect 8348 6500 8352 6556
rect 8352 6500 8408 6556
rect 8408 6500 8412 6556
rect 8348 6496 8412 6500
rect 8428 6556 8492 6560
rect 8428 6500 8432 6556
rect 8432 6500 8488 6556
rect 8488 6500 8492 6556
rect 8428 6496 8492 6500
rect 8508 6556 8572 6560
rect 8508 6500 8512 6556
rect 8512 6500 8568 6556
rect 8568 6500 8572 6556
rect 8508 6496 8572 6500
rect 8588 6556 8652 6560
rect 8588 6500 8592 6556
rect 8592 6500 8648 6556
rect 8648 6500 8652 6556
rect 8588 6496 8652 6500
rect 13278 6556 13342 6560
rect 13278 6500 13282 6556
rect 13282 6500 13338 6556
rect 13338 6500 13342 6556
rect 13278 6496 13342 6500
rect 13358 6556 13422 6560
rect 13358 6500 13362 6556
rect 13362 6500 13418 6556
rect 13418 6500 13422 6556
rect 13358 6496 13422 6500
rect 13438 6556 13502 6560
rect 13438 6500 13442 6556
rect 13442 6500 13498 6556
rect 13498 6500 13502 6556
rect 13438 6496 13502 6500
rect 13518 6556 13582 6560
rect 13518 6500 13522 6556
rect 13522 6500 13578 6556
rect 13578 6500 13582 6556
rect 13518 6496 13582 6500
rect 5882 6012 5946 6016
rect 5882 5956 5886 6012
rect 5886 5956 5942 6012
rect 5942 5956 5946 6012
rect 5882 5952 5946 5956
rect 5962 6012 6026 6016
rect 5962 5956 5966 6012
rect 5966 5956 6022 6012
rect 6022 5956 6026 6012
rect 5962 5952 6026 5956
rect 6042 6012 6106 6016
rect 6042 5956 6046 6012
rect 6046 5956 6102 6012
rect 6102 5956 6106 6012
rect 6042 5952 6106 5956
rect 6122 6012 6186 6016
rect 6122 5956 6126 6012
rect 6126 5956 6182 6012
rect 6182 5956 6186 6012
rect 6122 5952 6186 5956
rect 10813 6012 10877 6016
rect 10813 5956 10817 6012
rect 10817 5956 10873 6012
rect 10873 5956 10877 6012
rect 10813 5952 10877 5956
rect 10893 6012 10957 6016
rect 10893 5956 10897 6012
rect 10897 5956 10953 6012
rect 10953 5956 10957 6012
rect 10893 5952 10957 5956
rect 10973 6012 11037 6016
rect 10973 5956 10977 6012
rect 10977 5956 11033 6012
rect 11033 5956 11037 6012
rect 10973 5952 11037 5956
rect 11053 6012 11117 6016
rect 11053 5956 11057 6012
rect 11057 5956 11113 6012
rect 11113 5956 11117 6012
rect 11053 5952 11117 5956
rect 3417 5468 3481 5472
rect 3417 5412 3421 5468
rect 3421 5412 3477 5468
rect 3477 5412 3481 5468
rect 3417 5408 3481 5412
rect 3497 5468 3561 5472
rect 3497 5412 3501 5468
rect 3501 5412 3557 5468
rect 3557 5412 3561 5468
rect 3497 5408 3561 5412
rect 3577 5468 3641 5472
rect 3577 5412 3581 5468
rect 3581 5412 3637 5468
rect 3637 5412 3641 5468
rect 3577 5408 3641 5412
rect 3657 5468 3721 5472
rect 3657 5412 3661 5468
rect 3661 5412 3717 5468
rect 3717 5412 3721 5468
rect 3657 5408 3721 5412
rect 8348 5468 8412 5472
rect 8348 5412 8352 5468
rect 8352 5412 8408 5468
rect 8408 5412 8412 5468
rect 8348 5408 8412 5412
rect 8428 5468 8492 5472
rect 8428 5412 8432 5468
rect 8432 5412 8488 5468
rect 8488 5412 8492 5468
rect 8428 5408 8492 5412
rect 8508 5468 8572 5472
rect 8508 5412 8512 5468
rect 8512 5412 8568 5468
rect 8568 5412 8572 5468
rect 8508 5408 8572 5412
rect 8588 5468 8652 5472
rect 8588 5412 8592 5468
rect 8592 5412 8648 5468
rect 8648 5412 8652 5468
rect 8588 5408 8652 5412
rect 13278 5468 13342 5472
rect 13278 5412 13282 5468
rect 13282 5412 13338 5468
rect 13338 5412 13342 5468
rect 13278 5408 13342 5412
rect 13358 5468 13422 5472
rect 13358 5412 13362 5468
rect 13362 5412 13418 5468
rect 13418 5412 13422 5468
rect 13358 5408 13422 5412
rect 13438 5468 13502 5472
rect 13438 5412 13442 5468
rect 13442 5412 13498 5468
rect 13498 5412 13502 5468
rect 13438 5408 13502 5412
rect 13518 5468 13582 5472
rect 13518 5412 13522 5468
rect 13522 5412 13578 5468
rect 13578 5412 13582 5468
rect 13518 5408 13582 5412
rect 5882 4924 5946 4928
rect 5882 4868 5886 4924
rect 5886 4868 5942 4924
rect 5942 4868 5946 4924
rect 5882 4864 5946 4868
rect 5962 4924 6026 4928
rect 5962 4868 5966 4924
rect 5966 4868 6022 4924
rect 6022 4868 6026 4924
rect 5962 4864 6026 4868
rect 6042 4924 6106 4928
rect 6042 4868 6046 4924
rect 6046 4868 6102 4924
rect 6102 4868 6106 4924
rect 6042 4864 6106 4868
rect 6122 4924 6186 4928
rect 6122 4868 6126 4924
rect 6126 4868 6182 4924
rect 6182 4868 6186 4924
rect 6122 4864 6186 4868
rect 10813 4924 10877 4928
rect 10813 4868 10817 4924
rect 10817 4868 10873 4924
rect 10873 4868 10877 4924
rect 10813 4864 10877 4868
rect 10893 4924 10957 4928
rect 10893 4868 10897 4924
rect 10897 4868 10953 4924
rect 10953 4868 10957 4924
rect 10893 4864 10957 4868
rect 10973 4924 11037 4928
rect 10973 4868 10977 4924
rect 10977 4868 11033 4924
rect 11033 4868 11037 4924
rect 10973 4864 11037 4868
rect 11053 4924 11117 4928
rect 11053 4868 11057 4924
rect 11057 4868 11113 4924
rect 11113 4868 11117 4924
rect 11053 4864 11117 4868
rect 3417 4380 3481 4384
rect 3417 4324 3421 4380
rect 3421 4324 3477 4380
rect 3477 4324 3481 4380
rect 3417 4320 3481 4324
rect 3497 4380 3561 4384
rect 3497 4324 3501 4380
rect 3501 4324 3557 4380
rect 3557 4324 3561 4380
rect 3497 4320 3561 4324
rect 3577 4380 3641 4384
rect 3577 4324 3581 4380
rect 3581 4324 3637 4380
rect 3637 4324 3641 4380
rect 3577 4320 3641 4324
rect 3657 4380 3721 4384
rect 3657 4324 3661 4380
rect 3661 4324 3717 4380
rect 3717 4324 3721 4380
rect 3657 4320 3721 4324
rect 8348 4380 8412 4384
rect 8348 4324 8352 4380
rect 8352 4324 8408 4380
rect 8408 4324 8412 4380
rect 8348 4320 8412 4324
rect 8428 4380 8492 4384
rect 8428 4324 8432 4380
rect 8432 4324 8488 4380
rect 8488 4324 8492 4380
rect 8428 4320 8492 4324
rect 8508 4380 8572 4384
rect 8508 4324 8512 4380
rect 8512 4324 8568 4380
rect 8568 4324 8572 4380
rect 8508 4320 8572 4324
rect 8588 4380 8652 4384
rect 8588 4324 8592 4380
rect 8592 4324 8648 4380
rect 8648 4324 8652 4380
rect 8588 4320 8652 4324
rect 13278 4380 13342 4384
rect 13278 4324 13282 4380
rect 13282 4324 13338 4380
rect 13338 4324 13342 4380
rect 13278 4320 13342 4324
rect 13358 4380 13422 4384
rect 13358 4324 13362 4380
rect 13362 4324 13418 4380
rect 13418 4324 13422 4380
rect 13358 4320 13422 4324
rect 13438 4380 13502 4384
rect 13438 4324 13442 4380
rect 13442 4324 13498 4380
rect 13498 4324 13502 4380
rect 13438 4320 13502 4324
rect 13518 4380 13582 4384
rect 13518 4324 13522 4380
rect 13522 4324 13578 4380
rect 13578 4324 13582 4380
rect 13518 4320 13582 4324
rect 5882 3836 5946 3840
rect 5882 3780 5886 3836
rect 5886 3780 5942 3836
rect 5942 3780 5946 3836
rect 5882 3776 5946 3780
rect 5962 3836 6026 3840
rect 5962 3780 5966 3836
rect 5966 3780 6022 3836
rect 6022 3780 6026 3836
rect 5962 3776 6026 3780
rect 6042 3836 6106 3840
rect 6042 3780 6046 3836
rect 6046 3780 6102 3836
rect 6102 3780 6106 3836
rect 6042 3776 6106 3780
rect 6122 3836 6186 3840
rect 6122 3780 6126 3836
rect 6126 3780 6182 3836
rect 6182 3780 6186 3836
rect 6122 3776 6186 3780
rect 10813 3836 10877 3840
rect 10813 3780 10817 3836
rect 10817 3780 10873 3836
rect 10873 3780 10877 3836
rect 10813 3776 10877 3780
rect 10893 3836 10957 3840
rect 10893 3780 10897 3836
rect 10897 3780 10953 3836
rect 10953 3780 10957 3836
rect 10893 3776 10957 3780
rect 10973 3836 11037 3840
rect 10973 3780 10977 3836
rect 10977 3780 11033 3836
rect 11033 3780 11037 3836
rect 10973 3776 11037 3780
rect 11053 3836 11117 3840
rect 11053 3780 11057 3836
rect 11057 3780 11113 3836
rect 11113 3780 11117 3836
rect 11053 3776 11117 3780
rect 3417 3292 3481 3296
rect 3417 3236 3421 3292
rect 3421 3236 3477 3292
rect 3477 3236 3481 3292
rect 3417 3232 3481 3236
rect 3497 3292 3561 3296
rect 3497 3236 3501 3292
rect 3501 3236 3557 3292
rect 3557 3236 3561 3292
rect 3497 3232 3561 3236
rect 3577 3292 3641 3296
rect 3577 3236 3581 3292
rect 3581 3236 3637 3292
rect 3637 3236 3641 3292
rect 3577 3232 3641 3236
rect 3657 3292 3721 3296
rect 3657 3236 3661 3292
rect 3661 3236 3717 3292
rect 3717 3236 3721 3292
rect 3657 3232 3721 3236
rect 8348 3292 8412 3296
rect 8348 3236 8352 3292
rect 8352 3236 8408 3292
rect 8408 3236 8412 3292
rect 8348 3232 8412 3236
rect 8428 3292 8492 3296
rect 8428 3236 8432 3292
rect 8432 3236 8488 3292
rect 8488 3236 8492 3292
rect 8428 3232 8492 3236
rect 8508 3292 8572 3296
rect 8508 3236 8512 3292
rect 8512 3236 8568 3292
rect 8568 3236 8572 3292
rect 8508 3232 8572 3236
rect 8588 3292 8652 3296
rect 8588 3236 8592 3292
rect 8592 3236 8648 3292
rect 8648 3236 8652 3292
rect 8588 3232 8652 3236
rect 13278 3292 13342 3296
rect 13278 3236 13282 3292
rect 13282 3236 13338 3292
rect 13338 3236 13342 3292
rect 13278 3232 13342 3236
rect 13358 3292 13422 3296
rect 13358 3236 13362 3292
rect 13362 3236 13418 3292
rect 13418 3236 13422 3292
rect 13358 3232 13422 3236
rect 13438 3292 13502 3296
rect 13438 3236 13442 3292
rect 13442 3236 13498 3292
rect 13498 3236 13502 3292
rect 13438 3232 13502 3236
rect 13518 3292 13582 3296
rect 13518 3236 13522 3292
rect 13522 3236 13578 3292
rect 13578 3236 13582 3292
rect 13518 3232 13582 3236
rect 5882 2748 5946 2752
rect 5882 2692 5886 2748
rect 5886 2692 5942 2748
rect 5942 2692 5946 2748
rect 5882 2688 5946 2692
rect 5962 2748 6026 2752
rect 5962 2692 5966 2748
rect 5966 2692 6022 2748
rect 6022 2692 6026 2748
rect 5962 2688 6026 2692
rect 6042 2748 6106 2752
rect 6042 2692 6046 2748
rect 6046 2692 6102 2748
rect 6102 2692 6106 2748
rect 6042 2688 6106 2692
rect 6122 2748 6186 2752
rect 6122 2692 6126 2748
rect 6126 2692 6182 2748
rect 6182 2692 6186 2748
rect 6122 2688 6186 2692
rect 10813 2748 10877 2752
rect 10813 2692 10817 2748
rect 10817 2692 10873 2748
rect 10873 2692 10877 2748
rect 10813 2688 10877 2692
rect 10893 2748 10957 2752
rect 10893 2692 10897 2748
rect 10897 2692 10953 2748
rect 10953 2692 10957 2748
rect 10893 2688 10957 2692
rect 10973 2748 11037 2752
rect 10973 2692 10977 2748
rect 10977 2692 11033 2748
rect 11033 2692 11037 2748
rect 10973 2688 11037 2692
rect 11053 2748 11117 2752
rect 11053 2692 11057 2748
rect 11057 2692 11113 2748
rect 11113 2692 11117 2748
rect 11053 2688 11117 2692
rect 9628 2620 9692 2684
rect 3417 2204 3481 2208
rect 3417 2148 3421 2204
rect 3421 2148 3477 2204
rect 3477 2148 3481 2204
rect 3417 2144 3481 2148
rect 3497 2204 3561 2208
rect 3497 2148 3501 2204
rect 3501 2148 3557 2204
rect 3557 2148 3561 2204
rect 3497 2144 3561 2148
rect 3577 2204 3641 2208
rect 3577 2148 3581 2204
rect 3581 2148 3637 2204
rect 3637 2148 3641 2204
rect 3577 2144 3641 2148
rect 3657 2204 3721 2208
rect 3657 2148 3661 2204
rect 3661 2148 3717 2204
rect 3717 2148 3721 2204
rect 3657 2144 3721 2148
rect 8348 2204 8412 2208
rect 8348 2148 8352 2204
rect 8352 2148 8408 2204
rect 8408 2148 8412 2204
rect 8348 2144 8412 2148
rect 8428 2204 8492 2208
rect 8428 2148 8432 2204
rect 8432 2148 8488 2204
rect 8488 2148 8492 2204
rect 8428 2144 8492 2148
rect 8508 2204 8572 2208
rect 8508 2148 8512 2204
rect 8512 2148 8568 2204
rect 8568 2148 8572 2204
rect 8508 2144 8572 2148
rect 8588 2204 8652 2208
rect 8588 2148 8592 2204
rect 8592 2148 8648 2204
rect 8648 2148 8652 2204
rect 8588 2144 8652 2148
rect 13278 2204 13342 2208
rect 13278 2148 13282 2204
rect 13282 2148 13338 2204
rect 13338 2148 13342 2204
rect 13278 2144 13342 2148
rect 13358 2204 13422 2208
rect 13358 2148 13362 2204
rect 13362 2148 13418 2204
rect 13418 2148 13422 2204
rect 13358 2144 13422 2148
rect 13438 2204 13502 2208
rect 13438 2148 13442 2204
rect 13442 2148 13498 2204
rect 13498 2148 13502 2204
rect 13438 2144 13502 2148
rect 13518 2204 13582 2208
rect 13518 2148 13522 2204
rect 13522 2148 13578 2204
rect 13578 2148 13582 2204
rect 13518 2144 13582 2148
<< metal4 >>
rect 3409 17440 3729 17456
rect 3409 17376 3417 17440
rect 3481 17376 3497 17440
rect 3561 17376 3577 17440
rect 3641 17376 3657 17440
rect 3721 17376 3729 17440
rect 3409 16352 3729 17376
rect 3409 16288 3417 16352
rect 3481 16288 3497 16352
rect 3561 16288 3577 16352
rect 3641 16288 3657 16352
rect 3721 16288 3729 16352
rect 3409 15264 3729 16288
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 14176 3729 15200
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 13088 3729 14112
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 12000 3729 13024
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 10912 3729 11936
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 9824 3729 10848
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 8736 3729 9760
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 7648 3729 8672
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 6560 3729 7584
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 5472 3729 6496
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 4384 3729 5408
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 3296 3729 4320
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 2208 3729 3232
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2128 3729 2144
rect 5874 16896 6195 17456
rect 5874 16832 5882 16896
rect 5946 16832 5962 16896
rect 6026 16832 6042 16896
rect 6106 16832 6122 16896
rect 6186 16832 6195 16896
rect 5874 15808 6195 16832
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6195 15808
rect 5874 14720 6195 15744
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6195 14720
rect 5874 13632 6195 14656
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6195 13632
rect 5874 12544 6195 13568
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6195 12544
rect 5874 11456 6195 12480
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6195 11456
rect 5874 10368 6195 11392
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6195 10368
rect 5874 9280 6195 10304
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6195 9280
rect 5874 8192 6195 9216
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6195 8192
rect 5874 7104 6195 8128
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6195 7104
rect 5874 6016 6195 7040
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6195 6016
rect 5874 4928 6195 5952
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6195 4928
rect 5874 3840 6195 4864
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6195 3840
rect 5874 2752 6195 3776
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6195 2752
rect 5874 2128 6195 2688
rect 8340 17440 8660 17456
rect 8340 17376 8348 17440
rect 8412 17376 8428 17440
rect 8492 17376 8508 17440
rect 8572 17376 8588 17440
rect 8652 17376 8660 17440
rect 8340 16352 8660 17376
rect 8340 16288 8348 16352
rect 8412 16288 8428 16352
rect 8492 16288 8508 16352
rect 8572 16288 8588 16352
rect 8652 16288 8660 16352
rect 8340 15264 8660 16288
rect 10805 16896 11125 17456
rect 10805 16832 10813 16896
rect 10877 16832 10893 16896
rect 10957 16832 10973 16896
rect 11037 16832 11053 16896
rect 11117 16832 11125 16896
rect 9443 16148 9509 16149
rect 9443 16084 9444 16148
rect 9508 16084 9509 16148
rect 9443 16083 9509 16084
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 14176 8660 15200
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 13088 8660 14112
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 12000 8660 13024
rect 9446 12749 9506 16083
rect 10805 15808 11125 16832
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 14720 11125 15744
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 13632 11125 14656
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 9443 12748 9509 12749
rect 9443 12684 9444 12748
rect 9508 12684 9509 12748
rect 9443 12683 9509 12684
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 10912 8660 11936
rect 10805 12544 11125 13568
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 9443 11660 9509 11661
rect 9443 11596 9444 11660
rect 9508 11596 9509 11660
rect 9443 11595 9509 11596
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 9824 8660 10848
rect 9446 10301 9506 11595
rect 10805 11456 11125 12480
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 10368 11125 11392
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 9443 10300 9509 10301
rect 9443 10236 9444 10300
rect 9508 10236 9509 10300
rect 9443 10235 9509 10236
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 8736 8660 9760
rect 9811 9620 9877 9621
rect 9811 9556 9812 9620
rect 9876 9556 9877 9620
rect 9811 9555 9877 9556
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 7648 8660 8672
rect 9627 8260 9693 8261
rect 9627 8196 9628 8260
rect 9692 8196 9693 8260
rect 9627 8195 9693 8196
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 6560 8660 7584
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 5472 8660 6496
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 4384 8660 5408
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 3296 8660 4320
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 2208 8660 3232
rect 9630 2685 9690 8195
rect 9814 8125 9874 9555
rect 10805 9280 11125 10304
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 8192 11125 9216
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 9811 8124 9877 8125
rect 9811 8060 9812 8124
rect 9876 8060 9877 8124
rect 9811 8059 9877 8060
rect 10805 7104 11125 8128
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 6016 11125 7040
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 4928 11125 5952
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 3840 11125 4864
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 2752 11125 3776
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 9627 2684 9693 2685
rect 9627 2620 9628 2684
rect 9692 2620 9693 2684
rect 9627 2619 9693 2620
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2128 8660 2144
rect 10805 2128 11125 2688
rect 13270 17440 13590 17456
rect 13270 17376 13278 17440
rect 13342 17376 13358 17440
rect 13422 17376 13438 17440
rect 13502 17376 13518 17440
rect 13582 17376 13590 17440
rect 13270 16352 13590 17376
rect 13270 16288 13278 16352
rect 13342 16288 13358 16352
rect 13422 16288 13438 16352
rect 13502 16288 13518 16352
rect 13582 16288 13590 16352
rect 13270 15264 13590 16288
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 14176 13590 15200
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 13088 13590 14112
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 12000 13590 13024
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 10912 13590 11936
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 9824 13590 10848
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 8736 13590 9760
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 7648 13590 8672
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 6560 13590 7584
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 5472 13590 6496
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 4384 13590 5408
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 3296 13590 4320
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13270 2208 13590 3232
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2128 13590 2144
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608764939
transform -1 0 15824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608764939
transform -1 0 15824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608764939
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608764939
transform 1 0 15364 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_151
timestamp 1608764939
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_154
timestamp 1608764939
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_153
timestamp 1608764939
transform 1 0 15180 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_156
timestamp 1608764939
transform 1 0 15456 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608764939
transform 1 0 14168 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608764939
transform 1 0 13984 0 1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_26_138
timestamp 1608764939
transform 1 0 13800 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_134
timestamp 1608764939
transform 1 0 13432 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764939
transform 1 0 12328 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1608764939
transform 1 0 11040 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1608764939
transform 1 0 12604 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608764939
transform 1 0 12512 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_117
timestamp 1608764939
transform 1 0 11868 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_121
timestamp 1608764939
transform 1 0 12236 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1608764939
transform 1 0 11500 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_121
timestamp 1608764939
transform 1 0 12236 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1608764939
transform 1 0 9752 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1608764939
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1608764939
transform 1 0 10672 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608764939
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608764939
transform 1 0 9660 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_86
timestamp 1608764939
transform 1 0 9016 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_102
timestamp 1608764939
transform 1 0 10488 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_91
timestamp 1608764939
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_98
timestamp 1608764939
transform 1 0 10120 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1608764939
transform 1 0 6900 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1608764939
transform 1 0 8648 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764939
transform 1 0 6992 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1608764939
transform 1 0 8648 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1608764939
transform 1 0 7636 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_80
timestamp 1608764939
transform 1 0 8464 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_67
timestamp 1608764939
transform 1 0 7268 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_80
timestamp 1608764939
transform 1 0 8464 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1608764939
transform 1 0 5336 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1608764939
transform 1 0 5888 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764939
transform 1 0 5336 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608764939
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_45
timestamp 1608764939
transform 1 0 5244 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_62
timestamp 1608764939
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_44
timestamp 1608764939
transform 1 0 5152 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_50
timestamp 1608764939
transform 1 0 5704 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_56
timestamp 1608764939
transform 1 0 6256 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1608764939
transform 1 0 4784 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_39
timestamp 1608764939
transform 1 0 4692 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1608764939
transform 1 0 4324 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608764939
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608764939
transform 1 0 3956 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_32
timestamp 1608764939
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_32
timestamp 1608764939
transform 1 0 4048 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1608764939
transform 1 0 3404 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_25
timestamp 1608764939
transform 1 0 3404 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_23
timestamp 1608764939
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_29
timestamp 1608764939
transform 1 0 3772 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1608764939
transform 1 0 2852 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764939
transform 1 0 2852 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1608764939
transform 1 0 2116 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_9
timestamp 1608764939
transform 1 0 1932 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_15
timestamp 1608764939
transform 1 0 2484 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_9
timestamp 1608764939
transform 1 0 1932 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_17
timestamp 1608764939
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1608764939
transform 1 0 1564 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1608764939
transform 1 0 1564 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608764939
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608764939
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1608764939
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1608764939
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1608764939
transform 1 0 15088 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608764939
transform -1 0 15824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_150
timestamp 1608764939
transform 1 0 14904 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_155
timestamp 1608764939
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764939
transform 1 0 13432 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1608764939
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1608764939
transform 1 0 11684 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1608764939
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608764939
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1608764939
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1608764939
transform 1 0 11960 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764939
transform 1 0 10028 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_95
timestamp 1608764939
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1608764939
transform 1 0 7820 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764939
transform 1 0 8372 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_71
timestamp 1608764939
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_77
timestamp 1608764939
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1608764939
transform 1 0 5152 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1608764939
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1608764939
transform 1 0 5704 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608764939
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_43
timestamp 1608764939
transform 1 0 5060 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_48
timestamp 1608764939
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1608764939
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1608764939
transform 1 0 3404 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1608764939
transform 1 0 3956 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_23
timestamp 1608764939
transform 1 0 3220 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_29
timestamp 1608764939
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_35
timestamp 1608764939
transform 1 0 4324 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1608764939
transform 1 0 2300 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1608764939
transform 1 0 2852 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764939
transform 1 0 1564 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608764939
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1608764939
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1608764939
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_17
timestamp 1608764939
transform 1 0 2668 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608764939
transform -1 0 15824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608764939
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_148
timestamp 1608764939
transform 1 0 14720 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1608764939
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_154
timestamp 1608764939
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1608764939
transform 1 0 13892 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_137
timestamp 1608764939
transform 1 0 13708 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764939
transform 1 0 12236 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_113
timestamp 1608764939
transform 1 0 11500 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1608764939
transform 1 0 9016 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1608764939
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1608764939
transform 1 0 10672 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608764939
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1608764939
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1608764939
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_102
timestamp 1608764939
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1608764939
transform 1 0 6992 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1608764939
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_73
timestamp 1608764939
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1608764939
transform 1 0 6348 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_55
timestamp 1608764939
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_61
timestamp 1608764939
transform 1 0 6716 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764939
transform 1 0 4692 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608764939
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1608764939
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_32
timestamp 1608764939
transform 1 0 4048 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_38
timestamp 1608764939
transform 1 0 4600 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1608764939
transform 1 0 2208 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1608764939
transform 1 0 2944 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764939
transform 1 0 1472 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608764939
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1608764939
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_10
timestamp 1608764939
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_16
timestamp 1608764939
transform 1 0 2576 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608764939
transform -1 0 15824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_154
timestamp 1608764939
transform 1 0 15272 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1608764939
transform 1 0 13432 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1608764939
transform 1 0 14444 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_132
timestamp 1608764939
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_143
timestamp 1608764939
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1608764939
transform 1 0 11132 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1608764939
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608764939
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_107
timestamp 1608764939
transform 1 0 10948 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_118
timestamp 1608764939
transform 1 0 11960 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1608764939
transform 1 0 10120 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_96
timestamp 1608764939
transform 1 0 9936 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1608764939
transform 1 0 6992 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764939
transform 1 0 8464 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1608764939
transform 1 0 7452 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_67
timestamp 1608764939
transform 1 0 7268 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_78
timestamp 1608764939
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1608764939
transform 1 0 5336 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608764939
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608764939
transform 1 0 6348 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_44
timestamp 1608764939
transform 1 0 5152 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_55
timestamp 1608764939
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_60
timestamp 1608764939
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_62
timestamp 1608764939
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1608764939
transform 1 0 4324 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_33
timestamp 1608764939
transform 1 0 4140 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764939
transform 1 0 2668 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1608764939
transform 1 0 1656 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608764939
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1608764939
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_15
timestamp 1608764939
transform 1 0 2484 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608764939
transform -1 0 15824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608764939
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1608764939
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_154
timestamp 1608764939
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608764939
transform 1 0 13800 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_22_129
timestamp 1608764939
transform 1 0 12972 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_137
timestamp 1608764939
transform 1 0 13708 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764939
transform 1 0 11500 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_111
timestamp 1608764939
transform 1 0 11316 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764939
transform 1 0 9844 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608764939
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1608764939
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1608764939
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1608764939
transform 1 0 8556 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1608764939
transform 1 0 7544 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_68
timestamp 1608764939
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_79
timestamp 1608764939
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1608764939
transform 1 0 5796 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_49
timestamp 1608764939
transform 1 0 5612 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_60
timestamp 1608764939
transform 1 0 6624 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764939
transform 1 0 4140 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764939
transform 1 0 3128 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608764939
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_28
timestamp 1608764939
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_32
timestamp 1608764939
transform 1 0 4048 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764939
transform 1 0 1472 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608764939
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1608764939
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_20
timestamp 1608764939
transform 1 0 2944 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608764939
transform 1 0 14720 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608764939
transform -1 0 15824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_146
timestamp 1608764939
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_151
timestamp 1608764939
transform 1 0 14996 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764939
transform 1 0 13064 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_129
timestamp 1608764939
transform 1 0 12972 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1608764939
transform 1 0 11224 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608764939
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_107
timestamp 1608764939
transform 1 0 10948 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_119
timestamp 1608764939
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_123
timestamp 1608764939
transform 1 0 12420 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764939
transform 1 0 9016 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608764939
transform 1 0 10672 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_102
timestamp 1608764939
transform 1 0 10488 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_78
timestamp 1608764939
transform 1 0 8280 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1608764939
transform 1 0 4968 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764939
transform 1 0 6808 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1608764939
transform 1 0 5520 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608764939
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_45
timestamp 1608764939
transform 1 0 5244 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1608764939
transform 1 0 6348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1608764939
transform 1 0 3956 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_29
timestamp 1608764939
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_40
timestamp 1608764939
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1608764939
transform 1 0 2944 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1608764939
transform 1 0 1932 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608764939
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1608764939
transform 1 0 1380 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_18
timestamp 1608764939
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608764939
transform -1 0 15824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608764939
transform -1 0 15824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608764939
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_148
timestamp 1608764939
transform 1 0 14720 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_156
timestamp 1608764939
transform 1 0 15456 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_149
timestamp 1608764939
transform 1 0 14812 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1608764939
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1608764939
transform 1 0 12972 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1608764939
transform 1 0 13984 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1608764939
transform 1 0 13892 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_19_132
timestamp 1608764939
transform 1 0 13248 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_138
timestamp 1608764939
transform 1 0 13800 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_127
timestamp 1608764939
transform 1 0 12788 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1608764939
transform 1 0 13800 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1608764939
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1608764939
transform 1 0 11960 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1608764939
transform 1 0 10856 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608764939
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_115
timestamp 1608764939
transform 1 0 11684 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1608764939
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_116
timestamp 1608764939
transform 1 0 11776 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764939
transform 1 0 10304 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1608764939
transform 1 0 9844 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608764939
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608764939
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_91
timestamp 1608764939
transform 1 0 9476 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_104
timestamp 1608764939
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_86
timestamp 1608764939
transform 1 0 9016 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_93
timestamp 1608764939
transform 1 0 9660 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_99
timestamp 1608764939
transform 1 0 10212 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764939
transform 1 0 8004 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764939
transform 1 0 7544 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608764939
transform 1 0 7268 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_71
timestamp 1608764939
transform 1 0 7636 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_66
timestamp 1608764939
transform 1 0 7176 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1608764939
transform 1 0 5612 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1608764939
transform 1 0 5336 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1608764939
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608764939
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608764939
transform 1 0 6348 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_55
timestamp 1608764939
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1608764939
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_47
timestamp 1608764939
transform 1 0 5428 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_58
timestamp 1608764939
transform 1 0 6440 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764939
transform 1 0 3128 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1608764939
transform 1 0 4600 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608764939
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_38
timestamp 1608764939
transform 1 0 4600 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_26
timestamp 1608764939
transform 1 0 3496 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1608764939
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_32
timestamp 1608764939
transform 1 0 4048 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_20
timestamp 1608764939
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1608764939
transform 1 0 2116 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1608764939
transform 1 0 2668 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_15
timestamp 1608764939
transform 1 0 2484 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764939
transform 1 0 1380 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1608764939
transform 1 0 1656 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608764939
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608764939
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_9
timestamp 1608764939
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1608764939
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608764939
transform -1 0 15824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608764939
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1608764939
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1608764939
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1608764939
transform 1 0 14168 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1608764939
transform 1 0 13156 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_127
timestamp 1608764939
transform 1 0 12788 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_140
timestamp 1608764939
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1608764939
transform 1 0 12512 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764939
transform 1 0 10856 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_122
timestamp 1608764939
transform 1 0 12328 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1608764939
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608764939
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_89
timestamp 1608764939
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_102
timestamp 1608764939
transform 1 0 10488 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1608764939
transform 1 0 8188 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1608764939
transform 1 0 8464 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764939
transform 1 0 5060 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764939
transform 1 0 6716 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_59
timestamp 1608764939
transform 1 0 6532 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1608764939
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608764939
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608764939
transform 1 0 3680 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1608764939
transform 1 0 3404 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_41
timestamp 1608764939
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764939
transform 1 0 1932 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608764939
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1608764939
transform 1 0 1380 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1608764939
transform 1 0 14812 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608764939
transform -1 0 15824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_147
timestamp 1608764939
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1608764939
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00
timestamp 1608764939
transform 1 0 12788 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_139
timestamp 1608764939
transform 1 0 13892 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608764939
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1608764939
transform 1 0 11500 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1608764939
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_123
timestamp 1608764939
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1608764939
transform 1 0 9660 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1608764939
transform 1 0 10672 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_91
timestamp 1608764939
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_102
timestamp 1608764939
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1608764939
transform 1 0 6900 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1608764939
transform 1 0 8648 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1608764939
transform 1 0 7728 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_81
timestamp 1608764939
transform 1 0 8556 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1608764939
transform 1 0 5704 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608764939
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_47
timestamp 1608764939
transform 1 0 5428 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1608764939
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_62
timestamp 1608764939
transform 1 0 6808 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1608764939
transform 1 0 4600 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_35
timestamp 1608764939
transform 1 0 4324 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764939
transform 1 0 2852 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1608764939
transform 1 0 1840 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608764939
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1608764939
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1608764939
transform 1 0 1748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_17
timestamp 1608764939
transform 1 0 2668 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608764939
transform -1 0 15824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608764939
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1608764939
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1608764939
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_131
timestamp 1608764939
transform 1 0 13156 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_143
timestamp 1608764939
transform 1 0 14260 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764939
transform 1 0 11684 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_110
timestamp 1608764939
transform 1 0 11224 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_114
timestamp 1608764939
transform 1 0 11592 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1608764939
transform 1 0 10396 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608764939
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608764939
transform 1 0 10120 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1608764939
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_93
timestamp 1608764939
transform 1 0 9660 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_97
timestamp 1608764939
transform 1 0 10028 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1608764939
transform 1 0 7544 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1608764939
transform 1 0 8556 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_67
timestamp 1608764939
transform 1 0 7268 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_79
timestamp 1608764939
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764939
transform 1 0 5796 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_49
timestamp 1608764939
transform 1 0 5612 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764939
transform 1 0 3036 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1608764939
transform 1 0 4784 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764939
transform 1 0 4048 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608764939
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1608764939
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_38
timestamp 1608764939
transform 1 0 4600 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764939
transform 1 0 1380 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608764939
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_19
timestamp 1608764939
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608764939
transform -1 0 15824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_152
timestamp 1608764939
transform 1 0 15088 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_156
timestamp 1608764939
transform 1 0 15456 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1608764939
transform 1 0 14260 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_141
timestamp 1608764939
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764939
transform 1 0 12604 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608764939
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1608764939
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_123
timestamp 1608764939
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764939
transform 1 0 10672 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1608764939
transform 1 0 9660 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_15_87
timestamp 1608764939
transform 1 0 9108 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_102
timestamp 1608764939
transform 1 0 10488 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1608764939
transform 1 0 7176 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764939
transform 1 0 7636 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_69
timestamp 1608764939
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764939
transform 1 0 5888 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608764939
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_50
timestamp 1608764939
transform 1 0 5704 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_58
timestamp 1608764939
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1608764939
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764939
transform 1 0 4232 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1608764939
transform 1 0 3220 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_21
timestamp 1608764939
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_32
timestamp 1608764939
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764939
transform 1 0 1472 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1608764939
transform 1 0 2208 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608764939
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1608764939
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_10
timestamp 1608764939
transform 1 0 2024 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608764939
transform -1 0 15824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608764939
transform -1 0 15824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608764939
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_155
timestamp 1608764939
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_147
timestamp 1608764939
transform 1 0 14628 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_154
timestamp 1608764939
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1608764939
transform 1 0 14352 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1608764939
transform 1 0 13340 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1608764939
transform 1 0 13432 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1608764939
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_143
timestamp 1608764939
transform 1 0 14260 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_127
timestamp 1608764939
transform 1 0 12788 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_142
timestamp 1608764939
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1608764939
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1608764939
transform 1 0 11960 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1608764939
transform 1 0 11316 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608764939
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1608764939
transform 1 0 10948 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1608764939
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_112
timestamp 1608764939
transform 1 0 11408 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764939
transform 1 0 9936 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1608764939
transform 1 0 9292 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1608764939
transform 1 0 10120 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608764939
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_93
timestamp 1608764939
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1608764939
transform 1 0 7912 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1608764939
transform 1 0 8740 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608764939
transform 1 0 7452 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_13_68
timestamp 1608764939
transform 1 0 7360 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_66
timestamp 1608764939
transform 1 0 7176 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764939
transform 1 0 5704 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1608764939
transform 1 0 5888 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608764939
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608764939
transform 1 0 5428 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_45
timestamp 1608764939
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_50
timestamp 1608764939
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_62
timestamp 1608764939
transform 1 0 6808 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_45
timestamp 1608764939
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_49
timestamp 1608764939
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1608764939
transform 1 0 4416 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1608764939
transform 1 0 4416 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608764939
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_34
timestamp 1608764939
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_28
timestamp 1608764939
transform 1 0 3680 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1608764939
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764939
transform 1 0 2760 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1608764939
transform 1 0 2852 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_16
timestamp 1608764939
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_17
timestamp 1608764939
transform 1 0 2668 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1608764939
transform 1 0 1840 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1608764939
transform 1 0 1748 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608764939
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608764939
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1608764939
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1608764939
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1608764939
transform 1 0 1748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608764939
transform -1 0 15824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608764939
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1608764939
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1608764939
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1608764939
transform 1 0 13432 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_132
timestamp 1608764939
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_143
timestamp 1608764939
transform 1 0 14260 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1608764939
transform 1 0 12420 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_120
timestamp 1608764939
transform 1 0 12144 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764939
transform 1 0 10672 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1608764939
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608764939
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_89
timestamp 1608764939
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_102
timestamp 1608764939
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1608764939
transform 1 0 8464 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_76
timestamp 1608764939
transform 1 0 8096 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764939
transform 1 0 4968 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764939
transform 1 0 6624 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_58
timestamp 1608764939
transform 1 0 6440 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1608764939
transform 1 0 4508 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1608764939
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608764939
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1608764939
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_35
timestamp 1608764939
transform 1 0 4324 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_40
timestamp 1608764939
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764939
transform 1 0 2116 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764939
transform 1 0 1380 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608764939
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_9
timestamp 1608764939
transform 1 0 1932 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608764939
transform -1 0 15824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_155
timestamp 1608764939
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764939
transform 1 0 12788 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_11_143
timestamp 1608764939
transform 1 0 14260 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1608764939
transform 1 0 11592 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608764939
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_112
timestamp 1608764939
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1608764939
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1608764939
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_123
timestamp 1608764939
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764939
transform 1 0 9936 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608764939
transform 1 0 9660 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_90
timestamp 1608764939
transform 1 0 9384 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764939
transform 1 0 6900 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1608764939
transform 1 0 8556 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_79
timestamp 1608764939
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1608764939
transform 1 0 5704 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608764939
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_49
timestamp 1608764939
transform 1 0 5612 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1608764939
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_62
timestamp 1608764939
transform 1 0 6808 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1608764939
transform 1 0 4784 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1608764939
transform 1 0 3772 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_27
timestamp 1608764939
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_38
timestamp 1608764939
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1608764939
transform 1 0 2760 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1608764939
transform 1 0 1748 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608764939
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1608764939
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_16
timestamp 1608764939
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608764939
transform -1 0 15824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608764939
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_147
timestamp 1608764939
transform 1 0 14628 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_10_154
timestamp 1608764939
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1608764939
transform 1 0 12696 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_135
timestamp 1608764939
transform 1 0 13524 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1608764939
transform 1 0 11684 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_113
timestamp 1608764939
transform 1 0 11500 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_124
timestamp 1608764939
transform 1 0 12512 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1608764939
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1608764939
transform 1 0 10672 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608764939
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1608764939
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_102
timestamp 1608764939
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1608764939
transform 1 0 8556 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_71
timestamp 1608764939
transform 1 0 7636 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_79
timestamp 1608764939
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764939
transform 1 0 5152 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1608764939
transform 1 0 6808 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_42
timestamp 1608764939
transform 1 0 4968 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_60
timestamp 1608764939
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1608764939
transform 1 0 4140 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608764939
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1608764939
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_32
timestamp 1608764939
transform 1 0 4048 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1608764939
transform 1 0 2944 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764939
transform 1 0 1472 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764939
transform 1 0 2208 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608764939
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1608764939
transform 1 0 1380 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_10
timestamp 1608764939
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_18
timestamp 1608764939
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608764939
transform -1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_156
timestamp 1608764939
transform 1 0 15456 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_132
timestamp 1608764939
transform 1 0 13248 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_144
timestamp 1608764939
transform 1 0 14352 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1608764939
transform 1 0 11040 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1608764939
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608764939
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_106
timestamp 1608764939
transform 1 0 10856 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_117
timestamp 1608764939
transform 1 0 11868 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1608764939
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1608764939
transform 1 0 10028 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_94
timestamp 1608764939
transform 1 0 9752 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764939
transform 1 0 8280 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608764939
transform 1 0 7820 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_71
timestamp 1608764939
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_76
timestamp 1608764939
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1608764939
transform 1 0 5520 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1608764939
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608764939
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_46
timestamp 1608764939
transform 1 0 5336 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1608764939
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1608764939
transform 1 0 4508 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_35
timestamp 1608764939
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764939
transform 1 0 2852 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1608764939
transform 1 0 1840 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608764939
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1608764939
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1608764939
transform 1 0 1748 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_17
timestamp 1608764939
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608764939
transform -1 0 15824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608764939
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1608764939
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_154
timestamp 1608764939
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1608764939
transform 1 0 12880 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_126
timestamp 1608764939
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_137
timestamp 1608764939
transform 1 0 13708 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764939
transform 1 0 11224 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_8_107
timestamp 1608764939
transform 1 0 10948 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1608764939
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608764939
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608764939
transform 1 0 10672 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_88
timestamp 1608764939
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_102
timestamp 1608764939
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764939
transform 1 0 7728 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_70
timestamp 1608764939
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1608764939
transform 1 0 5980 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1608764939
transform 1 0 6716 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_49
timestamp 1608764939
transform 1 0 5612 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_57
timestamp 1608764939
transform 1 0 6348 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1608764939
transform 1 0 4784 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608764939
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608764939
transform 1 0 4508 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_22
timestamp 1608764939
transform 1 0 3128 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_30
timestamp 1608764939
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 1608764939
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_36
timestamp 1608764939
transform 1 0 4416 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764939
transform 1 0 1656 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608764939
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1608764939
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608764939
transform -1 0 15824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608764939
transform -1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608764939
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1608764939
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1608764939
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_150
timestamp 1608764939
transform 1 0 14904 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_156
timestamp 1608764939
transform 1 0 15456 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l4_in_0_
timestamp 1608764939
transform 1 0 12972 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764939
transform 1 0 14444 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_138
timestamp 1608764939
transform 1 0 13800 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_144
timestamp 1608764939
transform 1 0 14352 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_126
timestamp 1608764939
transform 1 0 12696 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_138
timestamp 1608764939
transform 1 0 13800 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1608764939
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1608764939
transform 1 0 11316 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608764939
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1608764939
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1608764939
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_107
timestamp 1608764939
transform 1 0 10948 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1608764939
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1608764939
transform 1 0 8924 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764939
transform 1 0 9476 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1608764939
transform 1 0 9936 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608764939
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_89
timestamp 1608764939
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_93
timestamp 1608764939
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_89
timestamp 1608764939
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1608764939
transform 1 0 6900 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1608764939
transform 1 0 8372 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1608764939
transform 1 0 7360 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1608764939
transform 1 0 8464 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_66
timestamp 1608764939
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_77
timestamp 1608764939
transform 1 0 8188 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_83
timestamp 1608764939
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_78
timestamp 1608764939
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764939
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764939
transform 1 0 5244 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1608764939
transform 1 0 5704 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608764939
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_61
timestamp 1608764939
transform 1 0 6716 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_46
timestamp 1608764939
transform 1 0 5336 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1608764939
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_41
timestamp 1608764939
transform 1 0 4876 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1608764939
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1608764939
transform 1 0 4508 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608764939
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_33
timestamp 1608764939
transform 1 0 4140 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1608764939
transform 1 0 3404 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1608764939
transform 1 0 3312 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_24
timestamp 1608764939
transform 1 0 3312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1608764939
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_22
timestamp 1608764939
transform 1 0 3128 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764939
transform 1 0 1656 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1608764939
transform 1 0 2116 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764939
transform 1 0 1380 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608764939
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608764939
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_9
timestamp 1608764939
transform 1 0 1932 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_20
timestamp 1608764939
transform 1 0 2944 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1608764939
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608764939
transform -1 0 15824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_150
timestamp 1608764939
transform 1 0 14904 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_156
timestamp 1608764939
transform 1 0 15456 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_3_
timestamp 1608764939
transform 1 0 14076 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_139
timestamp 1608764939
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764939
transform 1 0 12420 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608764939
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1608764939
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1608764939
transform 1 0 9936 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764939
transform 1 0 10672 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_94
timestamp 1608764939
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_100
timestamp 1608764939
transform 1 0 10304 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764939
transform 1 0 8280 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1608764939
transform 1 0 7268 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_65
timestamp 1608764939
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_76
timestamp 1608764939
transform 1 0 8096 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1608764939
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1608764939
transform 1 0 5704 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608764939
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_46
timestamp 1608764939
transform 1 0 5336 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1608764939
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1608764939
transform 1 0 3128 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764939
transform 1 0 3864 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_26
timestamp 1608764939
transform 1 0 3496 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1608764939
transform 1 0 1564 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1608764939
transform 1 0 2116 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608764939
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1608764939
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_9
timestamp 1608764939
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_20
timestamp 1608764939
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608764939
transform -1 0 15824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608764939
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1608764939
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1608764939
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_2_
timestamp 1608764939
transform 1 0 14168 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_140
timestamp 1608764939
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764939
transform 1 0 12512 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_4_115
timestamp 1608764939
transform 1 0 11684 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_123
timestamp 1608764939
transform 1 0 12420 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1608764939
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764939
transform 1 0 10212 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608764939
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1608764939
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_97
timestamp 1608764939
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1608764939
transform 1 0 8556 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1608764939
transform 1 0 7544 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_67
timestamp 1608764939
transform 1 0 7268 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_79
timestamp 1608764939
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1608764939
transform 1 0 5152 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764939
transform 1 0 5796 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_42
timestamp 1608764939
transform 1 0 4968 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_48
timestamp 1608764939
transform 1 0 5520 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1608764939
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1608764939
transform 1 0 4600 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608764939
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_28
timestamp 1608764939
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_36
timestamp 1608764939
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1608764939
transform 1 0 1840 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1608764939
transform 1 0 2852 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608764939
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1608764939
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1608764939
transform 1 0 1748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_17
timestamp 1608764939
transform 1 0 2668 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608764939
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_148
timestamp 1608764939
transform 1 0 14720 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_156
timestamp 1608764939
transform 1 0 15456 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1608764939
transform 1 0 14444 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_1_
timestamp 1608764939
transform 1 0 13432 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_132
timestamp 1608764939
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_143
timestamp 1608764939
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1608764939
transform 1 0 10764 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_0_
timestamp 1608764939
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_0_
timestamp 1608764939
transform 1 0 11316 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608764939
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_109
timestamp 1608764939
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1608764939
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1608764939
transform 1 0 9752 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608764939
transform 1 0 9476 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_89
timestamp 1608764939
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_103
timestamp 1608764939
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764939
transform 1 0 7820 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_3_66
timestamp 1608764939
transform 1 0 7176 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_72
timestamp 1608764939
transform 1 0 7728 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1608764939
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1608764939
transform 1 0 5704 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608764939
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_48
timestamp 1608764939
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1608764939
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1608764939
transform 1 0 4692 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_3_36
timestamp 1608764939
transform 1 0 4416 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764939
transform 1 0 2944 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764939
transform 1 0 1472 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764939
transform 1 0 2208 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608764939
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1608764939
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_10
timestamp 1608764939
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_18
timestamp 1608764939
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608764939
transform -1 0 15824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1608764939
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1608764939
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1608764939
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1608764939
transform 1 0 13432 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_132
timestamp 1608764939
transform 1 0 13248 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_143
timestamp 1608764939
transform 1 0 14260 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_0_
timestamp 1608764939
transform 1 0 12420 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_1_
timestamp 1608764939
transform 1 0 11408 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_2_105
timestamp 1608764939
transform 1 0 10764 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_111
timestamp 1608764939
transform 1 0 11316 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_121
timestamp 1608764939
transform 1 0 12236 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1608764939
transform 1 0 9936 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1608764939
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1608764939
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_93
timestamp 1608764939
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1608764939
transform 1 0 8556 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_2_74
timestamp 1608764939
transform 1 0 7912 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_80
timestamp 1608764939
transform 1 0 8464 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764939
transform 1 0 6440 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_2_51
timestamp 1608764939
transform 1 0 5796 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_57
timestamp 1608764939
transform 1 0 6348 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764939
transform 1 0 4324 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1608764939
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608764939
transform 1 0 3680 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_25
timestamp 1608764939
transform 1 0 3404 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_32
timestamp 1608764939
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1608764939
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764939
transform 1 0 1932 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608764939
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_7
timestamp 1608764939
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608764939
transform -1 0 15824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608764939
transform -1 0 15824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1608764939
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1608764939
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_155
timestamp 1608764939
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1608764939
transform 1 0 14720 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1608764939
transform 1 0 14812 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_146
timestamp 1608764939
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_152
timestamp 1608764939
transform 1 0 15088 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_148
timestamp 1608764939
transform 1 0 14720 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1608764939
transform 1 0 13616 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1608764939
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764939
transform 1 0 12880 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1608764939
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_140
timestamp 1608764939
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_126
timestamp 1608764939
transform 1 0 12696 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_144
timestamp 1608764939
transform 1 0 14352 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_1_
timestamp 1608764939
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1608764939
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1608764939
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1608764939
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1608764939
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_115
timestamp 1608764939
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_121
timestamp 1608764939
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1608764939
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_2_
timestamp 1608764939
transform 1 0 11316 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1608764939
transform 1 0 10856 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_1_108
timestamp 1608764939
transform 1 0 11040 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764939
transform 1 0 9568 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1608764939
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1608764939
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1608764939
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_103
timestamp 1608764939
transform 1 0 10580 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_90
timestamp 1608764939
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1608764939
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764939
transform 1 0 7912 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1608764939
transform 1 0 8648 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1608764939
transform 1 0 7636 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67
timestamp 1608764939
transform 1 0 7268 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80
timestamp 1608764939
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_71
timestamp 1608764939
transform 1 0 7636 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1608764939
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1608764939
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1608764939
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1608764939
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1608764939
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1608764939
transform 1 0 5244 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1608764939
transform 1 0 5704 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1608764939
transform 1 0 5428 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44
timestamp 1608764939
transform 1 0 5152 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_43
timestamp 1608764939
transform 1 0 5060 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_48
timestamp 1608764939
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1608764939
transform 1 0 4232 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1608764939
transform 1 0 4324 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1608764939
transform 1 0 3220 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1608764939
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26
timestamp 1608764939
transform 1 0 3496 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30
timestamp 1608764939
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp 1608764939
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_21
timestamp 1608764939
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_32
timestamp 1608764939
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764939
transform 1 0 2024 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1608764939
transform 1 0 2208 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1608764939
transform 1 0 1472 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764939
transform 1 0 1472 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608764939
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608764939
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3
timestamp 1608764939
transform 1 0 1380 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8
timestamp 1608764939
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3
timestamp 1608764939
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_10
timestamp 1608764939
transform 1 0 2024 0 1 2720
box -38 -48 222 592
<< labels >>
rlabel metal2 s 202 19200 258 20000 4 IO_ISOL_N
port 1 nsew
rlabel metal3 s 0 1368 800 1488 4 ccff_head
port 2 nsew
rlabel metal3 s 16200 1912 17000 2032 4 ccff_tail
port 3 nsew
rlabel metal2 s 8482 0 8538 800 4 chany_bottom_in[0]
port 4 nsew
rlabel metal2 s 12622 0 12678 800 4 chany_bottom_in[10]
port 5 nsew
rlabel metal2 s 12990 0 13046 800 4 chany_bottom_in[11]
port 6 nsew
rlabel metal2 s 13450 0 13506 800 4 chany_bottom_in[12]
port 7 nsew
rlabel metal2 s 13818 0 13874 800 4 chany_bottom_in[13]
port 8 nsew
rlabel metal2 s 14278 0 14334 800 4 chany_bottom_in[14]
port 9 nsew
rlabel metal2 s 14646 0 14702 800 4 chany_bottom_in[15]
port 10 nsew
rlabel metal2 s 15106 0 15162 800 4 chany_bottom_in[16]
port 11 nsew
rlabel metal2 s 15474 0 15530 800 4 chany_bottom_in[17]
port 12 nsew
rlabel metal2 s 15934 0 15990 800 4 chany_bottom_in[18]
port 13 nsew
rlabel metal2 s 16302 0 16358 800 4 chany_bottom_in[19]
port 14 nsew
rlabel metal2 s 8850 0 8906 800 4 chany_bottom_in[1]
port 15 nsew
rlabel metal2 s 9310 0 9366 800 4 chany_bottom_in[2]
port 16 nsew
rlabel metal2 s 9678 0 9734 800 4 chany_bottom_in[3]
port 17 nsew
rlabel metal2 s 10138 0 10194 800 4 chany_bottom_in[4]
port 18 nsew
rlabel metal2 s 10506 0 10562 800 4 chany_bottom_in[5]
port 19 nsew
rlabel metal2 s 10966 0 11022 800 4 chany_bottom_in[6]
port 20 nsew
rlabel metal2 s 11334 0 11390 800 4 chany_bottom_in[7]
port 21 nsew
rlabel metal2 s 11794 0 11850 800 4 chany_bottom_in[8]
port 22 nsew
rlabel metal2 s 12162 0 12218 800 4 chany_bottom_in[9]
port 23 nsew
rlabel metal2 s 202 0 258 800 4 chany_bottom_out[0]
port 24 nsew
rlabel metal2 s 4342 0 4398 800 4 chany_bottom_out[10]
port 25 nsew
rlabel metal2 s 4710 0 4766 800 4 chany_bottom_out[11]
port 26 nsew
rlabel metal2 s 5170 0 5226 800 4 chany_bottom_out[12]
port 27 nsew
rlabel metal2 s 5538 0 5594 800 4 chany_bottom_out[13]
port 28 nsew
rlabel metal2 s 5998 0 6054 800 4 chany_bottom_out[14]
port 29 nsew
rlabel metal2 s 6366 0 6422 800 4 chany_bottom_out[15]
port 30 nsew
rlabel metal2 s 6826 0 6882 800 4 chany_bottom_out[16]
port 31 nsew
rlabel metal2 s 7194 0 7250 800 4 chany_bottom_out[17]
port 32 nsew
rlabel metal2 s 7654 0 7710 800 4 chany_bottom_out[18]
port 33 nsew
rlabel metal2 s 8022 0 8078 800 4 chany_bottom_out[19]
port 34 nsew
rlabel metal2 s 570 0 626 800 4 chany_bottom_out[1]
port 35 nsew
rlabel metal2 s 1030 0 1086 800 4 chany_bottom_out[2]
port 36 nsew
rlabel metal2 s 1398 0 1454 800 4 chany_bottom_out[3]
port 37 nsew
rlabel metal2 s 1858 0 1914 800 4 chany_bottom_out[4]
port 38 nsew
rlabel metal2 s 2226 0 2282 800 4 chany_bottom_out[5]
port 39 nsew
rlabel metal2 s 2686 0 2742 800 4 chany_bottom_out[6]
port 40 nsew
rlabel metal2 s 3054 0 3110 800 4 chany_bottom_out[7]
port 41 nsew
rlabel metal2 s 3514 0 3570 800 4 chany_bottom_out[8]
port 42 nsew
rlabel metal2 s 3882 0 3938 800 4 chany_bottom_out[9]
port 43 nsew
rlabel metal2 s 8666 19200 8722 20000 4 chany_top_in[0]
port 44 nsew
rlabel metal2 s 12714 19200 12770 20000 4 chany_top_in[10]
port 45 nsew
rlabel metal2 s 13082 19200 13138 20000 4 chany_top_in[11]
port 46 nsew
rlabel metal2 s 13542 19200 13598 20000 4 chany_top_in[12]
port 47 nsew
rlabel metal2 s 13910 19200 13966 20000 4 chany_top_in[13]
port 48 nsew
rlabel metal2 s 14370 19200 14426 20000 4 chany_top_in[14]
port 49 nsew
rlabel metal2 s 14738 19200 14794 20000 4 chany_top_in[15]
port 50 nsew
rlabel metal2 s 15106 19200 15162 20000 4 chany_top_in[16]
port 51 nsew
rlabel metal2 s 15566 19200 15622 20000 4 chany_top_in[17]
port 52 nsew
rlabel metal2 s 15934 19200 15990 20000 4 chany_top_in[18]
port 53 nsew
rlabel metal2 s 16394 19200 16450 20000 4 chany_top_in[19]
port 54 nsew
rlabel metal2 s 9034 19200 9090 20000 4 chany_top_in[1]
port 55 nsew
rlabel metal2 s 9494 19200 9550 20000 4 chany_top_in[2]
port 56 nsew
rlabel metal2 s 9862 19200 9918 20000 4 chany_top_in[3]
port 57 nsew
rlabel metal2 s 10322 19200 10378 20000 4 chany_top_in[4]
port 58 nsew
rlabel metal2 s 10690 19200 10746 20000 4 chany_top_in[5]
port 59 nsew
rlabel metal2 s 11058 19200 11114 20000 4 chany_top_in[6]
port 60 nsew
rlabel metal2 s 11518 19200 11574 20000 4 chany_top_in[7]
port 61 nsew
rlabel metal2 s 11886 19200 11942 20000 4 chany_top_in[8]
port 62 nsew
rlabel metal2 s 12346 19200 12402 20000 4 chany_top_in[9]
port 63 nsew
rlabel metal2 s 570 19200 626 20000 4 chany_top_out[0]
port 64 nsew
rlabel metal2 s 4618 19200 4674 20000 4 chany_top_out[10]
port 65 nsew
rlabel metal2 s 4986 19200 5042 20000 4 chany_top_out[11]
port 66 nsew
rlabel metal2 s 5446 19200 5502 20000 4 chany_top_out[12]
port 67 nsew
rlabel metal2 s 5814 19200 5870 20000 4 chany_top_out[13]
port 68 nsew
rlabel metal2 s 6274 19200 6330 20000 4 chany_top_out[14]
port 69 nsew
rlabel metal2 s 6642 19200 6698 20000 4 chany_top_out[15]
port 70 nsew
rlabel metal2 s 7010 19200 7066 20000 4 chany_top_out[16]
port 71 nsew
rlabel metal2 s 7470 19200 7526 20000 4 chany_top_out[17]
port 72 nsew
rlabel metal2 s 7838 19200 7894 20000 4 chany_top_out[18]
port 73 nsew
rlabel metal2 s 8298 19200 8354 20000 4 chany_top_out[19]
port 74 nsew
rlabel metal2 s 938 19200 994 20000 4 chany_top_out[1]
port 75 nsew
rlabel metal2 s 1398 19200 1454 20000 4 chany_top_out[2]
port 76 nsew
rlabel metal2 s 1766 19200 1822 20000 4 chany_top_out[3]
port 77 nsew
rlabel metal2 s 2226 19200 2282 20000 4 chany_top_out[4]
port 78 nsew
rlabel metal2 s 2594 19200 2650 20000 4 chany_top_out[5]
port 79 nsew
rlabel metal2 s 2962 19200 3018 20000 4 chany_top_out[6]
port 80 nsew
rlabel metal2 s 3422 19200 3478 20000 4 chany_top_out[7]
port 81 nsew
rlabel metal2 s 3790 19200 3846 20000 4 chany_top_out[8]
port 82 nsew
rlabel metal2 s 4250 19200 4306 20000 4 chany_top_out[9]
port 83 nsew
rlabel metal3 s 16200 9800 17000 9920 4 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 84 nsew
rlabel metal3 s 16200 13880 17000 14000 4 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 85 nsew
rlabel metal3 s 16200 17824 17000 17944 4 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 86 nsew
rlabel metal3 s 0 3272 800 3392 4 left_grid_pin_16_
port 87 nsew
rlabel metal3 s 0 4224 800 4344 4 left_grid_pin_17_
port 88 nsew
rlabel metal3 s 0 5176 800 5296 4 left_grid_pin_18_
port 89 nsew
rlabel metal3 s 0 6128 800 6248 4 left_grid_pin_19_
port 90 nsew
rlabel metal3 s 0 7080 800 7200 4 left_grid_pin_20_
port 91 nsew
rlabel metal3 s 0 8032 800 8152 4 left_grid_pin_21_
port 92 nsew
rlabel metal3 s 0 8984 800 9104 4 left_grid_pin_22_
port 93 nsew
rlabel metal3 s 0 9936 800 10056 4 left_grid_pin_23_
port 94 nsew
rlabel metal3 s 0 10888 800 11008 4 left_grid_pin_24_
port 95 nsew
rlabel metal3 s 0 11840 800 11960 4 left_grid_pin_25_
port 96 nsew
rlabel metal3 s 0 12792 800 12912 4 left_grid_pin_26_
port 97 nsew
rlabel metal3 s 0 13744 800 13864 4 left_grid_pin_27_
port 98 nsew
rlabel metal3 s 0 14696 800 14816 4 left_grid_pin_28_
port 99 nsew
rlabel metal3 s 0 15648 800 15768 4 left_grid_pin_29_
port 100 nsew
rlabel metal3 s 0 16600 800 16720 4 left_grid_pin_30_
port 101 nsew
rlabel metal3 s 0 17552 800 17672 4 left_grid_pin_31_
port 102 nsew
rlabel metal3 s 0 18504 800 18624 4 left_width_0_height_0__pin_0_
port 103 nsew
rlabel metal3 s 0 416 800 536 4 left_width_0_height_0__pin_1_lower
port 104 nsew
rlabel metal3 s 0 19456 800 19576 4 left_width_0_height_0__pin_1_upper
port 105 nsew
rlabel metal2 s 16762 19200 16818 20000 4 prog_clk_0_N_out
port 106 nsew
rlabel metal2 s 16762 0 16818 800 4 prog_clk_0_S_out
port 107 nsew
rlabel metal3 s 0 2320 800 2440 4 prog_clk_0_W_in
port 108 nsew
rlabel metal3 s 16200 5856 17000 5976 4 right_grid_pin_0_
port 109 nsew
rlabel metal4 s 3409 2128 3729 17456 4 VPWR
port 110 nsew
rlabel metal4 s 5875 2128 6195 17456 4 VGND
port 111 nsew
<< properties >>
string FIXED_BBOX 0 0 17000 20000
string GDS_FILE /ef/openfpga/openlane/runs/cby_2__1_/results/magic/cby_2__1_.gds
string GDS_END 989412
string GDS_START 98316
<< end >>
