* NGSPICE file created from cbx_1__2_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxbp_1 abstract view
.subckt sky130_fd_sc_hd__dfxbp_1 D Q Q_N CLK VGND VNB VPB VPWR
.ends

.subckt cbx_1__2_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11]
+ chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16]
+ chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2]
+ chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7]
+ chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11]
+ chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16]
+ chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chanx_left_out[9] chanx_right_in[0] chanx_right_in[10] chanx_right_in[11]
+ chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16]
+ chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11]
+ chanx_right_out[12] chanx_right_out[13] chanx_right_out[14] chanx_right_out[15]
+ chanx_right_out[16] chanx_right_out[17] chanx_right_out[18] chanx_right_out[19]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9] prog_clk
+ top_grid_pin_0_ VPWR VGND
XFILLER_22_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0__S mux_bottom_ipin_0.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__04__A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12__A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07__A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_29_ chanx_right_in[7] chanx_left_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_4_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_0.mux_l4_in_0_/X top_grid_pin_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_3_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20__A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15__A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23__A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28_ chanx_right_in[8] chanx_left_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18__A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__31__A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__26__A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_1__S mux_bottom_ipin_0.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_27_ chanx_right_in[9] chanx_left_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__34__A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__29__A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__37__A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_26_ chanx_right_in[10] chanx_left_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A0 mux_bottom_ipin_0.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09_ chanx_left_in[7] chanx_right_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25_ chanx_right_in[11] chanx_left_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A1 mux_bottom_ipin_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08_ chanx_left_in[8] chanx_right_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_41_ chanx_left_in[15] chanx_right_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_14_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24_ chanx_right_in[12] chanx_left_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07_ chanx_left_in[9] chanx_right_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_25_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_40_ chanx_left_in[16] chanx_right_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23_ chanx_right_in[13] chanx_left_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A0 _01_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06_ chanx_left_in[10] chanx_right_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22_ chanx_right_in[14] chanx_left_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1 chanx_right_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05_ chanx_left_in[11] chanx_right_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_0.mux_l4_in_0__S ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_ipin_0.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21_ chanx_right_in[15] chanx_left_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_04_ chanx_left_in[12] chanx_right_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20_ chanx_right_in[16] chanx_left_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_03_ chanx_left_in[13] chanx_right_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_35_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_02_ chanx_left_in[14] chanx_right_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__02__A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1__S mux_bottom_ipin_0.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_01_ _01_/HI _01_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_2_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10__A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05__A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13__A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__08__A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21__A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16__A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24__A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19__A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__32__A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__27__A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__40__A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_2__S mux_bottom_ipin_0.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__35__A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__38__A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_0.mux_l2_in_3_ _01_/HI chanx_right_in[16] mux_bottom_ipin_0.mux_l2_in_2_/S
+ mux_bottom_ipin_0.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_ipin_0.mux_l4_in_0_ mux_bottom_ipin_0.mux_l3_in_1_/X mux_bottom_ipin_0.mux_l3_in_0_/X
+ ccff_tail mux_bottom_ipin_0.mux_l4_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_0.mux_l3_in_1_ mux_bottom_ipin_0.mux_l2_in_3_/X mux_bottom_ipin_0.mux_l2_in_2_/X
+ mux_bottom_ipin_0.mux_l3_in_1_/S mux_bottom_ipin_0.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_ipin_0.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_bottom_ipin_0.mux_l2_in_2_/S
+ mux_bottom_ipin_0.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_39_ chanx_left_in[17] chanx_right_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l3_in_0__S mux_bottom_ipin_0.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_ipin_0.mux_l3_in_0_ mux_bottom_ipin_0.mux_l2_in_1_/X mux_bottom_ipin_0.mux_l2_in_0_/X
+ mux_bottom_ipin_0.mux_l3_in_1_/S mux_bottom_ipin_0.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_0.mux_l2_in_1_ chanx_left_in[10] mux_bottom_ipin_0.mux_l1_in_2_/X
+ mux_bottom_ipin_0.mux_l2_in_2_/S mux_bottom_ipin_0.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A0 mux_bottom_ipin_0.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_38_ chanx_left_in[18] chanx_right_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_0.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_bottom_ipin_0.mux_l1_in_2_/S
+ mux_bottom_ipin_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A0 mux_bottom_ipin_0.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1 chanx_right_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_0.mux_l2_in_0_ mux_bottom_ipin_0.mux_l1_in_1_/X mux_bottom_ipin_0.mux_l1_in_0_/X
+ mux_bottom_ipin_0.mux_l2_in_2_/S mux_bottom_ipin_0.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A1 mux_bottom_ipin_0.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_37_ chanx_left_in[19] chanx_right_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_0.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_bottom_ipin_0.mux_l1_in_2_/S
+ mux_bottom_ipin_0.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A1 mux_bottom_ipin_0.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D ccff_head VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36_ chanx_right_in[0] chanx_left_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_9_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_0.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_0.mux_l1_in_2_/S
+ mux_bottom_ipin_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19_ chanx_right_in[17] chanx_left_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D mux_bottom_ipin_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_35_ chanx_right_in[1] chanx_left_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0__A mux_bottom_ipin_0.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18_ chanx_right_in[18] chanx_left_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_25_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_34_ chanx_right_in[2] chanx_left_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_ mux_bottom_ipin_0.mux_l3_in_1_/S ccff_tail
+ mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_22_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17_ chanx_right_in[19] chanx_left_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33_ chanx_right_in[3] chanx_left_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_ipin_0.mux_l2_in_2_/S mux_bottom_ipin_0.mux_l3_in_1_/S
+ mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16_ chanx_left_in[0] chanx_right_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__03__A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_ipin_0.mux_l1_in_2_/S mux_bottom_ipin_0.mux_l2_in_2_/S
+ mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_ipin_0.mux_l1_in_2__S mux_bottom_ipin_0.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_32_ chanx_right_in[4] chanx_left_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_13_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11__A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15_ chanx_left_in[1] chanx_right_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06__A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14__A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_ ccff_head mux_bottom_ipin_0.mux_l1_in_2_/S
+ mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA__09__A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31_ chanx_right_in[5] chanx_left_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_9_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14_ chanx_left_in[2] chanx_right_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22__A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17__A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__30__A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25__A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_30_ chanx_right_in[6] chanx_left_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_9_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13_ chanx_left_in[3] chanx_right_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_33_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0__S mux_bottom_ipin_0.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__33__A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__28__A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__41__A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_3__S mux_bottom_ipin_0.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__36__A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12_ chanx_left_in[4] chanx_right_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__39__A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11_ chanx_left_in[5] chanx_right_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A0 mux_bottom_ipin_0.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10_ chanx_left_in[6] chanx_right_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_0.mux_l3_in_1__S mux_bottom_ipin_0.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A1 mux_bottom_ipin_0.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A1 mux_bottom_ipin_0.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
.ends

