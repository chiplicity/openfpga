magic
tech EFS8A
magscale 1 2
timestamp 1602874135
<< locali >>
rect 4445 25347 4479 25449
rect 2881 25313 3042 25347
rect 4445 25313 4606 25347
rect 2881 25143 2915 25313
rect 15243 23137 15370 23171
rect 10051 22185 10057 22219
rect 10051 22117 10085 22185
rect 6595 22049 6630 22083
rect 17233 22049 17394 22083
rect 17233 21879 17267 22049
rect 9959 21335 9993 21403
rect 9959 21301 9965 21335
rect 15295 20247 15329 20315
rect 16773 17595 16807 17833
rect 13823 16745 13829 16779
rect 13823 16677 13857 16745
rect 17049 16031 17083 16133
rect 18383 15589 18429 15623
rect 16899 15521 16934 15555
rect 9499 13719 9533 13787
rect 9499 13685 9505 13719
rect 12535 13481 12541 13515
rect 12535 13413 12569 13481
rect 8855 12631 8889 12699
rect 8855 12597 8861 12631
rect 7935 11305 7941 11339
rect 10787 11305 10793 11339
rect 7935 11237 7969 11305
rect 10787 11237 10821 11305
rect 4813 10081 4974 10115
rect 4813 9911 4847 10081
rect 3387 9673 3525 9707
rect 16899 8993 16934 9027
rect 1547 8585 1685 8619
rect 12351 6953 12357 6987
rect 15663 6953 15669 6987
rect 12351 6885 12385 6953
rect 15663 6885 15697 6953
rect 15571 5015 15605 5083
rect 15571 4981 15577 5015
rect 12351 4777 12357 4811
rect 15663 4777 15669 4811
rect 12351 4709 12385 4777
rect 15663 4709 15697 4777
rect 5871 3961 6009 3995
rect 7757 2975 7791 3145
rect 7251 2601 7389 2635
<< viali >>
rect 4445 25449 4479 25483
rect 1476 25313 1510 25347
rect 5892 25313 5926 25347
rect 7389 25313 7423 25347
rect 8712 25313 8746 25347
rect 11564 25313 11598 25347
rect 13252 25313 13286 25347
rect 10057 25245 10091 25279
rect 7941 25177 7975 25211
rect 1547 25109 1581 25143
rect 2881 25109 2915 25143
rect 3111 25109 3145 25143
rect 4675 25109 4709 25143
rect 4997 25109 5031 25143
rect 5963 25109 5997 25143
rect 7205 25109 7239 25143
rect 8815 25109 8849 25143
rect 11667 25109 11701 25143
rect 13323 25109 13357 25143
rect 2053 24905 2087 24939
rect 4537 24905 4571 24939
rect 5917 24905 5951 24939
rect 11805 24905 11839 24939
rect 2421 24837 2455 24871
rect 13277 24837 13311 24871
rect 4721 24769 4755 24803
rect 4997 24769 5031 24803
rect 7205 24769 7239 24803
rect 7573 24769 7607 24803
rect 1409 24701 1443 24735
rect 3316 24701 3350 24735
rect 3801 24701 3835 24735
rect 8585 24701 8619 24735
rect 8769 24701 8803 24735
rect 10241 24701 10275 24735
rect 10793 24701 10827 24735
rect 11396 24701 11430 24735
rect 12173 24701 12207 24735
rect 12516 24701 12550 24735
rect 13001 24701 13035 24735
rect 13553 24701 13587 24735
rect 3065 24633 3099 24667
rect 4169 24633 4203 24667
rect 4813 24633 4847 24667
rect 7297 24633 7331 24667
rect 8677 24633 8711 24667
rect 11483 24633 11517 24667
rect 1593 24565 1627 24599
rect 3387 24565 3421 24599
rect 6285 24565 6319 24599
rect 6653 24565 6687 24599
rect 8217 24565 8251 24599
rect 10425 24565 10459 24599
rect 12587 24565 12621 24599
rect 13737 24565 13771 24599
rect 14105 24565 14139 24599
rect 1593 24361 1627 24395
rect 14289 24361 14323 24395
rect 21741 24361 21775 24395
rect 4721 24293 4755 24327
rect 6929 24293 6963 24327
rect 7021 24293 7055 24327
rect 7573 24293 7607 24327
rect 1409 24225 1443 24259
rect 2580 24225 2614 24259
rect 10701 24225 10735 24259
rect 11688 24225 11722 24259
rect 13645 24225 13679 24259
rect 21557 24225 21591 24259
rect 4629 24157 4663 24191
rect 7941 24157 7975 24191
rect 8401 24157 8435 24191
rect 10057 24157 10091 24191
rect 13829 24157 13863 24191
rect 14565 24157 14599 24191
rect 5181 24089 5215 24123
rect 2651 24021 2685 24055
rect 11759 24021 11793 24055
rect 1685 23817 1719 23851
rect 2237 23817 2271 23851
rect 2513 23817 2547 23851
rect 5181 23817 5215 23851
rect 6653 23817 6687 23851
rect 7113 23817 7147 23851
rect 9689 23817 9723 23851
rect 10057 23817 10091 23851
rect 11161 23817 11195 23851
rect 11713 23817 11747 23851
rect 13645 23817 13679 23851
rect 14105 23817 14139 23851
rect 19349 23817 19383 23851
rect 21557 23817 21591 23851
rect 24777 23817 24811 23851
rect 2973 23749 3007 23783
rect 4813 23749 4847 23783
rect 5549 23749 5583 23783
rect 14289 23749 14323 23783
rect 20453 23749 20487 23783
rect 3709 23681 3743 23715
rect 4261 23681 4295 23715
rect 5733 23681 5767 23715
rect 7665 23681 7699 23715
rect 10241 23681 10275 23715
rect 10701 23681 10735 23715
rect 16221 23681 16255 23715
rect 22293 23681 22327 23715
rect 2329 23613 2363 23647
rect 9204 23613 9238 23647
rect 12265 23613 12299 23647
rect 12725 23613 12759 23647
rect 14197 23613 14231 23647
rect 14473 23613 14507 23647
rect 15796 23613 15830 23647
rect 19165 23613 19199 23647
rect 19717 23613 19751 23647
rect 20269 23613 20303 23647
rect 20821 23613 20855 23647
rect 21373 23613 21407 23647
rect 21925 23613 21959 23647
rect 24593 23613 24627 23647
rect 25145 23613 25179 23647
rect 4353 23545 4387 23579
rect 7481 23545 7515 23579
rect 7757 23545 7791 23579
rect 8309 23545 8343 23579
rect 10333 23545 10367 23579
rect 15899 23545 15933 23579
rect 4077 23477 4111 23511
rect 9275 23477 9309 23511
rect 12909 23477 12943 23511
rect 14657 23477 14691 23511
rect 10149 23273 10183 23307
rect 13001 23273 13035 23307
rect 3157 23205 3191 23239
rect 4813 23205 4847 23239
rect 7757 23205 7791 23239
rect 10517 23205 10551 23239
rect 12081 23205 12115 23239
rect 3065 23137 3099 23171
rect 6628 23137 6662 23171
rect 14105 23137 14139 23171
rect 15209 23137 15243 23171
rect 1409 23069 1443 23103
rect 4721 23069 4755 23103
rect 4997 23069 5031 23103
rect 7665 23069 7699 23103
rect 8033 23069 8067 23103
rect 9505 23069 9539 23103
rect 10425 23069 10459 23103
rect 10701 23069 10735 23103
rect 11989 23069 12023 23103
rect 12265 23069 12299 23103
rect 13461 23069 13495 23103
rect 15439 23001 15473 23035
rect 4537 22933 4571 22967
rect 6699 22933 6733 22967
rect 14473 22933 14507 22967
rect 2513 22729 2547 22763
rect 3617 22729 3651 22763
rect 3847 22729 3881 22763
rect 6285 22729 6319 22763
rect 7757 22729 7791 22763
rect 8125 22729 8159 22763
rect 9781 22729 9815 22763
rect 11529 22729 11563 22763
rect 12265 22729 12299 22763
rect 13737 22729 13771 22763
rect 14105 22729 14139 22763
rect 22477 22729 22511 22763
rect 5641 22661 5675 22695
rect 12725 22661 12759 22695
rect 15945 22661 15979 22695
rect 10977 22593 11011 22627
rect 14657 22593 14691 22627
rect 1409 22525 1443 22559
rect 1961 22525 1995 22559
rect 2697 22525 2731 22559
rect 3744 22525 3778 22559
rect 4721 22525 4755 22559
rect 6837 22525 6871 22559
rect 8585 22525 8619 22559
rect 9321 22525 9355 22559
rect 12633 22525 12667 22559
rect 12909 22525 12943 22559
rect 14197 22525 14231 22559
rect 14289 22525 14323 22559
rect 14473 22525 14507 22559
rect 15761 22525 15795 22559
rect 16808 22525 16842 22559
rect 17233 22525 17267 22559
rect 22293 22525 22327 22559
rect 22845 22525 22879 22559
rect 4629 22457 4663 22491
rect 5083 22457 5117 22491
rect 6653 22457 6687 22491
rect 7199 22457 7233 22491
rect 9413 22457 9447 22491
rect 10057 22457 10091 22491
rect 10333 22457 10367 22491
rect 10425 22457 10459 22491
rect 11897 22457 11931 22491
rect 13369 22457 13403 22491
rect 16221 22457 16255 22491
rect 1593 22389 1627 22423
rect 2881 22389 2915 22423
rect 3249 22389 3283 22423
rect 4261 22389 4295 22423
rect 15301 22389 15335 22423
rect 16911 22389 16945 22423
rect 1593 22185 1627 22219
rect 5457 22185 5491 22219
rect 6699 22185 6733 22219
rect 7481 22185 7515 22219
rect 8493 22185 8527 22219
rect 10057 22185 10091 22219
rect 10977 22185 11011 22219
rect 14657 22185 14691 22219
rect 17463 22185 17497 22219
rect 4858 22117 4892 22151
rect 7935 22117 7969 22151
rect 12081 22117 12115 22151
rect 15485 22117 15519 22151
rect 1409 22049 1443 22083
rect 6561 22049 6595 22083
rect 11529 22049 11563 22083
rect 12633 22049 12667 22083
rect 12725 22049 12759 22083
rect 12909 22049 12943 22083
rect 14264 22049 14298 22083
rect 2513 21981 2547 22015
rect 4537 21981 4571 22015
rect 7573 21981 7607 22015
rect 9689 21981 9723 22015
rect 13369 21981 13403 22015
rect 13737 21981 13771 22015
rect 15393 21981 15427 22015
rect 15853 21981 15887 22015
rect 10609 21913 10643 21947
rect 2053 21845 2087 21879
rect 3249 21845 3283 21879
rect 4445 21845 4479 21879
rect 7021 21845 7055 21879
rect 9505 21845 9539 21879
rect 11713 21845 11747 21879
rect 14105 21845 14139 21879
rect 14335 21845 14369 21879
rect 17233 21845 17267 21879
rect 2513 21641 2547 21675
rect 4537 21641 4571 21675
rect 4997 21641 5031 21675
rect 8493 21641 8527 21675
rect 10517 21641 10551 21675
rect 12771 21641 12805 21675
rect 14657 21641 14691 21675
rect 15117 21641 15151 21675
rect 16221 21641 16255 21675
rect 24133 21641 24167 21675
rect 9505 21573 9539 21607
rect 10885 21573 10919 21607
rect 1501 21505 1535 21539
rect 13461 21505 13495 21539
rect 13737 21505 13771 21539
rect 15301 21505 15335 21539
rect 16589 21505 16623 21539
rect 4169 21437 4203 21471
rect 4813 21437 4847 21471
rect 7573 21437 7607 21471
rect 8585 21437 8619 21471
rect 9045 21437 9079 21471
rect 9597 21437 9631 21471
rect 11345 21437 11379 21471
rect 11805 21437 11839 21471
rect 12668 21437 12702 21471
rect 13093 21437 13127 21471
rect 16773 21437 16807 21471
rect 17233 21437 17267 21471
rect 23949 21437 23983 21471
rect 24501 21437 24535 21471
rect 1593 21369 1627 21403
rect 2145 21369 2179 21403
rect 3249 21369 3283 21403
rect 3341 21369 3375 21403
rect 3893 21369 3927 21403
rect 5825 21369 5859 21403
rect 8125 21369 8159 21403
rect 12173 21369 12207 21403
rect 13829 21369 13863 21403
rect 14381 21369 14415 21403
rect 15393 21369 15427 21403
rect 15945 21369 15979 21403
rect 17601 21369 17635 21403
rect 3065 21301 3099 21335
rect 6561 21301 6595 21335
rect 7113 21301 7147 21335
rect 7481 21301 7515 21335
rect 7757 21301 7791 21335
rect 8769 21301 8803 21335
rect 9965 21301 9999 21335
rect 11161 21301 11195 21335
rect 11529 21301 11563 21335
rect 16957 21301 16991 21335
rect 3801 21097 3835 21131
rect 5089 21097 5123 21131
rect 6101 21097 6135 21131
rect 6929 21097 6963 21131
rect 9781 21097 9815 21131
rect 13001 21097 13035 21131
rect 17463 21097 17497 21131
rect 2421 21029 2455 21063
rect 2973 21029 3007 21063
rect 4261 21029 4295 21063
rect 9505 21029 9539 21063
rect 13369 21029 13403 21063
rect 13829 21029 13863 21063
rect 15945 21029 15979 21063
rect 6653 20961 6687 20995
rect 7389 20961 7423 20995
rect 7665 20961 7699 20995
rect 8033 20961 8067 20995
rect 9689 20961 9723 20995
rect 10333 20961 10367 20995
rect 10517 20961 10551 20995
rect 10885 20961 10919 20995
rect 12081 20961 12115 20995
rect 17392 20961 17426 20995
rect 2145 20893 2179 20927
rect 2329 20893 2363 20927
rect 4169 20893 4203 20927
rect 4445 20893 4479 20927
rect 5641 20893 5675 20927
rect 11437 20893 11471 20927
rect 11989 20893 12023 20927
rect 13737 20893 13771 20927
rect 14381 20893 14415 20927
rect 15853 20893 15887 20927
rect 16405 20825 16439 20859
rect 1593 20757 1627 20791
rect 3249 20757 3283 20791
rect 6561 20757 6595 20791
rect 9045 20757 9079 20791
rect 15485 20757 15519 20791
rect 1547 20553 1581 20587
rect 12909 20553 12943 20587
rect 14841 20553 14875 20587
rect 15853 20553 15887 20587
rect 16129 20553 16163 20587
rect 16497 20553 16531 20587
rect 1961 20485 1995 20519
rect 3341 20485 3375 20519
rect 9229 20485 9263 20519
rect 18245 20485 18279 20519
rect 3985 20417 4019 20451
rect 4261 20417 4295 20451
rect 7297 20417 7331 20451
rect 11161 20417 11195 20451
rect 14105 20417 14139 20451
rect 1476 20349 1510 20383
rect 2421 20349 2455 20383
rect 4445 20349 4479 20383
rect 4905 20349 4939 20383
rect 5457 20349 5491 20383
rect 5641 20349 5675 20383
rect 7389 20349 7423 20383
rect 7849 20349 7883 20383
rect 8217 20349 8251 20383
rect 8769 20349 8803 20383
rect 9689 20349 9723 20383
rect 10425 20349 10459 20383
rect 10517 20349 10551 20383
rect 11069 20349 11103 20383
rect 14933 20349 14967 20383
rect 16716 20349 16750 20383
rect 17141 20349 17175 20383
rect 18061 20349 18095 20383
rect 19108 20349 19142 20383
rect 19533 20349 19567 20383
rect 2329 20281 2363 20315
rect 2783 20281 2817 20315
rect 6285 20281 6319 20315
rect 11437 20281 11471 20315
rect 13461 20281 13495 20315
rect 13553 20281 13587 20315
rect 4537 20213 4571 20247
rect 6653 20213 6687 20247
rect 7481 20213 7515 20247
rect 9597 20213 9631 20247
rect 12081 20213 12115 20247
rect 13277 20213 13311 20247
rect 14381 20213 14415 20247
rect 15295 20213 15329 20247
rect 16819 20213 16853 20247
rect 17509 20213 17543 20247
rect 18521 20213 18555 20247
rect 19211 20213 19245 20247
rect 6285 20009 6319 20043
rect 8309 20009 8343 20043
rect 11805 20009 11839 20043
rect 12541 20009 12575 20043
rect 14197 20009 14231 20043
rect 1593 19941 1627 19975
rect 4077 19941 4111 19975
rect 16405 19941 16439 19975
rect 2237 19873 2271 19907
rect 3893 19873 3927 19907
rect 4169 19873 4203 19907
rect 5733 19873 5767 19907
rect 6469 19873 6503 19907
rect 6837 19873 6871 19907
rect 7113 19873 7147 19907
rect 7573 19873 7607 19907
rect 8585 19873 8619 19907
rect 9965 19873 9999 19907
rect 10241 19873 10275 19907
rect 11621 19873 11655 19907
rect 13093 19873 13127 19907
rect 13369 19873 13403 19907
rect 17785 19873 17819 19907
rect 18797 19873 18831 19907
rect 9137 19805 9171 19839
rect 10701 19805 10735 19839
rect 13737 19805 13771 19839
rect 16313 19805 16347 19839
rect 10057 19737 10091 19771
rect 13185 19737 13219 19771
rect 16865 19737 16899 19771
rect 2697 19669 2731 19703
rect 2973 19669 3007 19703
rect 3433 19669 3467 19703
rect 5181 19669 5215 19703
rect 6009 19669 6043 19703
rect 7941 19669 7975 19703
rect 8769 19669 8803 19703
rect 9505 19669 9539 19703
rect 10977 19669 11011 19703
rect 11437 19669 11471 19703
rect 15025 19669 15059 19703
rect 15577 19669 15611 19703
rect 17969 19669 18003 19703
rect 18981 19669 19015 19703
rect 2421 19465 2455 19499
rect 2881 19465 2915 19499
rect 3985 19465 4019 19499
rect 4261 19465 4295 19499
rect 5917 19465 5951 19499
rect 10701 19465 10735 19499
rect 11805 19465 11839 19499
rect 13461 19465 13495 19499
rect 16405 19465 16439 19499
rect 16681 19465 16715 19499
rect 17509 19465 17543 19499
rect 6653 19397 6687 19431
rect 10885 19397 10919 19431
rect 17049 19397 17083 19431
rect 3065 19329 3099 19363
rect 9965 19329 9999 19363
rect 2053 19261 2087 19295
rect 4813 19261 4847 19295
rect 6285 19261 6319 19295
rect 7113 19261 7147 19295
rect 7389 19261 7423 19295
rect 7665 19261 7699 19295
rect 8217 19261 8251 19295
rect 9321 19261 9355 19295
rect 10793 19261 10827 19295
rect 11069 19261 11103 19295
rect 12173 19261 12207 19295
rect 12449 19261 12483 19295
rect 12541 19261 12575 19295
rect 12725 19261 12759 19295
rect 13185 19261 13219 19295
rect 14013 19261 14047 19295
rect 14841 19261 14875 19295
rect 15485 19261 15519 19295
rect 18061 19261 18095 19295
rect 18521 19261 18555 19295
rect 19073 19261 19107 19295
rect 3386 19193 3420 19227
rect 9045 19193 9079 19227
rect 11529 19193 11563 19227
rect 14565 19193 14599 19227
rect 15806 19193 15840 19227
rect 1685 19125 1719 19159
rect 4629 19125 4663 19159
rect 4997 19125 5031 19159
rect 5549 19125 5583 19159
rect 6929 19125 6963 19159
rect 8585 19125 8619 19159
rect 10241 19125 10275 19159
rect 13829 19125 13863 19159
rect 14197 19125 14231 19159
rect 15301 19125 15335 19159
rect 17785 19125 17819 19159
rect 18153 19125 18187 19159
rect 1593 18921 1627 18955
rect 3157 18921 3191 18955
rect 4215 18921 4249 18955
rect 5181 18921 5215 18955
rect 7205 18921 7239 18955
rect 16957 18921 16991 18955
rect 18153 18921 18187 18955
rect 2237 18853 2271 18887
rect 2789 18853 2823 18887
rect 4905 18853 4939 18887
rect 7573 18853 7607 18887
rect 8769 18853 8803 18887
rect 10793 18853 10827 18887
rect 15485 18853 15519 18887
rect 16037 18853 16071 18887
rect 4144 18785 4178 18819
rect 5089 18785 5123 18819
rect 5549 18785 5583 18819
rect 6009 18785 6043 18819
rect 6377 18785 6411 18819
rect 8217 18785 8251 18819
rect 9781 18785 9815 18819
rect 9873 18785 9907 18819
rect 10057 18785 10091 18819
rect 10517 18785 10551 18819
rect 11345 18785 11379 18819
rect 11621 18785 11655 18819
rect 13277 18785 13311 18819
rect 13645 18785 13679 18819
rect 17141 18785 17175 18819
rect 17417 18785 17451 18819
rect 18429 18785 18463 18819
rect 2145 18717 2179 18751
rect 9505 18717 9539 18751
rect 11805 18717 11839 18751
rect 13093 18717 13127 18751
rect 13921 18717 13955 18751
rect 14197 18717 14231 18751
rect 15393 18717 15427 18751
rect 4629 18649 4663 18683
rect 11437 18649 11471 18683
rect 12449 18649 12483 18683
rect 3433 18581 3467 18615
rect 3893 18581 3927 18615
rect 7941 18581 7975 18615
rect 9137 18581 9171 18615
rect 11253 18581 11287 18615
rect 16497 18581 16531 18615
rect 18613 18581 18647 18615
rect 2421 18377 2455 18411
rect 3157 18377 3191 18411
rect 4997 18377 5031 18411
rect 8217 18377 8251 18411
rect 9873 18377 9907 18411
rect 11345 18377 11379 18411
rect 11713 18377 11747 18411
rect 18429 18377 18463 18411
rect 4721 18309 4755 18343
rect 6285 18309 6319 18343
rect 8493 18309 8527 18343
rect 14841 18309 14875 18343
rect 15301 18309 15335 18343
rect 1501 18241 1535 18275
rect 2145 18241 2179 18275
rect 5917 18241 5951 18275
rect 6653 18241 6687 18275
rect 7849 18241 7883 18275
rect 8769 18241 8803 18275
rect 10609 18241 10643 18275
rect 13921 18241 13955 18275
rect 16497 18241 16531 18275
rect 16865 18241 16899 18275
rect 2881 18173 2915 18207
rect 3341 18173 3375 18207
rect 5825 18173 5859 18207
rect 7113 18173 7147 18207
rect 7205 18173 7239 18207
rect 7389 18173 7423 18207
rect 12265 18173 12299 18207
rect 12633 18173 12667 18207
rect 1593 18105 1627 18139
rect 3662 18105 3696 18139
rect 8861 18105 8895 18139
rect 9413 18105 9447 18139
rect 10333 18105 10367 18139
rect 10425 18105 10459 18139
rect 12449 18105 12483 18139
rect 13001 18105 13035 18139
rect 14242 18105 14276 18139
rect 16589 18105 16623 18139
rect 4261 18037 4295 18071
rect 13277 18037 13311 18071
rect 13829 18037 13863 18071
rect 15761 18037 15795 18071
rect 16313 18037 16347 18071
rect 17417 18037 17451 18071
rect 1685 17833 1719 17867
rect 3157 17833 3191 17867
rect 4261 17833 4295 17867
rect 5273 17833 5307 17867
rect 7205 17833 7239 17867
rect 8677 17833 8711 17867
rect 8953 17833 8987 17867
rect 9505 17833 9539 17867
rect 9873 17833 9907 17867
rect 11437 17833 11471 17867
rect 16681 17833 16715 17867
rect 16773 17833 16807 17867
rect 17049 17833 17083 17867
rect 2599 17765 2633 17799
rect 8078 17765 8112 17799
rect 11989 17765 12023 17799
rect 16082 17765 16116 17799
rect 4077 17697 4111 17731
rect 5457 17697 5491 17731
rect 5641 17697 5675 17731
rect 6009 17697 6043 17731
rect 6561 17697 6595 17731
rect 10241 17697 10275 17731
rect 12081 17697 12115 17731
rect 12633 17697 12667 17731
rect 13277 17697 13311 17731
rect 13645 17697 13679 17731
rect 14197 17697 14231 17731
rect 2237 17629 2271 17663
rect 7757 17629 7791 17663
rect 12817 17629 12851 17663
rect 14381 17629 14415 17663
rect 15761 17629 15795 17663
rect 17647 17765 17681 17799
rect 17544 17697 17578 17731
rect 18521 17697 18555 17731
rect 4629 17561 4663 17595
rect 16773 17561 16807 17595
rect 2053 17493 2087 17527
rect 3433 17493 3467 17527
rect 3893 17493 3927 17527
rect 5089 17493 5123 17527
rect 7481 17493 7515 17527
rect 10609 17493 10643 17527
rect 18705 17493 18739 17527
rect 2329 17289 2363 17323
rect 10149 17289 10183 17323
rect 13461 17289 13495 17323
rect 17049 17289 17083 17323
rect 18889 17289 18923 17323
rect 3985 17221 4019 17255
rect 14841 17221 14875 17255
rect 15209 17221 15243 17255
rect 16313 17221 16347 17255
rect 18245 17221 18279 17255
rect 4353 17153 4387 17187
rect 6653 17153 6687 17187
rect 10609 17153 10643 17187
rect 12265 17153 12299 17187
rect 15761 17153 15795 17187
rect 16681 17153 16715 17187
rect 1409 17085 1443 17119
rect 4721 17085 4755 17119
rect 4905 17085 4939 17119
rect 5273 17085 5307 17119
rect 5825 17085 5859 17119
rect 6837 17085 6871 17119
rect 7297 17085 7331 17119
rect 7849 17085 7883 17119
rect 8217 17085 8251 17119
rect 10701 17085 10735 17119
rect 10793 17085 10827 17119
rect 10977 17085 11011 17119
rect 12633 17085 12667 17119
rect 13921 17085 13955 17119
rect 18061 17085 18095 17119
rect 18521 17085 18555 17119
rect 2973 17017 3007 17051
rect 3065 17017 3099 17051
rect 3617 17017 3651 17051
rect 6285 17017 6319 17051
rect 8309 17017 8343 17051
rect 9229 17017 9263 17051
rect 9321 17017 9355 17051
rect 9873 17017 9907 17051
rect 12449 17017 12483 17051
rect 13001 17017 13035 17051
rect 14283 17017 14317 17051
rect 15853 17017 15887 17051
rect 1593 16949 1627 16983
rect 2789 16949 2823 16983
rect 4537 16949 4571 16983
rect 8585 16949 8619 16983
rect 9045 16949 9079 16983
rect 11161 16949 11195 16983
rect 11805 16949 11839 16983
rect 13829 16949 13863 16983
rect 15485 16949 15519 16983
rect 17509 16949 17543 16983
rect 2789 16745 2823 16779
rect 6469 16745 6503 16779
rect 8769 16745 8803 16779
rect 13829 16745 13863 16779
rect 16313 16745 16347 16779
rect 16865 16745 16899 16779
rect 3111 16677 3145 16711
rect 4169 16677 4203 16711
rect 4261 16677 4295 16711
rect 9873 16677 9907 16711
rect 10793 16677 10827 16711
rect 15485 16677 15519 16711
rect 16037 16677 16071 16711
rect 2053 16609 2087 16643
rect 3008 16609 3042 16643
rect 5676 16609 5710 16643
rect 6653 16609 6687 16643
rect 7113 16609 7147 16643
rect 7665 16609 7699 16643
rect 8033 16609 8067 16643
rect 11897 16609 11931 16643
rect 12357 16609 12391 16643
rect 13461 16609 13495 16643
rect 17877 16609 17911 16643
rect 4445 16541 4479 16575
rect 9137 16541 9171 16575
rect 9781 16541 9815 16575
rect 10057 16541 10091 16575
rect 12633 16541 12667 16575
rect 13001 16541 13035 16575
rect 15393 16541 15427 16575
rect 2421 16473 2455 16507
rect 3893 16473 3927 16507
rect 8033 16473 8067 16507
rect 11161 16473 11195 16507
rect 14657 16473 14691 16507
rect 18061 16473 18095 16507
rect 1685 16405 1719 16439
rect 3433 16405 3467 16439
rect 5181 16405 5215 16439
rect 5779 16405 5813 16439
rect 6193 16405 6227 16439
rect 8401 16405 8435 16439
rect 14381 16405 14415 16439
rect 4077 16201 4111 16235
rect 8861 16201 8895 16235
rect 11897 16201 11931 16235
rect 12725 16201 12759 16235
rect 14197 16201 14231 16235
rect 14657 16201 14691 16235
rect 15025 16201 15059 16235
rect 16957 16201 16991 16235
rect 18613 16201 18647 16235
rect 2881 16133 2915 16167
rect 6561 16133 6595 16167
rect 7113 16133 7147 16167
rect 15853 16133 15887 16167
rect 17049 16133 17083 16167
rect 17325 16133 17359 16167
rect 3065 16065 3099 16099
rect 4537 16065 4571 16099
rect 7665 16065 7699 16099
rect 9413 16065 9447 16099
rect 13921 16065 13955 16099
rect 4629 15997 4663 16031
rect 8585 15997 8619 16031
rect 9321 15997 9355 16031
rect 10057 15997 10091 16031
rect 10425 15997 10459 16031
rect 11161 15997 11195 16031
rect 13001 15997 13035 16031
rect 13185 15997 13219 16031
rect 13645 15997 13679 16031
rect 16773 15997 16807 16031
rect 17049 15997 17083 16031
rect 18061 15997 18095 16031
rect 18889 15997 18923 16031
rect 1501 15929 1535 15963
rect 1593 15929 1627 15963
rect 2145 15929 2179 15963
rect 3157 15929 3191 15963
rect 3709 15929 3743 15963
rect 6285 15929 6319 15963
rect 7481 15929 7515 15963
rect 7986 15929 8020 15963
rect 10885 15929 10919 15963
rect 10977 15929 11011 15963
rect 11529 15929 11563 15963
rect 15301 15929 15335 15963
rect 15393 15929 15427 15963
rect 2421 15861 2455 15895
rect 4445 15861 4479 15895
rect 5733 15861 5767 15895
rect 12173 15861 12207 15895
rect 16221 15861 16255 15895
rect 16589 15861 16623 15895
rect 18245 15861 18279 15895
rect 2513 15657 2547 15691
rect 3893 15657 3927 15691
rect 4629 15657 4663 15691
rect 5273 15657 5307 15691
rect 6929 15657 6963 15691
rect 7297 15657 7331 15691
rect 7757 15657 7791 15691
rect 9505 15657 9539 15691
rect 11713 15657 11747 15691
rect 13921 15657 13955 15691
rect 14289 15657 14323 15691
rect 15393 15657 15427 15691
rect 1685 15589 1719 15623
rect 2237 15589 2271 15623
rect 9873 15589 9907 15623
rect 12725 15589 12759 15623
rect 18429 15589 18463 15623
rect 4128 15521 4162 15555
rect 5457 15521 5491 15555
rect 5917 15521 5951 15555
rect 6193 15521 6227 15555
rect 6377 15521 6411 15555
rect 8309 15521 8343 15555
rect 8585 15521 8619 15555
rect 11529 15521 11563 15555
rect 14105 15521 14139 15555
rect 15301 15521 15335 15555
rect 15853 15521 15887 15555
rect 16865 15521 16899 15555
rect 18280 15521 18314 15555
rect 1593 15453 1627 15487
rect 4215 15453 4249 15487
rect 5089 15453 5123 15487
rect 8769 15453 8803 15487
rect 9781 15453 9815 15487
rect 10425 15453 10459 15487
rect 12633 15453 12667 15487
rect 13277 15453 13311 15487
rect 17003 15453 17037 15487
rect 3065 15317 3099 15351
rect 3525 15317 3559 15351
rect 12081 15317 12115 15351
rect 13645 15317 13679 15351
rect 2881 15113 2915 15147
rect 5733 15113 5767 15147
rect 8953 15113 8987 15147
rect 11161 15113 11195 15147
rect 12173 15113 12207 15147
rect 13277 15113 13311 15147
rect 14565 15113 14599 15147
rect 16129 15113 16163 15147
rect 18245 15113 18279 15147
rect 2145 15045 2179 15079
rect 4261 15045 4295 15079
rect 6009 15045 6043 15079
rect 15025 15045 15059 15079
rect 1593 14977 1627 15011
rect 2513 14977 2547 15011
rect 3065 14977 3099 15011
rect 4813 14977 4847 15011
rect 9873 14977 9907 15011
rect 11805 14977 11839 15011
rect 13645 14977 13679 15011
rect 14289 14977 14323 15011
rect 15209 14977 15243 15011
rect 16957 14977 16991 15011
rect 3985 14909 4019 14943
rect 7113 14909 7147 14943
rect 7297 14909 7331 14943
rect 7665 14909 7699 14943
rect 8125 14909 8159 14943
rect 11345 14909 11379 14943
rect 12449 14909 12483 14943
rect 12909 14909 12943 14943
rect 15853 14909 15887 14943
rect 17233 14909 17267 14943
rect 1685 14841 1719 14875
rect 3386 14841 3420 14875
rect 4629 14841 4663 14875
rect 5134 14841 5168 14875
rect 9965 14841 9999 14875
rect 10517 14841 10551 14875
rect 13746 14841 13780 14875
rect 15301 14841 15335 14875
rect 6653 14773 6687 14807
rect 7113 14773 7147 14807
rect 8585 14773 8619 14807
rect 9597 14773 9631 14807
rect 10793 14773 10827 14807
rect 11529 14773 11563 14807
rect 12633 14773 12667 14807
rect 16497 14773 16531 14807
rect 1685 14569 1719 14603
rect 2053 14569 2087 14603
rect 3157 14569 3191 14603
rect 5273 14569 5307 14603
rect 6929 14569 6963 14603
rect 7297 14569 7331 14603
rect 9045 14569 9079 14603
rect 9413 14569 9447 14603
rect 10793 14569 10827 14603
rect 12633 14569 12667 14603
rect 13001 14569 13035 14603
rect 14565 14569 14599 14603
rect 16221 14569 16255 14603
rect 2237 14501 2271 14535
rect 2329 14501 2363 14535
rect 2881 14501 2915 14535
rect 4629 14501 4663 14535
rect 5089 14501 5123 14535
rect 8125 14501 8159 14535
rect 8217 14501 8251 14535
rect 10235 14501 10269 14535
rect 11805 14501 11839 14535
rect 13277 14501 13311 14535
rect 13369 14501 13403 14535
rect 13921 14501 13955 14535
rect 15622 14501 15656 14535
rect 4169 14433 4203 14467
rect 5457 14433 5491 14467
rect 5917 14433 5951 14467
rect 6193 14433 6227 14467
rect 6561 14433 6595 14467
rect 7665 14433 7699 14467
rect 9873 14433 9907 14467
rect 15301 14433 15335 14467
rect 3893 14365 3927 14399
rect 8769 14365 8803 14399
rect 11713 14365 11747 14399
rect 12357 14365 12391 14399
rect 4353 14297 4387 14331
rect 14289 14229 14323 14263
rect 3249 14025 3283 14059
rect 3893 14025 3927 14059
rect 6193 14025 6227 14059
rect 6653 14025 6687 14059
rect 10425 14025 10459 14059
rect 10793 14025 10827 14059
rect 11805 14025 11839 14059
rect 13369 14025 13403 14059
rect 15117 14025 15151 14059
rect 16957 14025 16991 14059
rect 10057 13957 10091 13991
rect 15761 13957 15795 13991
rect 1593 13889 1627 13923
rect 2237 13889 2271 13923
rect 2881 13889 2915 13923
rect 12449 13889 12483 13923
rect 14105 13889 14139 13923
rect 15485 13889 15519 13923
rect 3065 13821 3099 13855
rect 4629 13821 4663 13855
rect 5181 13821 5215 13855
rect 5273 13821 5307 13855
rect 5825 13821 5859 13855
rect 7021 13821 7055 13855
rect 7297 13821 7331 13855
rect 7665 13821 7699 13855
rect 8033 13821 8067 13855
rect 9137 13821 9171 13855
rect 11069 13821 11103 13855
rect 14197 13821 14231 13855
rect 15945 13821 15979 13855
rect 16405 13821 16439 13855
rect 1685 13753 1719 13787
rect 4261 13753 4295 13787
rect 10885 13753 10919 13787
rect 12265 13753 12299 13787
rect 12811 13753 12845 13787
rect 13645 13753 13679 13787
rect 14518 13753 14552 13787
rect 2513 13685 2547 13719
rect 4537 13685 4571 13719
rect 6929 13685 6963 13719
rect 8677 13685 8711 13719
rect 8953 13685 8987 13719
rect 9505 13685 9539 13719
rect 11161 13685 11195 13719
rect 16037 13685 16071 13719
rect 1685 13481 1719 13515
rect 2513 13481 2547 13515
rect 3801 13481 3835 13515
rect 5273 13481 5307 13515
rect 6929 13481 6963 13515
rect 7665 13481 7699 13515
rect 7941 13481 7975 13515
rect 9137 13481 9171 13515
rect 9781 13481 9815 13515
rect 11621 13481 11655 13515
rect 11989 13481 12023 13515
rect 12541 13481 12575 13515
rect 13369 13481 13403 13515
rect 15393 13481 15427 13515
rect 16957 13481 16991 13515
rect 10885 13413 10919 13447
rect 2881 13345 2915 13379
rect 4112 13345 4146 13379
rect 5457 13345 5491 13379
rect 5641 13345 5675 13379
rect 6193 13345 6227 13379
rect 6561 13345 6595 13379
rect 7297 13345 7331 13379
rect 8125 13345 8159 13379
rect 8401 13345 8435 13379
rect 9873 13345 9907 13379
rect 10241 13345 10275 13379
rect 13093 13345 13127 13379
rect 13988 13345 14022 13379
rect 15577 13345 15611 13379
rect 15761 13345 15795 13379
rect 16313 13345 16347 13379
rect 16865 13345 16899 13379
rect 17325 13345 17359 13379
rect 3249 13277 3283 13311
rect 4629 13277 4663 13311
rect 12173 13277 12207 13311
rect 4215 13209 4249 13243
rect 1961 13141 1995 13175
rect 5089 13141 5123 13175
rect 13829 13141 13863 13175
rect 14059 13141 14093 13175
rect 15117 13141 15151 13175
rect 2973 12937 3007 12971
rect 3617 12937 3651 12971
rect 4905 12937 4939 12971
rect 5365 12937 5399 12971
rect 5917 12937 5951 12971
rect 8033 12937 8067 12971
rect 9413 12937 9447 12971
rect 10149 12937 10183 12971
rect 12265 12937 12299 12971
rect 14841 12937 14875 12971
rect 16865 12937 16899 12971
rect 9781 12869 9815 12903
rect 17233 12869 17267 12903
rect 2053 12801 2087 12835
rect 2513 12801 2547 12835
rect 3709 12801 3743 12835
rect 11529 12801 11563 12835
rect 12633 12801 12667 12835
rect 13185 12801 13219 12835
rect 15393 12801 15427 12835
rect 6653 12733 6687 12767
rect 7205 12733 7239 12767
rect 7481 12733 7515 12767
rect 7665 12733 7699 12767
rect 8493 12733 8527 12767
rect 10793 12733 10827 12767
rect 11345 12733 11379 12767
rect 1869 12665 1903 12699
rect 2145 12665 2179 12699
rect 4071 12665 4105 12699
rect 13277 12665 13311 12699
rect 13829 12665 13863 12699
rect 15485 12665 15519 12699
rect 16037 12665 16071 12699
rect 4629 12597 4663 12631
rect 5457 12597 5491 12631
rect 8309 12597 8343 12631
rect 8861 12597 8895 12631
rect 10701 12597 10735 12631
rect 14105 12597 14139 12631
rect 15209 12597 15243 12631
rect 16313 12597 16347 12631
rect 1409 12393 1443 12427
rect 1961 12393 1995 12427
rect 3801 12393 3835 12427
rect 4629 12393 4663 12427
rect 5089 12393 5123 12427
rect 7021 12393 7055 12427
rect 9045 12393 9079 12427
rect 13369 12393 13403 12427
rect 14933 12393 14967 12427
rect 17141 12393 17175 12427
rect 2237 12325 2271 12359
rect 2605 12325 2639 12359
rect 4215 12325 4249 12359
rect 5502 12325 5536 12359
rect 8170 12325 8204 12359
rect 10793 12325 10827 12359
rect 11345 12325 11379 12359
rect 13093 12325 13127 12359
rect 13829 12325 13863 12359
rect 14381 12325 14415 12359
rect 15663 12325 15697 12359
rect 4128 12257 4162 12291
rect 5181 12257 5215 12291
rect 7849 12257 7883 12291
rect 8769 12257 8803 12291
rect 12170 12257 12204 12291
rect 12357 12257 12391 12291
rect 15301 12257 15335 12291
rect 17325 12257 17359 12291
rect 17601 12257 17635 12291
rect 2513 12189 2547 12223
rect 3157 12189 3191 12223
rect 10701 12189 10735 12223
rect 12725 12189 12759 12223
rect 13737 12189 13771 12223
rect 6101 12053 6135 12087
rect 7757 12053 7791 12087
rect 16221 12053 16255 12087
rect 5089 11849 5123 11883
rect 8217 11849 8251 11883
rect 11161 11849 11195 11883
rect 11437 11849 11471 11883
rect 12173 11849 12207 11883
rect 13645 11849 13679 11883
rect 14657 11849 14691 11883
rect 15761 11849 15795 11883
rect 16037 11849 16071 11883
rect 16727 11849 16761 11883
rect 17417 11849 17451 11883
rect 4169 11781 4203 11815
rect 11805 11781 11839 11815
rect 16405 11781 16439 11815
rect 1593 11713 1627 11747
rect 3433 11713 3467 11747
rect 4721 11713 4755 11747
rect 5273 11713 5307 11747
rect 5549 11713 5583 11747
rect 9045 11713 9079 11747
rect 9689 11713 9723 11747
rect 10241 11713 10275 11747
rect 6653 11645 6687 11679
rect 6929 11645 6963 11679
rect 14841 11645 14875 11679
rect 16656 11645 16690 11679
rect 17049 11645 17083 11679
rect 1685 11577 1719 11611
rect 2237 11577 2271 11611
rect 3157 11577 3191 11611
rect 3249 11577 3283 11611
rect 5342 11577 5376 11611
rect 6837 11577 6871 11611
rect 8769 11577 8803 11611
rect 8861 11577 8895 11611
rect 10149 11577 10183 11611
rect 10603 11577 10637 11611
rect 12725 11577 12759 11611
rect 12817 11577 12851 11611
rect 13369 11577 13403 11611
rect 15162 11577 15196 11611
rect 2605 11509 2639 11543
rect 2973 11509 3007 11543
rect 7849 11509 7883 11543
rect 14105 11509 14139 11543
rect 17785 11509 17819 11543
rect 1685 11305 1719 11339
rect 3433 11305 3467 11339
rect 5273 11305 5307 11339
rect 6745 11305 6779 11339
rect 7941 11305 7975 11339
rect 8861 11305 8895 11339
rect 10241 11305 10275 11339
rect 10793 11305 10827 11339
rect 12541 11305 12575 11339
rect 14657 11305 14691 11339
rect 2237 11237 2271 11271
rect 4077 11237 4111 11271
rect 6146 11237 6180 11271
rect 12817 11237 12851 11271
rect 15485 11237 15519 11271
rect 16037 11237 16071 11271
rect 4721 11169 4755 11203
rect 5549 11169 5583 11203
rect 5825 11169 5859 11203
rect 7573 11169 7607 11203
rect 14264 11169 14298 11203
rect 2145 11101 2179 11135
rect 2789 11101 2823 11135
rect 3801 11101 3835 11135
rect 10425 11101 10459 11135
rect 12725 11101 12759 11135
rect 13369 11101 13403 11135
rect 15393 11101 15427 11135
rect 16865 11101 16899 11135
rect 3065 10965 3099 10999
rect 8493 10965 8527 10999
rect 9137 10965 9171 10999
rect 11345 10965 11379 10999
rect 11621 10965 11655 10999
rect 14335 10965 14369 10999
rect 4721 10761 4755 10795
rect 6193 10761 6227 10795
rect 6653 10761 6687 10795
rect 7113 10761 7147 10795
rect 10517 10761 10551 10795
rect 11805 10761 11839 10795
rect 14197 10761 14231 10795
rect 15393 10761 15427 10795
rect 15761 10761 15795 10795
rect 3157 10693 3191 10727
rect 7481 10693 7515 10727
rect 8309 10693 8343 10727
rect 11437 10693 11471 10727
rect 15991 10693 16025 10727
rect 2605 10625 2639 10659
rect 4169 10625 4203 10659
rect 9045 10625 9079 10659
rect 9321 10625 9355 10659
rect 9965 10625 9999 10659
rect 10885 10625 10919 10659
rect 12817 10625 12851 10659
rect 13829 10625 13863 10659
rect 14381 10625 14415 10659
rect 15920 10557 15954 10591
rect 16865 10557 16899 10591
rect 17325 10557 17359 10591
rect 1501 10489 1535 10523
rect 2697 10489 2731 10523
rect 3525 10489 3559 10523
rect 5273 10489 5307 10523
rect 5365 10489 5399 10523
rect 5917 10489 5951 10523
rect 7757 10489 7791 10523
rect 7849 10489 7883 10523
rect 9413 10489 9447 10523
rect 10977 10489 11011 10523
rect 12909 10489 12943 10523
rect 13461 10489 13495 10523
rect 14473 10489 14507 10523
rect 15025 10489 15059 10523
rect 16313 10489 16347 10523
rect 2053 10421 2087 10455
rect 5089 10421 5123 10455
rect 8677 10421 8711 10455
rect 12173 10421 12207 10455
rect 17049 10421 17083 10455
rect 2053 10217 2087 10251
rect 5043 10217 5077 10251
rect 9321 10217 9355 10251
rect 11345 10217 11379 10251
rect 12449 10217 12483 10251
rect 13093 10217 13127 10251
rect 13553 10217 13587 10251
rect 13737 10217 13771 10251
rect 16451 10217 16485 10251
rect 2881 10149 2915 10183
rect 6009 10149 6043 10183
rect 6101 10149 6135 10183
rect 7757 10149 7791 10183
rect 8217 10149 8251 10183
rect 8769 10149 8803 10183
rect 9873 10149 9907 10183
rect 15439 10149 15473 10183
rect 2237 10081 2271 10115
rect 11529 10081 11563 10115
rect 11805 10081 11839 10115
rect 12817 10081 12851 10115
rect 13645 10081 13679 10115
rect 14105 10081 14139 10115
rect 15352 10081 15386 10115
rect 16380 10081 16414 10115
rect 17325 10081 17359 10115
rect 6285 10013 6319 10047
rect 8125 10013 8159 10047
rect 9781 10013 9815 10047
rect 10057 10013 10091 10047
rect 5365 9945 5399 9979
rect 4813 9877 4847 9911
rect 10793 9877 10827 9911
rect 14657 9877 14691 9911
rect 17509 9877 17543 9911
rect 2145 9673 2179 9707
rect 2375 9673 2409 9707
rect 3525 9673 3559 9707
rect 6285 9673 6319 9707
rect 7205 9673 7239 9707
rect 10701 9673 10735 9707
rect 13645 9673 13679 9707
rect 17325 9673 17359 9707
rect 3801 9605 3835 9639
rect 6561 9605 6595 9639
rect 7849 9605 7883 9639
rect 8953 9605 8987 9639
rect 11805 9605 11839 9639
rect 2304 9469 2338 9503
rect 3316 9469 3350 9503
rect 4629 9469 4663 9503
rect 5273 9469 5307 9503
rect 7348 9469 7382 9503
rect 10793 9469 10827 9503
rect 11253 9469 11287 9503
rect 14381 9469 14415 9503
rect 16164 9469 16198 9503
rect 16957 9469 16991 9503
rect 18096 9469 18130 9503
rect 18521 9469 18555 9503
rect 5917 9401 5951 9435
rect 7435 9401 7469 9435
rect 8401 9401 8435 9435
rect 8493 9401 8527 9435
rect 9597 9401 9631 9435
rect 11529 9401 11563 9435
rect 12541 9401 12575 9435
rect 12633 9401 12667 9435
rect 13185 9401 13219 9435
rect 14702 9401 14736 9435
rect 16267 9401 16301 9435
rect 2789 9333 2823 9367
rect 4905 9333 4939 9367
rect 8125 9333 8159 9367
rect 10057 9333 10091 9367
rect 12265 9333 12299 9367
rect 14289 9333 14323 9367
rect 15301 9333 15335 9367
rect 15577 9333 15611 9367
rect 16681 9333 16715 9367
rect 18199 9333 18233 9367
rect 1823 9129 1857 9163
rect 2835 9129 2869 9163
rect 5135 9129 5169 9163
rect 7573 9129 7607 9163
rect 8125 9129 8159 9163
rect 9413 9129 9447 9163
rect 11345 9129 11379 9163
rect 13093 9129 13127 9163
rect 13737 9129 13771 9163
rect 6193 9061 6227 9095
rect 11891 9061 11925 9095
rect 15485 9061 15519 9095
rect 1752 8993 1786 9027
rect 2732 8993 2766 9027
rect 5064 8993 5098 9027
rect 8309 8993 8343 9027
rect 8585 8993 8619 9027
rect 10057 8993 10091 9027
rect 10425 8993 10459 9027
rect 11529 8993 11563 9027
rect 13553 8993 13587 9027
rect 14013 8993 14047 9027
rect 16865 8993 16899 9027
rect 6101 8925 6135 8959
rect 6377 8925 6411 8959
rect 7941 8925 7975 8959
rect 10701 8925 10735 8959
rect 15117 8925 15151 8959
rect 15393 8925 15427 8959
rect 12817 8857 12851 8891
rect 15945 8857 15979 8891
rect 9045 8789 9079 8823
rect 12449 8789 12483 8823
rect 14565 8789 14599 8823
rect 17003 8789 17037 8823
rect 1685 8585 1719 8619
rect 2559 8585 2593 8619
rect 2881 8585 2915 8619
rect 3341 8585 3375 8619
rect 5089 8585 5123 8619
rect 6561 8585 6595 8619
rect 7343 8585 7377 8619
rect 8033 8585 8067 8619
rect 9505 8585 9539 8619
rect 11069 8585 11103 8619
rect 16267 8585 16301 8619
rect 5871 8517 5905 8551
rect 13461 8517 13495 8551
rect 2329 8449 2363 8483
rect 8217 8449 8251 8483
rect 9873 8449 9907 8483
rect 11621 8449 11655 8483
rect 12541 8449 12575 8483
rect 13185 8449 13219 8483
rect 13921 8449 13955 8483
rect 1444 8381 1478 8415
rect 1869 8381 1903 8415
rect 2488 8381 2522 8415
rect 5800 8381 5834 8415
rect 6193 8381 6227 8415
rect 7240 8381 7274 8415
rect 7665 8381 7699 8415
rect 10241 8381 10275 8415
rect 10425 8381 10459 8415
rect 14381 8381 14415 8415
rect 16164 8381 16198 8415
rect 8538 8313 8572 8347
rect 12265 8313 12299 8347
rect 12633 8313 12667 8347
rect 14702 8313 14736 8347
rect 5549 8245 5583 8279
rect 9137 8245 9171 8279
rect 10057 8245 10091 8279
rect 14289 8245 14323 8279
rect 15301 8245 15335 8279
rect 15669 8245 15703 8279
rect 15945 8245 15979 8279
rect 16865 8245 16899 8279
rect 6009 8041 6043 8075
rect 6975 8041 7009 8075
rect 9505 8041 9539 8075
rect 11345 8041 11379 8075
rect 12357 8041 12391 8075
rect 12633 8041 12667 8075
rect 14841 8041 14875 8075
rect 8170 7973 8204 8007
rect 11799 7973 11833 8007
rect 15485 7973 15519 8007
rect 5825 7905 5859 7939
rect 6904 7905 6938 7939
rect 7849 7905 7883 7939
rect 9965 7905 9999 7939
rect 10333 7905 10367 7939
rect 11437 7905 11471 7939
rect 13277 7905 13311 7939
rect 13645 7905 13679 7939
rect 16900 7905 16934 7939
rect 9045 7837 9079 7871
rect 10609 7837 10643 7871
rect 13829 7837 13863 7871
rect 15393 7837 15427 7871
rect 17003 7837 17037 7871
rect 13001 7769 13035 7803
rect 15945 7769 15979 7803
rect 7297 7701 7331 7735
rect 7757 7701 7791 7735
rect 8769 7701 8803 7735
rect 14565 7701 14599 7735
rect 16405 7701 16439 7735
rect 5917 7497 5951 7531
rect 7159 7497 7193 7531
rect 9137 7497 9171 7531
rect 13461 7497 13495 7531
rect 13921 7497 13955 7531
rect 17141 7497 17175 7531
rect 10609 7429 10643 7463
rect 8125 7361 8159 7395
rect 16129 7361 16163 7395
rect 7056 7293 7090 7327
rect 7849 7293 7883 7327
rect 9873 7293 9907 7327
rect 10057 7293 10091 7327
rect 10977 7293 11011 7327
rect 11380 7293 11414 7327
rect 11805 7293 11839 7327
rect 12633 7293 12667 7327
rect 13001 7293 13035 7327
rect 14381 7293 14415 7327
rect 14473 7293 14507 7327
rect 15025 7293 15059 7327
rect 8217 7225 8251 7259
rect 8769 7225 8803 7259
rect 9505 7225 9539 7259
rect 15209 7225 15243 7259
rect 16221 7225 16255 7259
rect 16773 7225 16807 7259
rect 7481 7157 7515 7191
rect 9689 7157 9723 7191
rect 11483 7157 11517 7191
rect 12265 7157 12299 7191
rect 12541 7157 12575 7191
rect 15485 7157 15519 7191
rect 15945 7157 15979 7191
rect 7573 6953 7607 6987
rect 7941 6953 7975 6987
rect 11437 6953 11471 6987
rect 12357 6953 12391 6987
rect 15117 6953 15151 6987
rect 15669 6953 15703 6987
rect 16221 6953 16255 6987
rect 17141 6953 17175 6987
rect 8217 6885 8251 6919
rect 8769 6885 8803 6919
rect 9045 6885 9079 6919
rect 10010 6885 10044 6919
rect 7072 6817 7106 6851
rect 9505 6817 9539 6851
rect 9689 6817 9723 6851
rect 11989 6817 12023 6851
rect 15301 6817 15335 6851
rect 17049 6817 17083 6851
rect 17509 6817 17543 6851
rect 7159 6749 7193 6783
rect 8125 6749 8159 6783
rect 14197 6749 14231 6783
rect 10609 6613 10643 6647
rect 12909 6613 12943 6647
rect 6653 6409 6687 6443
rect 9505 6409 9539 6443
rect 10609 6409 10643 6443
rect 11253 6409 11287 6443
rect 12081 6409 12115 6443
rect 15945 6409 15979 6443
rect 17141 6409 17175 6443
rect 9045 6341 9079 6375
rect 8769 6273 8803 6307
rect 9689 6273 9723 6307
rect 10149 6273 10183 6307
rect 13185 6273 13219 6307
rect 14381 6273 14415 6307
rect 16221 6273 16255 6307
rect 16497 6273 16531 6307
rect 7021 6137 7055 6171
rect 7849 6137 7883 6171
rect 8125 6137 8159 6171
rect 8217 6137 8251 6171
rect 9781 6137 9815 6171
rect 11345 6137 11379 6171
rect 12541 6137 12575 6171
rect 12633 6137 12667 6171
rect 13461 6137 13495 6171
rect 14289 6137 14323 6171
rect 14743 6137 14777 6171
rect 16313 6137 16347 6171
rect 7481 6069 7515 6103
rect 15301 6069 15335 6103
rect 15577 6069 15611 6103
rect 17509 6069 17543 6103
rect 12633 5865 12667 5899
rect 14473 5865 14507 5899
rect 15117 5865 15151 5899
rect 16957 5865 16991 5899
rect 18521 5865 18555 5899
rect 8170 5797 8204 5831
rect 9873 5797 9907 5831
rect 11799 5797 11833 5831
rect 13369 5797 13403 5831
rect 6377 5729 6411 5763
rect 6745 5729 6779 5763
rect 7021 5729 7055 5763
rect 9137 5729 9171 5763
rect 11437 5729 11471 5763
rect 15301 5729 15335 5763
rect 15761 5729 15795 5763
rect 16865 5729 16899 5763
rect 17417 5729 17451 5763
rect 18429 5729 18463 5763
rect 18889 5729 18923 5763
rect 7389 5661 7423 5695
rect 7849 5661 7883 5695
rect 9781 5661 9815 5695
rect 10149 5661 10183 5695
rect 13277 5661 13311 5695
rect 15853 5661 15887 5695
rect 13829 5593 13863 5627
rect 7665 5525 7699 5559
rect 8769 5525 8803 5559
rect 12357 5525 12391 5559
rect 13001 5525 13035 5559
rect 16313 5525 16347 5559
rect 6377 5321 6411 5355
rect 7021 5321 7055 5355
rect 8585 5321 8619 5355
rect 8953 5321 8987 5355
rect 10333 5321 10367 5355
rect 12081 5321 12115 5355
rect 13737 5321 13771 5355
rect 16405 5321 16439 5355
rect 17417 5321 17451 5355
rect 17785 5321 17819 5355
rect 18521 5321 18555 5355
rect 18889 5321 18923 5355
rect 9137 5185 9171 5219
rect 13093 5185 13127 5219
rect 14381 5185 14415 5219
rect 15209 5185 15243 5219
rect 7481 5117 7515 5151
rect 7757 5117 7791 5151
rect 8033 5117 8067 5151
rect 10701 5117 10735 5151
rect 10952 5117 10986 5151
rect 17024 5117 17058 5151
rect 18096 5117 18130 5151
rect 8309 5049 8343 5083
rect 9458 5049 9492 5083
rect 11437 5049 11471 5083
rect 12817 5049 12851 5083
rect 12909 5049 12943 5083
rect 16773 5049 16807 5083
rect 10057 4981 10091 5015
rect 11023 4981 11057 5015
rect 11805 4981 11839 5015
rect 14657 4981 14691 5015
rect 15117 4981 15151 5015
rect 15577 4981 15611 5015
rect 16129 4981 16163 5015
rect 17095 4981 17129 5015
rect 18199 4981 18233 5015
rect 7665 4777 7699 4811
rect 8033 4777 8067 4811
rect 10609 4777 10643 4811
rect 12357 4777 12391 4811
rect 12909 4777 12943 4811
rect 13553 4777 13587 4811
rect 15669 4777 15703 4811
rect 16957 4777 16991 4811
rect 10010 4709 10044 4743
rect 17233 4709 17267 4743
rect 17785 4709 17819 4743
rect 6964 4641 6998 4675
rect 8217 4641 8251 4675
rect 8401 4641 8435 4675
rect 9689 4641 9723 4675
rect 13772 4641 13806 4675
rect 15301 4641 15335 4675
rect 11989 4573 12023 4607
rect 17141 4573 17175 4607
rect 7067 4437 7101 4471
rect 8953 4437 8987 4471
rect 10885 4437 10919 4471
rect 13185 4437 13219 4471
rect 13875 4437 13909 4471
rect 16221 4437 16255 4471
rect 6285 4233 6319 4267
rect 8769 4233 8803 4267
rect 10333 4233 10367 4267
rect 13737 4233 13771 4267
rect 14013 4233 14047 4267
rect 14657 4233 14691 4267
rect 16589 4233 16623 4267
rect 19211 4233 19245 4267
rect 6653 4165 6687 4199
rect 8401 4165 8435 4199
rect 17509 4165 17543 4199
rect 7481 4097 7515 4131
rect 9321 4097 9355 4131
rect 10609 4097 10643 4131
rect 10977 4097 11011 4131
rect 15209 4097 15243 4131
rect 17233 4097 17267 4131
rect 5800 4029 5834 4063
rect 12449 4029 12483 4063
rect 16748 4029 16782 4063
rect 18096 4029 18130 4063
rect 18521 4029 18555 4063
rect 19108 4029 19142 4063
rect 19533 4029 19567 4063
rect 6009 3961 6043 3995
rect 7573 3961 7607 3995
rect 8125 3961 8159 3995
rect 9045 3961 9079 3995
rect 9137 3961 9171 3995
rect 10701 3961 10735 3995
rect 11897 3961 11931 3995
rect 12265 3961 12299 3995
rect 12811 3961 12845 3995
rect 15301 3961 15335 3995
rect 15853 3961 15887 3995
rect 7021 3893 7055 3927
rect 9965 3893 9999 3927
rect 13369 3893 13403 3927
rect 15025 3893 15059 3927
rect 16129 3893 16163 3927
rect 16819 3893 16853 3927
rect 18199 3893 18233 3927
rect 5733 3689 5767 3723
rect 7573 3689 7607 3723
rect 9045 3689 9079 3723
rect 9873 3689 9907 3723
rect 13185 3689 13219 3723
rect 16773 3689 16807 3723
rect 8217 3621 8251 3655
rect 10701 3621 10735 3655
rect 11253 3621 11287 3655
rect 12265 3621 12299 3655
rect 13737 3621 13771 3655
rect 13829 3621 13863 3655
rect 15485 3621 15519 3655
rect 17049 3621 17083 3655
rect 17601 3621 17635 3655
rect 18613 3621 18647 3655
rect 5064 3553 5098 3587
rect 6076 3553 6110 3587
rect 7056 3553 7090 3587
rect 8125 3485 8159 3519
rect 8769 3485 8803 3519
rect 10425 3485 10459 3519
rect 10609 3485 10643 3519
rect 12173 3485 12207 3519
rect 14013 3485 14047 3519
rect 15393 3485 15427 3519
rect 15853 3485 15887 3519
rect 16957 3485 16991 3519
rect 18521 3485 18555 3519
rect 18797 3485 18831 3519
rect 5135 3417 5169 3451
rect 7159 3417 7193 3451
rect 7849 3417 7883 3451
rect 12725 3417 12759 3451
rect 17969 3417 18003 3451
rect 6147 3349 6181 3383
rect 6837 3349 6871 3383
rect 9413 3349 9447 3383
rect 14841 3349 14875 3383
rect 16405 3349 16439 3383
rect 4261 3145 4295 3179
rect 4859 3145 4893 3179
rect 7757 3145 7791 3179
rect 8033 3145 8067 3179
rect 8309 3145 8343 3179
rect 10333 3145 10367 3179
rect 11897 3145 11931 3179
rect 12265 3145 12299 3179
rect 13645 3145 13679 3179
rect 15853 3145 15887 3179
rect 17417 3145 17451 3179
rect 17877 3145 17911 3179
rect 18199 3145 18233 3179
rect 5871 3077 5905 3111
rect 6285 3009 6319 3043
rect 7021 3009 7055 3043
rect 7665 3009 7699 3043
rect 14013 3077 14047 3111
rect 16221 3077 16255 3111
rect 19211 3077 19245 3111
rect 20637 3077 20671 3111
rect 8861 3009 8895 3043
rect 11529 3009 11563 3043
rect 12817 3009 12851 3043
rect 16497 3009 16531 3043
rect 16773 3009 16807 3043
rect 18613 3009 18647 3043
rect 3760 2941 3794 2975
rect 4788 2941 4822 2975
rect 5800 2941 5834 2975
rect 7757 2941 7791 2975
rect 18128 2941 18162 2975
rect 19140 2941 19174 2975
rect 19533 2941 19567 2975
rect 20453 2941 20487 2975
rect 21005 2941 21039 2975
rect 23673 2941 23707 2975
rect 24225 2941 24259 2975
rect 3847 2873 3881 2907
rect 7113 2873 7147 2907
rect 8585 2873 8619 2907
rect 8686 2873 8720 2907
rect 9873 2873 9907 2907
rect 10885 2873 10919 2907
rect 10977 2873 11011 2907
rect 12541 2873 12575 2907
rect 12633 2873 12667 2907
rect 14933 2873 14967 2907
rect 15025 2873 15059 2907
rect 15577 2873 15611 2907
rect 16589 2873 16623 2907
rect 18889 2873 18923 2907
rect 5273 2805 5307 2839
rect 5641 2805 5675 2839
rect 6653 2805 6687 2839
rect 9505 2805 9539 2839
rect 10701 2805 10735 2839
rect 14749 2805 14783 2839
rect 23857 2805 23891 2839
rect 3111 2601 3145 2635
rect 5963 2601 5997 2635
rect 7389 2601 7423 2635
rect 10793 2601 10827 2635
rect 11989 2601 12023 2635
rect 12357 2601 12391 2635
rect 14105 2601 14139 2635
rect 14519 2601 14553 2635
rect 18613 2601 18647 2635
rect 21465 2601 21499 2635
rect 6377 2533 6411 2567
rect 8033 2533 8067 2567
rect 8309 2533 8343 2567
rect 8861 2533 8895 2567
rect 9505 2533 9539 2567
rect 11161 2533 11195 2567
rect 12725 2533 12759 2567
rect 12817 2533 12851 2567
rect 15301 2533 15335 2567
rect 15669 2533 15703 2567
rect 16589 2533 16623 2567
rect 16865 2533 16899 2567
rect 21833 2533 21867 2567
rect 3040 2465 3074 2499
rect 4880 2465 4914 2499
rect 5892 2465 5926 2499
rect 7180 2465 7214 2499
rect 9781 2465 9815 2499
rect 10333 2465 10367 2499
rect 14416 2465 14450 2499
rect 14841 2465 14875 2499
rect 17141 2465 17175 2499
rect 17693 2465 17727 2499
rect 18429 2465 18463 2499
rect 18981 2465 19015 2499
rect 19533 2465 19567 2499
rect 20085 2465 20119 2499
rect 21281 2465 21315 2499
rect 22385 2465 22419 2499
rect 22937 2465 22971 2499
rect 24593 2465 24627 2499
rect 25145 2465 25179 2499
rect 8217 2397 8251 2431
rect 9137 2397 9171 2431
rect 11069 2397 11103 2431
rect 11345 2397 11379 2431
rect 13001 2397 13035 2431
rect 15577 2397 15611 2431
rect 3525 2329 3559 2363
rect 7665 2329 7699 2363
rect 9965 2329 9999 2363
rect 16129 2329 16163 2363
rect 17325 2329 17359 2363
rect 19717 2329 19751 2363
rect 22569 2329 22603 2363
rect 24777 2329 24811 2363
rect 4951 2261 4985 2295
rect 5365 2261 5399 2295
rect 13645 2261 13679 2295
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 4433 25483 4491 25489
rect 4433 25449 4445 25483
rect 4479 25480 4491 25483
rect 4522 25480 4528 25492
rect 4479 25452 4528 25480
rect 4479 25449 4491 25452
rect 4433 25443 4491 25449
rect 4522 25440 4528 25452
rect 4580 25480 4586 25492
rect 5902 25480 5908 25492
rect 4580 25452 5908 25480
rect 4580 25440 4586 25452
rect 5902 25440 5908 25452
rect 5960 25440 5966 25492
rect 1464 25347 1522 25353
rect 1464 25313 1476 25347
rect 1510 25344 1522 25347
rect 2774 25344 2780 25356
rect 1510 25316 2780 25344
rect 1510 25313 1522 25316
rect 1464 25307 1522 25313
rect 2774 25304 2780 25316
rect 2832 25304 2838 25356
rect 5880 25347 5938 25353
rect 5880 25313 5892 25347
rect 5926 25344 5938 25347
rect 5994 25344 6000 25356
rect 5926 25316 6000 25344
rect 5926 25313 5938 25316
rect 5880 25307 5938 25313
rect 5994 25304 6000 25316
rect 6052 25344 6058 25356
rect 6730 25344 6736 25356
rect 6052 25316 6736 25344
rect 6052 25304 6058 25316
rect 6730 25304 6736 25316
rect 6788 25304 6794 25356
rect 7374 25344 7380 25356
rect 7335 25316 7380 25344
rect 7374 25304 7380 25316
rect 7432 25304 7438 25356
rect 8202 25304 8208 25356
rect 8260 25344 8266 25356
rect 8700 25347 8758 25353
rect 8700 25344 8712 25347
rect 8260 25316 8712 25344
rect 8260 25304 8266 25316
rect 8700 25313 8712 25316
rect 8746 25313 8758 25347
rect 8700 25307 8758 25313
rect 9122 25304 9128 25356
rect 9180 25344 9186 25356
rect 11552 25347 11610 25353
rect 11552 25344 11564 25347
rect 9180 25316 11564 25344
rect 9180 25304 9186 25316
rect 11552 25313 11564 25316
rect 11598 25344 11610 25347
rect 11698 25344 11704 25356
rect 11598 25316 11704 25344
rect 11598 25313 11610 25316
rect 11552 25307 11610 25313
rect 11698 25304 11704 25316
rect 11756 25304 11762 25356
rect 13240 25347 13298 25353
rect 13240 25313 13252 25347
rect 13286 25344 13298 25347
rect 13354 25344 13360 25356
rect 13286 25316 13360 25344
rect 13286 25313 13298 25316
rect 13240 25307 13298 25313
rect 13354 25304 13360 25316
rect 13412 25304 13418 25356
rect 10045 25279 10103 25285
rect 10045 25245 10057 25279
rect 10091 25276 10103 25279
rect 10134 25276 10140 25288
rect 10091 25248 10140 25276
rect 10091 25245 10103 25248
rect 10045 25239 10103 25245
rect 10134 25236 10140 25248
rect 10192 25236 10198 25288
rect 7006 25168 7012 25220
rect 7064 25208 7070 25220
rect 7929 25211 7987 25217
rect 7929 25208 7941 25211
rect 7064 25180 7941 25208
rect 7064 25168 7070 25180
rect 7929 25177 7941 25180
rect 7975 25177 7987 25211
rect 7929 25171 7987 25177
rect 1210 25100 1216 25152
rect 1268 25140 1274 25152
rect 1535 25143 1593 25149
rect 1535 25140 1547 25143
rect 1268 25112 1547 25140
rect 1268 25100 1274 25112
rect 1535 25109 1547 25112
rect 1581 25109 1593 25143
rect 2866 25140 2872 25152
rect 2827 25112 2872 25140
rect 1535 25103 1593 25109
rect 2866 25100 2872 25112
rect 2924 25100 2930 25152
rect 3099 25143 3157 25149
rect 3099 25109 3111 25143
rect 3145 25140 3157 25143
rect 3786 25140 3792 25152
rect 3145 25112 3792 25140
rect 3145 25109 3157 25112
rect 3099 25103 3157 25109
rect 3786 25100 3792 25112
rect 3844 25100 3850 25152
rect 4706 25149 4712 25152
rect 4663 25143 4712 25149
rect 4663 25140 4675 25143
rect 4619 25112 4675 25140
rect 4663 25109 4675 25112
rect 4709 25109 4712 25143
rect 4663 25103 4712 25109
rect 4706 25100 4712 25103
rect 4764 25140 4770 25152
rect 4985 25143 5043 25149
rect 4985 25140 4997 25143
rect 4764 25112 4997 25140
rect 4764 25100 4770 25112
rect 4985 25109 4997 25112
rect 5031 25109 5043 25143
rect 4985 25103 5043 25109
rect 5951 25143 6009 25149
rect 5951 25109 5963 25143
rect 5997 25140 6009 25143
rect 6914 25140 6920 25152
rect 5997 25112 6920 25140
rect 5997 25109 6009 25112
rect 5951 25103 6009 25109
rect 6914 25100 6920 25112
rect 6972 25100 6978 25152
rect 7190 25140 7196 25152
rect 7151 25112 7196 25140
rect 7190 25100 7196 25112
rect 7248 25100 7254 25152
rect 8018 25100 8024 25152
rect 8076 25140 8082 25152
rect 8803 25143 8861 25149
rect 8803 25140 8815 25143
rect 8076 25112 8815 25140
rect 8076 25100 8082 25112
rect 8803 25109 8815 25112
rect 8849 25109 8861 25143
rect 8803 25103 8861 25109
rect 11655 25143 11713 25149
rect 11655 25109 11667 25143
rect 11701 25140 11713 25143
rect 13170 25140 13176 25152
rect 11701 25112 13176 25140
rect 11701 25109 11713 25112
rect 11655 25103 11713 25109
rect 13170 25100 13176 25112
rect 13228 25100 13234 25152
rect 13311 25143 13369 25149
rect 13311 25109 13323 25143
rect 13357 25140 13369 25143
rect 13538 25140 13544 25152
rect 13357 25112 13544 25140
rect 13357 25109 13369 25112
rect 13311 25103 13369 25109
rect 13538 25100 13544 25112
rect 13596 25100 13602 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 2041 24939 2099 24945
rect 2041 24905 2053 24939
rect 2087 24936 2099 24939
rect 2774 24936 2780 24948
rect 2087 24908 2780 24936
rect 2087 24905 2099 24908
rect 2041 24899 2099 24905
rect 2774 24896 2780 24908
rect 2832 24896 2838 24948
rect 4522 24936 4528 24948
rect 4483 24908 4528 24936
rect 4522 24896 4528 24908
rect 4580 24896 4586 24948
rect 5905 24939 5963 24945
rect 5905 24905 5917 24939
rect 5951 24936 5963 24939
rect 5994 24936 6000 24948
rect 5951 24908 6000 24936
rect 5951 24905 5963 24908
rect 5905 24899 5963 24905
rect 5994 24896 6000 24908
rect 6052 24896 6058 24948
rect 11698 24896 11704 24948
rect 11756 24936 11762 24948
rect 11793 24939 11851 24945
rect 11793 24936 11805 24939
rect 11756 24908 11805 24936
rect 11756 24896 11762 24908
rect 11793 24905 11805 24908
rect 11839 24905 11851 24939
rect 11793 24899 11851 24905
rect 2409 24871 2467 24877
rect 2409 24837 2421 24871
rect 2455 24868 2467 24871
rect 8018 24868 8024 24880
rect 2455 24840 8024 24868
rect 2455 24837 2467 24840
rect 2409 24831 2467 24837
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24732 1455 24735
rect 2424 24732 2452 24831
rect 8018 24828 8024 24840
rect 8076 24828 8082 24880
rect 10686 24828 10692 24880
rect 10744 24868 10750 24880
rect 13265 24871 13323 24877
rect 13265 24868 13277 24871
rect 10744 24840 13277 24868
rect 10744 24828 10750 24840
rect 13265 24837 13277 24840
rect 13311 24868 13323 24871
rect 13354 24868 13360 24880
rect 13311 24840 13360 24868
rect 13311 24837 13323 24840
rect 13265 24831 13323 24837
rect 13354 24828 13360 24840
rect 13412 24828 13418 24880
rect 4706 24800 4712 24812
rect 4667 24772 4712 24800
rect 4706 24760 4712 24772
rect 4764 24760 4770 24812
rect 4982 24800 4988 24812
rect 4943 24772 4988 24800
rect 4982 24760 4988 24772
rect 5040 24760 5046 24812
rect 7006 24760 7012 24812
rect 7064 24800 7070 24812
rect 7193 24803 7251 24809
rect 7193 24800 7205 24803
rect 7064 24772 7205 24800
rect 7064 24760 7070 24772
rect 7193 24769 7205 24772
rect 7239 24769 7251 24803
rect 7558 24800 7564 24812
rect 7519 24772 7564 24800
rect 7193 24763 7251 24769
rect 7558 24760 7564 24772
rect 7616 24760 7622 24812
rect 1443 24704 2452 24732
rect 3304 24735 3362 24741
rect 1443 24701 1455 24704
rect 1397 24695 1455 24701
rect 3304 24701 3316 24735
rect 3350 24732 3362 24735
rect 3789 24735 3847 24741
rect 3789 24732 3801 24735
rect 3350 24704 3801 24732
rect 3350 24701 3362 24704
rect 3304 24695 3362 24701
rect 3789 24701 3801 24704
rect 3835 24732 3847 24735
rect 4522 24732 4528 24744
rect 3835 24704 4528 24732
rect 3835 24701 3847 24704
rect 3789 24695 3847 24701
rect 4522 24692 4528 24704
rect 4580 24692 4586 24744
rect 8570 24732 8576 24744
rect 8483 24704 8576 24732
rect 8570 24692 8576 24704
rect 8628 24732 8634 24744
rect 8757 24735 8815 24741
rect 8757 24732 8769 24735
rect 8628 24704 8769 24732
rect 8628 24692 8634 24704
rect 8757 24701 8769 24704
rect 8803 24701 8815 24735
rect 8757 24695 8815 24701
rect 8846 24692 8852 24744
rect 8904 24732 8910 24744
rect 10229 24735 10287 24741
rect 10229 24732 10241 24735
rect 8904 24704 10241 24732
rect 8904 24692 8910 24704
rect 10229 24701 10241 24704
rect 10275 24732 10287 24735
rect 10781 24735 10839 24741
rect 10781 24732 10793 24735
rect 10275 24704 10793 24732
rect 10275 24701 10287 24704
rect 10229 24695 10287 24701
rect 10781 24701 10793 24704
rect 10827 24701 10839 24735
rect 10781 24695 10839 24701
rect 11384 24735 11442 24741
rect 11384 24701 11396 24735
rect 11430 24732 11442 24735
rect 11790 24732 11796 24744
rect 11430 24704 11796 24732
rect 11430 24701 11442 24704
rect 11384 24695 11442 24701
rect 11790 24692 11796 24704
rect 11848 24732 11854 24744
rect 12161 24735 12219 24741
rect 12161 24732 12173 24735
rect 11848 24704 12173 24732
rect 11848 24692 11854 24704
rect 12161 24701 12173 24704
rect 12207 24701 12219 24735
rect 12161 24695 12219 24701
rect 12504 24735 12562 24741
rect 12504 24701 12516 24735
rect 12550 24732 12562 24735
rect 12989 24735 13047 24741
rect 12989 24732 13001 24735
rect 12550 24704 13001 24732
rect 12550 24701 12562 24704
rect 12504 24695 12562 24701
rect 12989 24701 13001 24704
rect 13035 24732 13047 24735
rect 13541 24735 13599 24741
rect 13541 24732 13553 24735
rect 13035 24704 13553 24732
rect 13035 24701 13047 24704
rect 12989 24695 13047 24701
rect 13541 24701 13553 24704
rect 13587 24732 13599 24735
rect 13587 24704 14136 24732
rect 13587 24701 13599 24704
rect 13541 24695 13599 24701
rect 2866 24624 2872 24676
rect 2924 24664 2930 24676
rect 3053 24667 3111 24673
rect 3053 24664 3065 24667
rect 2924 24636 3065 24664
rect 2924 24624 2930 24636
rect 3053 24633 3065 24636
rect 3099 24664 3111 24667
rect 4157 24667 4215 24673
rect 3099 24636 3556 24664
rect 3099 24633 3111 24636
rect 3053 24627 3111 24633
rect 1578 24596 1584 24608
rect 1539 24568 1584 24596
rect 1578 24556 1584 24568
rect 1636 24556 1642 24608
rect 2406 24556 2412 24608
rect 2464 24596 2470 24608
rect 3375 24599 3433 24605
rect 3375 24596 3387 24599
rect 2464 24568 3387 24596
rect 2464 24556 2470 24568
rect 3375 24565 3387 24568
rect 3421 24565 3433 24599
rect 3528 24596 3556 24636
rect 4157 24633 4169 24667
rect 4203 24664 4215 24667
rect 4798 24664 4804 24676
rect 4203 24636 4804 24664
rect 4203 24633 4215 24636
rect 4157 24627 4215 24633
rect 4798 24624 4804 24636
rect 4856 24624 4862 24676
rect 7285 24667 7343 24673
rect 7285 24633 7297 24667
rect 7331 24664 7343 24667
rect 7374 24664 7380 24676
rect 7331 24636 7380 24664
rect 7331 24633 7343 24636
rect 7285 24627 7343 24633
rect 4338 24596 4344 24608
rect 3528 24568 4344 24596
rect 3375 24559 3433 24565
rect 4338 24556 4344 24568
rect 4396 24596 4402 24608
rect 5350 24596 5356 24608
rect 4396 24568 5356 24596
rect 4396 24556 4402 24568
rect 5350 24556 5356 24568
rect 5408 24556 5414 24608
rect 6273 24599 6331 24605
rect 6273 24565 6285 24599
rect 6319 24596 6331 24599
rect 6641 24599 6699 24605
rect 6641 24596 6653 24599
rect 6319 24568 6653 24596
rect 6319 24565 6331 24568
rect 6273 24559 6331 24565
rect 6641 24565 6653 24568
rect 6687 24596 6699 24599
rect 7300 24596 7328 24627
rect 7374 24624 7380 24636
rect 7432 24624 7438 24676
rect 7926 24624 7932 24676
rect 7984 24664 7990 24676
rect 8665 24667 8723 24673
rect 8665 24664 8677 24667
rect 7984 24636 8677 24664
rect 7984 24624 7990 24636
rect 8665 24633 8677 24636
rect 8711 24633 8723 24667
rect 8665 24627 8723 24633
rect 11471 24667 11529 24673
rect 11471 24633 11483 24667
rect 11517 24664 11529 24667
rect 11974 24664 11980 24676
rect 11517 24636 11980 24664
rect 11517 24633 11529 24636
rect 11471 24627 11529 24633
rect 11974 24624 11980 24636
rect 12032 24624 12038 24676
rect 14108 24608 14136 24704
rect 8202 24596 8208 24608
rect 6687 24568 7328 24596
rect 8163 24568 8208 24596
rect 6687 24565 6699 24568
rect 6641 24559 6699 24565
rect 8202 24556 8208 24568
rect 8260 24556 8266 24608
rect 10413 24599 10471 24605
rect 10413 24565 10425 24599
rect 10459 24596 10471 24599
rect 10686 24596 10692 24608
rect 10459 24568 10692 24596
rect 10459 24565 10471 24568
rect 10413 24559 10471 24565
rect 10686 24556 10692 24568
rect 10744 24556 10750 24608
rect 12250 24556 12256 24608
rect 12308 24596 12314 24608
rect 12575 24599 12633 24605
rect 12575 24596 12587 24599
rect 12308 24568 12587 24596
rect 12308 24556 12314 24568
rect 12575 24565 12587 24568
rect 12621 24565 12633 24599
rect 13722 24596 13728 24608
rect 13683 24568 13728 24596
rect 12575 24559 12633 24565
rect 13722 24556 13728 24568
rect 13780 24556 13786 24608
rect 14090 24596 14096 24608
rect 14051 24568 14096 24596
rect 14090 24556 14096 24568
rect 14148 24556 14154 24608
rect 14458 24556 14464 24608
rect 14516 24596 14522 24608
rect 17954 24596 17960 24608
rect 14516 24568 17960 24596
rect 14516 24556 14522 24568
rect 17954 24556 17960 24568
rect 18012 24556 18018 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1486 24352 1492 24404
rect 1544 24392 1550 24404
rect 1581 24395 1639 24401
rect 1581 24392 1593 24395
rect 1544 24364 1593 24392
rect 1544 24352 1550 24364
rect 1581 24361 1593 24364
rect 1627 24361 1639 24395
rect 14274 24392 14280 24404
rect 14187 24364 14280 24392
rect 1581 24355 1639 24361
rect 14274 24352 14280 24364
rect 14332 24392 14338 24404
rect 18690 24392 18696 24404
rect 14332 24364 18696 24392
rect 14332 24352 14338 24364
rect 18690 24352 18696 24364
rect 18748 24352 18754 24404
rect 21729 24395 21787 24401
rect 21729 24361 21741 24395
rect 21775 24392 21787 24395
rect 23474 24392 23480 24404
rect 21775 24364 23480 24392
rect 21775 24361 21787 24364
rect 21729 24355 21787 24361
rect 23474 24352 23480 24364
rect 23532 24352 23538 24404
rect 4706 24324 4712 24336
rect 4667 24296 4712 24324
rect 4706 24284 4712 24296
rect 4764 24284 4770 24336
rect 6914 24324 6920 24336
rect 6875 24296 6920 24324
rect 6914 24284 6920 24296
rect 6972 24284 6978 24336
rect 7009 24327 7067 24333
rect 7009 24293 7021 24327
rect 7055 24324 7067 24327
rect 7190 24324 7196 24336
rect 7055 24296 7196 24324
rect 7055 24293 7067 24296
rect 7009 24287 7067 24293
rect 7190 24284 7196 24296
rect 7248 24284 7254 24336
rect 7558 24324 7564 24336
rect 7519 24296 7564 24324
rect 7558 24284 7564 24296
rect 7616 24284 7622 24336
rect 8202 24284 8208 24336
rect 8260 24324 8266 24336
rect 10594 24324 10600 24336
rect 8260 24296 10600 24324
rect 8260 24284 8266 24296
rect 10594 24284 10600 24296
rect 10652 24284 10658 24336
rect 1397 24259 1455 24265
rect 1397 24225 1409 24259
rect 1443 24256 1455 24259
rect 1670 24256 1676 24268
rect 1443 24228 1676 24256
rect 1443 24225 1455 24228
rect 1397 24219 1455 24225
rect 1670 24216 1676 24228
rect 1728 24216 1734 24268
rect 2568 24259 2626 24265
rect 2568 24225 2580 24259
rect 2614 24256 2626 24259
rect 2958 24256 2964 24268
rect 2614 24228 2964 24256
rect 2614 24225 2626 24228
rect 2568 24219 2626 24225
rect 2958 24216 2964 24228
rect 3016 24216 3022 24268
rect 10686 24256 10692 24268
rect 10647 24228 10692 24256
rect 10686 24216 10692 24228
rect 10744 24216 10750 24268
rect 11698 24265 11704 24268
rect 11676 24259 11704 24265
rect 11676 24256 11688 24259
rect 11611 24228 11688 24256
rect 11676 24225 11688 24228
rect 11756 24256 11762 24268
rect 12342 24256 12348 24268
rect 11756 24228 12348 24256
rect 11676 24219 11704 24225
rect 11698 24216 11704 24219
rect 11756 24216 11762 24228
rect 12342 24216 12348 24228
rect 12400 24216 12406 24268
rect 13630 24256 13636 24268
rect 13591 24228 13636 24256
rect 13630 24216 13636 24228
rect 13688 24256 13694 24268
rect 14734 24256 14740 24268
rect 13688 24228 14740 24256
rect 13688 24216 13694 24228
rect 14734 24216 14740 24228
rect 14792 24216 14798 24268
rect 20714 24216 20720 24268
rect 20772 24256 20778 24268
rect 21545 24259 21603 24265
rect 21545 24256 21557 24259
rect 20772 24228 21557 24256
rect 20772 24216 20778 24228
rect 21545 24225 21557 24228
rect 21591 24225 21603 24259
rect 21545 24219 21603 24225
rect 4617 24191 4675 24197
rect 4617 24157 4629 24191
rect 4663 24188 4675 24191
rect 4982 24188 4988 24200
rect 4663 24160 4988 24188
rect 4663 24157 4675 24160
rect 4617 24151 4675 24157
rect 4982 24148 4988 24160
rect 5040 24148 5046 24200
rect 7650 24148 7656 24200
rect 7708 24188 7714 24200
rect 7929 24191 7987 24197
rect 7929 24188 7941 24191
rect 7708 24160 7941 24188
rect 7708 24148 7714 24160
rect 7929 24157 7941 24160
rect 7975 24188 7987 24191
rect 8389 24191 8447 24197
rect 8389 24188 8401 24191
rect 7975 24160 8401 24188
rect 7975 24157 7987 24160
rect 7929 24151 7987 24157
rect 8389 24157 8401 24160
rect 8435 24157 8447 24191
rect 10042 24188 10048 24200
rect 10003 24160 10048 24188
rect 8389 24151 8447 24157
rect 10042 24148 10048 24160
rect 10100 24148 10106 24200
rect 13817 24191 13875 24197
rect 13817 24157 13829 24191
rect 13863 24188 13875 24191
rect 14182 24188 14188 24200
rect 13863 24160 14188 24188
rect 13863 24157 13875 24160
rect 13817 24151 13875 24157
rect 14182 24148 14188 24160
rect 14240 24188 14246 24200
rect 14553 24191 14611 24197
rect 14553 24188 14565 24191
rect 14240 24160 14565 24188
rect 14240 24148 14246 24160
rect 14553 24157 14565 24160
rect 14599 24157 14611 24191
rect 14553 24151 14611 24157
rect 4522 24080 4528 24132
rect 4580 24120 4586 24132
rect 5169 24123 5227 24129
rect 5169 24120 5181 24123
rect 4580 24092 5181 24120
rect 4580 24080 4586 24092
rect 5169 24089 5181 24092
rect 5215 24089 5227 24123
rect 5169 24083 5227 24089
rect 1670 24012 1676 24064
rect 1728 24052 1734 24064
rect 2639 24055 2697 24061
rect 2639 24052 2651 24055
rect 1728 24024 2651 24052
rect 1728 24012 1734 24024
rect 2639 24021 2651 24024
rect 2685 24021 2697 24055
rect 2639 24015 2697 24021
rect 10226 24012 10232 24064
rect 10284 24052 10290 24064
rect 11747 24055 11805 24061
rect 11747 24052 11759 24055
rect 10284 24024 11759 24052
rect 10284 24012 10290 24024
rect 11747 24021 11759 24024
rect 11793 24021 11805 24055
rect 11747 24015 11805 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1670 23848 1676 23860
rect 1631 23820 1676 23848
rect 1670 23808 1676 23820
rect 1728 23808 1734 23860
rect 2225 23851 2283 23857
rect 2225 23817 2237 23851
rect 2271 23848 2283 23851
rect 2406 23848 2412 23860
rect 2271 23820 2412 23848
rect 2271 23817 2283 23820
rect 2225 23811 2283 23817
rect 2332 23653 2360 23820
rect 2406 23808 2412 23820
rect 2464 23808 2470 23860
rect 2498 23808 2504 23860
rect 2556 23848 2562 23860
rect 2556 23820 2601 23848
rect 2556 23808 2562 23820
rect 4706 23808 4712 23860
rect 4764 23848 4770 23860
rect 5169 23851 5227 23857
rect 5169 23848 5181 23851
rect 4764 23820 5181 23848
rect 4764 23808 4770 23820
rect 5169 23817 5181 23820
rect 5215 23848 5227 23851
rect 5442 23848 5448 23860
rect 5215 23820 5448 23848
rect 5215 23817 5227 23820
rect 5169 23811 5227 23817
rect 5442 23808 5448 23820
rect 5500 23808 5506 23860
rect 6641 23851 6699 23857
rect 6641 23817 6653 23851
rect 6687 23848 6699 23851
rect 6914 23848 6920 23860
rect 6687 23820 6920 23848
rect 6687 23817 6699 23820
rect 6641 23811 6699 23817
rect 6914 23808 6920 23820
rect 6972 23808 6978 23860
rect 7101 23851 7159 23857
rect 7101 23817 7113 23851
rect 7147 23848 7159 23851
rect 7190 23848 7196 23860
rect 7147 23820 7196 23848
rect 7147 23817 7159 23820
rect 7101 23811 7159 23817
rect 7190 23808 7196 23820
rect 7248 23808 7254 23860
rect 9674 23848 9680 23860
rect 9635 23820 9680 23848
rect 9674 23808 9680 23820
rect 9732 23808 9738 23860
rect 10042 23848 10048 23860
rect 10003 23820 10048 23848
rect 10042 23808 10048 23820
rect 10100 23808 10106 23860
rect 10686 23808 10692 23860
rect 10744 23848 10750 23860
rect 11149 23851 11207 23857
rect 11149 23848 11161 23851
rect 10744 23820 11161 23848
rect 10744 23808 10750 23820
rect 11149 23817 11161 23820
rect 11195 23817 11207 23851
rect 11698 23848 11704 23860
rect 11659 23820 11704 23848
rect 11149 23811 11207 23817
rect 11698 23808 11704 23820
rect 11756 23808 11762 23860
rect 13630 23848 13636 23860
rect 13591 23820 13636 23848
rect 13630 23808 13636 23820
rect 13688 23808 13694 23860
rect 14093 23851 14151 23857
rect 14093 23817 14105 23851
rect 14139 23848 14151 23851
rect 14458 23848 14464 23860
rect 14139 23820 14464 23848
rect 14139 23817 14151 23820
rect 14093 23811 14151 23817
rect 14458 23808 14464 23820
rect 14516 23808 14522 23860
rect 19337 23851 19395 23857
rect 19337 23817 19349 23851
rect 19383 23848 19395 23851
rect 21082 23848 21088 23860
rect 19383 23820 21088 23848
rect 19383 23817 19395 23820
rect 19337 23811 19395 23817
rect 21082 23808 21088 23820
rect 21140 23808 21146 23860
rect 21545 23851 21603 23857
rect 21545 23817 21557 23851
rect 21591 23848 21603 23851
rect 22738 23848 22744 23860
rect 21591 23820 22744 23848
rect 21591 23817 21603 23820
rect 21545 23811 21603 23817
rect 22738 23808 22744 23820
rect 22796 23808 22802 23860
rect 24765 23851 24823 23857
rect 24765 23817 24777 23851
rect 24811 23848 24823 23851
rect 27522 23848 27528 23860
rect 24811 23820 27528 23848
rect 24811 23817 24823 23820
rect 24765 23811 24823 23817
rect 27522 23808 27528 23820
rect 27580 23808 27586 23860
rect 2958 23780 2964 23792
rect 2871 23752 2964 23780
rect 2958 23740 2964 23752
rect 3016 23780 3022 23792
rect 4430 23780 4436 23792
rect 3016 23752 4436 23780
rect 3016 23740 3022 23752
rect 4430 23740 4436 23752
rect 4488 23740 4494 23792
rect 4522 23740 4528 23792
rect 4580 23780 4586 23792
rect 4801 23783 4859 23789
rect 4801 23780 4813 23783
rect 4580 23752 4813 23780
rect 4580 23740 4586 23752
rect 4801 23749 4813 23752
rect 4847 23749 4859 23783
rect 4801 23743 4859 23749
rect 4982 23740 4988 23792
rect 5040 23780 5046 23792
rect 5537 23783 5595 23789
rect 5537 23780 5549 23783
rect 5040 23752 5549 23780
rect 5040 23740 5046 23752
rect 5537 23749 5549 23752
rect 5583 23749 5595 23783
rect 5537 23743 5595 23749
rect 9766 23740 9772 23792
rect 9824 23780 9830 23792
rect 10134 23780 10140 23792
rect 9824 23752 10140 23780
rect 9824 23740 9830 23752
rect 10134 23740 10140 23752
rect 10192 23780 10198 23792
rect 14274 23780 14280 23792
rect 10192 23752 10272 23780
rect 10192 23740 10198 23752
rect 3697 23715 3755 23721
rect 3697 23681 3709 23715
rect 3743 23712 3755 23715
rect 4249 23715 4307 23721
rect 4249 23712 4261 23715
rect 3743 23684 4261 23712
rect 3743 23681 3755 23684
rect 3697 23675 3755 23681
rect 4249 23681 4261 23684
rect 4295 23712 4307 23715
rect 5721 23715 5779 23721
rect 5721 23712 5733 23715
rect 4295 23684 5733 23712
rect 4295 23681 4307 23684
rect 4249 23675 4307 23681
rect 5721 23681 5733 23684
rect 5767 23681 5779 23715
rect 7650 23712 7656 23724
rect 7611 23684 7656 23712
rect 5721 23675 5779 23681
rect 7650 23672 7656 23684
rect 7708 23672 7714 23724
rect 10244 23721 10272 23752
rect 13786 23752 14280 23780
rect 10229 23715 10287 23721
rect 10229 23681 10241 23715
rect 10275 23681 10287 23715
rect 10686 23712 10692 23724
rect 10647 23684 10692 23712
rect 10229 23675 10287 23681
rect 10686 23672 10692 23684
rect 10744 23672 10750 23724
rect 2317 23647 2375 23653
rect 2317 23613 2329 23647
rect 2363 23613 2375 23647
rect 2317 23607 2375 23613
rect 9192 23647 9250 23653
rect 9192 23613 9204 23647
rect 9238 23644 9250 23647
rect 9674 23644 9680 23656
rect 9238 23616 9680 23644
rect 9238 23613 9250 23616
rect 9192 23607 9250 23613
rect 9674 23604 9680 23616
rect 9732 23604 9738 23656
rect 12253 23647 12311 23653
rect 12253 23613 12265 23647
rect 12299 23644 12311 23647
rect 12342 23644 12348 23656
rect 12299 23616 12348 23644
rect 12299 23613 12311 23616
rect 12253 23607 12311 23613
rect 12342 23604 12348 23616
rect 12400 23644 12406 23656
rect 12713 23647 12771 23653
rect 12713 23644 12725 23647
rect 12400 23616 12725 23644
rect 12400 23604 12406 23616
rect 12713 23613 12725 23616
rect 12759 23644 12771 23647
rect 13786 23644 13814 23752
rect 14274 23740 14280 23752
rect 14332 23740 14338 23792
rect 20441 23783 20499 23789
rect 20441 23749 20453 23783
rect 20487 23780 20499 23783
rect 21634 23780 21640 23792
rect 20487 23752 21640 23780
rect 20487 23749 20499 23752
rect 20441 23743 20499 23749
rect 21634 23740 21640 23752
rect 21692 23740 21698 23792
rect 13906 23672 13912 23724
rect 13964 23712 13970 23724
rect 16209 23715 16267 23721
rect 16209 23712 16221 23715
rect 13964 23684 16221 23712
rect 13964 23672 13970 23684
rect 14182 23644 14188 23656
rect 12759 23616 13814 23644
rect 14143 23616 14188 23644
rect 12759 23613 12771 23616
rect 12713 23607 12771 23613
rect 14182 23604 14188 23616
rect 14240 23604 14246 23656
rect 14458 23644 14464 23656
rect 14419 23616 14464 23644
rect 14458 23604 14464 23616
rect 14516 23604 14522 23656
rect 15799 23653 15827 23684
rect 16209 23681 16221 23684
rect 16255 23681 16267 23715
rect 16209 23675 16267 23681
rect 20714 23672 20720 23724
rect 20772 23712 20778 23724
rect 22281 23715 22339 23721
rect 22281 23712 22293 23715
rect 20772 23684 22293 23712
rect 20772 23672 20778 23684
rect 22281 23681 22293 23684
rect 22327 23681 22339 23715
rect 22281 23675 22339 23681
rect 15784 23647 15842 23653
rect 15784 23613 15796 23647
rect 15830 23613 15842 23647
rect 15784 23607 15842 23613
rect 18414 23604 18420 23656
rect 18472 23644 18478 23656
rect 19153 23647 19211 23653
rect 19153 23644 19165 23647
rect 18472 23616 19165 23644
rect 18472 23604 18478 23616
rect 19153 23613 19165 23616
rect 19199 23644 19211 23647
rect 19705 23647 19763 23653
rect 19705 23644 19717 23647
rect 19199 23616 19717 23644
rect 19199 23613 19211 23616
rect 19153 23607 19211 23613
rect 19705 23613 19717 23616
rect 19751 23613 19763 23647
rect 20254 23644 20260 23656
rect 20167 23616 20260 23644
rect 19705 23607 19763 23613
rect 20254 23604 20260 23616
rect 20312 23644 20318 23656
rect 20809 23647 20867 23653
rect 20809 23644 20821 23647
rect 20312 23616 20821 23644
rect 20312 23604 20318 23616
rect 20809 23613 20821 23616
rect 20855 23613 20867 23647
rect 21358 23644 21364 23656
rect 21271 23616 21364 23644
rect 20809 23607 20867 23613
rect 21358 23604 21364 23616
rect 21416 23644 21422 23656
rect 21913 23647 21971 23653
rect 21913 23644 21925 23647
rect 21416 23616 21925 23644
rect 21416 23604 21422 23616
rect 21913 23613 21925 23616
rect 21959 23613 21971 23647
rect 21913 23607 21971 23613
rect 23474 23604 23480 23656
rect 23532 23644 23538 23656
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 23532 23616 24593 23644
rect 23532 23604 23538 23616
rect 24581 23613 24593 23616
rect 24627 23644 24639 23647
rect 25133 23647 25191 23653
rect 25133 23644 25145 23647
rect 24627 23616 25145 23644
rect 24627 23613 24639 23616
rect 24581 23607 24639 23613
rect 25133 23613 25145 23616
rect 25179 23613 25191 23647
rect 25133 23607 25191 23613
rect 4341 23579 4399 23585
rect 4341 23545 4353 23579
rect 4387 23545 4399 23579
rect 4341 23539 4399 23545
rect 7469 23579 7527 23585
rect 7469 23545 7481 23579
rect 7515 23576 7527 23579
rect 7745 23579 7803 23585
rect 7745 23576 7757 23579
rect 7515 23548 7757 23576
rect 7515 23545 7527 23548
rect 7469 23539 7527 23545
rect 7745 23545 7757 23548
rect 7791 23576 7803 23579
rect 7926 23576 7932 23588
rect 7791 23548 7932 23576
rect 7791 23545 7803 23548
rect 7745 23539 7803 23545
rect 3970 23468 3976 23520
rect 4028 23508 4034 23520
rect 4065 23511 4123 23517
rect 4065 23508 4077 23511
rect 4028 23480 4077 23508
rect 4028 23468 4034 23480
rect 4065 23477 4077 23480
rect 4111 23508 4123 23511
rect 4356 23508 4384 23539
rect 7926 23536 7932 23548
rect 7984 23536 7990 23588
rect 8297 23579 8355 23585
rect 8297 23545 8309 23579
rect 8343 23545 8355 23579
rect 8297 23539 8355 23545
rect 10321 23579 10379 23585
rect 10321 23545 10333 23579
rect 10367 23545 10379 23579
rect 10321 23539 10379 23545
rect 13786 23548 14228 23576
rect 4111 23480 4384 23508
rect 4111 23477 4123 23480
rect 4065 23471 4123 23477
rect 4430 23468 4436 23520
rect 4488 23508 4494 23520
rect 8018 23508 8024 23520
rect 4488 23480 8024 23508
rect 4488 23468 4494 23480
rect 8018 23468 8024 23480
rect 8076 23508 8082 23520
rect 8312 23508 8340 23539
rect 8076 23480 8340 23508
rect 9263 23511 9321 23517
rect 8076 23468 8082 23480
rect 9263 23477 9275 23511
rect 9309 23508 9321 23511
rect 9398 23508 9404 23520
rect 9309 23480 9404 23508
rect 9309 23477 9321 23480
rect 9263 23471 9321 23477
rect 9398 23468 9404 23480
rect 9456 23468 9462 23520
rect 10042 23468 10048 23520
rect 10100 23508 10106 23520
rect 10336 23508 10364 23539
rect 10100 23480 10364 23508
rect 10100 23468 10106 23480
rect 12710 23468 12716 23520
rect 12768 23508 12774 23520
rect 12897 23511 12955 23517
rect 12897 23508 12909 23511
rect 12768 23480 12909 23508
rect 12768 23468 12774 23480
rect 12897 23477 12909 23480
rect 12943 23477 12955 23511
rect 12897 23471 12955 23477
rect 12986 23468 12992 23520
rect 13044 23508 13050 23520
rect 13786 23508 13814 23548
rect 13044 23480 13814 23508
rect 14200 23508 14228 23548
rect 14550 23536 14556 23588
rect 14608 23576 14614 23588
rect 15887 23579 15945 23585
rect 15887 23576 15899 23579
rect 14608 23548 15899 23576
rect 14608 23536 14614 23548
rect 15887 23545 15899 23548
rect 15933 23545 15945 23579
rect 15887 23539 15945 23545
rect 14645 23511 14703 23517
rect 14645 23508 14657 23511
rect 14200 23480 14657 23508
rect 13044 23468 13050 23480
rect 14645 23477 14657 23480
rect 14691 23477 14703 23511
rect 14645 23471 14703 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 5442 23304 5448 23316
rect 3068 23276 5448 23304
rect 2498 23128 2504 23180
rect 2556 23168 2562 23180
rect 3068 23177 3096 23276
rect 5442 23264 5448 23276
rect 5500 23264 5506 23316
rect 9674 23264 9680 23316
rect 9732 23304 9738 23316
rect 10137 23307 10195 23313
rect 10137 23304 10149 23307
rect 9732 23276 10149 23304
rect 9732 23264 9738 23276
rect 10137 23273 10149 23276
rect 10183 23273 10195 23307
rect 10137 23267 10195 23273
rect 12618 23264 12624 23316
rect 12676 23304 12682 23316
rect 12989 23307 13047 23313
rect 12989 23304 13001 23307
rect 12676 23276 13001 23304
rect 12676 23264 12682 23276
rect 12989 23273 13001 23276
rect 13035 23304 13047 23307
rect 14182 23304 14188 23316
rect 13035 23276 14188 23304
rect 13035 23273 13047 23276
rect 12989 23267 13047 23273
rect 14182 23264 14188 23276
rect 14240 23264 14246 23316
rect 3145 23239 3203 23245
rect 3145 23205 3157 23239
rect 3191 23236 3203 23239
rect 3970 23236 3976 23248
rect 3191 23208 3976 23236
rect 3191 23205 3203 23208
rect 3145 23199 3203 23205
rect 3970 23196 3976 23208
rect 4028 23196 4034 23248
rect 4522 23196 4528 23248
rect 4580 23236 4586 23248
rect 4801 23239 4859 23245
rect 4801 23236 4813 23239
rect 4580 23208 4813 23236
rect 4580 23196 4586 23208
rect 4801 23205 4813 23208
rect 4847 23205 4859 23239
rect 4801 23199 4859 23205
rect 7745 23239 7803 23245
rect 7745 23205 7757 23239
rect 7791 23236 7803 23239
rect 8110 23236 8116 23248
rect 7791 23208 8116 23236
rect 7791 23205 7803 23208
rect 7745 23199 7803 23205
rect 8110 23196 8116 23208
rect 8168 23236 8174 23248
rect 8570 23236 8576 23248
rect 8168 23208 8576 23236
rect 8168 23196 8174 23208
rect 8570 23196 8576 23208
rect 8628 23196 8634 23248
rect 10505 23239 10563 23245
rect 10505 23205 10517 23239
rect 10551 23236 10563 23239
rect 10778 23236 10784 23248
rect 10551 23208 10784 23236
rect 10551 23205 10563 23208
rect 10505 23199 10563 23205
rect 10778 23196 10784 23208
rect 10836 23196 10842 23248
rect 11514 23196 11520 23248
rect 11572 23236 11578 23248
rect 12069 23239 12127 23245
rect 12069 23236 12081 23239
rect 11572 23208 12081 23236
rect 11572 23196 11578 23208
rect 12069 23205 12081 23208
rect 12115 23205 12127 23239
rect 12069 23199 12127 23205
rect 3053 23171 3111 23177
rect 3053 23168 3065 23171
rect 2556 23140 3065 23168
rect 2556 23128 2562 23140
rect 3053 23137 3065 23140
rect 3099 23137 3111 23171
rect 3053 23131 3111 23137
rect 6270 23128 6276 23180
rect 6328 23168 6334 23180
rect 6616 23171 6674 23177
rect 6616 23168 6628 23171
rect 6328 23140 6628 23168
rect 6328 23128 6334 23140
rect 6616 23137 6628 23140
rect 6662 23168 6674 23171
rect 7282 23168 7288 23180
rect 6662 23140 7288 23168
rect 6662 23137 6674 23140
rect 6616 23131 6674 23137
rect 7282 23128 7288 23140
rect 7340 23128 7346 23180
rect 14093 23171 14151 23177
rect 14093 23137 14105 23171
rect 14139 23168 14151 23171
rect 14458 23168 14464 23180
rect 14139 23140 14464 23168
rect 14139 23137 14151 23140
rect 14093 23131 14151 23137
rect 14458 23128 14464 23140
rect 14516 23128 14522 23180
rect 15197 23171 15255 23177
rect 15197 23137 15209 23171
rect 15243 23168 15255 23171
rect 15286 23168 15292 23180
rect 15243 23140 15292 23168
rect 15243 23137 15255 23140
rect 15197 23131 15255 23137
rect 15286 23128 15292 23140
rect 15344 23128 15350 23180
rect 1397 23103 1455 23109
rect 1397 23069 1409 23103
rect 1443 23100 1455 23103
rect 1486 23100 1492 23112
rect 1443 23072 1492 23100
rect 1443 23069 1455 23072
rect 1397 23063 1455 23069
rect 1486 23060 1492 23072
rect 1544 23060 1550 23112
rect 4706 23100 4712 23112
rect 4667 23072 4712 23100
rect 4706 23060 4712 23072
rect 4764 23060 4770 23112
rect 4982 23100 4988 23112
rect 4943 23072 4988 23100
rect 4982 23060 4988 23072
rect 5040 23060 5046 23112
rect 7466 23060 7472 23112
rect 7524 23100 7530 23112
rect 7653 23103 7711 23109
rect 7653 23100 7665 23103
rect 7524 23072 7665 23100
rect 7524 23060 7530 23072
rect 7653 23069 7665 23072
rect 7699 23069 7711 23103
rect 8018 23100 8024 23112
rect 7979 23072 8024 23100
rect 7653 23063 7711 23069
rect 8018 23060 8024 23072
rect 8076 23060 8082 23112
rect 9493 23103 9551 23109
rect 9493 23069 9505 23103
rect 9539 23100 9551 23103
rect 10410 23100 10416 23112
rect 9539 23072 10416 23100
rect 9539 23069 9551 23072
rect 9493 23063 9551 23069
rect 10410 23060 10416 23072
rect 10468 23060 10474 23112
rect 10686 23100 10692 23112
rect 10647 23072 10692 23100
rect 10686 23060 10692 23072
rect 10744 23060 10750 23112
rect 11977 23103 12035 23109
rect 11977 23069 11989 23103
rect 12023 23069 12035 23103
rect 12250 23100 12256 23112
rect 12211 23072 12256 23100
rect 11977 23063 12035 23069
rect 11992 23032 12020 23063
rect 12250 23060 12256 23072
rect 12308 23060 12314 23112
rect 12894 23060 12900 23112
rect 12952 23100 12958 23112
rect 13449 23103 13507 23109
rect 13449 23100 13461 23103
rect 12952 23072 13461 23100
rect 12952 23060 12958 23072
rect 13449 23069 13461 23072
rect 13495 23069 13507 23103
rect 13449 23063 13507 23069
rect 12066 23032 12072 23044
rect 11979 23004 12072 23032
rect 12066 22992 12072 23004
rect 12124 23032 12130 23044
rect 15427 23035 15485 23041
rect 15427 23032 15439 23035
rect 12124 23004 15439 23032
rect 12124 22992 12130 23004
rect 15427 23001 15439 23004
rect 15473 23001 15485 23035
rect 15427 22995 15485 23001
rect 4522 22964 4528 22976
rect 4483 22936 4528 22964
rect 4522 22924 4528 22936
rect 4580 22924 4586 22976
rect 6687 22967 6745 22973
rect 6687 22933 6699 22967
rect 6733 22964 6745 22967
rect 7926 22964 7932 22976
rect 6733 22936 7932 22964
rect 6733 22933 6745 22936
rect 6687 22927 6745 22933
rect 7926 22924 7932 22936
rect 7984 22924 7990 22976
rect 8570 22924 8576 22976
rect 8628 22964 8634 22976
rect 12986 22964 12992 22976
rect 8628 22936 12992 22964
rect 8628 22924 8634 22936
rect 12986 22924 12992 22936
rect 13044 22924 13050 22976
rect 14182 22924 14188 22976
rect 14240 22964 14246 22976
rect 14461 22967 14519 22973
rect 14461 22964 14473 22967
rect 14240 22936 14473 22964
rect 14240 22924 14246 22936
rect 14461 22933 14473 22936
rect 14507 22933 14519 22967
rect 14461 22927 14519 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 2498 22760 2504 22772
rect 2459 22732 2504 22760
rect 2498 22720 2504 22732
rect 2556 22720 2562 22772
rect 3605 22763 3663 22769
rect 3605 22729 3617 22763
rect 3651 22760 3663 22763
rect 3835 22763 3893 22769
rect 3835 22760 3847 22763
rect 3651 22732 3847 22760
rect 3651 22729 3663 22732
rect 3605 22723 3663 22729
rect 3835 22729 3847 22732
rect 3881 22760 3893 22763
rect 4706 22760 4712 22772
rect 3881 22732 4712 22760
rect 3881 22729 3893 22732
rect 3835 22723 3893 22729
rect 4706 22720 4712 22732
rect 4764 22720 4770 22772
rect 6270 22760 6276 22772
rect 6231 22732 6276 22760
rect 6270 22720 6276 22732
rect 6328 22720 6334 22772
rect 7374 22720 7380 22772
rect 7432 22760 7438 22772
rect 7745 22763 7803 22769
rect 7745 22760 7757 22763
rect 7432 22732 7757 22760
rect 7432 22720 7438 22732
rect 7745 22729 7757 22732
rect 7791 22729 7803 22763
rect 8110 22760 8116 22772
rect 8071 22732 8116 22760
rect 7745 22723 7803 22729
rect 8110 22720 8116 22732
rect 8168 22720 8174 22772
rect 9769 22763 9827 22769
rect 9769 22729 9781 22763
rect 9815 22760 9827 22763
rect 10778 22760 10784 22772
rect 9815 22732 10784 22760
rect 9815 22729 9827 22732
rect 9769 22723 9827 22729
rect 10778 22720 10784 22732
rect 10836 22720 10842 22772
rect 11514 22760 11520 22772
rect 11475 22732 11520 22760
rect 11514 22720 11520 22732
rect 11572 22720 11578 22772
rect 12253 22763 12311 22769
rect 12253 22729 12265 22763
rect 12299 22760 12311 22763
rect 12342 22760 12348 22772
rect 12299 22732 12348 22760
rect 12299 22729 12311 22732
rect 12253 22723 12311 22729
rect 12342 22720 12348 22732
rect 12400 22760 12406 22772
rect 13725 22763 13783 22769
rect 12400 22732 12756 22760
rect 12400 22720 12406 22732
rect 4522 22652 4528 22704
rect 4580 22692 4586 22704
rect 12728 22701 12756 22732
rect 13725 22729 13737 22763
rect 13771 22760 13783 22763
rect 14093 22763 14151 22769
rect 14093 22760 14105 22763
rect 13771 22732 14105 22760
rect 13771 22729 13783 22732
rect 13725 22723 13783 22729
rect 14093 22729 14105 22732
rect 14139 22760 14151 22763
rect 14458 22760 14464 22772
rect 14139 22732 14464 22760
rect 14139 22729 14151 22732
rect 14093 22723 14151 22729
rect 14458 22720 14464 22732
rect 14516 22720 14522 22772
rect 22465 22763 22523 22769
rect 22465 22729 22477 22763
rect 22511 22760 22523 22763
rect 23934 22760 23940 22772
rect 22511 22732 23940 22760
rect 22511 22729 22523 22732
rect 22465 22723 22523 22729
rect 23934 22720 23940 22732
rect 23992 22720 23998 22772
rect 5629 22695 5687 22701
rect 5629 22692 5641 22695
rect 4580 22664 5641 22692
rect 4580 22652 4586 22664
rect 5629 22661 5641 22664
rect 5675 22661 5687 22695
rect 5629 22655 5687 22661
rect 12713 22695 12771 22701
rect 12713 22661 12725 22695
rect 12759 22661 12771 22695
rect 12713 22655 12771 22661
rect 12802 22652 12808 22704
rect 12860 22692 12866 22704
rect 14274 22692 14280 22704
rect 12860 22664 14280 22692
rect 12860 22652 12866 22664
rect 14274 22652 14280 22664
rect 14332 22652 14338 22704
rect 14734 22652 14740 22704
rect 14792 22692 14798 22704
rect 15933 22695 15991 22701
rect 15933 22692 15945 22695
rect 14792 22664 15945 22692
rect 14792 22652 14798 22664
rect 15933 22661 15945 22664
rect 15979 22661 15991 22695
rect 15933 22655 15991 22661
rect 1118 22584 1124 22636
rect 1176 22624 1182 22636
rect 1176 22596 3775 22624
rect 1176 22584 1182 22596
rect 1394 22556 1400 22568
rect 1355 22528 1400 22556
rect 1394 22516 1400 22528
rect 1452 22556 1458 22568
rect 1949 22559 2007 22565
rect 1949 22556 1961 22559
rect 1452 22528 1961 22556
rect 1452 22516 1458 22528
rect 1949 22525 1961 22528
rect 1995 22525 2007 22559
rect 1949 22519 2007 22525
rect 2685 22559 2743 22565
rect 2685 22525 2697 22559
rect 2731 22556 2743 22559
rect 3418 22556 3424 22568
rect 2731 22528 3424 22556
rect 2731 22525 2743 22528
rect 2685 22519 2743 22525
rect 3418 22516 3424 22528
rect 3476 22516 3482 22568
rect 3747 22565 3775 22596
rect 10410 22584 10416 22636
rect 10468 22624 10474 22636
rect 10965 22627 11023 22633
rect 10965 22624 10977 22627
rect 10468 22596 10977 22624
rect 10468 22584 10474 22596
rect 10965 22593 10977 22596
rect 11011 22624 11023 22627
rect 12250 22624 12256 22636
rect 11011 22596 12256 22624
rect 11011 22593 11023 22596
rect 10965 22587 11023 22593
rect 12250 22584 12256 22596
rect 12308 22584 12314 22636
rect 13446 22584 13452 22636
rect 13504 22624 13510 22636
rect 14645 22627 14703 22633
rect 14645 22624 14657 22627
rect 13504 22596 14657 22624
rect 13504 22584 13510 22596
rect 14645 22593 14657 22596
rect 14691 22593 14703 22627
rect 14645 22587 14703 22593
rect 3732 22559 3790 22565
rect 3732 22525 3744 22559
rect 3778 22556 3790 22559
rect 4246 22556 4252 22568
rect 3778 22528 4252 22556
rect 3778 22525 3790 22528
rect 3732 22519 3790 22525
rect 4246 22516 4252 22528
rect 4304 22516 4310 22568
rect 4706 22556 4712 22568
rect 4667 22528 4712 22556
rect 4706 22516 4712 22528
rect 4764 22516 4770 22568
rect 6825 22559 6883 22565
rect 6825 22525 6837 22559
rect 6871 22556 6883 22559
rect 6914 22556 6920 22568
rect 6871 22528 6920 22556
rect 6871 22525 6883 22528
rect 6825 22519 6883 22525
rect 6914 22516 6920 22528
rect 6972 22516 6978 22568
rect 8573 22559 8631 22565
rect 8573 22525 8585 22559
rect 8619 22556 8631 22559
rect 9306 22556 9312 22568
rect 8619 22528 9312 22556
rect 8619 22525 8631 22528
rect 8573 22519 8631 22525
rect 9306 22516 9312 22528
rect 9364 22516 9370 22568
rect 12618 22556 12624 22568
rect 12579 22528 12624 22556
rect 12618 22516 12624 22528
rect 12676 22516 12682 22568
rect 12894 22556 12900 22568
rect 12855 22528 12900 22556
rect 12894 22516 12900 22528
rect 12952 22516 12958 22568
rect 14182 22556 14188 22568
rect 14143 22528 14188 22556
rect 14182 22516 14188 22528
rect 14240 22516 14246 22568
rect 14274 22516 14280 22568
rect 14332 22556 14338 22568
rect 14458 22556 14464 22568
rect 14332 22528 14377 22556
rect 14419 22528 14464 22556
rect 14332 22516 14338 22528
rect 14458 22516 14464 22528
rect 14516 22516 14522 22568
rect 15749 22559 15807 22565
rect 15749 22525 15761 22559
rect 15795 22525 15807 22559
rect 15749 22519 15807 22525
rect 4338 22488 4344 22500
rect 3068 22460 4344 22488
rect 106 22380 112 22432
rect 164 22420 170 22432
rect 1581 22423 1639 22429
rect 1581 22420 1593 22423
rect 164 22392 1593 22420
rect 164 22380 170 22392
rect 1581 22389 1593 22392
rect 1627 22389 1639 22423
rect 1581 22383 1639 22389
rect 2869 22423 2927 22429
rect 2869 22389 2881 22423
rect 2915 22420 2927 22423
rect 3068 22420 3096 22460
rect 4338 22448 4344 22460
rect 4396 22448 4402 22500
rect 4430 22448 4436 22500
rect 4488 22488 4494 22500
rect 4617 22491 4675 22497
rect 4617 22488 4629 22491
rect 4488 22460 4629 22488
rect 4488 22448 4494 22460
rect 4617 22457 4629 22460
rect 4663 22488 4675 22491
rect 5071 22491 5129 22497
rect 5071 22488 5083 22491
rect 4663 22460 5083 22488
rect 4663 22457 4675 22460
rect 4617 22451 4675 22457
rect 5071 22457 5083 22460
rect 5117 22488 5129 22491
rect 6641 22491 6699 22497
rect 6641 22488 6653 22491
rect 5117 22460 6653 22488
rect 5117 22457 5129 22460
rect 5071 22451 5129 22457
rect 6641 22457 6653 22460
rect 6687 22488 6699 22491
rect 7187 22491 7245 22497
rect 7187 22488 7199 22491
rect 6687 22460 7199 22488
rect 6687 22457 6699 22460
rect 6641 22451 6699 22457
rect 7187 22457 7199 22460
rect 7233 22488 7245 22491
rect 8018 22488 8024 22500
rect 7233 22460 8024 22488
rect 7233 22457 7245 22460
rect 7187 22451 7245 22457
rect 8018 22448 8024 22460
rect 8076 22448 8082 22500
rect 9401 22491 9459 22497
rect 9401 22457 9413 22491
rect 9447 22488 9459 22491
rect 10045 22491 10103 22497
rect 10045 22488 10057 22491
rect 9447 22460 10057 22488
rect 9447 22457 9459 22460
rect 9401 22451 9459 22457
rect 10045 22457 10057 22460
rect 10091 22457 10103 22491
rect 10045 22451 10103 22457
rect 2915 22392 3096 22420
rect 3237 22423 3295 22429
rect 2915 22389 2927 22392
rect 2869 22383 2927 22389
rect 3237 22389 3249 22423
rect 3283 22420 3295 22423
rect 3418 22420 3424 22432
rect 3283 22392 3424 22420
rect 3283 22389 3295 22392
rect 3237 22383 3295 22389
rect 3418 22380 3424 22392
rect 3476 22380 3482 22432
rect 4246 22420 4252 22432
rect 4159 22392 4252 22420
rect 4246 22380 4252 22392
rect 4304 22420 4310 22432
rect 6086 22420 6092 22432
rect 4304 22392 6092 22420
rect 4304 22380 4310 22392
rect 6086 22380 6092 22392
rect 6144 22380 6150 22432
rect 10060 22420 10088 22451
rect 10134 22448 10140 22500
rect 10192 22488 10198 22500
rect 10321 22491 10379 22497
rect 10321 22488 10333 22491
rect 10192 22460 10333 22488
rect 10192 22448 10198 22460
rect 10321 22457 10333 22460
rect 10367 22457 10379 22491
rect 10321 22451 10379 22457
rect 10413 22491 10471 22497
rect 10413 22457 10425 22491
rect 10459 22457 10471 22491
rect 10413 22451 10471 22457
rect 11885 22491 11943 22497
rect 11885 22457 11897 22491
rect 11931 22488 11943 22491
rect 12912 22488 12940 22516
rect 11931 22460 12940 22488
rect 13357 22491 13415 22497
rect 11931 22457 11943 22460
rect 11885 22451 11943 22457
rect 13357 22457 13369 22491
rect 13403 22488 13415 22491
rect 15764 22488 15792 22519
rect 16390 22516 16396 22568
rect 16448 22556 16454 22568
rect 16796 22559 16854 22565
rect 16796 22556 16808 22559
rect 16448 22528 16808 22556
rect 16448 22516 16454 22528
rect 16796 22525 16808 22528
rect 16842 22556 16854 22559
rect 17221 22559 17279 22565
rect 17221 22556 17233 22559
rect 16842 22528 17233 22556
rect 16842 22525 16854 22528
rect 16796 22519 16854 22525
rect 17221 22525 17233 22528
rect 17267 22525 17279 22559
rect 22278 22556 22284 22568
rect 22239 22528 22284 22556
rect 17221 22519 17279 22525
rect 22278 22516 22284 22528
rect 22336 22556 22342 22568
rect 22833 22559 22891 22565
rect 22833 22556 22845 22559
rect 22336 22528 22845 22556
rect 22336 22516 22342 22528
rect 22833 22525 22845 22528
rect 22879 22525 22891 22559
rect 22833 22519 22891 22525
rect 16209 22491 16267 22497
rect 16209 22488 16221 22491
rect 13403 22460 16221 22488
rect 13403 22457 13415 22460
rect 13357 22451 13415 22457
rect 16209 22457 16221 22460
rect 16255 22457 16267 22491
rect 16209 22451 16267 22457
rect 10428 22420 10456 22451
rect 15286 22420 15292 22432
rect 10060 22392 10456 22420
rect 15247 22392 15292 22420
rect 15286 22380 15292 22392
rect 15344 22380 15350 22432
rect 16022 22380 16028 22432
rect 16080 22420 16086 22432
rect 16899 22423 16957 22429
rect 16899 22420 16911 22423
rect 16080 22392 16911 22420
rect 16080 22380 16086 22392
rect 16899 22389 16911 22392
rect 16945 22389 16957 22423
rect 16899 22383 16957 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1578 22216 1584 22228
rect 1539 22188 1584 22216
rect 1578 22176 1584 22188
rect 1636 22176 1642 22228
rect 5442 22216 5448 22228
rect 5403 22188 5448 22216
rect 5442 22176 5448 22188
rect 5500 22176 5506 22228
rect 6687 22219 6745 22225
rect 6687 22185 6699 22219
rect 6733 22216 6745 22219
rect 7006 22216 7012 22228
rect 6733 22188 7012 22216
rect 6733 22185 6745 22188
rect 6687 22179 6745 22185
rect 7006 22176 7012 22188
rect 7064 22176 7070 22228
rect 7466 22216 7472 22228
rect 7427 22188 7472 22216
rect 7466 22176 7472 22188
rect 7524 22176 7530 22228
rect 8110 22176 8116 22228
rect 8168 22216 8174 22228
rect 8481 22219 8539 22225
rect 8481 22216 8493 22219
rect 8168 22188 8493 22216
rect 8168 22176 8174 22188
rect 8481 22185 8493 22188
rect 8527 22185 8539 22219
rect 8481 22179 8539 22185
rect 9950 22176 9956 22228
rect 10008 22216 10014 22228
rect 10045 22219 10103 22225
rect 10045 22216 10057 22219
rect 10008 22188 10057 22216
rect 10008 22176 10014 22188
rect 10045 22185 10057 22188
rect 10091 22185 10103 22219
rect 10045 22179 10103 22185
rect 10134 22176 10140 22228
rect 10192 22216 10198 22228
rect 10965 22219 11023 22225
rect 10965 22216 10977 22219
rect 10192 22188 10977 22216
rect 10192 22176 10198 22188
rect 10965 22185 10977 22188
rect 11011 22216 11023 22219
rect 12158 22216 12164 22228
rect 11011 22188 12164 22216
rect 11011 22185 11023 22188
rect 10965 22179 11023 22185
rect 12158 22176 12164 22188
rect 12216 22176 12222 22228
rect 14274 22176 14280 22228
rect 14332 22216 14338 22228
rect 14645 22219 14703 22225
rect 14645 22216 14657 22219
rect 14332 22188 14657 22216
rect 14332 22176 14338 22188
rect 14645 22185 14657 22188
rect 14691 22185 14703 22219
rect 14645 22179 14703 22185
rect 17451 22219 17509 22225
rect 17451 22185 17463 22219
rect 17497 22216 17509 22219
rect 22278 22216 22284 22228
rect 17497 22188 22284 22216
rect 17497 22185 17509 22188
rect 17451 22179 17509 22185
rect 22278 22176 22284 22188
rect 22336 22176 22342 22228
rect 4430 22108 4436 22160
rect 4488 22148 4494 22160
rect 4846 22151 4904 22157
rect 4846 22148 4858 22151
rect 4488 22120 4858 22148
rect 4488 22108 4494 22120
rect 4846 22117 4858 22120
rect 4892 22117 4904 22151
rect 4846 22111 4904 22117
rect 7923 22151 7981 22157
rect 7923 22117 7935 22151
rect 7969 22148 7981 22151
rect 8018 22148 8024 22160
rect 7969 22120 8024 22148
rect 7969 22117 7981 22120
rect 7923 22111 7981 22117
rect 8018 22108 8024 22120
rect 8076 22108 8082 22160
rect 12066 22148 12072 22160
rect 12027 22120 12072 22148
rect 12066 22108 12072 22120
rect 12124 22108 12130 22160
rect 15194 22108 15200 22160
rect 15252 22148 15258 22160
rect 15473 22151 15531 22157
rect 15473 22148 15485 22151
rect 15252 22120 15485 22148
rect 15252 22108 15258 22120
rect 15473 22117 15485 22120
rect 15519 22117 15531 22151
rect 15473 22111 15531 22117
rect 1397 22083 1455 22089
rect 1397 22049 1409 22083
rect 1443 22080 1455 22083
rect 2038 22080 2044 22092
rect 1443 22052 2044 22080
rect 1443 22049 1455 22052
rect 1397 22043 1455 22049
rect 2038 22040 2044 22052
rect 2096 22040 2102 22092
rect 2314 22040 2320 22092
rect 2372 22080 2378 22092
rect 6546 22080 6552 22092
rect 2372 22052 6552 22080
rect 2372 22040 2378 22052
rect 6546 22040 6552 22052
rect 6604 22040 6610 22092
rect 11238 22040 11244 22092
rect 11296 22080 11302 22092
rect 11517 22083 11575 22089
rect 11517 22080 11529 22083
rect 11296 22052 11529 22080
rect 11296 22040 11302 22052
rect 11517 22049 11529 22052
rect 11563 22049 11575 22083
rect 12618 22080 12624 22092
rect 12579 22052 12624 22080
rect 11517 22043 11575 22049
rect 12618 22040 12624 22052
rect 12676 22040 12682 22092
rect 12710 22040 12716 22092
rect 12768 22080 12774 22092
rect 12894 22080 12900 22092
rect 12768 22052 12813 22080
rect 12855 22052 12900 22080
rect 12768 22040 12774 22052
rect 12894 22040 12900 22052
rect 12952 22040 12958 22092
rect 13078 22040 13084 22092
rect 13136 22080 13142 22092
rect 14252 22083 14310 22089
rect 14252 22080 14264 22083
rect 13136 22052 14264 22080
rect 13136 22040 13142 22052
rect 14252 22049 14264 22052
rect 14298 22080 14310 22083
rect 14642 22080 14648 22092
rect 14298 22052 14648 22080
rect 14298 22049 14310 22052
rect 14252 22043 14310 22049
rect 14642 22040 14648 22052
rect 14700 22040 14706 22092
rect 2498 22012 2504 22024
rect 2459 21984 2504 22012
rect 2498 21972 2504 21984
rect 2556 21972 2562 22024
rect 4525 22015 4583 22021
rect 4525 21981 4537 22015
rect 4571 22012 4583 22015
rect 4614 22012 4620 22024
rect 4571 21984 4620 22012
rect 4571 21981 4583 21984
rect 4525 21975 4583 21981
rect 4614 21972 4620 21984
rect 4672 21972 4678 22024
rect 7282 21972 7288 22024
rect 7340 22012 7346 22024
rect 7561 22015 7619 22021
rect 7561 22012 7573 22015
rect 7340 21984 7573 22012
rect 7340 21972 7346 21984
rect 7561 21981 7573 21984
rect 7607 21981 7619 22015
rect 7561 21975 7619 21981
rect 9677 22015 9735 22021
rect 9677 21981 9689 22015
rect 9723 22012 9735 22015
rect 11146 22012 11152 22024
rect 9723 21984 11152 22012
rect 9723 21981 9735 21984
rect 9677 21975 9735 21981
rect 11146 21972 11152 21984
rect 11204 21972 11210 22024
rect 13354 22012 13360 22024
rect 13315 21984 13360 22012
rect 13354 21972 13360 21984
rect 13412 21972 13418 22024
rect 13725 22015 13783 22021
rect 13725 21981 13737 22015
rect 13771 22012 13783 22015
rect 13814 22012 13820 22024
rect 13771 21984 13820 22012
rect 13771 21981 13783 21984
rect 13725 21975 13783 21981
rect 13814 21972 13820 21984
rect 13872 21972 13878 22024
rect 14458 21972 14464 22024
rect 14516 22012 14522 22024
rect 15378 22012 15384 22024
rect 14516 21984 15384 22012
rect 14516 21972 14522 21984
rect 15378 21972 15384 21984
rect 15436 21972 15442 22024
rect 15838 22012 15844 22024
rect 15799 21984 15844 22012
rect 15838 21972 15844 21984
rect 15896 21972 15902 22024
rect 9306 21904 9312 21956
rect 9364 21944 9370 21956
rect 10597 21947 10655 21953
rect 10597 21944 10609 21947
rect 9364 21916 10609 21944
rect 9364 21904 9370 21916
rect 10597 21913 10609 21916
rect 10643 21944 10655 21947
rect 11514 21944 11520 21956
rect 10643 21916 11520 21944
rect 10643 21913 10655 21916
rect 10597 21907 10655 21913
rect 11514 21904 11520 21916
rect 11572 21904 11578 21956
rect 2038 21876 2044 21888
rect 1999 21848 2044 21876
rect 2038 21836 2044 21848
rect 2096 21836 2102 21888
rect 3234 21876 3240 21888
rect 3195 21848 3240 21876
rect 3234 21836 3240 21848
rect 3292 21836 3298 21888
rect 4433 21879 4491 21885
rect 4433 21845 4445 21879
rect 4479 21876 4491 21879
rect 4706 21876 4712 21888
rect 4479 21848 4712 21876
rect 4479 21845 4491 21848
rect 4433 21839 4491 21845
rect 4706 21836 4712 21848
rect 4764 21876 4770 21888
rect 6270 21876 6276 21888
rect 4764 21848 6276 21876
rect 4764 21836 4770 21848
rect 6270 21836 6276 21848
rect 6328 21836 6334 21888
rect 6914 21836 6920 21888
rect 6972 21876 6978 21888
rect 7009 21879 7067 21885
rect 7009 21876 7021 21879
rect 6972 21848 7021 21876
rect 6972 21836 6978 21848
rect 7009 21845 7021 21848
rect 7055 21845 7067 21879
rect 7009 21839 7067 21845
rect 9493 21879 9551 21885
rect 9493 21845 9505 21879
rect 9539 21876 9551 21879
rect 9766 21876 9772 21888
rect 9539 21848 9772 21876
rect 9539 21845 9551 21848
rect 9493 21839 9551 21845
rect 9766 21836 9772 21848
rect 9824 21836 9830 21888
rect 11698 21876 11704 21888
rect 11659 21848 11704 21876
rect 11698 21836 11704 21848
rect 11756 21836 11762 21888
rect 13722 21836 13728 21888
rect 13780 21876 13786 21888
rect 14093 21879 14151 21885
rect 14093 21876 14105 21879
rect 13780 21848 14105 21876
rect 13780 21836 13786 21848
rect 14093 21845 14105 21848
rect 14139 21876 14151 21879
rect 14323 21879 14381 21885
rect 14323 21876 14335 21879
rect 14139 21848 14335 21876
rect 14139 21845 14151 21848
rect 14093 21839 14151 21845
rect 14323 21845 14335 21848
rect 14369 21845 14381 21879
rect 14323 21839 14381 21845
rect 16850 21836 16856 21888
rect 16908 21876 16914 21888
rect 17221 21879 17279 21885
rect 17221 21876 17233 21879
rect 16908 21848 17233 21876
rect 16908 21836 16914 21848
rect 17221 21845 17233 21848
rect 17267 21845 17279 21879
rect 17221 21839 17279 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 2498 21672 2504 21684
rect 2459 21644 2504 21672
rect 2498 21632 2504 21644
rect 2556 21632 2562 21684
rect 4430 21632 4436 21684
rect 4488 21672 4494 21684
rect 4525 21675 4583 21681
rect 4525 21672 4537 21675
rect 4488 21644 4537 21672
rect 4488 21632 4494 21644
rect 4525 21641 4537 21644
rect 4571 21641 4583 21675
rect 4525 21635 4583 21641
rect 4798 21632 4804 21684
rect 4856 21672 4862 21684
rect 4985 21675 5043 21681
rect 4985 21672 4997 21675
rect 4856 21644 4997 21672
rect 4856 21632 4862 21644
rect 4985 21641 4997 21644
rect 5031 21641 5043 21675
rect 4985 21635 5043 21641
rect 8481 21675 8539 21681
rect 8481 21641 8493 21675
rect 8527 21672 8539 21675
rect 8570 21672 8576 21684
rect 8527 21644 8576 21672
rect 8527 21641 8539 21644
rect 8481 21635 8539 21641
rect 1489 21539 1547 21545
rect 1489 21505 1501 21539
rect 1535 21536 1547 21539
rect 2516 21536 2544 21632
rect 8496 21604 8524 21635
rect 8570 21632 8576 21644
rect 8628 21632 8634 21684
rect 10505 21675 10563 21681
rect 10505 21641 10517 21675
rect 10551 21672 10563 21675
rect 10778 21672 10784 21684
rect 10551 21644 10784 21672
rect 10551 21641 10563 21644
rect 10505 21635 10563 21641
rect 10778 21632 10784 21644
rect 10836 21632 10842 21684
rect 12759 21675 12817 21681
rect 12759 21641 12771 21675
rect 12805 21672 12817 21675
rect 14458 21672 14464 21684
rect 12805 21644 14464 21672
rect 12805 21641 12817 21644
rect 12759 21635 12817 21641
rect 14458 21632 14464 21644
rect 14516 21632 14522 21684
rect 14642 21672 14648 21684
rect 14603 21644 14648 21672
rect 14642 21632 14648 21644
rect 14700 21632 14706 21684
rect 14826 21632 14832 21684
rect 14884 21672 14890 21684
rect 15105 21675 15163 21681
rect 15105 21672 15117 21675
rect 14884 21644 15117 21672
rect 14884 21632 14890 21644
rect 15105 21641 15117 21644
rect 15151 21672 15163 21675
rect 15286 21672 15292 21684
rect 15151 21644 15292 21672
rect 15151 21641 15163 21644
rect 15105 21635 15163 21641
rect 15286 21632 15292 21644
rect 15344 21632 15350 21684
rect 15378 21632 15384 21684
rect 15436 21672 15442 21684
rect 16209 21675 16267 21681
rect 16209 21672 16221 21675
rect 15436 21644 16221 21672
rect 15436 21632 15442 21644
rect 16209 21641 16221 21644
rect 16255 21641 16267 21675
rect 16209 21635 16267 21641
rect 24121 21675 24179 21681
rect 24121 21641 24133 21675
rect 24167 21672 24179 21675
rect 25866 21672 25872 21684
rect 24167 21644 25872 21672
rect 24167 21641 24179 21644
rect 24121 21635 24179 21641
rect 25866 21632 25872 21644
rect 25924 21632 25930 21684
rect 1535 21508 2544 21536
rect 7576 21576 8524 21604
rect 9493 21607 9551 21613
rect 1535 21505 1547 21508
rect 1489 21499 1547 21505
rect 4157 21471 4215 21477
rect 4157 21437 4169 21471
rect 4203 21468 4215 21471
rect 4522 21468 4528 21480
rect 4203 21440 4528 21468
rect 4203 21437 4215 21440
rect 4157 21431 4215 21437
rect 4522 21428 4528 21440
rect 4580 21468 4586 21480
rect 7576 21477 7604 21576
rect 9493 21573 9505 21607
rect 9539 21604 9551 21607
rect 9950 21604 9956 21616
rect 9539 21576 9956 21604
rect 9539 21573 9551 21576
rect 9493 21567 9551 21573
rect 9950 21564 9956 21576
rect 10008 21604 10014 21616
rect 10873 21607 10931 21613
rect 10873 21604 10885 21607
rect 10008 21576 10885 21604
rect 10008 21564 10014 21576
rect 10873 21573 10885 21576
rect 10919 21573 10931 21607
rect 10873 21567 10931 21573
rect 12618 21564 12624 21616
rect 12676 21564 12682 21616
rect 13354 21564 13360 21616
rect 13412 21604 13418 21616
rect 13412 21576 16804 21604
rect 13412 21564 13418 21576
rect 8478 21496 8484 21548
rect 8536 21536 8542 21548
rect 12636 21536 12664 21564
rect 13449 21539 13507 21545
rect 13449 21536 13461 21539
rect 8536 21508 12525 21536
rect 12636 21508 13461 21536
rect 8536 21496 8542 21508
rect 4801 21471 4859 21477
rect 4801 21468 4813 21471
rect 4580 21440 4813 21468
rect 4580 21428 4586 21440
rect 4801 21437 4813 21440
rect 4847 21437 4859 21471
rect 4801 21431 4859 21437
rect 7561 21471 7619 21477
rect 7561 21437 7573 21471
rect 7607 21437 7619 21471
rect 7561 21431 7619 21437
rect 8573 21471 8631 21477
rect 8573 21437 8585 21471
rect 8619 21468 8631 21471
rect 9033 21471 9091 21477
rect 9033 21468 9045 21471
rect 8619 21440 9045 21468
rect 8619 21437 8631 21440
rect 8573 21431 8631 21437
rect 9033 21437 9045 21440
rect 9079 21468 9091 21471
rect 9490 21468 9496 21480
rect 9079 21440 9496 21468
rect 9079 21437 9091 21440
rect 9033 21431 9091 21437
rect 9490 21428 9496 21440
rect 9548 21428 9554 21480
rect 9585 21471 9643 21477
rect 9585 21437 9597 21471
rect 9631 21468 9643 21471
rect 9766 21468 9772 21480
rect 9631 21440 9772 21468
rect 9631 21437 9643 21440
rect 9585 21431 9643 21437
rect 9766 21428 9772 21440
rect 9824 21428 9830 21480
rect 11333 21471 11391 21477
rect 11333 21437 11345 21471
rect 11379 21468 11391 21471
rect 11790 21468 11796 21480
rect 11379 21440 11796 21468
rect 11379 21437 11391 21440
rect 11333 21431 11391 21437
rect 11790 21428 11796 21440
rect 11848 21428 11854 21480
rect 12497 21468 12525 21508
rect 13449 21505 13461 21508
rect 13495 21505 13507 21539
rect 13722 21536 13728 21548
rect 13683 21508 13728 21536
rect 13449 21499 13507 21505
rect 13722 21496 13728 21508
rect 13780 21496 13786 21548
rect 15289 21539 15347 21545
rect 15289 21505 15301 21539
rect 15335 21536 15347 21539
rect 16574 21536 16580 21548
rect 15335 21508 16580 21536
rect 15335 21505 15347 21508
rect 15289 21499 15347 21505
rect 16574 21496 16580 21508
rect 16632 21496 16638 21548
rect 16776 21477 16804 21576
rect 12656 21471 12714 21477
rect 12656 21468 12668 21471
rect 12497 21440 12668 21468
rect 12656 21437 12668 21440
rect 12702 21468 12714 21471
rect 13081 21471 13139 21477
rect 13081 21468 13093 21471
rect 12702 21440 13093 21468
rect 12702 21437 12714 21440
rect 12656 21431 12714 21437
rect 13081 21437 13093 21440
rect 13127 21437 13139 21471
rect 13081 21431 13139 21437
rect 16761 21471 16819 21477
rect 16761 21437 16773 21471
rect 16807 21468 16819 21471
rect 17221 21471 17279 21477
rect 17221 21468 17233 21471
rect 16807 21440 17233 21468
rect 16807 21437 16819 21440
rect 16761 21431 16819 21437
rect 17221 21437 17233 21440
rect 17267 21437 17279 21471
rect 23934 21468 23940 21480
rect 23895 21440 23940 21468
rect 17221 21431 17279 21437
rect 23934 21428 23940 21440
rect 23992 21468 23998 21480
rect 24489 21471 24547 21477
rect 24489 21468 24501 21471
rect 23992 21440 24501 21468
rect 23992 21428 23998 21440
rect 24489 21437 24501 21440
rect 24535 21437 24547 21471
rect 24489 21431 24547 21437
rect 1578 21360 1584 21412
rect 1636 21400 1642 21412
rect 2133 21403 2191 21409
rect 1636 21372 1681 21400
rect 1636 21360 1642 21372
rect 2133 21369 2145 21403
rect 2179 21400 2191 21403
rect 2958 21400 2964 21412
rect 2179 21372 2964 21400
rect 2179 21369 2191 21372
rect 2133 21363 2191 21369
rect 2958 21360 2964 21372
rect 3016 21360 3022 21412
rect 3234 21400 3240 21412
rect 3195 21372 3240 21400
rect 3234 21360 3240 21372
rect 3292 21360 3298 21412
rect 3326 21360 3332 21412
rect 3384 21400 3390 21412
rect 3881 21403 3939 21409
rect 3384 21372 3429 21400
rect 3384 21360 3390 21372
rect 3881 21369 3893 21403
rect 3927 21400 3939 21403
rect 4246 21400 4252 21412
rect 3927 21372 4252 21400
rect 3927 21369 3939 21372
rect 3881 21363 3939 21369
rect 4246 21360 4252 21372
rect 4304 21360 4310 21412
rect 4614 21360 4620 21412
rect 4672 21400 4678 21412
rect 5813 21403 5871 21409
rect 5813 21400 5825 21403
rect 4672 21372 5825 21400
rect 4672 21360 4678 21372
rect 5813 21369 5825 21372
rect 5859 21400 5871 21403
rect 6638 21400 6644 21412
rect 5859 21372 6644 21400
rect 5859 21369 5871 21372
rect 5813 21363 5871 21369
rect 6638 21360 6644 21372
rect 6696 21360 6702 21412
rect 8018 21360 8024 21412
rect 8076 21400 8082 21412
rect 8113 21403 8171 21409
rect 8113 21400 8125 21403
rect 8076 21372 8125 21400
rect 8076 21360 8082 21372
rect 8113 21369 8125 21372
rect 8159 21400 8171 21403
rect 8159 21372 9996 21400
rect 8159 21369 8171 21372
rect 8113 21363 8171 21369
rect 3053 21335 3111 21341
rect 3053 21301 3065 21335
rect 3099 21332 3111 21335
rect 3344 21332 3372 21360
rect 9968 21344 9996 21372
rect 11238 21360 11244 21412
rect 11296 21400 11302 21412
rect 12161 21403 12219 21409
rect 12161 21400 12173 21403
rect 11296 21372 12173 21400
rect 11296 21360 11302 21372
rect 12161 21369 12173 21372
rect 12207 21369 12219 21403
rect 12161 21363 12219 21369
rect 13814 21360 13820 21412
rect 13872 21400 13878 21412
rect 14366 21400 14372 21412
rect 13872 21372 13917 21400
rect 14327 21372 14372 21400
rect 13872 21360 13878 21372
rect 14366 21360 14372 21372
rect 14424 21360 14430 21412
rect 15378 21400 15384 21412
rect 15339 21372 15384 21400
rect 15378 21360 15384 21372
rect 15436 21360 15442 21412
rect 15654 21360 15660 21412
rect 15712 21400 15718 21412
rect 15933 21403 15991 21409
rect 15933 21400 15945 21403
rect 15712 21372 15945 21400
rect 15712 21360 15718 21372
rect 15933 21369 15945 21372
rect 15979 21369 15991 21403
rect 15933 21363 15991 21369
rect 16850 21360 16856 21412
rect 16908 21400 16914 21412
rect 17589 21403 17647 21409
rect 17589 21400 17601 21403
rect 16908 21372 17601 21400
rect 16908 21360 16914 21372
rect 17589 21369 17601 21372
rect 17635 21369 17647 21403
rect 17589 21363 17647 21369
rect 3099 21304 3372 21332
rect 3099 21301 3111 21304
rect 3053 21295 3111 21301
rect 3510 21292 3516 21344
rect 3568 21332 3574 21344
rect 4430 21332 4436 21344
rect 3568 21304 4436 21332
rect 3568 21292 3574 21304
rect 4430 21292 4436 21304
rect 4488 21292 4494 21344
rect 6546 21332 6552 21344
rect 6507 21304 6552 21332
rect 6546 21292 6552 21304
rect 6604 21292 6610 21344
rect 7101 21335 7159 21341
rect 7101 21301 7113 21335
rect 7147 21332 7159 21335
rect 7282 21332 7288 21344
rect 7147 21304 7288 21332
rect 7147 21301 7159 21304
rect 7101 21295 7159 21301
rect 7282 21292 7288 21304
rect 7340 21292 7346 21344
rect 7466 21332 7472 21344
rect 7427 21304 7472 21332
rect 7466 21292 7472 21304
rect 7524 21292 7530 21344
rect 7742 21332 7748 21344
rect 7703 21304 7748 21332
rect 7742 21292 7748 21304
rect 7800 21292 7806 21344
rect 8757 21335 8815 21341
rect 8757 21301 8769 21335
rect 8803 21332 8815 21335
rect 9122 21332 9128 21344
rect 8803 21304 9128 21332
rect 8803 21301 8815 21304
rect 8757 21295 8815 21301
rect 9122 21292 9128 21304
rect 9180 21292 9186 21344
rect 9950 21332 9956 21344
rect 9911 21304 9956 21332
rect 9950 21292 9956 21304
rect 10008 21292 10014 21344
rect 11146 21332 11152 21344
rect 11107 21304 11152 21332
rect 11146 21292 11152 21304
rect 11204 21292 11210 21344
rect 11514 21332 11520 21344
rect 11475 21304 11520 21332
rect 11514 21292 11520 21304
rect 11572 21292 11578 21344
rect 13832 21332 13860 21360
rect 14642 21332 14648 21344
rect 13832 21304 14648 21332
rect 14642 21292 14648 21304
rect 14700 21292 14706 21344
rect 16942 21332 16948 21344
rect 16903 21304 16948 21332
rect 16942 21292 16948 21304
rect 17000 21292 17006 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 3786 21128 3792 21140
rect 3747 21100 3792 21128
rect 3786 21088 3792 21100
rect 3844 21088 3850 21140
rect 4338 21088 4344 21140
rect 4396 21128 4402 21140
rect 5077 21131 5135 21137
rect 5077 21128 5089 21131
rect 4396 21100 5089 21128
rect 4396 21088 4402 21100
rect 5077 21097 5089 21100
rect 5123 21128 5135 21131
rect 6089 21131 6147 21137
rect 6089 21128 6101 21131
rect 5123 21100 6101 21128
rect 5123 21097 5135 21100
rect 5077 21091 5135 21097
rect 6089 21097 6101 21100
rect 6135 21097 6147 21131
rect 6914 21128 6920 21140
rect 6875 21100 6920 21128
rect 6089 21091 6147 21097
rect 2406 21060 2412 21072
rect 2367 21032 2412 21060
rect 2406 21020 2412 21032
rect 2464 21020 2470 21072
rect 2958 21060 2964 21072
rect 2919 21032 2964 21060
rect 2958 21020 2964 21032
rect 3016 21020 3022 21072
rect 4154 21020 4160 21072
rect 4212 21060 4218 21072
rect 4249 21063 4307 21069
rect 4249 21060 4261 21063
rect 4212 21032 4261 21060
rect 4212 21020 4218 21032
rect 4249 21029 4261 21032
rect 4295 21029 4307 21063
rect 4249 21023 4307 21029
rect 6104 20992 6132 21091
rect 6914 21088 6920 21100
rect 6972 21088 6978 21140
rect 9766 21128 9772 21140
rect 9727 21100 9772 21128
rect 9766 21088 9772 21100
rect 9824 21088 9830 21140
rect 12894 21088 12900 21140
rect 12952 21128 12958 21140
rect 12989 21131 13047 21137
rect 12989 21128 13001 21131
rect 12952 21100 13001 21128
rect 12952 21088 12958 21100
rect 12989 21097 13001 21100
rect 13035 21097 13047 21131
rect 12989 21091 13047 21097
rect 16574 21088 16580 21140
rect 16632 21128 16638 21140
rect 17451 21131 17509 21137
rect 17451 21128 17463 21131
rect 16632 21100 17463 21128
rect 16632 21088 16638 21100
rect 17451 21097 17463 21100
rect 17497 21097 17509 21131
rect 17451 21091 17509 21097
rect 9122 21060 9128 21072
rect 8036 21032 9128 21060
rect 6641 20995 6699 21001
rect 6641 20992 6653 20995
rect 6104 20964 6653 20992
rect 6641 20961 6653 20964
rect 6687 20992 6699 20995
rect 7006 20992 7012 21004
rect 6687 20964 7012 20992
rect 6687 20961 6699 20964
rect 6641 20955 6699 20961
rect 7006 20952 7012 20964
rect 7064 20952 7070 21004
rect 7377 20995 7435 21001
rect 7377 20961 7389 20995
rect 7423 20992 7435 20995
rect 7466 20992 7472 21004
rect 7423 20964 7472 20992
rect 7423 20961 7435 20964
rect 7377 20955 7435 20961
rect 7466 20952 7472 20964
rect 7524 20952 7530 21004
rect 7650 20992 7656 21004
rect 7611 20964 7656 20992
rect 7650 20952 7656 20964
rect 7708 20952 7714 21004
rect 8036 21001 8064 21032
rect 9122 21020 9128 21032
rect 9180 21020 9186 21072
rect 9214 21020 9220 21072
rect 9272 21060 9278 21072
rect 9493 21063 9551 21069
rect 9493 21060 9505 21063
rect 9272 21032 9505 21060
rect 9272 21020 9278 21032
rect 9493 21029 9505 21032
rect 9539 21060 9551 21063
rect 9539 21032 10364 21060
rect 9539 21029 9551 21032
rect 9493 21023 9551 21029
rect 10336 21004 10364 21032
rect 12710 21020 12716 21072
rect 12768 21060 12774 21072
rect 13357 21063 13415 21069
rect 13357 21060 13369 21063
rect 12768 21032 13369 21060
rect 12768 21020 12774 21032
rect 13357 21029 13369 21032
rect 13403 21029 13415 21063
rect 13357 21023 13415 21029
rect 13817 21063 13875 21069
rect 13817 21029 13829 21063
rect 13863 21060 13875 21063
rect 14182 21060 14188 21072
rect 13863 21032 14188 21060
rect 13863 21029 13875 21032
rect 13817 21023 13875 21029
rect 14182 21020 14188 21032
rect 14240 21020 14246 21072
rect 15930 21060 15936 21072
rect 15891 21032 15936 21060
rect 15930 21020 15936 21032
rect 15988 21020 15994 21072
rect 8021 20995 8079 21001
rect 8021 20961 8033 20995
rect 8067 20961 8079 20995
rect 8021 20955 8079 20961
rect 9030 20952 9036 21004
rect 9088 20992 9094 21004
rect 9677 20995 9735 21001
rect 9677 20992 9689 20995
rect 9088 20964 9689 20992
rect 9088 20952 9094 20964
rect 9677 20961 9689 20964
rect 9723 20961 9735 20995
rect 10318 20992 10324 21004
rect 10279 20964 10324 20992
rect 9677 20955 9735 20961
rect 2133 20927 2191 20933
rect 2133 20893 2145 20927
rect 2179 20924 2191 20927
rect 2317 20927 2375 20933
rect 2317 20924 2329 20927
rect 2179 20896 2329 20924
rect 2179 20893 2191 20896
rect 2133 20887 2191 20893
rect 2317 20893 2329 20896
rect 2363 20924 2375 20927
rect 2363 20896 3004 20924
rect 2363 20893 2375 20896
rect 2317 20887 2375 20893
rect 2976 20856 3004 20896
rect 3786 20884 3792 20936
rect 3844 20924 3850 20936
rect 4157 20927 4215 20933
rect 4157 20924 4169 20927
rect 3844 20896 4169 20924
rect 3844 20884 3850 20896
rect 4157 20893 4169 20896
rect 4203 20893 4215 20927
rect 4157 20887 4215 20893
rect 4246 20884 4252 20936
rect 4304 20924 4310 20936
rect 4433 20927 4491 20933
rect 4433 20924 4445 20927
rect 4304 20896 4445 20924
rect 4304 20884 4310 20896
rect 4433 20893 4445 20896
rect 4479 20893 4491 20927
rect 4433 20887 4491 20893
rect 5629 20927 5687 20933
rect 5629 20893 5641 20927
rect 5675 20924 5687 20927
rect 8478 20924 8484 20936
rect 5675 20896 8484 20924
rect 5675 20893 5687 20896
rect 5629 20887 5687 20893
rect 8478 20884 8484 20896
rect 8536 20884 8542 20936
rect 9692 20924 9720 20955
rect 10318 20952 10324 20964
rect 10376 20952 10382 21004
rect 10502 20992 10508 21004
rect 10463 20964 10508 20992
rect 10502 20952 10508 20964
rect 10560 20952 10566 21004
rect 10778 20952 10784 21004
rect 10836 20992 10842 21004
rect 10873 20995 10931 21001
rect 10873 20992 10885 20995
rect 10836 20964 10885 20992
rect 10836 20952 10842 20964
rect 10873 20961 10885 20964
rect 10919 20992 10931 20995
rect 11514 20992 11520 21004
rect 10919 20964 11520 20992
rect 10919 20961 10931 20964
rect 10873 20955 10931 20961
rect 11514 20952 11520 20964
rect 11572 20952 11578 21004
rect 12066 20992 12072 21004
rect 12027 20964 12072 20992
rect 12066 20952 12072 20964
rect 12124 20952 12130 21004
rect 17380 20995 17438 21001
rect 17380 20961 17392 20995
rect 17426 20992 17438 20995
rect 17494 20992 17500 21004
rect 17426 20964 17500 20992
rect 17426 20961 17438 20964
rect 17380 20955 17438 20961
rect 17494 20952 17500 20964
rect 17552 20952 17558 21004
rect 11425 20927 11483 20933
rect 11425 20924 11437 20927
rect 9692 20896 11437 20924
rect 11425 20893 11437 20896
rect 11471 20893 11483 20927
rect 11425 20887 11483 20893
rect 11606 20884 11612 20936
rect 11664 20924 11670 20936
rect 11977 20927 12035 20933
rect 11977 20924 11989 20927
rect 11664 20896 11989 20924
rect 11664 20884 11670 20896
rect 11977 20893 11989 20896
rect 12023 20893 12035 20927
rect 11977 20887 12035 20893
rect 13538 20884 13544 20936
rect 13596 20924 13602 20936
rect 13725 20927 13783 20933
rect 13725 20924 13737 20927
rect 13596 20896 13737 20924
rect 13596 20884 13602 20896
rect 13725 20893 13737 20896
rect 13771 20893 13783 20927
rect 14366 20924 14372 20936
rect 14279 20896 14372 20924
rect 13725 20887 13783 20893
rect 14366 20884 14372 20896
rect 14424 20924 14430 20936
rect 15838 20924 15844 20936
rect 14424 20896 15844 20924
rect 14424 20884 14430 20896
rect 15838 20884 15844 20896
rect 15896 20924 15902 20936
rect 16482 20924 16488 20936
rect 15896 20896 16488 20924
rect 15896 20884 15902 20896
rect 16482 20884 16488 20896
rect 16540 20884 16546 20936
rect 4264 20856 4292 20884
rect 2976 20828 4292 20856
rect 11698 20816 11704 20868
rect 11756 20856 11762 20868
rect 16393 20859 16451 20865
rect 11756 20828 13584 20856
rect 11756 20816 11762 20828
rect 1578 20788 1584 20800
rect 1539 20760 1584 20788
rect 1578 20748 1584 20760
rect 1636 20748 1642 20800
rect 1670 20748 1676 20800
rect 1728 20788 1734 20800
rect 2774 20788 2780 20800
rect 1728 20760 2780 20788
rect 1728 20748 1734 20760
rect 2774 20748 2780 20760
rect 2832 20788 2838 20800
rect 3237 20791 3295 20797
rect 3237 20788 3249 20791
rect 2832 20760 3249 20788
rect 2832 20748 2838 20760
rect 3237 20757 3249 20760
rect 3283 20757 3295 20791
rect 3237 20751 3295 20757
rect 6549 20791 6607 20797
rect 6549 20757 6561 20791
rect 6595 20788 6607 20791
rect 6822 20788 6828 20800
rect 6595 20760 6828 20788
rect 6595 20757 6607 20760
rect 6549 20751 6607 20757
rect 6822 20748 6828 20760
rect 6880 20748 6886 20800
rect 9030 20788 9036 20800
rect 8991 20760 9036 20788
rect 9030 20748 9036 20760
rect 9088 20748 9094 20800
rect 13556 20788 13584 20828
rect 16393 20825 16405 20859
rect 16439 20856 16451 20859
rect 16850 20856 16856 20868
rect 16439 20828 16856 20856
rect 16439 20825 16451 20828
rect 16393 20819 16451 20825
rect 16850 20816 16856 20828
rect 16908 20816 16914 20868
rect 13998 20788 14004 20800
rect 13556 20760 14004 20788
rect 13998 20748 14004 20760
rect 14056 20748 14062 20800
rect 14366 20748 14372 20800
rect 14424 20788 14430 20800
rect 15378 20788 15384 20800
rect 14424 20760 15384 20788
rect 14424 20748 14430 20760
rect 15378 20748 15384 20760
rect 15436 20788 15442 20800
rect 15473 20791 15531 20797
rect 15473 20788 15485 20791
rect 15436 20760 15485 20788
rect 15436 20748 15442 20760
rect 15473 20757 15485 20760
rect 15519 20757 15531 20791
rect 15473 20751 15531 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1394 20544 1400 20596
rect 1452 20584 1458 20596
rect 1535 20587 1593 20593
rect 1535 20584 1547 20587
rect 1452 20556 1547 20584
rect 1452 20544 1458 20556
rect 1535 20553 1547 20556
rect 1581 20553 1593 20587
rect 1535 20547 1593 20553
rect 10410 20544 10416 20596
rect 10468 20584 10474 20596
rect 12897 20587 12955 20593
rect 10468 20556 10640 20584
rect 10468 20544 10474 20556
rect 1949 20519 2007 20525
rect 1949 20485 1961 20519
rect 1995 20516 2007 20519
rect 2222 20516 2228 20528
rect 1995 20488 2228 20516
rect 1995 20485 2007 20488
rect 1949 20479 2007 20485
rect 2222 20476 2228 20488
rect 2280 20516 2286 20528
rect 2406 20516 2412 20528
rect 2280 20488 2412 20516
rect 2280 20476 2286 20488
rect 2406 20476 2412 20488
rect 2464 20516 2470 20528
rect 3329 20519 3387 20525
rect 3329 20516 3341 20519
rect 2464 20488 3341 20516
rect 2464 20476 2470 20488
rect 3329 20485 3341 20488
rect 3375 20485 3387 20519
rect 3329 20479 3387 20485
rect 4126 20488 5488 20516
rect 3973 20451 4031 20457
rect 3973 20417 3985 20451
rect 4019 20448 4031 20451
rect 4126 20448 4154 20488
rect 4019 20420 4154 20448
rect 4249 20451 4307 20457
rect 4019 20417 4031 20420
rect 3973 20411 4031 20417
rect 4249 20417 4261 20451
rect 4295 20448 4307 20451
rect 4295 20420 4936 20448
rect 4295 20417 4307 20420
rect 4249 20411 4307 20417
rect 4908 20392 4936 20420
rect 5460 20392 5488 20488
rect 7742 20476 7748 20528
rect 7800 20516 7806 20528
rect 9217 20519 9275 20525
rect 9217 20516 9229 20519
rect 7800 20488 9229 20516
rect 7800 20476 7806 20488
rect 9217 20485 9229 20488
rect 9263 20516 9275 20519
rect 10502 20516 10508 20528
rect 9263 20488 10508 20516
rect 9263 20485 9275 20488
rect 9217 20479 9275 20485
rect 10502 20476 10508 20488
rect 10560 20476 10566 20528
rect 10612 20516 10640 20556
rect 12897 20553 12909 20587
rect 12943 20584 12955 20587
rect 13538 20584 13544 20596
rect 12943 20556 13544 20584
rect 12943 20553 12955 20556
rect 12897 20547 12955 20553
rect 13538 20544 13544 20556
rect 13596 20544 13602 20596
rect 14829 20587 14887 20593
rect 14829 20553 14841 20587
rect 14875 20584 14887 20587
rect 15286 20584 15292 20596
rect 14875 20556 15292 20584
rect 14875 20553 14887 20556
rect 14829 20547 14887 20553
rect 15286 20544 15292 20556
rect 15344 20544 15350 20596
rect 15841 20587 15899 20593
rect 15841 20553 15853 20587
rect 15887 20584 15899 20587
rect 15930 20584 15936 20596
rect 15887 20556 15936 20584
rect 15887 20553 15899 20556
rect 15841 20547 15899 20553
rect 15930 20544 15936 20556
rect 15988 20584 15994 20596
rect 16117 20587 16175 20593
rect 16117 20584 16129 20587
rect 15988 20556 16129 20584
rect 15988 20544 15994 20556
rect 16117 20553 16129 20556
rect 16163 20553 16175 20587
rect 16482 20584 16488 20596
rect 16443 20556 16488 20584
rect 16117 20547 16175 20553
rect 16482 20544 16488 20556
rect 16540 20544 16546 20596
rect 18233 20519 18291 20525
rect 18233 20516 18245 20519
rect 10612 20488 18245 20516
rect 18233 20485 18245 20488
rect 18279 20485 18291 20519
rect 18233 20479 18291 20485
rect 7285 20451 7343 20457
rect 7285 20417 7297 20451
rect 7331 20448 7343 20451
rect 7331 20420 8800 20448
rect 7331 20417 7343 20420
rect 7285 20411 7343 20417
rect 1464 20383 1522 20389
rect 1464 20349 1476 20383
rect 1510 20380 1522 20383
rect 1670 20380 1676 20392
rect 1510 20352 1676 20380
rect 1510 20349 1522 20352
rect 1464 20343 1522 20349
rect 1670 20340 1676 20352
rect 1728 20340 1734 20392
rect 2409 20383 2467 20389
rect 2409 20349 2421 20383
rect 2455 20380 2467 20383
rect 2590 20380 2596 20392
rect 2455 20352 2596 20380
rect 2455 20349 2467 20352
rect 2409 20343 2467 20349
rect 2590 20340 2596 20352
rect 2648 20340 2654 20392
rect 4338 20340 4344 20392
rect 4396 20380 4402 20392
rect 4433 20383 4491 20389
rect 4433 20380 4445 20383
rect 4396 20352 4445 20380
rect 4396 20340 4402 20352
rect 4433 20349 4445 20352
rect 4479 20349 4491 20383
rect 4890 20380 4896 20392
rect 4803 20352 4896 20380
rect 4433 20343 4491 20349
rect 4890 20340 4896 20352
rect 4948 20340 4954 20392
rect 5442 20380 5448 20392
rect 5403 20352 5448 20380
rect 5442 20340 5448 20352
rect 5500 20340 5506 20392
rect 5629 20383 5687 20389
rect 5629 20349 5641 20383
rect 5675 20349 5687 20383
rect 5629 20343 5687 20349
rect 2317 20315 2375 20321
rect 2317 20281 2329 20315
rect 2363 20312 2375 20315
rect 2771 20315 2829 20321
rect 2771 20312 2783 20315
rect 2363 20284 2783 20312
rect 2363 20281 2375 20284
rect 2317 20275 2375 20281
rect 2771 20281 2783 20284
rect 2817 20312 2829 20315
rect 2866 20312 2872 20324
rect 2817 20284 2872 20312
rect 2817 20281 2829 20284
rect 2771 20275 2829 20281
rect 2866 20272 2872 20284
rect 2924 20312 2930 20324
rect 3510 20312 3516 20324
rect 2924 20284 3516 20312
rect 2924 20272 2930 20284
rect 3510 20272 3516 20284
rect 3568 20272 3574 20324
rect 4522 20244 4528 20256
rect 4483 20216 4528 20244
rect 4522 20204 4528 20216
rect 4580 20204 4586 20256
rect 5258 20204 5264 20256
rect 5316 20244 5322 20256
rect 5644 20244 5672 20343
rect 7006 20340 7012 20392
rect 7064 20380 7070 20392
rect 7377 20383 7435 20389
rect 7377 20380 7389 20383
rect 7064 20352 7389 20380
rect 7064 20340 7070 20352
rect 7377 20349 7389 20352
rect 7423 20349 7435 20383
rect 7377 20343 7435 20349
rect 7466 20340 7472 20392
rect 7524 20380 7530 20392
rect 7837 20383 7895 20389
rect 7837 20380 7849 20383
rect 7524 20352 7849 20380
rect 7524 20340 7530 20352
rect 7837 20349 7849 20352
rect 7883 20349 7895 20383
rect 8202 20380 8208 20392
rect 8163 20352 8208 20380
rect 7837 20343 7895 20349
rect 8202 20340 8208 20352
rect 8260 20340 8266 20392
rect 8772 20389 8800 20420
rect 9030 20408 9036 20460
rect 9088 20448 9094 20460
rect 9088 20420 9720 20448
rect 9088 20408 9094 20420
rect 9692 20389 9720 20420
rect 8757 20383 8815 20389
rect 8757 20349 8769 20383
rect 8803 20380 8815 20383
rect 9677 20383 9735 20389
rect 8803 20352 9628 20380
rect 8803 20349 8815 20352
rect 8757 20343 8815 20349
rect 6273 20315 6331 20321
rect 6273 20281 6285 20315
rect 6319 20312 6331 20315
rect 7650 20312 7656 20324
rect 6319 20284 7656 20312
rect 6319 20281 6331 20284
rect 6273 20275 6331 20281
rect 7650 20272 7656 20284
rect 7708 20312 7714 20324
rect 8220 20312 8248 20340
rect 7708 20284 8248 20312
rect 7708 20272 7714 20284
rect 5316 20216 5672 20244
rect 6641 20247 6699 20253
rect 5316 20204 5322 20216
rect 6641 20213 6653 20247
rect 6687 20244 6699 20247
rect 6730 20244 6736 20256
rect 6687 20216 6736 20244
rect 6687 20213 6699 20216
rect 6641 20207 6699 20213
rect 6730 20204 6736 20216
rect 6788 20204 6794 20256
rect 7282 20204 7288 20256
rect 7340 20244 7346 20256
rect 9600 20253 9628 20352
rect 9677 20349 9689 20383
rect 9723 20349 9735 20383
rect 10410 20380 10416 20392
rect 10371 20352 10416 20380
rect 9677 20343 9735 20349
rect 10410 20340 10416 20352
rect 10468 20340 10474 20392
rect 10520 20389 10548 20476
rect 11146 20448 11152 20460
rect 11107 20420 11152 20448
rect 11146 20408 11152 20420
rect 11204 20408 11210 20460
rect 14093 20451 14151 20457
rect 14093 20417 14105 20451
rect 14139 20448 14151 20451
rect 15654 20448 15660 20460
rect 14139 20420 15660 20448
rect 14139 20417 14151 20420
rect 14093 20411 14151 20417
rect 15654 20408 15660 20420
rect 15712 20408 15718 20460
rect 21358 20448 21364 20460
rect 17144 20420 21364 20448
rect 10505 20383 10563 20389
rect 10505 20349 10517 20383
rect 10551 20380 10563 20383
rect 10962 20380 10968 20392
rect 10551 20352 10968 20380
rect 10551 20349 10563 20352
rect 10505 20343 10563 20349
rect 10962 20340 10968 20352
rect 11020 20340 11026 20392
rect 11057 20383 11115 20389
rect 11057 20349 11069 20383
rect 11103 20380 11115 20383
rect 11330 20380 11336 20392
rect 11103 20352 11336 20380
rect 11103 20349 11115 20352
rect 11057 20343 11115 20349
rect 11330 20340 11336 20352
rect 11388 20340 11394 20392
rect 14921 20383 14979 20389
rect 14921 20349 14933 20383
rect 14967 20380 14979 20383
rect 15378 20380 15384 20392
rect 14967 20352 15384 20380
rect 14967 20349 14979 20352
rect 14921 20343 14979 20349
rect 15378 20340 15384 20352
rect 15436 20340 15442 20392
rect 15930 20340 15936 20392
rect 15988 20380 15994 20392
rect 17144 20389 17172 20420
rect 21358 20408 21364 20420
rect 21416 20408 21422 20460
rect 16704 20383 16762 20389
rect 16704 20380 16716 20383
rect 15988 20352 16716 20380
rect 15988 20340 15994 20352
rect 16704 20349 16716 20352
rect 16750 20380 16762 20383
rect 17129 20383 17187 20389
rect 17129 20380 17141 20383
rect 16750 20352 17141 20380
rect 16750 20349 16762 20352
rect 16704 20343 16762 20349
rect 17129 20349 17141 20352
rect 17175 20349 17187 20383
rect 17129 20343 17187 20349
rect 18049 20383 18107 20389
rect 18049 20349 18061 20383
rect 18095 20380 18107 20383
rect 18506 20380 18512 20392
rect 18095 20352 18512 20380
rect 18095 20349 18107 20352
rect 18049 20343 18107 20349
rect 18506 20340 18512 20352
rect 18564 20340 18570 20392
rect 19096 20383 19154 20389
rect 19096 20380 19108 20383
rect 19076 20349 19108 20380
rect 19142 20380 19154 20383
rect 19521 20383 19579 20389
rect 19521 20380 19533 20383
rect 19142 20352 19533 20380
rect 19142 20349 19154 20352
rect 19076 20343 19154 20349
rect 19521 20349 19533 20352
rect 19567 20380 19579 20383
rect 23934 20380 23940 20392
rect 19567 20352 23940 20380
rect 19567 20349 19579 20352
rect 19521 20343 19579 20349
rect 10980 20312 11008 20340
rect 11425 20315 11483 20321
rect 11425 20312 11437 20315
rect 10980 20284 11437 20312
rect 11425 20281 11437 20284
rect 11471 20281 11483 20315
rect 13446 20312 13452 20324
rect 13407 20284 13452 20312
rect 11425 20275 11483 20281
rect 13446 20272 13452 20284
rect 13504 20272 13510 20324
rect 13541 20315 13599 20321
rect 13541 20281 13553 20315
rect 13587 20312 13599 20315
rect 14826 20312 14832 20324
rect 13587 20284 14832 20312
rect 13587 20281 13599 20284
rect 13541 20275 13599 20281
rect 7469 20247 7527 20253
rect 7469 20244 7481 20247
rect 7340 20216 7481 20244
rect 7340 20204 7346 20216
rect 7469 20213 7481 20216
rect 7515 20213 7527 20247
rect 7469 20207 7527 20213
rect 9585 20247 9643 20253
rect 9585 20213 9597 20247
rect 9631 20244 9643 20247
rect 9858 20244 9864 20256
rect 9631 20216 9864 20244
rect 9631 20213 9643 20216
rect 9585 20207 9643 20213
rect 9858 20204 9864 20216
rect 9916 20204 9922 20256
rect 12066 20244 12072 20256
rect 12027 20216 12072 20244
rect 12066 20204 12072 20216
rect 12124 20204 12130 20256
rect 13265 20247 13323 20253
rect 13265 20213 13277 20247
rect 13311 20244 13323 20247
rect 13556 20244 13584 20275
rect 14826 20272 14832 20284
rect 14884 20272 14890 20324
rect 19076 20312 19104 20343
rect 23934 20340 23940 20352
rect 23992 20340 23998 20392
rect 17512 20284 19104 20312
rect 17512 20256 17540 20284
rect 14366 20244 14372 20256
rect 13311 20216 13584 20244
rect 14327 20216 14372 20244
rect 13311 20213 13323 20216
rect 13265 20207 13323 20213
rect 14366 20204 14372 20216
rect 14424 20204 14430 20256
rect 15280 20244 15286 20256
rect 15241 20216 15286 20244
rect 15280 20204 15286 20216
rect 15338 20204 15344 20256
rect 16574 20204 16580 20256
rect 16632 20244 16638 20256
rect 16807 20247 16865 20253
rect 16807 20244 16819 20247
rect 16632 20216 16819 20244
rect 16632 20204 16638 20216
rect 16807 20213 16819 20216
rect 16853 20213 16865 20247
rect 17494 20244 17500 20256
rect 17455 20216 17500 20244
rect 16807 20207 16865 20213
rect 17494 20204 17500 20216
rect 17552 20204 17558 20256
rect 18506 20244 18512 20256
rect 18467 20216 18512 20244
rect 18506 20204 18512 20216
rect 18564 20204 18570 20256
rect 18598 20204 18604 20256
rect 18656 20244 18662 20256
rect 19199 20247 19257 20253
rect 19199 20244 19211 20247
rect 18656 20216 19211 20244
rect 18656 20204 18662 20216
rect 19199 20213 19211 20216
rect 19245 20213 19257 20247
rect 19199 20207 19257 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 3418 20000 3424 20052
rect 3476 20040 3482 20052
rect 6270 20040 6276 20052
rect 3476 20012 5764 20040
rect 6231 20012 6276 20040
rect 3476 20000 3482 20012
rect 1578 19972 1584 19984
rect 1539 19944 1584 19972
rect 1578 19932 1584 19944
rect 1636 19932 1642 19984
rect 3326 19932 3332 19984
rect 3384 19972 3390 19984
rect 4065 19975 4123 19981
rect 4065 19972 4077 19975
rect 3384 19944 4077 19972
rect 3384 19932 3390 19944
rect 4065 19941 4077 19944
rect 4111 19941 4123 19975
rect 4065 19935 4123 19941
rect 2222 19904 2228 19916
rect 2183 19876 2228 19904
rect 2222 19864 2228 19876
rect 2280 19864 2286 19916
rect 3881 19907 3939 19913
rect 3881 19873 3893 19907
rect 3927 19904 3939 19907
rect 4154 19904 4160 19916
rect 3927 19876 4160 19904
rect 3927 19873 3939 19876
rect 3881 19867 3939 19873
rect 4154 19864 4160 19876
rect 4212 19904 4218 19916
rect 5736 19913 5764 20012
rect 6270 20000 6276 20012
rect 6328 20000 6334 20052
rect 7006 20000 7012 20052
rect 7064 20040 7070 20052
rect 8297 20043 8355 20049
rect 8297 20040 8309 20043
rect 7064 20012 8309 20040
rect 7064 20000 7070 20012
rect 8297 20009 8309 20012
rect 8343 20040 8355 20043
rect 9030 20040 9036 20052
rect 8343 20012 9036 20040
rect 8343 20009 8355 20012
rect 8297 20003 8355 20009
rect 9030 20000 9036 20012
rect 9088 20000 9094 20052
rect 11790 20040 11796 20052
rect 11751 20012 11796 20040
rect 11790 20000 11796 20012
rect 11848 20040 11854 20052
rect 12434 20040 12440 20052
rect 11848 20012 12440 20040
rect 11848 20000 11854 20012
rect 12434 20000 12440 20012
rect 12492 20040 12498 20052
rect 12529 20043 12587 20049
rect 12529 20040 12541 20043
rect 12492 20012 12541 20040
rect 12492 20000 12498 20012
rect 12529 20009 12541 20012
rect 12575 20009 12587 20043
rect 12529 20003 12587 20009
rect 13446 20000 13452 20052
rect 13504 20040 13510 20052
rect 14185 20043 14243 20049
rect 14185 20040 14197 20043
rect 13504 20012 14197 20040
rect 13504 20000 13510 20012
rect 14185 20009 14197 20012
rect 14231 20040 14243 20043
rect 16574 20040 16580 20052
rect 14231 20012 16580 20040
rect 14231 20009 14243 20012
rect 14185 20003 14243 20009
rect 16574 20000 16580 20012
rect 16632 20000 16638 20052
rect 6730 19932 6736 19984
rect 6788 19972 6794 19984
rect 9122 19972 9128 19984
rect 6788 19944 9128 19972
rect 6788 19932 6794 19944
rect 5721 19907 5779 19913
rect 4212 19876 4257 19904
rect 4212 19864 4218 19876
rect 5721 19873 5733 19907
rect 5767 19904 5779 19907
rect 6454 19904 6460 19916
rect 5767 19876 6460 19904
rect 5767 19873 5779 19876
rect 5721 19867 5779 19873
rect 6454 19864 6460 19876
rect 6512 19864 6518 19916
rect 6822 19904 6828 19916
rect 6783 19876 6828 19904
rect 6822 19864 6828 19876
rect 6880 19864 6886 19916
rect 7576 19913 7604 19944
rect 9122 19932 9128 19944
rect 9180 19932 9186 19984
rect 9490 19932 9496 19984
rect 9548 19972 9554 19984
rect 9548 19944 11652 19972
rect 9548 19932 9554 19944
rect 7101 19907 7159 19913
rect 7101 19873 7113 19907
rect 7147 19873 7159 19907
rect 7101 19867 7159 19873
rect 7561 19907 7619 19913
rect 7561 19873 7573 19907
rect 7607 19873 7619 19907
rect 8570 19904 8576 19916
rect 8531 19876 8576 19904
rect 7561 19867 7619 19873
rect 7116 19836 7144 19867
rect 8570 19864 8576 19876
rect 8628 19864 8634 19916
rect 9858 19864 9864 19916
rect 9916 19904 9922 19916
rect 9953 19907 10011 19913
rect 9953 19904 9965 19907
rect 9916 19876 9965 19904
rect 9916 19864 9922 19876
rect 9953 19873 9965 19876
rect 9999 19873 10011 19907
rect 9953 19867 10011 19873
rect 10134 19864 10140 19916
rect 10192 19904 10198 19916
rect 11624 19913 11652 19944
rect 12066 19932 12072 19984
rect 12124 19972 12130 19984
rect 16390 19972 16396 19984
rect 12124 19944 13400 19972
rect 16351 19944 16396 19972
rect 12124 19932 12130 19944
rect 10229 19907 10287 19913
rect 10229 19904 10241 19907
rect 10192 19876 10241 19904
rect 10192 19864 10198 19876
rect 10229 19873 10241 19876
rect 10275 19873 10287 19907
rect 10229 19867 10287 19873
rect 11609 19907 11667 19913
rect 11609 19873 11621 19907
rect 11655 19904 11667 19907
rect 11790 19904 11796 19916
rect 11655 19876 11796 19904
rect 11655 19873 11667 19876
rect 11609 19867 11667 19873
rect 11790 19864 11796 19876
rect 11848 19904 11854 19916
rect 13081 19907 13139 19913
rect 13081 19904 13093 19907
rect 11848 19876 13093 19904
rect 11848 19864 11854 19876
rect 13081 19873 13093 19876
rect 13127 19904 13139 19907
rect 13262 19904 13268 19916
rect 13127 19876 13268 19904
rect 13127 19873 13139 19876
rect 13081 19867 13139 19873
rect 13262 19864 13268 19876
rect 13320 19864 13326 19916
rect 13372 19913 13400 19944
rect 16390 19932 16396 19944
rect 16448 19932 16454 19984
rect 13357 19907 13415 19913
rect 13357 19873 13369 19907
rect 13403 19904 13415 19907
rect 13998 19904 14004 19916
rect 13403 19876 14004 19904
rect 13403 19873 13415 19876
rect 13357 19867 13415 19873
rect 13998 19864 14004 19876
rect 14056 19904 14062 19916
rect 16114 19904 16120 19916
rect 14056 19876 16120 19904
rect 14056 19864 14062 19876
rect 16114 19864 16120 19876
rect 16172 19864 16178 19916
rect 17770 19904 17776 19916
rect 17731 19876 17776 19904
rect 17770 19864 17776 19876
rect 17828 19864 17834 19916
rect 18782 19904 18788 19916
rect 18743 19876 18788 19904
rect 18782 19864 18788 19876
rect 18840 19864 18846 19916
rect 7282 19836 7288 19848
rect 6012 19808 7288 19836
rect 2682 19700 2688 19712
rect 2643 19672 2688 19700
rect 2682 19660 2688 19672
rect 2740 19660 2746 19712
rect 2958 19700 2964 19712
rect 2919 19672 2964 19700
rect 2958 19660 2964 19672
rect 3016 19660 3022 19712
rect 3421 19703 3479 19709
rect 3421 19669 3433 19703
rect 3467 19700 3479 19703
rect 3602 19700 3608 19712
rect 3467 19672 3608 19700
rect 3467 19669 3479 19672
rect 3421 19663 3479 19669
rect 3602 19660 3608 19672
rect 3660 19660 3666 19712
rect 5169 19703 5227 19709
rect 5169 19669 5181 19703
rect 5215 19700 5227 19703
rect 5258 19700 5264 19712
rect 5215 19672 5264 19700
rect 5215 19669 5227 19672
rect 5169 19663 5227 19669
rect 5258 19660 5264 19672
rect 5316 19660 5322 19712
rect 5534 19660 5540 19712
rect 5592 19700 5598 19712
rect 6012 19709 6040 19808
rect 7282 19796 7288 19808
rect 7340 19796 7346 19848
rect 9125 19839 9183 19845
rect 9125 19805 9137 19839
rect 9171 19836 9183 19839
rect 9214 19836 9220 19848
rect 9171 19808 9220 19836
rect 9171 19805 9183 19808
rect 9125 19799 9183 19805
rect 9214 19796 9220 19808
rect 9272 19796 9278 19848
rect 10686 19836 10692 19848
rect 10647 19808 10692 19836
rect 10686 19796 10692 19808
rect 10744 19796 10750 19848
rect 13722 19836 13728 19848
rect 13683 19808 13728 19836
rect 13722 19796 13728 19808
rect 13780 19796 13786 19848
rect 15654 19796 15660 19848
rect 15712 19836 15718 19848
rect 16022 19836 16028 19848
rect 15712 19808 16028 19836
rect 15712 19796 15718 19808
rect 16022 19796 16028 19808
rect 16080 19836 16086 19848
rect 16301 19839 16359 19845
rect 16301 19836 16313 19839
rect 16080 19808 16313 19836
rect 16080 19796 16086 19808
rect 16301 19805 16313 19808
rect 16347 19805 16359 19839
rect 18506 19836 18512 19848
rect 16301 19799 16359 19805
rect 16408 19808 18512 19836
rect 9950 19728 9956 19780
rect 10008 19768 10014 19780
rect 10045 19771 10103 19777
rect 10045 19768 10057 19771
rect 10008 19740 10057 19768
rect 10008 19728 10014 19740
rect 10045 19737 10057 19740
rect 10091 19737 10103 19771
rect 10045 19731 10103 19737
rect 12526 19728 12532 19780
rect 12584 19768 12590 19780
rect 13173 19771 13231 19777
rect 13173 19768 13185 19771
rect 12584 19740 13185 19768
rect 12584 19728 12590 19740
rect 13173 19737 13185 19740
rect 13219 19737 13231 19771
rect 16408 19768 16436 19808
rect 18506 19796 18512 19808
rect 18564 19796 18570 19848
rect 16850 19768 16856 19780
rect 13173 19731 13231 19737
rect 13786 19740 16436 19768
rect 16811 19740 16856 19768
rect 5997 19703 6055 19709
rect 5997 19700 6009 19703
rect 5592 19672 6009 19700
rect 5592 19660 5598 19672
rect 5997 19669 6009 19672
rect 6043 19669 6055 19703
rect 5997 19663 6055 19669
rect 7650 19660 7656 19712
rect 7708 19700 7714 19712
rect 7929 19703 7987 19709
rect 7929 19700 7941 19703
rect 7708 19672 7941 19700
rect 7708 19660 7714 19672
rect 7929 19669 7941 19672
rect 7975 19700 7987 19703
rect 8202 19700 8208 19712
rect 7975 19672 8208 19700
rect 7975 19669 7987 19672
rect 7929 19663 7987 19669
rect 8202 19660 8208 19672
rect 8260 19660 8266 19712
rect 8662 19660 8668 19712
rect 8720 19700 8726 19712
rect 8757 19703 8815 19709
rect 8757 19700 8769 19703
rect 8720 19672 8769 19700
rect 8720 19660 8726 19672
rect 8757 19669 8769 19672
rect 8803 19669 8815 19703
rect 8757 19663 8815 19669
rect 9122 19660 9128 19712
rect 9180 19700 9186 19712
rect 9493 19703 9551 19709
rect 9493 19700 9505 19703
rect 9180 19672 9505 19700
rect 9180 19660 9186 19672
rect 9493 19669 9505 19672
rect 9539 19700 9551 19703
rect 9766 19700 9772 19712
rect 9539 19672 9772 19700
rect 9539 19669 9551 19672
rect 9493 19663 9551 19669
rect 9766 19660 9772 19672
rect 9824 19660 9830 19712
rect 10962 19700 10968 19712
rect 10923 19672 10968 19700
rect 10962 19660 10968 19672
rect 11020 19660 11026 19712
rect 11422 19700 11428 19712
rect 11335 19672 11428 19700
rect 11422 19660 11428 19672
rect 11480 19700 11486 19712
rect 13786 19700 13814 19740
rect 16850 19728 16856 19740
rect 16908 19728 16914 19780
rect 11480 19672 13814 19700
rect 15013 19703 15071 19709
rect 11480 19660 11486 19672
rect 15013 19669 15025 19703
rect 15059 19700 15071 19703
rect 15378 19700 15384 19712
rect 15059 19672 15384 19700
rect 15059 19669 15071 19672
rect 15013 19663 15071 19669
rect 15378 19660 15384 19672
rect 15436 19660 15442 19712
rect 15562 19700 15568 19712
rect 15523 19672 15568 19700
rect 15562 19660 15568 19672
rect 15620 19660 15626 19712
rect 15838 19660 15844 19712
rect 15896 19700 15902 19712
rect 17957 19703 18015 19709
rect 17957 19700 17969 19703
rect 15896 19672 17969 19700
rect 15896 19660 15902 19672
rect 17957 19669 17969 19672
rect 18003 19669 18015 19703
rect 18966 19700 18972 19712
rect 18927 19672 18972 19700
rect 17957 19663 18015 19669
rect 18966 19660 18972 19672
rect 19024 19660 19030 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 2222 19456 2228 19508
rect 2280 19496 2286 19508
rect 2409 19499 2467 19505
rect 2409 19496 2421 19499
rect 2280 19468 2421 19496
rect 2280 19456 2286 19468
rect 2409 19465 2421 19468
rect 2455 19465 2467 19499
rect 2866 19496 2872 19508
rect 2827 19468 2872 19496
rect 2409 19459 2467 19465
rect 2866 19456 2872 19468
rect 2924 19456 2930 19508
rect 3973 19499 4031 19505
rect 3973 19465 3985 19499
rect 4019 19496 4031 19499
rect 4154 19496 4160 19508
rect 4019 19468 4160 19496
rect 4019 19465 4031 19468
rect 3973 19459 4031 19465
rect 4154 19456 4160 19468
rect 4212 19496 4218 19508
rect 4249 19499 4307 19505
rect 4249 19496 4261 19499
rect 4212 19468 4261 19496
rect 4212 19456 4218 19468
rect 4249 19465 4261 19468
rect 4295 19465 4307 19499
rect 4249 19459 4307 19465
rect 5905 19499 5963 19505
rect 5905 19465 5917 19499
rect 5951 19496 5963 19499
rect 6822 19496 6828 19508
rect 5951 19468 6828 19496
rect 5951 19465 5963 19468
rect 5905 19459 5963 19465
rect 6822 19456 6828 19468
rect 6880 19496 6886 19508
rect 7466 19496 7472 19508
rect 6880 19468 7472 19496
rect 6880 19456 6886 19468
rect 7466 19456 7472 19468
rect 7524 19456 7530 19508
rect 9858 19456 9864 19508
rect 9916 19496 9922 19508
rect 10689 19499 10747 19505
rect 10689 19496 10701 19499
rect 9916 19468 10701 19496
rect 9916 19456 9922 19468
rect 10689 19465 10701 19468
rect 10735 19496 10747 19499
rect 10778 19496 10784 19508
rect 10735 19468 10784 19496
rect 10735 19465 10747 19468
rect 10689 19459 10747 19465
rect 10778 19456 10784 19468
rect 10836 19456 10842 19508
rect 11790 19496 11796 19508
rect 11751 19468 11796 19496
rect 11790 19456 11796 19468
rect 11848 19456 11854 19508
rect 13262 19456 13268 19508
rect 13320 19496 13326 19508
rect 13449 19499 13507 19505
rect 13449 19496 13461 19499
rect 13320 19468 13461 19496
rect 13320 19456 13326 19468
rect 13449 19465 13461 19468
rect 13495 19496 13507 19499
rect 15470 19496 15476 19508
rect 13495 19468 15476 19496
rect 13495 19465 13507 19468
rect 13449 19459 13507 19465
rect 15470 19456 15476 19468
rect 15528 19456 15534 19508
rect 16390 19496 16396 19508
rect 16351 19468 16396 19496
rect 16390 19456 16396 19468
rect 16448 19496 16454 19508
rect 16669 19499 16727 19505
rect 16669 19496 16681 19499
rect 16448 19468 16681 19496
rect 16448 19456 16454 19468
rect 16669 19465 16681 19468
rect 16715 19465 16727 19499
rect 16669 19459 16727 19465
rect 17497 19499 17555 19505
rect 17497 19465 17509 19499
rect 17543 19496 17555 19499
rect 17770 19496 17776 19508
rect 17543 19468 17776 19496
rect 17543 19465 17555 19468
rect 17497 19459 17555 19465
rect 6641 19431 6699 19437
rect 6641 19397 6653 19431
rect 6687 19428 6699 19431
rect 9876 19428 9904 19456
rect 10870 19428 10876 19440
rect 6687 19400 7788 19428
rect 6687 19397 6699 19400
rect 6641 19391 6699 19397
rect 3053 19363 3111 19369
rect 3053 19329 3065 19363
rect 3099 19360 3111 19363
rect 3142 19360 3148 19372
rect 3099 19332 3148 19360
rect 3099 19329 3111 19332
rect 3053 19323 3111 19329
rect 3142 19320 3148 19332
rect 3200 19360 3206 19372
rect 4522 19360 4528 19372
rect 3200 19332 4528 19360
rect 3200 19320 3206 19332
rect 4522 19320 4528 19332
rect 4580 19320 4586 19372
rect 6454 19320 6460 19372
rect 6512 19360 6518 19372
rect 7558 19360 7564 19372
rect 6512 19332 7564 19360
rect 6512 19320 6518 19332
rect 2041 19295 2099 19301
rect 2041 19261 2053 19295
rect 2087 19292 2099 19295
rect 2222 19292 2228 19304
rect 2087 19264 2228 19292
rect 2087 19261 2099 19264
rect 2041 19255 2099 19261
rect 2222 19252 2228 19264
rect 2280 19292 2286 19304
rect 2958 19292 2964 19304
rect 2280 19264 2964 19292
rect 2280 19252 2286 19264
rect 2958 19252 2964 19264
rect 3016 19252 3022 19304
rect 4801 19295 4859 19301
rect 4801 19292 4813 19295
rect 4632 19264 4813 19292
rect 2866 19184 2872 19236
rect 2924 19224 2930 19236
rect 3374 19227 3432 19233
rect 3374 19224 3386 19227
rect 2924 19196 3386 19224
rect 2924 19184 2930 19196
rect 3374 19193 3386 19196
rect 3420 19193 3432 19227
rect 3374 19187 3432 19193
rect 4632 19168 4660 19264
rect 4801 19261 4813 19264
rect 4847 19261 4859 19295
rect 4801 19255 4859 19261
rect 6273 19295 6331 19301
rect 6273 19261 6285 19295
rect 6319 19292 6331 19295
rect 6730 19292 6736 19304
rect 6319 19264 6736 19292
rect 6319 19261 6331 19264
rect 6273 19255 6331 19261
rect 6730 19252 6736 19264
rect 6788 19252 6794 19304
rect 7116 19301 7144 19332
rect 7558 19320 7564 19332
rect 7616 19320 7622 19372
rect 7760 19304 7788 19400
rect 9232 19400 9904 19428
rect 10783 19400 10876 19428
rect 7101 19295 7159 19301
rect 7101 19261 7113 19295
rect 7147 19261 7159 19295
rect 7374 19292 7380 19304
rect 7335 19264 7380 19292
rect 7101 19255 7159 19261
rect 7374 19252 7380 19264
rect 7432 19252 7438 19304
rect 7653 19295 7711 19301
rect 7653 19292 7665 19295
rect 7576 19264 7665 19292
rect 7282 19184 7288 19236
rect 7340 19224 7346 19236
rect 7576 19224 7604 19264
rect 7653 19261 7665 19264
rect 7699 19261 7711 19295
rect 7653 19255 7711 19261
rect 7742 19252 7748 19304
rect 7800 19292 7806 19304
rect 8205 19295 8263 19301
rect 8205 19292 8217 19295
rect 7800 19264 8217 19292
rect 7800 19252 7806 19264
rect 8205 19261 8217 19264
rect 8251 19292 8263 19295
rect 9232 19292 9260 19400
rect 10870 19388 10876 19400
rect 10928 19428 10934 19440
rect 11422 19428 11428 19440
rect 10928 19400 11428 19428
rect 10928 19388 10934 19400
rect 11422 19388 11428 19400
rect 11480 19388 11486 19440
rect 16022 19388 16028 19440
rect 16080 19428 16086 19440
rect 17037 19431 17095 19437
rect 17037 19428 17049 19431
rect 16080 19400 17049 19428
rect 16080 19388 16086 19400
rect 17037 19397 17049 19400
rect 17083 19397 17095 19431
rect 17037 19391 17095 19397
rect 9950 19360 9956 19372
rect 9911 19332 9956 19360
rect 9950 19320 9956 19332
rect 10008 19320 10014 19372
rect 12176 19332 12756 19360
rect 8251 19264 9260 19292
rect 9309 19295 9367 19301
rect 8251 19261 8263 19264
rect 8205 19255 8263 19261
rect 9309 19261 9321 19295
rect 9355 19261 9367 19295
rect 9309 19255 9367 19261
rect 10781 19295 10839 19301
rect 10781 19261 10793 19295
rect 10827 19292 10839 19295
rect 10962 19292 10968 19304
rect 10827 19264 10968 19292
rect 10827 19261 10839 19264
rect 10781 19255 10839 19261
rect 9033 19227 9091 19233
rect 9033 19224 9045 19227
rect 7340 19196 7604 19224
rect 7760 19196 9045 19224
rect 7340 19184 7346 19196
rect 1670 19156 1676 19168
rect 1631 19128 1676 19156
rect 1670 19116 1676 19128
rect 1728 19116 1734 19168
rect 4614 19156 4620 19168
rect 4575 19128 4620 19156
rect 4614 19116 4620 19128
rect 4672 19116 4678 19168
rect 4982 19156 4988 19168
rect 4943 19128 4988 19156
rect 4982 19116 4988 19128
rect 5040 19116 5046 19168
rect 5534 19156 5540 19168
rect 5495 19128 5540 19156
rect 5534 19116 5540 19128
rect 5592 19116 5598 19168
rect 6638 19116 6644 19168
rect 6696 19156 6702 19168
rect 6917 19159 6975 19165
rect 6917 19156 6929 19159
rect 6696 19128 6929 19156
rect 6696 19116 6702 19128
rect 6917 19125 6929 19128
rect 6963 19125 6975 19159
rect 6917 19119 6975 19125
rect 7190 19116 7196 19168
rect 7248 19156 7254 19168
rect 7760 19156 7788 19196
rect 9033 19193 9045 19196
rect 9079 19224 9091 19227
rect 9324 19224 9352 19255
rect 10962 19252 10968 19264
rect 11020 19252 11026 19304
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 12066 19292 12072 19304
rect 11112 19264 11157 19292
rect 11440 19264 12072 19292
rect 11112 19252 11118 19264
rect 9858 19224 9864 19236
rect 9079 19196 9864 19224
rect 9079 19193 9091 19196
rect 9033 19187 9091 19193
rect 9858 19184 9864 19196
rect 9916 19184 9922 19236
rect 11440 19224 11468 19264
rect 12066 19252 12072 19264
rect 12124 19292 12130 19304
rect 12176 19301 12204 19332
rect 12161 19295 12219 19301
rect 12161 19292 12173 19295
rect 12124 19264 12173 19292
rect 12124 19252 12130 19264
rect 12161 19261 12173 19264
rect 12207 19261 12219 19295
rect 12434 19292 12440 19304
rect 12395 19264 12440 19292
rect 12161 19255 12219 19261
rect 12434 19252 12440 19264
rect 12492 19252 12498 19304
rect 12526 19252 12532 19304
rect 12584 19292 12590 19304
rect 12728 19301 12756 19332
rect 13722 19320 13728 19372
rect 13780 19360 13786 19372
rect 17512 19360 17540 19459
rect 17770 19456 17776 19468
rect 17828 19456 17834 19508
rect 13780 19332 17540 19360
rect 13780 19320 13786 19332
rect 17770 19320 17776 19372
rect 17828 19360 17834 19372
rect 17828 19332 18092 19360
rect 17828 19320 17834 19332
rect 12713 19295 12771 19301
rect 12584 19264 12629 19292
rect 12584 19252 12590 19264
rect 12713 19261 12725 19295
rect 12759 19261 12771 19295
rect 12713 19255 12771 19261
rect 13173 19295 13231 19301
rect 13173 19261 13185 19295
rect 13219 19292 13231 19295
rect 14001 19295 14059 19301
rect 14001 19292 14013 19295
rect 13219 19264 14013 19292
rect 13219 19261 13231 19264
rect 13173 19255 13231 19261
rect 14001 19261 14013 19264
rect 14047 19292 14059 19295
rect 14829 19295 14887 19301
rect 14829 19292 14841 19295
rect 14047 19264 14841 19292
rect 14047 19261 14059 19264
rect 14001 19255 14059 19261
rect 14829 19261 14841 19264
rect 14875 19261 14887 19295
rect 14829 19255 14887 19261
rect 15473 19295 15531 19301
rect 15473 19261 15485 19295
rect 15519 19292 15531 19295
rect 15562 19292 15568 19304
rect 15519 19264 15568 19292
rect 15519 19261 15531 19264
rect 15473 19255 15531 19261
rect 15562 19252 15568 19264
rect 15620 19292 15626 19304
rect 18064 19301 18092 19332
rect 18049 19295 18107 19301
rect 15620 19264 17908 19292
rect 15620 19252 15626 19264
rect 10244 19196 11468 19224
rect 11517 19227 11575 19233
rect 7248 19128 7788 19156
rect 7248 19116 7254 19128
rect 7834 19116 7840 19168
rect 7892 19156 7898 19168
rect 8570 19156 8576 19168
rect 7892 19128 8576 19156
rect 7892 19116 7898 19128
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 10134 19116 10140 19168
rect 10192 19156 10198 19168
rect 10244 19165 10272 19196
rect 11517 19193 11529 19227
rect 11563 19224 11575 19227
rect 12250 19224 12256 19236
rect 11563 19196 12256 19224
rect 11563 19193 11575 19196
rect 11517 19187 11575 19193
rect 12250 19184 12256 19196
rect 12308 19184 12314 19236
rect 14458 19184 14464 19236
rect 14516 19224 14522 19236
rect 14553 19227 14611 19233
rect 14553 19224 14565 19227
rect 14516 19196 14565 19224
rect 14516 19184 14522 19196
rect 14553 19193 14565 19196
rect 14599 19224 14611 19227
rect 14599 19196 15516 19224
rect 14599 19193 14611 19196
rect 14553 19187 14611 19193
rect 10229 19159 10287 19165
rect 10229 19156 10241 19159
rect 10192 19128 10241 19156
rect 10192 19116 10198 19128
rect 10229 19125 10241 19128
rect 10275 19125 10287 19159
rect 10229 19119 10287 19125
rect 13817 19159 13875 19165
rect 13817 19125 13829 19159
rect 13863 19156 13875 19159
rect 13998 19156 14004 19168
rect 13863 19128 14004 19156
rect 13863 19125 13875 19128
rect 13817 19119 13875 19125
rect 13998 19116 14004 19128
rect 14056 19116 14062 19168
rect 14182 19156 14188 19168
rect 14143 19128 14188 19156
rect 14182 19116 14188 19128
rect 14240 19116 14246 19168
rect 15286 19156 15292 19168
rect 15247 19128 15292 19156
rect 15286 19116 15292 19128
rect 15344 19116 15350 19168
rect 15488 19156 15516 19196
rect 15654 19184 15660 19236
rect 15712 19224 15718 19236
rect 15794 19227 15852 19233
rect 15794 19224 15806 19227
rect 15712 19196 15806 19224
rect 15712 19184 15718 19196
rect 15794 19193 15806 19196
rect 15840 19193 15852 19227
rect 15794 19187 15852 19193
rect 16758 19156 16764 19168
rect 15488 19128 16764 19156
rect 16758 19116 16764 19128
rect 16816 19116 16822 19168
rect 17770 19156 17776 19168
rect 17731 19128 17776 19156
rect 17770 19116 17776 19128
rect 17828 19116 17834 19168
rect 17880 19156 17908 19264
rect 18049 19261 18061 19295
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 18138 19252 18144 19304
rect 18196 19292 18202 19304
rect 18509 19295 18567 19301
rect 18509 19292 18521 19295
rect 18196 19264 18521 19292
rect 18196 19252 18202 19264
rect 18509 19261 18521 19264
rect 18555 19261 18567 19295
rect 18509 19255 18567 19261
rect 18782 19252 18788 19304
rect 18840 19292 18846 19304
rect 19061 19295 19119 19301
rect 19061 19292 19073 19295
rect 18840 19264 19073 19292
rect 18840 19252 18846 19264
rect 19061 19261 19073 19264
rect 19107 19261 19119 19295
rect 19061 19255 19119 19261
rect 18141 19159 18199 19165
rect 18141 19156 18153 19159
rect 17880 19128 18153 19156
rect 18141 19125 18153 19128
rect 18187 19125 18199 19159
rect 18141 19119 18199 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1486 18912 1492 18964
rect 1544 18952 1550 18964
rect 1581 18955 1639 18961
rect 1581 18952 1593 18955
rect 1544 18924 1593 18952
rect 1544 18912 1550 18924
rect 1581 18921 1593 18924
rect 1627 18921 1639 18955
rect 3142 18952 3148 18964
rect 3103 18924 3148 18952
rect 1581 18915 1639 18921
rect 3142 18912 3148 18924
rect 3200 18912 3206 18964
rect 4203 18955 4261 18961
rect 4203 18921 4215 18955
rect 4249 18952 4261 18955
rect 4614 18952 4620 18964
rect 4249 18924 4620 18952
rect 4249 18921 4261 18924
rect 4203 18915 4261 18921
rect 4614 18912 4620 18924
rect 4672 18912 4678 18964
rect 5166 18952 5172 18964
rect 5127 18924 5172 18952
rect 5166 18912 5172 18924
rect 5224 18912 5230 18964
rect 7098 18912 7104 18964
rect 7156 18952 7162 18964
rect 7193 18955 7251 18961
rect 7193 18952 7205 18955
rect 7156 18924 7205 18952
rect 7156 18912 7162 18924
rect 7193 18921 7205 18924
rect 7239 18952 7251 18955
rect 7742 18952 7748 18964
rect 7239 18924 7748 18952
rect 7239 18921 7251 18924
rect 7193 18915 7251 18921
rect 7742 18912 7748 18924
rect 7800 18912 7806 18964
rect 10870 18952 10876 18964
rect 7944 18924 10876 18952
rect 2222 18884 2228 18896
rect 2183 18856 2228 18884
rect 2222 18844 2228 18856
rect 2280 18844 2286 18896
rect 2774 18884 2780 18896
rect 2735 18856 2780 18884
rect 2774 18844 2780 18856
rect 2832 18844 2838 18896
rect 4338 18844 4344 18896
rect 4396 18884 4402 18896
rect 4893 18887 4951 18893
rect 4893 18884 4905 18887
rect 4396 18856 4905 18884
rect 4396 18844 4402 18856
rect 4893 18853 4905 18856
rect 4939 18884 4951 18887
rect 4939 18856 5120 18884
rect 4939 18853 4951 18856
rect 4893 18847 4951 18853
rect 5092 18825 5120 18856
rect 7466 18844 7472 18896
rect 7524 18884 7530 18896
rect 7561 18887 7619 18893
rect 7561 18884 7573 18887
rect 7524 18856 7573 18884
rect 7524 18844 7530 18856
rect 7561 18853 7573 18856
rect 7607 18884 7619 18887
rect 7944 18884 7972 18924
rect 10870 18912 10876 18924
rect 10928 18912 10934 18964
rect 15378 18912 15384 18964
rect 15436 18952 15442 18964
rect 16945 18955 17003 18961
rect 16945 18952 16957 18955
rect 15436 18924 16957 18952
rect 15436 18912 15442 18924
rect 16945 18921 16957 18924
rect 16991 18921 17003 18955
rect 18138 18952 18144 18964
rect 18099 18924 18144 18952
rect 16945 18915 17003 18921
rect 18138 18912 18144 18924
rect 18196 18912 18202 18964
rect 7607 18856 7972 18884
rect 8757 18887 8815 18893
rect 7607 18853 7619 18856
rect 7561 18847 7619 18853
rect 8757 18853 8769 18887
rect 8803 18884 8815 18887
rect 10410 18884 10416 18896
rect 8803 18856 10416 18884
rect 8803 18853 8815 18856
rect 8757 18847 8815 18853
rect 10410 18844 10416 18856
rect 10468 18884 10474 18896
rect 10781 18887 10839 18893
rect 10781 18884 10793 18887
rect 10468 18856 10793 18884
rect 10468 18844 10474 18856
rect 10781 18853 10793 18856
rect 10827 18853 10839 18887
rect 10781 18847 10839 18853
rect 14642 18844 14648 18896
rect 14700 18884 14706 18896
rect 15473 18887 15531 18893
rect 15473 18884 15485 18887
rect 14700 18856 15485 18884
rect 14700 18844 14706 18856
rect 15473 18853 15485 18856
rect 15519 18853 15531 18887
rect 16022 18884 16028 18896
rect 15983 18856 16028 18884
rect 15473 18847 15531 18853
rect 16022 18844 16028 18856
rect 16080 18844 16086 18896
rect 4132 18819 4190 18825
rect 4132 18785 4144 18819
rect 4178 18816 4190 18819
rect 5077 18819 5135 18825
rect 4178 18788 4660 18816
rect 4178 18785 4190 18788
rect 4132 18779 4190 18785
rect 2133 18751 2191 18757
rect 2133 18717 2145 18751
rect 2179 18748 2191 18751
rect 3602 18748 3608 18760
rect 2179 18720 3608 18748
rect 2179 18717 2191 18720
rect 2133 18711 2191 18717
rect 3602 18708 3608 18720
rect 3660 18708 3666 18760
rect 4632 18689 4660 18788
rect 5077 18785 5089 18819
rect 5123 18785 5135 18819
rect 5077 18779 5135 18785
rect 5537 18819 5595 18825
rect 5537 18785 5549 18819
rect 5583 18785 5595 18819
rect 5994 18816 6000 18828
rect 5955 18788 6000 18816
rect 5537 18779 5595 18785
rect 4890 18708 4896 18760
rect 4948 18748 4954 18760
rect 5552 18748 5580 18779
rect 5994 18776 6000 18788
rect 6052 18776 6058 18828
rect 6362 18816 6368 18828
rect 6323 18788 6368 18816
rect 6362 18776 6368 18788
rect 6420 18776 6426 18828
rect 8202 18816 8208 18828
rect 8163 18788 8208 18816
rect 8202 18776 8208 18788
rect 8260 18776 8266 18828
rect 9766 18816 9772 18828
rect 9727 18788 9772 18816
rect 9766 18776 9772 18788
rect 9824 18776 9830 18828
rect 9861 18819 9919 18825
rect 9861 18785 9873 18819
rect 9907 18816 9919 18819
rect 9950 18816 9956 18828
rect 9907 18788 9956 18816
rect 9907 18785 9919 18788
rect 9861 18779 9919 18785
rect 9950 18776 9956 18788
rect 10008 18776 10014 18828
rect 10045 18819 10103 18825
rect 10045 18785 10057 18819
rect 10091 18816 10103 18819
rect 10134 18816 10140 18828
rect 10091 18788 10140 18816
rect 10091 18785 10103 18788
rect 10045 18779 10103 18785
rect 10134 18776 10140 18788
rect 10192 18776 10198 18828
rect 10505 18819 10563 18825
rect 10505 18785 10517 18819
rect 10551 18816 10563 18819
rect 11238 18816 11244 18828
rect 10551 18788 11244 18816
rect 10551 18785 10563 18788
rect 10505 18779 10563 18785
rect 11238 18776 11244 18788
rect 11296 18776 11302 18828
rect 11330 18776 11336 18828
rect 11388 18816 11394 18828
rect 11606 18816 11612 18828
rect 11388 18788 11433 18816
rect 11567 18788 11612 18816
rect 11388 18776 11394 18788
rect 11606 18776 11612 18788
rect 11664 18776 11670 18828
rect 13262 18816 13268 18828
rect 13223 18788 13268 18816
rect 13262 18776 13268 18788
rect 13320 18776 13326 18828
rect 13633 18819 13691 18825
rect 13633 18816 13645 18819
rect 13464 18788 13645 18816
rect 9306 18748 9312 18760
rect 4948 18720 9312 18748
rect 4948 18708 4954 18720
rect 9306 18708 9312 18720
rect 9364 18708 9370 18760
rect 9490 18748 9496 18760
rect 9403 18720 9496 18748
rect 9490 18708 9496 18720
rect 9548 18748 9554 18760
rect 11790 18748 11796 18760
rect 9548 18720 9720 18748
rect 11751 18720 11796 18748
rect 9548 18708 9554 18720
rect 4617 18683 4675 18689
rect 4617 18649 4629 18683
rect 4663 18680 4675 18683
rect 9030 18680 9036 18692
rect 4663 18652 9036 18680
rect 4663 18649 4675 18652
rect 4617 18643 4675 18649
rect 9030 18640 9036 18652
rect 9088 18640 9094 18692
rect 2958 18572 2964 18624
rect 3016 18612 3022 18624
rect 3421 18615 3479 18621
rect 3421 18612 3433 18615
rect 3016 18584 3433 18612
rect 3016 18572 3022 18584
rect 3421 18581 3433 18584
rect 3467 18581 3479 18615
rect 3878 18612 3884 18624
rect 3839 18584 3884 18612
rect 3421 18575 3479 18581
rect 3878 18572 3884 18584
rect 3936 18572 3942 18624
rect 7558 18572 7564 18624
rect 7616 18612 7622 18624
rect 7929 18615 7987 18621
rect 7929 18612 7941 18615
rect 7616 18584 7941 18612
rect 7616 18572 7622 18584
rect 7929 18581 7941 18584
rect 7975 18612 7987 18615
rect 8018 18612 8024 18624
rect 7975 18584 8024 18612
rect 7975 18581 7987 18584
rect 7929 18575 7987 18581
rect 8018 18572 8024 18584
rect 8076 18572 8082 18624
rect 9122 18612 9128 18624
rect 9083 18584 9128 18612
rect 9122 18572 9128 18584
rect 9180 18572 9186 18624
rect 9692 18612 9720 18720
rect 11790 18708 11796 18720
rect 11848 18708 11854 18760
rect 13081 18751 13139 18757
rect 13081 18717 13093 18751
rect 13127 18748 13139 18751
rect 13464 18748 13492 18788
rect 13633 18785 13645 18788
rect 13679 18816 13691 18819
rect 13722 18816 13728 18828
rect 13679 18788 13728 18816
rect 13679 18785 13691 18788
rect 13633 18779 13691 18785
rect 13722 18776 13728 18788
rect 13780 18776 13786 18828
rect 17129 18819 17187 18825
rect 17129 18785 17141 18819
rect 17175 18816 17187 18819
rect 17218 18816 17224 18828
rect 17175 18788 17224 18816
rect 17175 18785 17187 18788
rect 17129 18779 17187 18785
rect 17218 18776 17224 18788
rect 17276 18776 17282 18828
rect 17402 18816 17408 18828
rect 17315 18788 17408 18816
rect 17402 18776 17408 18788
rect 17460 18816 17466 18828
rect 18156 18816 18184 18912
rect 17460 18788 18184 18816
rect 17460 18776 17466 18788
rect 18322 18776 18328 18828
rect 18380 18816 18386 18828
rect 18417 18819 18475 18825
rect 18417 18816 18429 18819
rect 18380 18788 18429 18816
rect 18380 18776 18386 18788
rect 18417 18785 18429 18788
rect 18463 18785 18475 18819
rect 18417 18779 18475 18785
rect 13906 18748 13912 18760
rect 13127 18720 13492 18748
rect 13819 18720 13912 18748
rect 13127 18717 13139 18720
rect 13081 18711 13139 18717
rect 13906 18708 13912 18720
rect 13964 18748 13970 18760
rect 14185 18751 14243 18757
rect 14185 18748 14197 18751
rect 13964 18720 14197 18748
rect 13964 18708 13970 18720
rect 14185 18717 14197 18720
rect 14231 18717 14243 18751
rect 15378 18748 15384 18760
rect 15339 18720 15384 18748
rect 14185 18711 14243 18717
rect 15378 18708 15384 18720
rect 15436 18708 15442 18760
rect 9858 18640 9864 18692
rect 9916 18680 9922 18692
rect 11330 18680 11336 18692
rect 9916 18652 11336 18680
rect 9916 18640 9922 18652
rect 11330 18640 11336 18652
rect 11388 18680 11394 18692
rect 11425 18683 11483 18689
rect 11425 18680 11437 18683
rect 11388 18652 11437 18680
rect 11388 18640 11394 18652
rect 11425 18649 11437 18652
rect 11471 18680 11483 18683
rect 12437 18683 12495 18689
rect 12437 18680 12449 18683
rect 11471 18652 12449 18680
rect 11471 18649 11483 18652
rect 11425 18643 11483 18649
rect 12437 18649 12449 18652
rect 12483 18680 12495 18683
rect 12526 18680 12532 18692
rect 12483 18652 12532 18680
rect 12483 18649 12495 18652
rect 12437 18643 12495 18649
rect 12526 18640 12532 18652
rect 12584 18680 12590 18692
rect 14458 18680 14464 18692
rect 12584 18652 14464 18680
rect 12584 18640 12590 18652
rect 14458 18640 14464 18652
rect 14516 18640 14522 18692
rect 9950 18612 9956 18624
rect 9692 18584 9956 18612
rect 9950 18572 9956 18584
rect 10008 18572 10014 18624
rect 11054 18572 11060 18624
rect 11112 18612 11118 18624
rect 11241 18615 11299 18621
rect 11241 18612 11253 18615
rect 11112 18584 11253 18612
rect 11112 18572 11118 18584
rect 11241 18581 11253 18584
rect 11287 18612 11299 18615
rect 16298 18612 16304 18624
rect 11287 18584 16304 18612
rect 11287 18581 11299 18584
rect 11241 18575 11299 18581
rect 16298 18572 16304 18584
rect 16356 18572 16362 18624
rect 16482 18612 16488 18624
rect 16443 18584 16488 18612
rect 16482 18572 16488 18584
rect 16540 18572 16546 18624
rect 18598 18612 18604 18624
rect 18559 18584 18604 18612
rect 18598 18572 18604 18584
rect 18656 18572 18662 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 2222 18368 2228 18420
rect 2280 18408 2286 18420
rect 2409 18411 2467 18417
rect 2409 18408 2421 18411
rect 2280 18380 2421 18408
rect 2280 18368 2286 18380
rect 2409 18377 2421 18380
rect 2455 18377 2467 18411
rect 2409 18371 2467 18377
rect 2866 18368 2872 18420
rect 2924 18408 2930 18420
rect 3145 18411 3203 18417
rect 3145 18408 3157 18411
rect 2924 18380 3157 18408
rect 2924 18368 2930 18380
rect 3145 18377 3157 18380
rect 3191 18377 3203 18411
rect 3145 18371 3203 18377
rect 1486 18272 1492 18284
rect 1447 18244 1492 18272
rect 1486 18232 1492 18244
rect 1544 18232 1550 18284
rect 2133 18275 2191 18281
rect 2133 18241 2145 18275
rect 2179 18272 2191 18275
rect 2774 18272 2780 18284
rect 2179 18244 2780 18272
rect 2179 18241 2191 18244
rect 2133 18235 2191 18241
rect 2774 18232 2780 18244
rect 2832 18232 2838 18284
rect 3160 18272 3188 18371
rect 4890 18368 4896 18420
rect 4948 18408 4954 18420
rect 4985 18411 5043 18417
rect 4985 18408 4997 18411
rect 4948 18380 4997 18408
rect 4948 18368 4954 18380
rect 4985 18377 4997 18380
rect 5031 18377 5043 18411
rect 5994 18408 6000 18420
rect 4985 18371 5043 18377
rect 5092 18380 6000 18408
rect 4709 18343 4767 18349
rect 4709 18309 4721 18343
rect 4755 18340 4767 18343
rect 5092 18340 5120 18380
rect 5994 18368 6000 18380
rect 6052 18368 6058 18420
rect 8202 18408 8208 18420
rect 8163 18380 8208 18408
rect 8202 18368 8208 18380
rect 8260 18408 8266 18420
rect 8846 18408 8852 18420
rect 8260 18380 8852 18408
rect 8260 18368 8266 18380
rect 8846 18368 8852 18380
rect 8904 18368 8910 18420
rect 9861 18411 9919 18417
rect 9861 18377 9873 18411
rect 9907 18408 9919 18411
rect 10134 18408 10140 18420
rect 9907 18380 10140 18408
rect 9907 18377 9919 18380
rect 9861 18371 9919 18377
rect 10134 18368 10140 18380
rect 10192 18368 10198 18420
rect 11330 18408 11336 18420
rect 11291 18380 11336 18408
rect 11330 18368 11336 18380
rect 11388 18368 11394 18420
rect 11422 18368 11428 18420
rect 11480 18408 11486 18420
rect 11701 18411 11759 18417
rect 11701 18408 11713 18411
rect 11480 18380 11713 18408
rect 11480 18368 11486 18380
rect 11701 18377 11713 18380
rect 11747 18377 11759 18411
rect 11701 18371 11759 18377
rect 18322 18368 18328 18420
rect 18380 18408 18386 18420
rect 18417 18411 18475 18417
rect 18417 18408 18429 18411
rect 18380 18380 18429 18408
rect 18380 18368 18386 18380
rect 18417 18377 18429 18380
rect 18463 18377 18475 18411
rect 18417 18371 18475 18377
rect 6270 18340 6276 18352
rect 4755 18312 5120 18340
rect 5828 18312 6276 18340
rect 4755 18309 4767 18312
rect 4709 18303 4767 18309
rect 5000 18284 5028 18312
rect 3160 18244 3693 18272
rect 2869 18207 2927 18213
rect 2869 18173 2881 18207
rect 2915 18204 2927 18207
rect 3326 18204 3332 18216
rect 2915 18176 3332 18204
rect 2915 18173 2927 18176
rect 2869 18167 2927 18173
rect 3326 18164 3332 18176
rect 3384 18164 3390 18216
rect 1581 18139 1639 18145
rect 1581 18105 1593 18139
rect 1627 18136 1639 18139
rect 1670 18136 1676 18148
rect 1627 18108 1676 18136
rect 1627 18105 1639 18108
rect 1581 18099 1639 18105
rect 1670 18096 1676 18108
rect 1728 18096 1734 18148
rect 3665 18145 3693 18244
rect 4982 18232 4988 18284
rect 5040 18232 5046 18284
rect 5442 18164 5448 18216
rect 5500 18204 5506 18216
rect 5828 18213 5856 18312
rect 6270 18300 6276 18312
rect 6328 18300 6334 18352
rect 8478 18340 8484 18352
rect 8439 18312 8484 18340
rect 8478 18300 8484 18312
rect 8536 18340 8542 18352
rect 10318 18340 10324 18352
rect 8536 18312 10324 18340
rect 8536 18300 8542 18312
rect 10318 18300 10324 18312
rect 10376 18300 10382 18352
rect 14642 18300 14648 18352
rect 14700 18340 14706 18352
rect 14829 18343 14887 18349
rect 14829 18340 14841 18343
rect 14700 18312 14841 18340
rect 14700 18300 14706 18312
rect 14829 18309 14841 18312
rect 14875 18340 14887 18343
rect 15289 18343 15347 18349
rect 15289 18340 15301 18343
rect 14875 18312 15301 18340
rect 14875 18309 14887 18312
rect 14829 18303 14887 18309
rect 15289 18309 15301 18312
rect 15335 18340 15347 18343
rect 15562 18340 15568 18352
rect 15335 18312 15568 18340
rect 15335 18309 15347 18312
rect 15289 18303 15347 18309
rect 15562 18300 15568 18312
rect 15620 18300 15626 18352
rect 5905 18275 5963 18281
rect 5905 18241 5917 18275
rect 5951 18272 5963 18275
rect 6454 18272 6460 18284
rect 5951 18244 6460 18272
rect 5951 18241 5963 18244
rect 5905 18235 5963 18241
rect 6454 18232 6460 18244
rect 6512 18232 6518 18284
rect 6641 18275 6699 18281
rect 6641 18241 6653 18275
rect 6687 18272 6699 18275
rect 7834 18272 7840 18284
rect 6687 18244 7420 18272
rect 7795 18244 7840 18272
rect 6687 18241 6699 18244
rect 6641 18235 6699 18241
rect 5813 18207 5871 18213
rect 5813 18204 5825 18207
rect 5500 18176 5825 18204
rect 5500 18164 5506 18176
rect 5813 18173 5825 18176
rect 5859 18173 5871 18207
rect 7098 18204 7104 18216
rect 7059 18176 7104 18204
rect 5813 18167 5871 18173
rect 7098 18164 7104 18176
rect 7156 18164 7162 18216
rect 7190 18164 7196 18216
rect 7248 18204 7254 18216
rect 7392 18213 7420 18244
rect 7834 18232 7840 18244
rect 7892 18232 7898 18284
rect 8757 18275 8815 18281
rect 8757 18241 8769 18275
rect 8803 18272 8815 18275
rect 9122 18272 9128 18284
rect 8803 18244 9128 18272
rect 8803 18241 8815 18244
rect 8757 18235 8815 18241
rect 9122 18232 9128 18244
rect 9180 18272 9186 18284
rect 10042 18272 10048 18284
rect 9180 18244 10048 18272
rect 9180 18232 9186 18244
rect 10042 18232 10048 18244
rect 10100 18232 10106 18284
rect 10597 18275 10655 18281
rect 10597 18272 10609 18275
rect 10152 18244 10609 18272
rect 7377 18207 7435 18213
rect 7248 18176 7293 18204
rect 7248 18164 7254 18176
rect 7377 18173 7389 18207
rect 7423 18204 7435 18207
rect 7423 18176 8616 18204
rect 7423 18173 7435 18176
rect 7377 18167 7435 18173
rect 3650 18139 3708 18145
rect 3650 18105 3662 18139
rect 3696 18105 3708 18139
rect 3650 18099 3708 18105
rect 4249 18071 4307 18077
rect 4249 18037 4261 18071
rect 4295 18068 4307 18071
rect 4338 18068 4344 18080
rect 4295 18040 4344 18068
rect 4295 18037 4307 18040
rect 4249 18031 4307 18037
rect 4338 18028 4344 18040
rect 4396 18028 4402 18080
rect 8588 18068 8616 18176
rect 8846 18096 8852 18148
rect 8904 18136 8910 18148
rect 8904 18108 8949 18136
rect 8904 18096 8910 18108
rect 9030 18096 9036 18148
rect 9088 18136 9094 18148
rect 9401 18139 9459 18145
rect 9401 18136 9413 18139
rect 9088 18108 9413 18136
rect 9088 18096 9094 18108
rect 9401 18105 9413 18108
rect 9447 18136 9459 18139
rect 10152 18136 10180 18244
rect 10597 18241 10609 18244
rect 10643 18241 10655 18275
rect 13906 18272 13912 18284
rect 13867 18244 13912 18272
rect 10597 18235 10655 18241
rect 13906 18232 13912 18244
rect 13964 18232 13970 18284
rect 16482 18272 16488 18284
rect 16443 18244 16488 18272
rect 16482 18232 16488 18244
rect 16540 18232 16546 18284
rect 16850 18272 16856 18284
rect 16811 18244 16856 18272
rect 16850 18232 16856 18244
rect 16908 18232 16914 18284
rect 12253 18207 12311 18213
rect 12253 18173 12265 18207
rect 12299 18204 12311 18207
rect 12618 18204 12624 18216
rect 12299 18176 12624 18204
rect 12299 18173 12311 18176
rect 12253 18167 12311 18173
rect 12618 18164 12624 18176
rect 12676 18164 12682 18216
rect 16114 18204 16120 18216
rect 13280 18176 16120 18204
rect 10318 18136 10324 18148
rect 9447 18108 10180 18136
rect 10279 18108 10324 18136
rect 9447 18105 9459 18108
rect 9401 18099 9459 18105
rect 10318 18096 10324 18108
rect 10376 18096 10382 18148
rect 10410 18096 10416 18148
rect 10468 18136 10474 18148
rect 11606 18136 11612 18148
rect 10468 18108 10513 18136
rect 10888 18108 11612 18136
rect 10468 18096 10474 18108
rect 10888 18068 10916 18108
rect 11606 18096 11612 18108
rect 11664 18096 11670 18148
rect 12437 18139 12495 18145
rect 12437 18105 12449 18139
rect 12483 18105 12495 18139
rect 12437 18099 12495 18105
rect 8588 18040 10916 18068
rect 11514 18028 11520 18080
rect 11572 18068 11578 18080
rect 12452 18068 12480 18099
rect 12894 18096 12900 18148
rect 12952 18136 12958 18148
rect 12989 18139 13047 18145
rect 12989 18136 13001 18139
rect 12952 18108 13001 18136
rect 12952 18096 12958 18108
rect 12989 18105 13001 18108
rect 13035 18105 13047 18139
rect 12989 18099 13047 18105
rect 13280 18077 13308 18176
rect 16114 18164 16120 18176
rect 16172 18164 16178 18216
rect 14230 18139 14288 18145
rect 14230 18136 14242 18139
rect 14016 18108 14242 18136
rect 14016 18080 14044 18108
rect 14230 18105 14242 18108
rect 14276 18105 14288 18139
rect 14230 18099 14288 18105
rect 16577 18139 16635 18145
rect 16577 18105 16589 18139
rect 16623 18105 16635 18139
rect 16577 18099 16635 18105
rect 13265 18071 13323 18077
rect 13265 18068 13277 18071
rect 11572 18040 13277 18068
rect 11572 18028 11578 18040
rect 13265 18037 13277 18040
rect 13311 18037 13323 18071
rect 13265 18031 13323 18037
rect 13817 18071 13875 18077
rect 13817 18037 13829 18071
rect 13863 18068 13875 18071
rect 13998 18068 14004 18080
rect 13863 18040 14004 18068
rect 13863 18037 13875 18040
rect 13817 18031 13875 18037
rect 13998 18028 14004 18040
rect 14056 18028 14062 18080
rect 15378 18028 15384 18080
rect 15436 18068 15442 18080
rect 15749 18071 15807 18077
rect 15749 18068 15761 18071
rect 15436 18040 15761 18068
rect 15436 18028 15442 18040
rect 15749 18037 15761 18040
rect 15795 18068 15807 18071
rect 16206 18068 16212 18080
rect 15795 18040 16212 18068
rect 15795 18037 15807 18040
rect 15749 18031 15807 18037
rect 16206 18028 16212 18040
rect 16264 18028 16270 18080
rect 16301 18071 16359 18077
rect 16301 18037 16313 18071
rect 16347 18068 16359 18071
rect 16592 18068 16620 18099
rect 16666 18068 16672 18080
rect 16347 18040 16672 18068
rect 16347 18037 16359 18040
rect 16301 18031 16359 18037
rect 16666 18028 16672 18040
rect 16724 18028 16730 18080
rect 17310 18028 17316 18080
rect 17368 18068 17374 18080
rect 17405 18071 17463 18077
rect 17405 18068 17417 18071
rect 17368 18040 17417 18068
rect 17368 18028 17374 18040
rect 17405 18037 17417 18040
rect 17451 18037 17463 18071
rect 17405 18031 17463 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1670 17864 1676 17876
rect 1631 17836 1676 17864
rect 1670 17824 1676 17836
rect 1728 17824 1734 17876
rect 2222 17824 2228 17876
rect 2280 17864 2286 17876
rect 3145 17867 3203 17873
rect 3145 17864 3157 17867
rect 2280 17836 3157 17864
rect 2280 17824 2286 17836
rect 3145 17833 3157 17836
rect 3191 17833 3203 17867
rect 3145 17827 3203 17833
rect 3326 17824 3332 17876
rect 3384 17864 3390 17876
rect 4246 17864 4252 17876
rect 3384 17836 4154 17864
rect 4207 17836 4252 17864
rect 3384 17824 3390 17836
rect 2587 17799 2645 17805
rect 2587 17765 2599 17799
rect 2633 17796 2645 17799
rect 2866 17796 2872 17808
rect 2633 17768 2872 17796
rect 2633 17765 2645 17768
rect 2587 17759 2645 17765
rect 2866 17756 2872 17768
rect 2924 17756 2930 17808
rect 4126 17796 4154 17836
rect 4246 17824 4252 17836
rect 4304 17824 4310 17876
rect 5261 17867 5319 17873
rect 5261 17864 5273 17867
rect 4540 17836 5273 17864
rect 4540 17796 4568 17836
rect 5261 17833 5273 17836
rect 5307 17833 5319 17867
rect 7190 17864 7196 17876
rect 7151 17836 7196 17864
rect 5261 17827 5319 17833
rect 7190 17824 7196 17836
rect 7248 17824 7254 17876
rect 8665 17867 8723 17873
rect 8665 17833 8677 17867
rect 8711 17864 8723 17867
rect 8846 17864 8852 17876
rect 8711 17836 8852 17864
rect 8711 17833 8723 17836
rect 8665 17827 8723 17833
rect 8846 17824 8852 17836
rect 8904 17864 8910 17876
rect 8941 17867 8999 17873
rect 8941 17864 8953 17867
rect 8904 17836 8953 17864
rect 8904 17824 8910 17836
rect 8941 17833 8953 17836
rect 8987 17833 8999 17867
rect 9490 17864 9496 17876
rect 9451 17836 9496 17864
rect 8941 17827 8999 17833
rect 9490 17824 9496 17836
rect 9548 17824 9554 17876
rect 9766 17824 9772 17876
rect 9824 17864 9830 17876
rect 9861 17867 9919 17873
rect 9861 17864 9873 17867
rect 9824 17836 9873 17864
rect 9824 17824 9830 17836
rect 9861 17833 9873 17836
rect 9907 17833 9919 17867
rect 9861 17827 9919 17833
rect 11425 17867 11483 17873
rect 11425 17833 11437 17867
rect 11471 17864 11483 17867
rect 11606 17864 11612 17876
rect 11471 17836 11612 17864
rect 11471 17833 11483 17836
rect 11425 17827 11483 17833
rect 11606 17824 11612 17836
rect 11664 17824 11670 17876
rect 14182 17864 14188 17876
rect 11900 17836 14188 17864
rect 4126 17768 4568 17796
rect 5166 17756 5172 17808
rect 5224 17796 5230 17808
rect 5534 17796 5540 17808
rect 5224 17768 5540 17796
rect 5224 17756 5230 17768
rect 5534 17756 5540 17768
rect 5592 17796 5598 17808
rect 5592 17768 6040 17796
rect 5592 17756 5598 17768
rect 4065 17731 4123 17737
rect 4065 17728 4077 17731
rect 3436 17700 4077 17728
rect 2225 17663 2283 17669
rect 2225 17629 2237 17663
rect 2271 17660 2283 17663
rect 2774 17660 2780 17672
rect 2271 17632 2780 17660
rect 2271 17629 2283 17632
rect 2225 17623 2283 17629
rect 2774 17620 2780 17632
rect 2832 17620 2838 17672
rect 2041 17527 2099 17533
rect 2041 17493 2053 17527
rect 2087 17524 2099 17527
rect 2130 17524 2136 17536
rect 2087 17496 2136 17524
rect 2087 17493 2099 17496
rect 2041 17487 2099 17493
rect 2130 17484 2136 17496
rect 2188 17484 2194 17536
rect 3326 17484 3332 17536
rect 3384 17524 3390 17536
rect 3436 17533 3464 17700
rect 4065 17697 4077 17700
rect 4111 17697 4123 17731
rect 4065 17691 4123 17697
rect 5445 17731 5503 17737
rect 5445 17697 5457 17731
rect 5491 17697 5503 17731
rect 5626 17728 5632 17740
rect 5587 17700 5632 17728
rect 5445 17691 5503 17697
rect 4706 17620 4712 17672
rect 4764 17660 4770 17672
rect 5460 17660 5488 17691
rect 5626 17688 5632 17700
rect 5684 17688 5690 17740
rect 6012 17737 6040 17768
rect 7466 17756 7472 17808
rect 7524 17796 7530 17808
rect 8066 17799 8124 17805
rect 8066 17796 8078 17799
rect 7524 17768 8078 17796
rect 7524 17756 7530 17768
rect 8066 17765 8078 17768
rect 8112 17765 8124 17799
rect 8066 17759 8124 17765
rect 5997 17731 6055 17737
rect 5997 17697 6009 17731
rect 6043 17697 6055 17731
rect 6546 17728 6552 17740
rect 6459 17700 6552 17728
rect 5997 17691 6055 17697
rect 6546 17688 6552 17700
rect 6604 17728 6610 17740
rect 8202 17728 8208 17740
rect 6604 17700 8208 17728
rect 6604 17688 6610 17700
rect 8202 17688 8208 17700
rect 8260 17688 8266 17740
rect 9306 17688 9312 17740
rect 9364 17728 9370 17740
rect 10134 17728 10140 17740
rect 9364 17700 10140 17728
rect 9364 17688 9370 17700
rect 10134 17688 10140 17700
rect 10192 17728 10198 17740
rect 10229 17731 10287 17737
rect 10229 17728 10241 17731
rect 10192 17700 10241 17728
rect 10192 17688 10198 17700
rect 10229 17697 10241 17700
rect 10275 17728 10287 17731
rect 11514 17728 11520 17740
rect 10275 17700 11520 17728
rect 10275 17697 10287 17700
rect 10229 17691 10287 17697
rect 11514 17688 11520 17700
rect 11572 17688 11578 17740
rect 11698 17688 11704 17740
rect 11756 17728 11762 17740
rect 11900 17728 11928 17836
rect 14182 17824 14188 17836
rect 14240 17824 14246 17876
rect 16666 17864 16672 17876
rect 16627 17836 16672 17864
rect 16666 17824 16672 17836
rect 16724 17824 16730 17876
rect 16761 17867 16819 17873
rect 16761 17833 16773 17867
rect 16807 17864 16819 17867
rect 17037 17867 17095 17873
rect 17037 17864 17049 17867
rect 16807 17836 17049 17864
rect 16807 17833 16819 17836
rect 16761 17827 16819 17833
rect 17037 17833 17049 17836
rect 17083 17864 17095 17867
rect 17402 17864 17408 17876
rect 17083 17836 17408 17864
rect 17083 17833 17095 17836
rect 17037 17827 17095 17833
rect 17402 17824 17408 17836
rect 17460 17824 17466 17876
rect 11977 17799 12035 17805
rect 11977 17765 11989 17799
rect 12023 17796 12035 17799
rect 12710 17796 12716 17808
rect 12023 17768 12716 17796
rect 12023 17765 12035 17768
rect 11977 17759 12035 17765
rect 12636 17737 12664 17768
rect 12710 17756 12716 17768
rect 12768 17796 12774 17808
rect 12768 17768 13768 17796
rect 12768 17756 12774 17768
rect 13740 17740 13768 17768
rect 15470 17756 15476 17808
rect 15528 17796 15534 17808
rect 16070 17799 16128 17805
rect 16070 17796 16082 17799
rect 15528 17768 16082 17796
rect 15528 17756 15534 17768
rect 16070 17765 16082 17768
rect 16116 17765 16128 17799
rect 16070 17759 16128 17765
rect 16206 17756 16212 17808
rect 16264 17796 16270 17808
rect 17635 17799 17693 17805
rect 17635 17796 17647 17799
rect 16264 17768 17647 17796
rect 16264 17756 16270 17768
rect 17635 17765 17647 17768
rect 17681 17765 17693 17799
rect 17635 17759 17693 17765
rect 12069 17731 12127 17737
rect 12069 17728 12081 17731
rect 11756 17700 12081 17728
rect 11756 17688 11762 17700
rect 12069 17697 12081 17700
rect 12115 17697 12127 17731
rect 12069 17691 12127 17697
rect 12621 17731 12679 17737
rect 12621 17697 12633 17731
rect 12667 17697 12679 17731
rect 13262 17728 13268 17740
rect 13223 17700 13268 17728
rect 12621 17691 12679 17697
rect 13262 17688 13268 17700
rect 13320 17688 13326 17740
rect 13630 17728 13636 17740
rect 13591 17700 13636 17728
rect 13630 17688 13636 17700
rect 13688 17688 13694 17740
rect 13722 17688 13728 17740
rect 13780 17728 13786 17740
rect 14185 17731 14243 17737
rect 14185 17728 14197 17731
rect 13780 17700 14197 17728
rect 13780 17688 13786 17700
rect 14185 17697 14197 17700
rect 14231 17697 14243 17731
rect 14185 17691 14243 17697
rect 7745 17663 7803 17669
rect 4764 17632 6868 17660
rect 4764 17620 4770 17632
rect 4617 17595 4675 17601
rect 4617 17561 4629 17595
rect 4663 17592 4675 17595
rect 5258 17592 5264 17604
rect 4663 17564 5264 17592
rect 4663 17561 4675 17564
rect 4617 17555 4675 17561
rect 5258 17552 5264 17564
rect 5316 17592 5322 17604
rect 6546 17592 6552 17604
rect 5316 17564 6552 17592
rect 5316 17552 5322 17564
rect 6546 17552 6552 17564
rect 6604 17552 6610 17604
rect 6840 17536 6868 17632
rect 7745 17629 7757 17663
rect 7791 17660 7803 17663
rect 8294 17660 8300 17672
rect 7791 17632 8300 17660
rect 7791 17629 7803 17632
rect 7745 17623 7803 17629
rect 8294 17620 8300 17632
rect 8352 17620 8358 17672
rect 12802 17660 12808 17672
rect 12763 17632 12808 17660
rect 12802 17620 12808 17632
rect 12860 17620 12866 17672
rect 14200 17592 14228 17691
rect 17402 17688 17408 17740
rect 17460 17728 17466 17740
rect 17532 17731 17590 17737
rect 17532 17728 17544 17731
rect 17460 17700 17544 17728
rect 17460 17688 17466 17700
rect 17532 17697 17544 17700
rect 17578 17697 17590 17731
rect 17532 17691 17590 17697
rect 18509 17731 18567 17737
rect 18509 17697 18521 17731
rect 18555 17697 18567 17731
rect 18509 17691 18567 17697
rect 14369 17663 14427 17669
rect 14369 17629 14381 17663
rect 14415 17660 14427 17663
rect 15749 17663 15807 17669
rect 15749 17660 15761 17663
rect 14415 17632 15761 17660
rect 14415 17629 14427 17632
rect 14369 17623 14427 17629
rect 15749 17629 15761 17632
rect 15795 17660 15807 17663
rect 17034 17660 17040 17672
rect 15795 17632 17040 17660
rect 15795 17629 15807 17632
rect 15749 17623 15807 17629
rect 17034 17620 17040 17632
rect 17092 17620 17098 17672
rect 18322 17620 18328 17672
rect 18380 17660 18386 17672
rect 18516 17660 18544 17691
rect 18380 17632 18544 17660
rect 18380 17620 18386 17632
rect 15286 17592 15292 17604
rect 14200 17564 15292 17592
rect 15286 17552 15292 17564
rect 15344 17592 15350 17604
rect 16761 17595 16819 17601
rect 16761 17592 16773 17595
rect 15344 17564 16773 17592
rect 15344 17552 15350 17564
rect 16761 17561 16773 17564
rect 16807 17561 16819 17595
rect 16761 17555 16819 17561
rect 3421 17527 3479 17533
rect 3421 17524 3433 17527
rect 3384 17496 3433 17524
rect 3384 17484 3390 17496
rect 3421 17493 3433 17496
rect 3467 17493 3479 17527
rect 3421 17487 3479 17493
rect 3881 17527 3939 17533
rect 3881 17493 3893 17527
rect 3927 17524 3939 17527
rect 4890 17524 4896 17536
rect 3927 17496 4896 17524
rect 3927 17493 3939 17496
rect 3881 17487 3939 17493
rect 4890 17484 4896 17496
rect 4948 17484 4954 17536
rect 5077 17527 5135 17533
rect 5077 17493 5089 17527
rect 5123 17524 5135 17527
rect 5534 17524 5540 17536
rect 5123 17496 5540 17524
rect 5123 17493 5135 17496
rect 5077 17487 5135 17493
rect 5534 17484 5540 17496
rect 5592 17484 5598 17536
rect 6822 17484 6828 17536
rect 6880 17524 6886 17536
rect 7469 17527 7527 17533
rect 7469 17524 7481 17527
rect 6880 17496 7481 17524
rect 6880 17484 6886 17496
rect 7469 17493 7481 17496
rect 7515 17493 7527 17527
rect 7469 17487 7527 17493
rect 10597 17527 10655 17533
rect 10597 17493 10609 17527
rect 10643 17524 10655 17527
rect 10778 17524 10784 17536
rect 10643 17496 10784 17524
rect 10643 17493 10655 17496
rect 10597 17487 10655 17493
rect 10778 17484 10784 17496
rect 10836 17484 10842 17536
rect 13262 17484 13268 17536
rect 13320 17524 13326 17536
rect 15838 17524 15844 17536
rect 13320 17496 15844 17524
rect 13320 17484 13326 17496
rect 15838 17484 15844 17496
rect 15896 17484 15902 17536
rect 18690 17524 18696 17536
rect 18651 17496 18696 17524
rect 18690 17484 18696 17496
rect 18748 17484 18754 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 2317 17323 2375 17329
rect 2317 17289 2329 17323
rect 2363 17320 2375 17323
rect 2682 17320 2688 17332
rect 2363 17292 2688 17320
rect 2363 17289 2375 17292
rect 2317 17283 2375 17289
rect 2682 17280 2688 17292
rect 2740 17320 2746 17332
rect 2866 17320 2872 17332
rect 2740 17292 2872 17320
rect 2740 17280 2746 17292
rect 2866 17280 2872 17292
rect 2924 17280 2930 17332
rect 10134 17320 10140 17332
rect 10095 17292 10140 17320
rect 10134 17280 10140 17292
rect 10192 17280 10198 17332
rect 13078 17280 13084 17332
rect 13136 17320 13142 17332
rect 13449 17323 13507 17329
rect 13449 17320 13461 17323
rect 13136 17292 13461 17320
rect 13136 17280 13142 17292
rect 13449 17289 13461 17292
rect 13495 17320 13507 17323
rect 13630 17320 13636 17332
rect 13495 17292 13636 17320
rect 13495 17289 13507 17292
rect 13449 17283 13507 17289
rect 13630 17280 13636 17292
rect 13688 17280 13694 17332
rect 13814 17280 13820 17332
rect 13872 17320 13878 17332
rect 17034 17320 17040 17332
rect 13872 17292 16942 17320
rect 16995 17292 17040 17320
rect 13872 17280 13878 17292
rect 3973 17255 4031 17261
rect 3973 17221 3985 17255
rect 4019 17252 4031 17255
rect 4614 17252 4620 17264
rect 4019 17224 4620 17252
rect 4019 17221 4031 17224
rect 3973 17215 4031 17221
rect 4614 17212 4620 17224
rect 4672 17252 4678 17264
rect 5534 17252 5540 17264
rect 4672 17224 5540 17252
rect 4672 17212 4678 17224
rect 5534 17212 5540 17224
rect 5592 17212 5598 17264
rect 14826 17252 14832 17264
rect 14787 17224 14832 17252
rect 14826 17212 14832 17224
rect 14884 17212 14890 17264
rect 15197 17255 15255 17261
rect 15197 17221 15209 17255
rect 15243 17252 15255 17255
rect 15286 17252 15292 17264
rect 15243 17224 15292 17252
rect 15243 17221 15255 17224
rect 15197 17215 15255 17221
rect 15286 17212 15292 17224
rect 15344 17212 15350 17264
rect 16301 17255 16359 17261
rect 16301 17221 16313 17255
rect 16347 17252 16359 17255
rect 16482 17252 16488 17264
rect 16347 17224 16488 17252
rect 16347 17221 16359 17224
rect 16301 17215 16359 17221
rect 16482 17212 16488 17224
rect 16540 17212 16546 17264
rect 16914 17252 16942 17292
rect 17034 17280 17040 17292
rect 17092 17280 17098 17332
rect 18322 17280 18328 17332
rect 18380 17320 18386 17332
rect 18877 17323 18935 17329
rect 18877 17320 18889 17323
rect 18380 17292 18889 17320
rect 18380 17280 18386 17292
rect 18877 17289 18889 17292
rect 18923 17289 18935 17323
rect 18877 17283 18935 17289
rect 18233 17255 18291 17261
rect 16914 17224 18000 17252
rect 4341 17187 4399 17193
rect 4341 17153 4353 17187
rect 4387 17184 4399 17187
rect 6641 17187 6699 17193
rect 4387 17156 5304 17184
rect 4387 17153 4399 17156
rect 4341 17147 4399 17153
rect 5276 17128 5304 17156
rect 6641 17153 6653 17187
rect 6687 17184 6699 17187
rect 10597 17187 10655 17193
rect 6687 17156 9904 17184
rect 6687 17153 6699 17156
rect 6641 17147 6699 17153
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 2130 17116 2136 17128
rect 1443 17088 2136 17116
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 2130 17076 2136 17088
rect 2188 17076 2194 17128
rect 4706 17116 4712 17128
rect 4667 17088 4712 17116
rect 4706 17076 4712 17088
rect 4764 17076 4770 17128
rect 4890 17116 4896 17128
rect 4851 17088 4896 17116
rect 4890 17076 4896 17088
rect 4948 17076 4954 17128
rect 5258 17076 5264 17128
rect 5316 17116 5322 17128
rect 5316 17088 5361 17116
rect 5316 17076 5322 17088
rect 5534 17076 5540 17128
rect 5592 17116 5598 17128
rect 5813 17119 5871 17125
rect 5813 17116 5825 17119
rect 5592 17088 5825 17116
rect 5592 17076 5598 17088
rect 5813 17085 5825 17088
rect 5859 17116 5871 17119
rect 6822 17116 6828 17128
rect 5859 17088 6316 17116
rect 6783 17088 6828 17116
rect 5859 17085 5871 17088
rect 5813 17079 5871 17085
rect 2958 17048 2964 17060
rect 2919 17020 2964 17048
rect 2958 17008 2964 17020
rect 3016 17008 3022 17060
rect 3053 17051 3111 17057
rect 3053 17017 3065 17051
rect 3099 17017 3111 17051
rect 3602 17048 3608 17060
rect 3563 17020 3608 17048
rect 3053 17011 3111 17017
rect 106 16940 112 16992
rect 164 16980 170 16992
rect 1581 16983 1639 16989
rect 1581 16980 1593 16983
rect 164 16952 1593 16980
rect 164 16940 170 16952
rect 1581 16949 1593 16952
rect 1627 16949 1639 16983
rect 1581 16943 1639 16949
rect 2777 16983 2835 16989
rect 2777 16949 2789 16983
rect 2823 16980 2835 16983
rect 3068 16980 3096 17011
rect 3602 17008 3608 17020
rect 3660 17008 3666 17060
rect 6288 17057 6316 17088
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 7282 17116 7288 17128
rect 7243 17088 7288 17116
rect 7282 17076 7288 17088
rect 7340 17076 7346 17128
rect 7650 17076 7656 17128
rect 7708 17116 7714 17128
rect 7852 17125 7880 17156
rect 7837 17119 7895 17125
rect 7837 17116 7849 17119
rect 7708 17088 7849 17116
rect 7708 17076 7714 17088
rect 7837 17085 7849 17088
rect 7883 17085 7895 17119
rect 8202 17116 8208 17128
rect 7837 17079 7895 17085
rect 7944 17088 8208 17116
rect 6273 17051 6331 17057
rect 6273 17017 6285 17051
rect 6319 17048 6331 17051
rect 6362 17048 6368 17060
rect 6319 17020 6368 17048
rect 6319 17017 6331 17020
rect 6273 17011 6331 17017
rect 6362 17008 6368 17020
rect 6420 17048 6426 17060
rect 7944 17048 7972 17088
rect 8202 17076 8208 17088
rect 8260 17076 8266 17128
rect 9876 17116 9904 17156
rect 10597 17153 10609 17187
rect 10643 17184 10655 17187
rect 10643 17156 11008 17184
rect 10643 17153 10655 17156
rect 10597 17147 10655 17153
rect 10689 17119 10747 17125
rect 10689 17116 10701 17119
rect 9876 17088 10701 17116
rect 10689 17085 10701 17088
rect 10735 17085 10747 17119
rect 10689 17079 10747 17085
rect 8294 17048 8300 17060
rect 6420 17020 7972 17048
rect 8255 17020 8300 17048
rect 6420 17008 6426 17020
rect 8294 17008 8300 17020
rect 8352 17008 8358 17060
rect 9214 17048 9220 17060
rect 9175 17020 9220 17048
rect 9214 17008 9220 17020
rect 9272 17008 9278 17060
rect 9309 17051 9367 17057
rect 9309 17017 9321 17051
rect 9355 17048 9367 17051
rect 9398 17048 9404 17060
rect 9355 17020 9404 17048
rect 9355 17017 9367 17020
rect 9309 17011 9367 17017
rect 3510 16980 3516 16992
rect 2823 16952 3516 16980
rect 2823 16949 2835 16952
rect 2777 16943 2835 16949
rect 3510 16940 3516 16952
rect 3568 16940 3574 16992
rect 4522 16980 4528 16992
rect 4483 16952 4528 16980
rect 4522 16940 4528 16952
rect 4580 16940 4586 16992
rect 7466 16940 7472 16992
rect 7524 16980 7530 16992
rect 8573 16983 8631 16989
rect 8573 16980 8585 16983
rect 7524 16952 8585 16980
rect 7524 16940 7530 16952
rect 8573 16949 8585 16952
rect 8619 16949 8631 16983
rect 8573 16943 8631 16949
rect 9033 16983 9091 16989
rect 9033 16949 9045 16983
rect 9079 16980 9091 16983
rect 9324 16980 9352 17011
rect 9398 17008 9404 17020
rect 9456 17008 9462 17060
rect 9861 17051 9919 17057
rect 9861 17017 9873 17051
rect 9907 17048 9919 17051
rect 10042 17048 10048 17060
rect 9907 17020 10048 17048
rect 9907 17017 9919 17020
rect 9861 17011 9919 17017
rect 10042 17008 10048 17020
rect 10100 17008 10106 17060
rect 10704 17048 10732 17079
rect 10778 17076 10784 17128
rect 10836 17116 10842 17128
rect 10980 17125 11008 17156
rect 11882 17144 11888 17196
rect 11940 17184 11946 17196
rect 12253 17187 12311 17193
rect 12253 17184 12265 17187
rect 11940 17156 12265 17184
rect 11940 17144 11946 17156
rect 12253 17153 12265 17156
rect 12299 17184 12311 17187
rect 12299 17156 12664 17184
rect 12299 17153 12311 17156
rect 12253 17147 12311 17153
rect 10965 17119 11023 17125
rect 10836 17088 10881 17116
rect 10836 17076 10842 17088
rect 10965 17085 10977 17119
rect 11011 17116 11023 17119
rect 12526 17116 12532 17128
rect 11011 17088 12532 17116
rect 11011 17085 11023 17088
rect 10965 17079 11023 17085
rect 12526 17076 12532 17088
rect 12584 17076 12590 17128
rect 12636 17125 12664 17156
rect 13722 17144 13728 17196
rect 13780 17184 13786 17196
rect 13998 17184 14004 17196
rect 13780 17156 14004 17184
rect 13780 17144 13786 17156
rect 13998 17144 14004 17156
rect 14056 17184 14062 17196
rect 15749 17187 15807 17193
rect 14056 17156 14314 17184
rect 14056 17144 14062 17156
rect 12621 17119 12679 17125
rect 12621 17085 12633 17119
rect 12667 17116 12679 17119
rect 12894 17116 12900 17128
rect 12667 17088 12900 17116
rect 12667 17085 12679 17088
rect 12621 17079 12679 17085
rect 12894 17076 12900 17088
rect 12952 17076 12958 17128
rect 13906 17116 13912 17128
rect 13867 17088 13912 17116
rect 13906 17076 13912 17088
rect 13964 17076 13970 17128
rect 11054 17048 11060 17060
rect 10704 17020 11060 17048
rect 11054 17008 11060 17020
rect 11112 17008 11118 17060
rect 12434 17048 12440 17060
rect 12395 17020 12440 17048
rect 12434 17008 12440 17020
rect 12492 17008 12498 17060
rect 12989 17051 13047 17057
rect 12989 17017 13001 17051
rect 13035 17048 13047 17051
rect 13998 17048 14004 17060
rect 13035 17020 14004 17048
rect 13035 17017 13047 17020
rect 12989 17011 13047 17017
rect 13998 17008 14004 17020
rect 14056 17008 14062 17060
rect 14286 17057 14314 17156
rect 15749 17153 15761 17187
rect 15795 17184 15807 17187
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 15795 17156 16681 17184
rect 15795 17153 15807 17156
rect 15749 17147 15807 17153
rect 16669 17153 16681 17156
rect 16715 17184 16727 17187
rect 16850 17184 16856 17196
rect 16715 17156 16856 17184
rect 16715 17153 16727 17156
rect 16669 17147 16727 17153
rect 16850 17144 16856 17156
rect 16908 17144 16914 17196
rect 17972 17116 18000 17224
rect 18233 17221 18245 17255
rect 18279 17252 18291 17255
rect 18506 17252 18512 17264
rect 18279 17224 18512 17252
rect 18279 17221 18291 17224
rect 18233 17215 18291 17221
rect 18506 17212 18512 17224
rect 18564 17212 18570 17264
rect 18049 17119 18107 17125
rect 18049 17116 18061 17119
rect 17972 17088 18061 17116
rect 18049 17085 18061 17088
rect 18095 17116 18107 17119
rect 18509 17119 18567 17125
rect 18509 17116 18521 17119
rect 18095 17088 18521 17116
rect 18095 17085 18107 17088
rect 18049 17079 18107 17085
rect 18509 17085 18521 17088
rect 18555 17085 18567 17119
rect 18509 17079 18567 17085
rect 14271 17051 14329 17057
rect 14271 17017 14283 17051
rect 14317 17017 14329 17051
rect 14271 17011 14329 17017
rect 11146 16980 11152 16992
rect 9079 16952 9352 16980
rect 11107 16952 11152 16980
rect 9079 16949 9091 16952
rect 9033 16943 9091 16949
rect 11146 16940 11152 16952
rect 11204 16940 11210 16992
rect 11698 16940 11704 16992
rect 11756 16980 11762 16992
rect 11793 16983 11851 16989
rect 11793 16980 11805 16983
rect 11756 16952 11805 16980
rect 11756 16940 11762 16952
rect 11793 16949 11805 16952
rect 11839 16949 11851 16983
rect 11793 16943 11851 16949
rect 13817 16983 13875 16989
rect 13817 16949 13829 16983
rect 13863 16980 13875 16983
rect 14286 16980 14314 17011
rect 15562 17008 15568 17060
rect 15620 17048 15626 17060
rect 15841 17051 15899 17057
rect 15841 17048 15853 17051
rect 15620 17020 15853 17048
rect 15620 17008 15626 17020
rect 15841 17017 15853 17020
rect 15887 17017 15899 17051
rect 15841 17011 15899 17017
rect 14458 16980 14464 16992
rect 13863 16952 14464 16980
rect 13863 16949 13875 16952
rect 13817 16943 13875 16949
rect 14458 16940 14464 16952
rect 14516 16980 14522 16992
rect 15470 16980 15476 16992
rect 14516 16952 15476 16980
rect 14516 16940 14522 16952
rect 15470 16940 15476 16952
rect 15528 16940 15534 16992
rect 17402 16940 17408 16992
rect 17460 16980 17466 16992
rect 17497 16983 17555 16989
rect 17497 16980 17509 16983
rect 17460 16952 17509 16980
rect 17460 16940 17466 16952
rect 17497 16949 17509 16952
rect 17543 16949 17555 16983
rect 17497 16943 17555 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 2774 16776 2780 16788
rect 2735 16748 2780 16776
rect 2774 16736 2780 16748
rect 2832 16776 2838 16788
rect 4522 16776 4528 16788
rect 2832 16748 4528 16776
rect 2832 16736 2838 16748
rect 4522 16736 4528 16748
rect 4580 16736 4586 16788
rect 4890 16736 4896 16788
rect 4948 16776 4954 16788
rect 6457 16779 6515 16785
rect 6457 16776 6469 16779
rect 4948 16748 6469 16776
rect 4948 16736 4954 16748
rect 6457 16745 6469 16748
rect 6503 16745 6515 16779
rect 6457 16739 6515 16745
rect 3099 16711 3157 16717
rect 3099 16677 3111 16711
rect 3145 16708 3157 16711
rect 3878 16708 3884 16720
rect 3145 16680 3884 16708
rect 3145 16677 3157 16680
rect 3099 16671 3157 16677
rect 3878 16668 3884 16680
rect 3936 16708 3942 16720
rect 4157 16711 4215 16717
rect 4157 16708 4169 16711
rect 3936 16680 4169 16708
rect 3936 16668 3942 16680
rect 4157 16677 4169 16680
rect 4203 16677 4215 16711
rect 4157 16671 4215 16677
rect 4249 16711 4307 16717
rect 4249 16677 4261 16711
rect 4295 16708 4307 16711
rect 4338 16708 4344 16720
rect 4295 16680 4344 16708
rect 4295 16677 4307 16680
rect 4249 16671 4307 16677
rect 4338 16668 4344 16680
rect 4396 16668 4402 16720
rect 6472 16708 6500 16739
rect 8294 16736 8300 16788
rect 8352 16776 8358 16788
rect 8757 16779 8815 16785
rect 8757 16776 8769 16779
rect 8352 16748 8769 16776
rect 8352 16736 8358 16748
rect 8757 16745 8769 16748
rect 8803 16745 8815 16779
rect 8757 16739 8815 16745
rect 13722 16736 13728 16788
rect 13780 16776 13786 16788
rect 13817 16779 13875 16785
rect 13817 16776 13829 16779
rect 13780 16748 13829 16776
rect 13780 16736 13786 16748
rect 13817 16745 13829 16748
rect 13863 16745 13875 16779
rect 13817 16739 13875 16745
rect 15562 16736 15568 16788
rect 15620 16776 15626 16788
rect 16301 16779 16359 16785
rect 16301 16776 16313 16779
rect 15620 16748 16313 16776
rect 15620 16736 15626 16748
rect 16301 16745 16313 16748
rect 16347 16745 16359 16779
rect 16850 16776 16856 16788
rect 16811 16748 16856 16776
rect 16301 16739 16359 16745
rect 16850 16736 16856 16748
rect 16908 16736 16914 16788
rect 7282 16708 7288 16720
rect 6472 16680 7288 16708
rect 2038 16640 2044 16652
rect 1999 16612 2044 16640
rect 2038 16600 2044 16612
rect 2096 16600 2102 16652
rect 2866 16600 2872 16652
rect 2924 16640 2930 16652
rect 2996 16643 3054 16649
rect 2996 16640 3008 16643
rect 2924 16612 3008 16640
rect 2924 16600 2930 16612
rect 2996 16609 3008 16612
rect 3042 16609 3054 16643
rect 2996 16603 3054 16609
rect 5534 16600 5540 16652
rect 5592 16640 5598 16652
rect 5664 16643 5722 16649
rect 5664 16640 5676 16643
rect 5592 16612 5676 16640
rect 5592 16600 5598 16612
rect 5664 16609 5676 16612
rect 5710 16609 5722 16643
rect 5664 16603 5722 16609
rect 6178 16600 6184 16652
rect 6236 16640 6242 16652
rect 6641 16643 6699 16649
rect 6641 16640 6653 16643
rect 6236 16612 6653 16640
rect 6236 16600 6242 16612
rect 6641 16609 6653 16612
rect 6687 16640 6699 16643
rect 6822 16640 6828 16652
rect 6687 16612 6828 16640
rect 6687 16609 6699 16612
rect 6641 16603 6699 16609
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 7116 16649 7144 16680
rect 7282 16668 7288 16680
rect 7340 16668 7346 16720
rect 9858 16708 9864 16720
rect 9819 16680 9864 16708
rect 9858 16668 9864 16680
rect 9916 16668 9922 16720
rect 10781 16711 10839 16717
rect 10781 16677 10793 16711
rect 10827 16708 10839 16711
rect 11054 16708 11060 16720
rect 10827 16680 11060 16708
rect 10827 16677 10839 16680
rect 10781 16671 10839 16677
rect 11054 16668 11060 16680
rect 11112 16708 11118 16720
rect 11112 16680 12480 16708
rect 11112 16668 11118 16680
rect 12452 16652 12480 16680
rect 14366 16668 14372 16720
rect 14424 16708 14430 16720
rect 15473 16711 15531 16717
rect 15473 16708 15485 16711
rect 14424 16680 15485 16708
rect 14424 16668 14430 16680
rect 15473 16677 15485 16680
rect 15519 16677 15531 16711
rect 15473 16671 15531 16677
rect 15838 16668 15844 16720
rect 15896 16708 15902 16720
rect 16025 16711 16083 16717
rect 16025 16708 16037 16711
rect 15896 16680 16037 16708
rect 15896 16668 15902 16680
rect 16025 16677 16037 16680
rect 16071 16708 16083 16711
rect 16482 16708 16488 16720
rect 16071 16680 16488 16708
rect 16071 16677 16083 16680
rect 16025 16671 16083 16677
rect 16482 16668 16488 16680
rect 16540 16668 16546 16720
rect 7101 16643 7159 16649
rect 7101 16609 7113 16643
rect 7147 16609 7159 16643
rect 7650 16640 7656 16652
rect 7611 16612 7656 16640
rect 7101 16603 7159 16609
rect 7650 16600 7656 16612
rect 7708 16600 7714 16652
rect 8021 16643 8079 16649
rect 8021 16609 8033 16643
rect 8067 16640 8079 16643
rect 8110 16640 8116 16652
rect 8067 16612 8116 16640
rect 8067 16609 8079 16612
rect 8021 16603 8079 16609
rect 8110 16600 8116 16612
rect 8168 16600 8174 16652
rect 11698 16600 11704 16652
rect 11756 16640 11762 16652
rect 11885 16643 11943 16649
rect 11885 16640 11897 16643
rect 11756 16612 11897 16640
rect 11756 16600 11762 16612
rect 11885 16609 11897 16612
rect 11931 16609 11943 16643
rect 12342 16640 12348 16652
rect 12303 16612 12348 16640
rect 11885 16603 11943 16609
rect 12342 16600 12348 16612
rect 12400 16600 12406 16652
rect 12434 16600 12440 16652
rect 12492 16640 12498 16652
rect 12492 16612 12756 16640
rect 12492 16600 12498 16612
rect 3602 16532 3608 16584
rect 3660 16572 3666 16584
rect 4433 16575 4491 16581
rect 4433 16572 4445 16575
rect 3660 16544 4445 16572
rect 3660 16532 3666 16544
rect 4433 16541 4445 16544
rect 4479 16541 4491 16575
rect 4433 16535 4491 16541
rect 7190 16532 7196 16584
rect 7248 16572 7254 16584
rect 9125 16575 9183 16581
rect 9125 16572 9137 16575
rect 7248 16544 9137 16572
rect 7248 16532 7254 16544
rect 9125 16541 9137 16544
rect 9171 16572 9183 16575
rect 9214 16572 9220 16584
rect 9171 16544 9220 16572
rect 9171 16541 9183 16544
rect 9125 16535 9183 16541
rect 9214 16532 9220 16544
rect 9272 16532 9278 16584
rect 9766 16572 9772 16584
rect 9727 16544 9772 16572
rect 9766 16532 9772 16544
rect 9824 16532 9830 16584
rect 10042 16572 10048 16584
rect 10003 16544 10048 16572
rect 10042 16532 10048 16544
rect 10100 16532 10106 16584
rect 12618 16572 12624 16584
rect 12579 16544 12624 16572
rect 12618 16532 12624 16544
rect 12676 16532 12682 16584
rect 12728 16572 12756 16612
rect 12802 16600 12808 16652
rect 12860 16640 12866 16652
rect 13446 16640 13452 16652
rect 12860 16612 13452 16640
rect 12860 16600 12866 16612
rect 13446 16600 13452 16612
rect 13504 16600 13510 16652
rect 16114 16600 16120 16652
rect 16172 16640 16178 16652
rect 17865 16643 17923 16649
rect 17865 16640 17877 16643
rect 16172 16612 17877 16640
rect 16172 16600 16178 16612
rect 17865 16609 17877 16612
rect 17911 16640 17923 16643
rect 18598 16640 18604 16652
rect 17911 16612 18604 16640
rect 17911 16609 17923 16612
rect 17865 16603 17923 16609
rect 18598 16600 18604 16612
rect 18656 16600 18662 16652
rect 12989 16575 13047 16581
rect 12989 16572 13001 16575
rect 12728 16544 13001 16572
rect 12989 16541 13001 16544
rect 13035 16572 13047 16575
rect 14734 16572 14740 16584
rect 13035 16544 14740 16572
rect 13035 16541 13047 16544
rect 12989 16535 13047 16541
rect 14734 16532 14740 16544
rect 14792 16532 14798 16584
rect 15381 16575 15439 16581
rect 15381 16541 15393 16575
rect 15427 16572 15439 16575
rect 16574 16572 16580 16584
rect 15427 16544 16580 16572
rect 15427 16541 15439 16544
rect 15381 16535 15439 16541
rect 16574 16532 16580 16544
rect 16632 16532 16638 16584
rect 1486 16464 1492 16516
rect 1544 16504 1550 16516
rect 2409 16507 2467 16513
rect 2409 16504 2421 16507
rect 1544 16476 2421 16504
rect 1544 16464 1550 16476
rect 2409 16473 2421 16476
rect 2455 16473 2467 16507
rect 2409 16467 2467 16473
rect 3881 16507 3939 16513
rect 3881 16473 3893 16507
rect 3927 16504 3939 16507
rect 4706 16504 4712 16516
rect 3927 16476 4712 16504
rect 3927 16473 3939 16476
rect 3881 16467 3939 16473
rect 4706 16464 4712 16476
rect 4764 16464 4770 16516
rect 8018 16504 8024 16516
rect 7979 16476 8024 16504
rect 8018 16464 8024 16476
rect 8076 16464 8082 16516
rect 10778 16464 10784 16516
rect 10836 16504 10842 16516
rect 11149 16507 11207 16513
rect 11149 16504 11161 16507
rect 10836 16476 11161 16504
rect 10836 16464 10842 16476
rect 11149 16473 11161 16476
rect 11195 16504 11207 16507
rect 13814 16504 13820 16516
rect 11195 16476 13820 16504
rect 11195 16473 11207 16476
rect 11149 16467 11207 16473
rect 13814 16464 13820 16476
rect 13872 16464 13878 16516
rect 13906 16464 13912 16516
rect 13964 16504 13970 16516
rect 14645 16507 14703 16513
rect 14645 16504 14657 16507
rect 13964 16476 14657 16504
rect 13964 16464 13970 16476
rect 14645 16473 14657 16476
rect 14691 16473 14703 16507
rect 14645 16467 14703 16473
rect 16022 16464 16028 16516
rect 16080 16504 16086 16516
rect 18049 16507 18107 16513
rect 18049 16504 18061 16507
rect 16080 16476 18061 16504
rect 16080 16464 16086 16476
rect 18049 16473 18061 16476
rect 18095 16473 18107 16507
rect 18049 16467 18107 16473
rect 1670 16436 1676 16448
rect 1631 16408 1676 16436
rect 1670 16396 1676 16408
rect 1728 16396 1734 16448
rect 3418 16436 3424 16448
rect 3379 16408 3424 16436
rect 3418 16396 3424 16408
rect 3476 16396 3482 16448
rect 5166 16436 5172 16448
rect 5127 16408 5172 16436
rect 5166 16396 5172 16408
rect 5224 16396 5230 16448
rect 5767 16439 5825 16445
rect 5767 16405 5779 16439
rect 5813 16436 5825 16439
rect 5994 16436 6000 16448
rect 5813 16408 6000 16436
rect 5813 16405 5825 16408
rect 5767 16399 5825 16405
rect 5994 16396 6000 16408
rect 6052 16396 6058 16448
rect 6178 16436 6184 16448
rect 6139 16408 6184 16436
rect 6178 16396 6184 16408
rect 6236 16396 6242 16448
rect 7282 16396 7288 16448
rect 7340 16436 7346 16448
rect 8386 16436 8392 16448
rect 7340 16408 8392 16436
rect 7340 16396 7346 16408
rect 8386 16396 8392 16408
rect 8444 16396 8450 16448
rect 14366 16436 14372 16448
rect 14327 16408 14372 16436
rect 14366 16396 14372 16408
rect 14424 16396 14430 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 4065 16235 4123 16241
rect 4065 16201 4077 16235
rect 4111 16232 4123 16235
rect 4338 16232 4344 16244
rect 4111 16204 4344 16232
rect 4111 16201 4123 16204
rect 4065 16195 4123 16201
rect 4338 16192 4344 16204
rect 4396 16192 4402 16244
rect 5994 16192 6000 16244
rect 6052 16232 6058 16244
rect 8849 16235 8907 16241
rect 8849 16232 8861 16235
rect 6052 16204 8861 16232
rect 6052 16192 6058 16204
rect 8849 16201 8861 16204
rect 8895 16232 8907 16235
rect 9766 16232 9772 16244
rect 8895 16204 9772 16232
rect 8895 16201 8907 16204
rect 8849 16195 8907 16201
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 11882 16232 11888 16244
rect 11843 16204 11888 16232
rect 11882 16192 11888 16204
rect 11940 16192 11946 16244
rect 12710 16232 12716 16244
rect 12671 16204 12716 16232
rect 12710 16192 12716 16204
rect 12768 16192 12774 16244
rect 13722 16192 13728 16244
rect 13780 16232 13786 16244
rect 14185 16235 14243 16241
rect 14185 16232 14197 16235
rect 13780 16204 14197 16232
rect 13780 16192 13786 16204
rect 14185 16201 14197 16204
rect 14231 16201 14243 16235
rect 14185 16195 14243 16201
rect 14366 16192 14372 16244
rect 14424 16232 14430 16244
rect 14645 16235 14703 16241
rect 14645 16232 14657 16235
rect 14424 16204 14657 16232
rect 14424 16192 14430 16204
rect 14645 16201 14657 16204
rect 14691 16201 14703 16235
rect 14645 16195 14703 16201
rect 14826 16192 14832 16244
rect 14884 16232 14890 16244
rect 15013 16235 15071 16241
rect 15013 16232 15025 16235
rect 14884 16204 15025 16232
rect 14884 16192 14890 16204
rect 15013 16201 15025 16204
rect 15059 16232 15071 16235
rect 15378 16232 15384 16244
rect 15059 16204 15384 16232
rect 15059 16201 15071 16204
rect 15013 16195 15071 16201
rect 15378 16192 15384 16204
rect 15436 16192 15442 16244
rect 16298 16192 16304 16244
rect 16356 16232 16362 16244
rect 16945 16235 17003 16241
rect 16945 16232 16957 16235
rect 16356 16204 16957 16232
rect 16356 16192 16362 16204
rect 16945 16201 16957 16204
rect 16991 16201 17003 16235
rect 18598 16232 18604 16244
rect 18511 16204 18604 16232
rect 16945 16195 17003 16201
rect 18598 16192 18604 16204
rect 18656 16232 18662 16244
rect 19518 16232 19524 16244
rect 18656 16204 19524 16232
rect 18656 16192 18662 16204
rect 19518 16192 19524 16204
rect 19576 16192 19582 16244
rect 2866 16164 2872 16176
rect 2779 16136 2872 16164
rect 2866 16124 2872 16136
rect 2924 16164 2930 16176
rect 3878 16164 3884 16176
rect 2924 16136 3884 16164
rect 2924 16124 2930 16136
rect 3878 16124 3884 16136
rect 3936 16164 3942 16176
rect 5074 16164 5080 16176
rect 3936 16136 5080 16164
rect 3936 16124 3942 16136
rect 5074 16124 5080 16136
rect 5132 16124 5138 16176
rect 6546 16164 6552 16176
rect 6507 16136 6552 16164
rect 6546 16124 6552 16136
rect 6604 16124 6610 16176
rect 7101 16167 7159 16173
rect 7101 16133 7113 16167
rect 7147 16164 7159 16167
rect 7558 16164 7564 16176
rect 7147 16136 7564 16164
rect 7147 16133 7159 16136
rect 7101 16127 7159 16133
rect 7558 16124 7564 16136
rect 7616 16124 7622 16176
rect 3053 16099 3111 16105
rect 3053 16065 3065 16099
rect 3099 16096 3111 16099
rect 3418 16096 3424 16108
rect 3099 16068 3424 16096
rect 3099 16065 3111 16068
rect 3053 16059 3111 16065
rect 3418 16056 3424 16068
rect 3476 16056 3482 16108
rect 3510 16056 3516 16108
rect 3568 16096 3574 16108
rect 4525 16099 4583 16105
rect 4525 16096 4537 16099
rect 3568 16068 4537 16096
rect 3568 16056 3574 16068
rect 4525 16065 4537 16068
rect 4571 16065 4583 16099
rect 4525 16059 4583 16065
rect 7653 16099 7711 16105
rect 7653 16065 7665 16099
rect 7699 16096 7711 16099
rect 8018 16096 8024 16108
rect 7699 16068 8024 16096
rect 7699 16065 7711 16068
rect 7653 16059 7711 16065
rect 8018 16056 8024 16068
rect 8076 16056 8082 16108
rect 9398 16096 9404 16108
rect 9359 16068 9404 16096
rect 9398 16056 9404 16068
rect 9456 16056 9462 16108
rect 11054 16056 11060 16108
rect 11112 16096 11118 16108
rect 12728 16096 12756 16192
rect 15838 16164 15844 16176
rect 15799 16136 15844 16164
rect 15838 16124 15844 16136
rect 15896 16124 15902 16176
rect 17037 16167 17095 16173
rect 17037 16133 17049 16167
rect 17083 16164 17095 16167
rect 17313 16167 17371 16173
rect 17313 16164 17325 16167
rect 17083 16136 17325 16164
rect 17083 16133 17095 16136
rect 17037 16127 17095 16133
rect 17313 16133 17325 16136
rect 17359 16164 17371 16167
rect 19978 16164 19984 16176
rect 17359 16136 19984 16164
rect 17359 16133 17371 16136
rect 17313 16127 17371 16133
rect 19978 16124 19984 16136
rect 20036 16124 20042 16176
rect 13906 16096 13912 16108
rect 11112 16068 12664 16096
rect 12728 16068 13676 16096
rect 13867 16068 13912 16096
rect 11112 16056 11118 16068
rect 4338 15988 4344 16040
rect 4396 16028 4402 16040
rect 4617 16031 4675 16037
rect 4617 16028 4629 16031
rect 4396 16000 4629 16028
rect 4396 15988 4402 16000
rect 4617 15997 4629 16000
rect 4663 15997 4675 16031
rect 4617 15991 4675 15997
rect 8573 16031 8631 16037
rect 8573 15997 8585 16031
rect 8619 16028 8631 16031
rect 9309 16031 9367 16037
rect 9309 16028 9321 16031
rect 8619 16000 9321 16028
rect 8619 15997 8631 16000
rect 8573 15991 8631 15997
rect 9309 15997 9321 16000
rect 9355 16028 9367 16031
rect 9858 16028 9864 16040
rect 9355 16000 9864 16028
rect 9355 15997 9367 16000
rect 9309 15991 9367 15997
rect 9858 15988 9864 16000
rect 9916 16028 9922 16040
rect 10045 16031 10103 16037
rect 10045 16028 10057 16031
rect 9916 16000 10057 16028
rect 9916 15988 9922 16000
rect 10045 15997 10057 16000
rect 10091 16028 10103 16031
rect 10413 16031 10471 16037
rect 10413 16028 10425 16031
rect 10091 16000 10425 16028
rect 10091 15997 10103 16000
rect 10045 15991 10103 15997
rect 10413 15997 10425 16000
rect 10459 15997 10471 16031
rect 10413 15991 10471 15997
rect 11149 16031 11207 16037
rect 11149 15997 11161 16031
rect 11195 16028 11207 16031
rect 11882 16028 11888 16040
rect 11195 16000 11888 16028
rect 11195 15997 11207 16000
rect 11149 15991 11207 15997
rect 11882 15988 11888 16000
rect 11940 15988 11946 16040
rect 12636 16028 12664 16068
rect 12989 16031 13047 16037
rect 12989 16028 13001 16031
rect 12636 16000 13001 16028
rect 12989 15997 13001 16000
rect 13035 16028 13047 16031
rect 13173 16031 13231 16037
rect 13173 16028 13185 16031
rect 13035 16000 13185 16028
rect 13035 15997 13047 16000
rect 12989 15991 13047 15997
rect 13173 15997 13185 16000
rect 13219 16028 13231 16031
rect 13262 16028 13268 16040
rect 13219 16000 13268 16028
rect 13219 15997 13231 16000
rect 13173 15991 13231 15997
rect 13262 15988 13268 16000
rect 13320 15988 13326 16040
rect 13648 16037 13676 16068
rect 13906 16056 13912 16068
rect 13964 16056 13970 16108
rect 15120 16068 18092 16096
rect 13633 16031 13691 16037
rect 13633 15997 13645 16031
rect 13679 16028 13691 16031
rect 14274 16028 14280 16040
rect 13679 16000 14280 16028
rect 13679 15997 13691 16000
rect 13633 15991 13691 15997
rect 14274 15988 14280 16000
rect 14332 15988 14338 16040
rect 1486 15960 1492 15972
rect 1447 15932 1492 15960
rect 1486 15920 1492 15932
rect 1544 15920 1550 15972
rect 1581 15963 1639 15969
rect 1581 15929 1593 15963
rect 1627 15960 1639 15963
rect 1670 15960 1676 15972
rect 1627 15932 1676 15960
rect 1627 15929 1639 15932
rect 1581 15923 1639 15929
rect 1670 15920 1676 15932
rect 1728 15920 1734 15972
rect 2133 15963 2191 15969
rect 2133 15929 2145 15963
rect 2179 15960 2191 15963
rect 2222 15960 2228 15972
rect 2179 15932 2228 15960
rect 2179 15929 2191 15932
rect 2133 15923 2191 15929
rect 2222 15920 2228 15932
rect 2280 15920 2286 15972
rect 3145 15963 3203 15969
rect 3145 15929 3157 15963
rect 3191 15960 3203 15963
rect 3510 15960 3516 15972
rect 3191 15932 3516 15960
rect 3191 15929 3203 15932
rect 3145 15923 3203 15929
rect 3510 15920 3516 15932
rect 3568 15920 3574 15972
rect 3694 15960 3700 15972
rect 3655 15932 3700 15960
rect 3694 15920 3700 15932
rect 3752 15920 3758 15972
rect 4798 15920 4804 15972
rect 4856 15960 4862 15972
rect 4856 15932 5764 15960
rect 4856 15920 4862 15932
rect 1688 15892 1716 15920
rect 5736 15904 5764 15932
rect 6178 15920 6184 15972
rect 6236 15960 6242 15972
rect 6273 15963 6331 15969
rect 6273 15960 6285 15963
rect 6236 15932 6285 15960
rect 6236 15920 6242 15932
rect 6273 15929 6285 15932
rect 6319 15960 6331 15963
rect 7098 15960 7104 15972
rect 6319 15932 7104 15960
rect 6319 15929 6331 15932
rect 6273 15923 6331 15929
rect 7098 15920 7104 15932
rect 7156 15920 7162 15972
rect 7466 15960 7472 15972
rect 7427 15932 7472 15960
rect 7466 15920 7472 15932
rect 7524 15960 7530 15972
rect 7974 15963 8032 15969
rect 7974 15960 7986 15963
rect 7524 15932 7986 15960
rect 7524 15920 7530 15932
rect 7974 15929 7986 15932
rect 8020 15929 8032 15963
rect 7974 15923 8032 15929
rect 10873 15963 10931 15969
rect 10873 15929 10885 15963
rect 10919 15960 10931 15963
rect 10965 15963 11023 15969
rect 10965 15960 10977 15963
rect 10919 15932 10977 15960
rect 10919 15929 10931 15932
rect 10873 15923 10931 15929
rect 10965 15929 10977 15932
rect 11011 15929 11023 15963
rect 11514 15960 11520 15972
rect 11475 15932 11520 15960
rect 10965 15923 11023 15929
rect 2409 15895 2467 15901
rect 2409 15892 2421 15895
rect 1688 15864 2421 15892
rect 2409 15861 2421 15864
rect 2455 15861 2467 15895
rect 2409 15855 2467 15861
rect 4433 15895 4491 15901
rect 4433 15861 4445 15895
rect 4479 15892 4491 15895
rect 5258 15892 5264 15904
rect 4479 15864 5264 15892
rect 4479 15861 4491 15864
rect 4433 15855 4491 15861
rect 5258 15852 5264 15864
rect 5316 15852 5322 15904
rect 5718 15892 5724 15904
rect 5679 15864 5724 15892
rect 5718 15852 5724 15864
rect 5776 15852 5782 15904
rect 5902 15852 5908 15904
rect 5960 15892 5966 15904
rect 9122 15892 9128 15904
rect 5960 15864 9128 15892
rect 5960 15852 5966 15864
rect 9122 15852 9128 15864
rect 9180 15852 9186 15904
rect 10980 15892 11008 15923
rect 11514 15920 11520 15932
rect 11572 15920 11578 15972
rect 13538 15960 13544 15972
rect 11624 15932 13544 15960
rect 11624 15892 11652 15932
rect 13538 15920 13544 15932
rect 13596 15960 13602 15972
rect 15120 15960 15148 16068
rect 16758 16028 16764 16040
rect 16671 16000 16764 16028
rect 16758 15988 16764 16000
rect 16816 16028 16822 16040
rect 18064 16037 18092 16068
rect 17037 16031 17095 16037
rect 17037 16028 17049 16031
rect 16816 16000 17049 16028
rect 16816 15988 16822 16000
rect 17037 15997 17049 16000
rect 17083 15997 17095 16031
rect 17037 15991 17095 15997
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 16028 18107 16031
rect 18877 16031 18935 16037
rect 18877 16028 18889 16031
rect 18095 16000 18889 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 18877 15997 18889 16000
rect 18923 15997 18935 16031
rect 18877 15991 18935 15997
rect 13596 15932 15148 15960
rect 15289 15963 15347 15969
rect 13596 15920 13602 15932
rect 15289 15929 15301 15963
rect 15335 15929 15347 15963
rect 15289 15923 15347 15929
rect 10980 15864 11652 15892
rect 11698 15852 11704 15904
rect 11756 15892 11762 15904
rect 12161 15895 12219 15901
rect 12161 15892 12173 15895
rect 11756 15864 12173 15892
rect 11756 15852 11762 15864
rect 12161 15861 12173 15864
rect 12207 15861 12219 15895
rect 15304 15892 15332 15923
rect 15378 15920 15384 15972
rect 15436 15960 15442 15972
rect 15436 15932 15481 15960
rect 15436 15920 15442 15932
rect 15562 15892 15568 15904
rect 15304 15864 15568 15892
rect 12161 15855 12219 15861
rect 15562 15852 15568 15864
rect 15620 15892 15626 15904
rect 16209 15895 16267 15901
rect 16209 15892 16221 15895
rect 15620 15864 16221 15892
rect 15620 15852 15626 15864
rect 16209 15861 16221 15864
rect 16255 15861 16267 15895
rect 16574 15892 16580 15904
rect 16535 15864 16580 15892
rect 16209 15855 16267 15861
rect 16574 15852 16580 15864
rect 16632 15852 16638 15904
rect 18230 15892 18236 15904
rect 18191 15864 18236 15892
rect 18230 15852 18236 15864
rect 18288 15852 18294 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 2038 15648 2044 15700
rect 2096 15688 2102 15700
rect 2501 15691 2559 15697
rect 2501 15688 2513 15691
rect 2096 15660 2513 15688
rect 2096 15648 2102 15660
rect 2501 15657 2513 15660
rect 2547 15657 2559 15691
rect 2501 15651 2559 15657
rect 3881 15691 3939 15697
rect 3881 15657 3893 15691
rect 3927 15688 3939 15691
rect 4338 15688 4344 15700
rect 3927 15660 4344 15688
rect 3927 15657 3939 15660
rect 3881 15651 3939 15657
rect 4338 15648 4344 15660
rect 4396 15648 4402 15700
rect 4614 15688 4620 15700
rect 4575 15660 4620 15688
rect 4614 15648 4620 15660
rect 4672 15648 4678 15700
rect 5258 15688 5264 15700
rect 5219 15660 5264 15688
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 6546 15648 6552 15700
rect 6604 15688 6610 15700
rect 6917 15691 6975 15697
rect 6917 15688 6929 15691
rect 6604 15660 6929 15688
rect 6604 15648 6610 15660
rect 6917 15657 6929 15660
rect 6963 15657 6975 15691
rect 7282 15688 7288 15700
rect 7243 15660 7288 15688
rect 6917 15651 6975 15657
rect 7282 15648 7288 15660
rect 7340 15648 7346 15700
rect 7745 15691 7803 15697
rect 7745 15657 7757 15691
rect 7791 15688 7803 15691
rect 8018 15688 8024 15700
rect 7791 15660 8024 15688
rect 7791 15657 7803 15660
rect 7745 15651 7803 15657
rect 8018 15648 8024 15660
rect 8076 15648 8082 15700
rect 9493 15691 9551 15697
rect 9493 15657 9505 15691
rect 9539 15688 9551 15691
rect 9950 15688 9956 15700
rect 9539 15660 9956 15688
rect 9539 15657 9551 15660
rect 9493 15651 9551 15657
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 11238 15648 11244 15700
rect 11296 15688 11302 15700
rect 11701 15691 11759 15697
rect 11701 15688 11713 15691
rect 11296 15660 11713 15688
rect 11296 15648 11302 15660
rect 11701 15657 11713 15660
rect 11747 15688 11759 15691
rect 13354 15688 13360 15700
rect 11747 15660 13360 15688
rect 11747 15657 11759 15660
rect 11701 15651 11759 15657
rect 13354 15648 13360 15660
rect 13412 15648 13418 15700
rect 13446 15648 13452 15700
rect 13504 15688 13510 15700
rect 13909 15691 13967 15697
rect 13909 15688 13921 15691
rect 13504 15660 13921 15688
rect 13504 15648 13510 15660
rect 13909 15657 13921 15660
rect 13955 15657 13967 15691
rect 14274 15688 14280 15700
rect 14235 15660 14280 15688
rect 13909 15651 13967 15657
rect 14274 15648 14280 15660
rect 14332 15648 14338 15700
rect 15378 15688 15384 15700
rect 15339 15660 15384 15688
rect 15378 15648 15384 15660
rect 15436 15648 15442 15700
rect 1670 15620 1676 15632
rect 1631 15592 1676 15620
rect 1670 15580 1676 15592
rect 1728 15580 1734 15632
rect 2225 15623 2283 15629
rect 2225 15589 2237 15623
rect 2271 15620 2283 15623
rect 2314 15620 2320 15632
rect 2271 15592 2320 15620
rect 2271 15589 2283 15592
rect 2225 15583 2283 15589
rect 2314 15580 2320 15592
rect 2372 15620 2378 15632
rect 3418 15620 3424 15632
rect 2372 15592 3424 15620
rect 2372 15580 2378 15592
rect 3418 15580 3424 15592
rect 3476 15580 3482 15632
rect 4246 15620 4252 15632
rect 4131 15592 4252 15620
rect 4131 15561 4159 15592
rect 4246 15580 4252 15592
rect 4304 15620 4310 15632
rect 8754 15620 8760 15632
rect 4304 15592 8760 15620
rect 4304 15580 4310 15592
rect 8754 15580 8760 15592
rect 8812 15580 8818 15632
rect 9582 15580 9588 15632
rect 9640 15620 9646 15632
rect 9861 15623 9919 15629
rect 9861 15620 9873 15623
rect 9640 15592 9873 15620
rect 9640 15580 9646 15592
rect 9861 15589 9873 15592
rect 9907 15589 9919 15623
rect 12710 15620 12716 15632
rect 12671 15592 12716 15620
rect 9861 15583 9919 15589
rect 12710 15580 12716 15592
rect 12768 15580 12774 15632
rect 18414 15620 18420 15632
rect 18375 15592 18420 15620
rect 18414 15580 18420 15592
rect 18472 15580 18478 15632
rect 4116 15555 4174 15561
rect 4116 15521 4128 15555
rect 4162 15521 4174 15555
rect 5442 15552 5448 15564
rect 5403 15524 5448 15552
rect 4116 15515 4174 15521
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 5902 15552 5908 15564
rect 5863 15524 5908 15552
rect 5902 15512 5908 15524
rect 5960 15512 5966 15564
rect 6178 15552 6184 15564
rect 6139 15524 6184 15552
rect 6178 15512 6184 15524
rect 6236 15512 6242 15564
rect 6362 15552 6368 15564
rect 6323 15524 6368 15552
rect 6362 15512 6368 15524
rect 6420 15512 6426 15564
rect 8294 15552 8300 15564
rect 8255 15524 8300 15552
rect 8294 15512 8300 15524
rect 8352 15512 8358 15564
rect 8573 15555 8631 15561
rect 8573 15521 8585 15555
rect 8619 15552 8631 15555
rect 8662 15552 8668 15564
rect 8619 15524 8668 15552
rect 8619 15521 8631 15524
rect 8573 15515 8631 15521
rect 8662 15512 8668 15524
rect 8720 15512 8726 15564
rect 11517 15555 11575 15561
rect 11517 15521 11529 15555
rect 11563 15552 11575 15555
rect 11790 15552 11796 15564
rect 11563 15524 11796 15552
rect 11563 15521 11575 15524
rect 11517 15515 11575 15521
rect 11790 15512 11796 15524
rect 11848 15512 11854 15564
rect 13998 15512 14004 15564
rect 14056 15552 14062 15564
rect 14093 15555 14151 15561
rect 14093 15552 14105 15555
rect 14056 15524 14105 15552
rect 14056 15512 14062 15524
rect 14093 15521 14105 15524
rect 14139 15521 14151 15555
rect 14093 15515 14151 15521
rect 14734 15512 14740 15564
rect 14792 15552 14798 15564
rect 15289 15555 15347 15561
rect 15289 15552 15301 15555
rect 14792 15524 15301 15552
rect 14792 15512 14798 15524
rect 15289 15521 15301 15524
rect 15335 15521 15347 15555
rect 15838 15552 15844 15564
rect 15799 15524 15844 15552
rect 15289 15515 15347 15521
rect 15838 15512 15844 15524
rect 15896 15512 15902 15564
rect 16850 15552 16856 15564
rect 16811 15524 16856 15552
rect 16850 15512 16856 15524
rect 16908 15512 16914 15564
rect 18138 15512 18144 15564
rect 18196 15552 18202 15564
rect 18268 15555 18326 15561
rect 18268 15552 18280 15555
rect 18196 15524 18280 15552
rect 18196 15512 18202 15524
rect 18268 15521 18280 15524
rect 18314 15521 18326 15555
rect 18268 15515 18326 15521
rect 1210 15444 1216 15496
rect 1268 15484 1274 15496
rect 1581 15487 1639 15493
rect 1581 15484 1593 15487
rect 1268 15456 1593 15484
rect 1268 15444 1274 15456
rect 1581 15453 1593 15456
rect 1627 15484 1639 15487
rect 2774 15484 2780 15496
rect 1627 15456 2780 15484
rect 1627 15453 1639 15456
rect 1581 15447 1639 15453
rect 2774 15444 2780 15456
rect 2832 15444 2838 15496
rect 2958 15444 2964 15496
rect 3016 15484 3022 15496
rect 4203 15487 4261 15493
rect 4203 15484 4215 15487
rect 3016 15456 4215 15484
rect 3016 15444 3022 15456
rect 4203 15453 4215 15456
rect 4249 15453 4261 15487
rect 4203 15447 4261 15453
rect 5077 15487 5135 15493
rect 5077 15453 5089 15487
rect 5123 15484 5135 15487
rect 5166 15484 5172 15496
rect 5123 15456 5172 15484
rect 5123 15453 5135 15456
rect 5077 15447 5135 15453
rect 5166 15444 5172 15456
rect 5224 15484 5230 15496
rect 6196 15484 6224 15512
rect 5224 15456 6224 15484
rect 8757 15487 8815 15493
rect 5224 15444 5230 15456
rect 8757 15453 8769 15487
rect 8803 15484 8815 15487
rect 9398 15484 9404 15496
rect 8803 15456 9404 15484
rect 8803 15453 8815 15456
rect 8757 15447 8815 15453
rect 9398 15444 9404 15456
rect 9456 15444 9462 15496
rect 9490 15444 9496 15496
rect 9548 15484 9554 15496
rect 9769 15487 9827 15493
rect 9769 15484 9781 15487
rect 9548 15456 9781 15484
rect 9548 15444 9554 15456
rect 9769 15453 9781 15456
rect 9815 15453 9827 15487
rect 9769 15447 9827 15453
rect 10413 15487 10471 15493
rect 10413 15453 10425 15487
rect 10459 15484 10471 15487
rect 10502 15484 10508 15496
rect 10459 15456 10508 15484
rect 10459 15453 10471 15456
rect 10413 15447 10471 15453
rect 10502 15444 10508 15456
rect 10560 15444 10566 15496
rect 11974 15444 11980 15496
rect 12032 15484 12038 15496
rect 12621 15487 12679 15493
rect 12621 15484 12633 15487
rect 12032 15456 12633 15484
rect 12032 15444 12038 15456
rect 12621 15453 12633 15456
rect 12667 15484 12679 15487
rect 12986 15484 12992 15496
rect 12667 15456 12992 15484
rect 12667 15453 12679 15456
rect 12621 15447 12679 15453
rect 12986 15444 12992 15456
rect 13044 15444 13050 15496
rect 13265 15487 13323 15493
rect 13265 15453 13277 15487
rect 13311 15484 13323 15487
rect 13906 15484 13912 15496
rect 13311 15456 13912 15484
rect 13311 15453 13323 15456
rect 13265 15447 13323 15453
rect 13906 15444 13912 15456
rect 13964 15444 13970 15496
rect 16991 15487 17049 15493
rect 16991 15453 17003 15487
rect 17037 15484 17049 15487
rect 17218 15484 17224 15496
rect 17037 15456 17224 15484
rect 17037 15453 17049 15456
rect 16991 15447 17049 15453
rect 17218 15444 17224 15456
rect 17276 15444 17282 15496
rect 6086 15376 6092 15428
rect 6144 15416 6150 15428
rect 10778 15416 10784 15428
rect 6144 15388 10784 15416
rect 6144 15376 6150 15388
rect 10778 15376 10784 15388
rect 10836 15376 10842 15428
rect 12250 15376 12256 15428
rect 12308 15416 12314 15428
rect 12308 15388 13854 15416
rect 12308 15376 12314 15388
rect 3050 15348 3056 15360
rect 3011 15320 3056 15348
rect 3050 15308 3056 15320
rect 3108 15308 3114 15360
rect 3510 15348 3516 15360
rect 3471 15320 3516 15348
rect 3510 15308 3516 15320
rect 3568 15348 3574 15360
rect 4522 15348 4528 15360
rect 3568 15320 4528 15348
rect 3568 15308 3574 15320
rect 4522 15308 4528 15320
rect 4580 15308 4586 15360
rect 12069 15351 12127 15357
rect 12069 15317 12081 15351
rect 12115 15348 12127 15351
rect 12342 15348 12348 15360
rect 12115 15320 12348 15348
rect 12115 15317 12127 15320
rect 12069 15311 12127 15317
rect 12342 15308 12348 15320
rect 12400 15308 12406 15360
rect 13630 15348 13636 15360
rect 13591 15320 13636 15348
rect 13630 15308 13636 15320
rect 13688 15308 13694 15360
rect 13826 15348 13854 15388
rect 17218 15348 17224 15360
rect 13826 15320 17224 15348
rect 17218 15308 17224 15320
rect 17276 15308 17282 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 2682 15104 2688 15156
rect 2740 15144 2746 15156
rect 2869 15147 2927 15153
rect 2869 15144 2881 15147
rect 2740 15116 2881 15144
rect 2740 15104 2746 15116
rect 2869 15113 2881 15116
rect 2915 15113 2927 15147
rect 2869 15107 2927 15113
rect 4522 15104 4528 15156
rect 4580 15144 4586 15156
rect 5721 15147 5779 15153
rect 5721 15144 5733 15147
rect 4580 15116 5733 15144
rect 4580 15104 4586 15116
rect 5721 15113 5733 15116
rect 5767 15113 5779 15147
rect 5721 15107 5779 15113
rect 8662 15104 8668 15156
rect 8720 15144 8726 15156
rect 8941 15147 8999 15153
rect 8941 15144 8953 15147
rect 8720 15116 8953 15144
rect 8720 15104 8726 15116
rect 8941 15113 8953 15116
rect 8987 15144 8999 15147
rect 9030 15144 9036 15156
rect 8987 15116 9036 15144
rect 8987 15113 8999 15116
rect 8941 15107 8999 15113
rect 9030 15104 9036 15116
rect 9088 15104 9094 15156
rect 9490 15104 9496 15156
rect 9548 15144 9554 15156
rect 11149 15147 11207 15153
rect 11149 15144 11161 15147
rect 9548 15116 11161 15144
rect 9548 15104 9554 15116
rect 11149 15113 11161 15116
rect 11195 15113 11207 15147
rect 11149 15107 11207 15113
rect 11790 15104 11796 15156
rect 11848 15144 11854 15156
rect 12161 15147 12219 15153
rect 12161 15144 12173 15147
rect 11848 15116 12173 15144
rect 11848 15104 11854 15116
rect 12161 15113 12173 15116
rect 12207 15113 12219 15147
rect 12161 15107 12219 15113
rect 12710 15104 12716 15156
rect 12768 15144 12774 15156
rect 13265 15147 13323 15153
rect 13265 15144 13277 15147
rect 12768 15116 13277 15144
rect 12768 15104 12774 15116
rect 13265 15113 13277 15116
rect 13311 15144 13323 15147
rect 13354 15144 13360 15156
rect 13311 15116 13360 15144
rect 13311 15113 13323 15116
rect 13265 15107 13323 15113
rect 13354 15104 13360 15116
rect 13412 15104 13418 15156
rect 13998 15104 14004 15156
rect 14056 15144 14062 15156
rect 14553 15147 14611 15153
rect 14553 15144 14565 15147
rect 14056 15116 14565 15144
rect 14056 15104 14062 15116
rect 14553 15113 14565 15116
rect 14599 15113 14611 15147
rect 14553 15107 14611 15113
rect 14734 15104 14740 15156
rect 14792 15144 14798 15156
rect 16117 15147 16175 15153
rect 16117 15144 16129 15147
rect 14792 15116 16129 15144
rect 14792 15104 14798 15116
rect 16117 15113 16129 15116
rect 16163 15144 16175 15147
rect 17310 15144 17316 15156
rect 16163 15116 17316 15144
rect 16163 15113 16175 15116
rect 16117 15107 16175 15113
rect 17310 15104 17316 15116
rect 17368 15104 17374 15156
rect 18138 15104 18144 15156
rect 18196 15144 18202 15156
rect 18233 15147 18291 15153
rect 18233 15144 18245 15147
rect 18196 15116 18245 15144
rect 18196 15104 18202 15116
rect 18233 15113 18245 15116
rect 18279 15113 18291 15147
rect 18233 15107 18291 15113
rect 2133 15079 2191 15085
rect 2133 15045 2145 15079
rect 2179 15076 2191 15079
rect 2314 15076 2320 15088
rect 2179 15048 2320 15076
rect 2179 15045 2191 15048
rect 2133 15039 2191 15045
rect 2314 15036 2320 15048
rect 2372 15036 2378 15088
rect 4246 15076 4252 15088
rect 4207 15048 4252 15076
rect 4246 15036 4252 15048
rect 4304 15036 4310 15088
rect 5442 15036 5448 15088
rect 5500 15076 5506 15088
rect 5997 15079 6055 15085
rect 5997 15076 6009 15079
rect 5500 15048 6009 15076
rect 5500 15036 5506 15048
rect 5997 15045 6009 15048
rect 6043 15045 6055 15079
rect 5997 15039 6055 15045
rect 12342 15036 12348 15088
rect 12400 15076 12406 15088
rect 15013 15079 15071 15085
rect 15013 15076 15025 15079
rect 12400 15048 15025 15076
rect 12400 15036 12406 15048
rect 15013 15045 15025 15048
rect 15059 15076 15071 15079
rect 15838 15076 15844 15088
rect 15059 15048 15844 15076
rect 15059 15045 15071 15048
rect 15013 15039 15071 15045
rect 15838 15036 15844 15048
rect 15896 15036 15902 15088
rect 1578 15008 1584 15020
rect 1491 14980 1584 15008
rect 1578 14968 1584 14980
rect 1636 15008 1642 15020
rect 2501 15011 2559 15017
rect 2501 15008 2513 15011
rect 1636 14980 2513 15008
rect 1636 14968 1642 14980
rect 2501 14977 2513 14980
rect 2547 14977 2559 15011
rect 3050 15008 3056 15020
rect 3011 14980 3056 15008
rect 2501 14971 2559 14977
rect 3050 14968 3056 14980
rect 3108 15008 3114 15020
rect 4706 15008 4712 15020
rect 3108 14980 4712 15008
rect 3108 14968 3114 14980
rect 4706 14968 4712 14980
rect 4764 14968 4770 15020
rect 4801 15011 4859 15017
rect 4801 14977 4813 15011
rect 4847 15008 4859 15011
rect 5258 15008 5264 15020
rect 4847 14980 5264 15008
rect 4847 14977 4859 14980
rect 4801 14971 4859 14977
rect 5258 14968 5264 14980
rect 5316 14968 5322 15020
rect 6730 14968 6736 15020
rect 6788 15008 6794 15020
rect 9861 15011 9919 15017
rect 6788 14980 7696 15008
rect 6788 14968 6794 14980
rect 3973 14943 4031 14949
rect 3973 14940 3985 14943
rect 2332 14912 3985 14940
rect 1673 14875 1731 14881
rect 1673 14841 1685 14875
rect 1719 14872 1731 14875
rect 2038 14872 2044 14884
rect 1719 14844 2044 14872
rect 1719 14841 1731 14844
rect 1673 14835 1731 14841
rect 2038 14832 2044 14844
rect 2096 14872 2102 14884
rect 2332 14872 2360 14912
rect 3973 14909 3985 14912
rect 4019 14909 4031 14943
rect 7098 14940 7104 14952
rect 7059 14912 7104 14940
rect 3973 14903 4031 14909
rect 7098 14900 7104 14912
rect 7156 14900 7162 14952
rect 7282 14940 7288 14952
rect 7243 14912 7288 14940
rect 7282 14900 7288 14912
rect 7340 14900 7346 14952
rect 7668 14949 7696 14980
rect 9861 14977 9873 15011
rect 9907 15008 9919 15011
rect 9950 15008 9956 15020
rect 9907 14980 9956 15008
rect 9907 14977 9919 14980
rect 9861 14971 9919 14977
rect 9950 14968 9956 14980
rect 10008 14968 10014 15020
rect 11793 15011 11851 15017
rect 11793 15008 11805 15011
rect 11348 14980 11805 15008
rect 7653 14943 7711 14949
rect 7653 14909 7665 14943
rect 7699 14909 7711 14943
rect 8110 14940 8116 14952
rect 8071 14912 8116 14940
rect 7653 14903 7711 14909
rect 8110 14900 8116 14912
rect 8168 14900 8174 14952
rect 10686 14900 10692 14952
rect 10744 14940 10750 14952
rect 11348 14949 11376 14980
rect 11793 14977 11805 14980
rect 11839 14977 11851 15011
rect 11793 14971 11851 14977
rect 13633 15011 13691 15017
rect 13633 14977 13645 15011
rect 13679 15008 13691 15011
rect 13722 15008 13728 15020
rect 13679 14980 13728 15008
rect 13679 14977 13691 14980
rect 13633 14971 13691 14977
rect 13722 14968 13728 14980
rect 13780 14968 13786 15020
rect 13906 14968 13912 15020
rect 13964 15008 13970 15020
rect 14277 15011 14335 15017
rect 14277 15008 14289 15011
rect 13964 14980 14289 15008
rect 13964 14968 13970 14980
rect 14277 14977 14289 14980
rect 14323 15008 14335 15011
rect 15197 15011 15255 15017
rect 15197 15008 15209 15011
rect 14323 14980 15209 15008
rect 14323 14977 14335 14980
rect 14277 14971 14335 14977
rect 15197 14977 15209 14980
rect 15243 15008 15255 15011
rect 16945 15011 17003 15017
rect 16945 15008 16957 15011
rect 15243 14980 16957 15008
rect 15243 14977 15255 14980
rect 15197 14971 15255 14977
rect 16945 14977 16957 14980
rect 16991 14977 17003 15011
rect 16945 14971 17003 14977
rect 11333 14943 11391 14949
rect 11333 14940 11345 14943
rect 10744 14912 11345 14940
rect 10744 14900 10750 14912
rect 11333 14909 11345 14912
rect 11379 14909 11391 14943
rect 11333 14903 11391 14909
rect 11514 14900 11520 14952
rect 11572 14940 11578 14952
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 11572 14912 12449 14940
rect 11572 14900 11578 14912
rect 12437 14909 12449 14912
rect 12483 14940 12495 14943
rect 12897 14943 12955 14949
rect 12897 14940 12909 14943
rect 12483 14912 12909 14940
rect 12483 14909 12495 14912
rect 12437 14903 12495 14909
rect 12897 14909 12909 14912
rect 12943 14909 12955 14943
rect 12897 14903 12955 14909
rect 15841 14943 15899 14949
rect 15841 14909 15853 14943
rect 15887 14940 15899 14943
rect 16022 14940 16028 14952
rect 15887 14912 16028 14940
rect 15887 14909 15899 14912
rect 15841 14903 15899 14909
rect 16022 14900 16028 14912
rect 16080 14940 16086 14952
rect 16850 14940 16856 14952
rect 16080 14912 16856 14940
rect 16080 14900 16086 14912
rect 16850 14900 16856 14912
rect 16908 14940 16914 14952
rect 17221 14943 17279 14949
rect 17221 14940 17233 14943
rect 16908 14912 17233 14940
rect 16908 14900 16914 14912
rect 17221 14909 17233 14912
rect 17267 14909 17279 14943
rect 17221 14903 17279 14909
rect 2096 14844 2360 14872
rect 2096 14832 2102 14844
rect 2682 14832 2688 14884
rect 2740 14872 2746 14884
rect 3374 14875 3432 14881
rect 3374 14872 3386 14875
rect 2740 14844 3386 14872
rect 2740 14832 2746 14844
rect 3374 14841 3386 14844
rect 3420 14872 3432 14875
rect 3602 14872 3608 14884
rect 3420 14844 3608 14872
rect 3420 14841 3432 14844
rect 3374 14835 3432 14841
rect 3602 14832 3608 14844
rect 3660 14872 3666 14884
rect 4617 14875 4675 14881
rect 4617 14872 4629 14875
rect 3660 14844 4629 14872
rect 3660 14832 3666 14844
rect 4617 14841 4629 14844
rect 4663 14872 4675 14875
rect 5122 14875 5180 14881
rect 5122 14872 5134 14875
rect 4663 14844 5134 14872
rect 4663 14841 4675 14844
rect 4617 14835 4675 14841
rect 5122 14841 5134 14844
rect 5168 14872 5180 14875
rect 7466 14872 7472 14884
rect 5168 14844 7472 14872
rect 5168 14841 5180 14844
rect 5122 14835 5180 14841
rect 7466 14832 7472 14844
rect 7524 14832 7530 14884
rect 9953 14875 10011 14881
rect 9953 14841 9965 14875
rect 9999 14841 10011 14875
rect 10502 14872 10508 14884
rect 10415 14844 10508 14872
rect 9953 14835 10011 14841
rect 6641 14807 6699 14813
rect 6641 14773 6653 14807
rect 6687 14804 6699 14807
rect 6730 14804 6736 14816
rect 6687 14776 6736 14804
rect 6687 14773 6699 14776
rect 6641 14767 6699 14773
rect 6730 14764 6736 14776
rect 6788 14764 6794 14816
rect 7098 14804 7104 14816
rect 7059 14776 7104 14804
rect 7098 14764 7104 14776
rect 7156 14764 7162 14816
rect 8294 14764 8300 14816
rect 8352 14804 8358 14816
rect 8573 14807 8631 14813
rect 8573 14804 8585 14807
rect 8352 14776 8585 14804
rect 8352 14764 8358 14776
rect 8573 14773 8585 14776
rect 8619 14773 8631 14807
rect 9582 14804 9588 14816
rect 9543 14776 9588 14804
rect 8573 14767 8631 14773
rect 9582 14764 9588 14776
rect 9640 14764 9646 14816
rect 9674 14764 9680 14816
rect 9732 14804 9738 14816
rect 9968 14804 9996 14835
rect 10502 14832 10508 14844
rect 10560 14872 10566 14884
rect 11974 14872 11980 14884
rect 10560 14844 11980 14872
rect 10560 14832 10566 14844
rect 11974 14832 11980 14844
rect 12032 14832 12038 14884
rect 13630 14832 13636 14884
rect 13688 14872 13694 14884
rect 13734 14875 13792 14881
rect 13734 14872 13746 14875
rect 13688 14844 13746 14872
rect 13688 14832 13694 14844
rect 13734 14841 13746 14844
rect 13780 14872 13792 14875
rect 14826 14872 14832 14884
rect 13780 14844 14832 14872
rect 13780 14841 13792 14844
rect 13734 14835 13792 14841
rect 14826 14832 14832 14844
rect 14884 14832 14890 14884
rect 15289 14875 15347 14881
rect 15289 14841 15301 14875
rect 15335 14841 15347 14875
rect 15289 14835 15347 14841
rect 15948 14844 16252 14872
rect 10781 14807 10839 14813
rect 10781 14804 10793 14807
rect 9732 14776 10793 14804
rect 9732 14764 9738 14776
rect 10781 14773 10793 14776
rect 10827 14773 10839 14807
rect 11514 14804 11520 14816
rect 11475 14776 11520 14804
rect 10781 14767 10839 14773
rect 11514 14764 11520 14776
rect 11572 14764 11578 14816
rect 12342 14764 12348 14816
rect 12400 14804 12406 14816
rect 12621 14807 12679 14813
rect 12621 14804 12633 14807
rect 12400 14776 12633 14804
rect 12400 14764 12406 14776
rect 12621 14773 12633 14776
rect 12667 14773 12679 14807
rect 15304 14804 15332 14835
rect 15948 14804 15976 14844
rect 16224 14816 16252 14844
rect 15304 14776 15976 14804
rect 12621 14767 12679 14773
rect 16206 14764 16212 14816
rect 16264 14804 16270 14816
rect 16485 14807 16543 14813
rect 16485 14804 16497 14807
rect 16264 14776 16497 14804
rect 16264 14764 16270 14776
rect 16485 14773 16497 14776
rect 16531 14773 16543 14807
rect 16485 14767 16543 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1670 14600 1676 14612
rect 1631 14572 1676 14600
rect 1670 14560 1676 14572
rect 1728 14560 1734 14612
rect 2038 14600 2044 14612
rect 1999 14572 2044 14600
rect 2038 14560 2044 14572
rect 2096 14560 2102 14612
rect 2774 14560 2780 14612
rect 2832 14600 2838 14612
rect 3145 14603 3203 14609
rect 3145 14600 3157 14603
rect 2832 14572 3157 14600
rect 2832 14560 2838 14572
rect 3145 14569 3157 14572
rect 3191 14569 3203 14603
rect 3145 14563 3203 14569
rect 4706 14560 4712 14612
rect 4764 14600 4770 14612
rect 5261 14603 5319 14609
rect 5261 14600 5273 14603
rect 4764 14572 5273 14600
rect 4764 14560 4770 14572
rect 5261 14569 5273 14572
rect 5307 14569 5319 14603
rect 5261 14563 5319 14569
rect 6362 14560 6368 14612
rect 6420 14600 6426 14612
rect 6822 14600 6828 14612
rect 6420 14572 6828 14600
rect 6420 14560 6426 14572
rect 6822 14560 6828 14572
rect 6880 14600 6886 14612
rect 6917 14603 6975 14609
rect 6917 14600 6929 14603
rect 6880 14572 6929 14600
rect 6880 14560 6886 14572
rect 6917 14569 6929 14572
rect 6963 14569 6975 14603
rect 6917 14563 6975 14569
rect 7006 14560 7012 14612
rect 7064 14600 7070 14612
rect 7285 14603 7343 14609
rect 7285 14600 7297 14603
rect 7064 14572 7297 14600
rect 7064 14560 7070 14572
rect 7285 14569 7297 14572
rect 7331 14569 7343 14603
rect 9033 14603 9091 14609
rect 9033 14600 9045 14603
rect 7285 14563 7343 14569
rect 8128 14572 9045 14600
rect 2222 14532 2228 14544
rect 2183 14504 2228 14532
rect 2222 14492 2228 14504
rect 2280 14492 2286 14544
rect 2317 14535 2375 14541
rect 2317 14501 2329 14535
rect 2363 14532 2375 14535
rect 2498 14532 2504 14544
rect 2363 14504 2504 14532
rect 2363 14501 2375 14504
rect 2317 14495 2375 14501
rect 2498 14492 2504 14504
rect 2556 14492 2562 14544
rect 2869 14535 2927 14541
rect 2869 14501 2881 14535
rect 2915 14532 2927 14535
rect 3234 14532 3240 14544
rect 2915 14504 3240 14532
rect 2915 14501 2927 14504
rect 2869 14495 2927 14501
rect 3234 14492 3240 14504
rect 3292 14532 3298 14544
rect 3694 14532 3700 14544
rect 3292 14504 3700 14532
rect 3292 14492 3298 14504
rect 3694 14492 3700 14504
rect 3752 14492 3758 14544
rect 4617 14535 4675 14541
rect 4617 14501 4629 14535
rect 4663 14532 4675 14535
rect 5077 14535 5135 14541
rect 5077 14532 5089 14535
rect 4663 14504 5089 14532
rect 4663 14501 4675 14504
rect 4617 14495 4675 14501
rect 5077 14501 5089 14504
rect 5123 14532 5135 14535
rect 5166 14532 5172 14544
rect 5123 14504 5172 14532
rect 5123 14501 5135 14504
rect 5077 14495 5135 14501
rect 5166 14492 5172 14504
rect 5224 14532 5230 14544
rect 5224 14504 5948 14532
rect 5224 14492 5230 14504
rect 4157 14467 4215 14473
rect 4157 14433 4169 14467
rect 4203 14464 4215 14467
rect 4246 14464 4252 14476
rect 4203 14436 4252 14464
rect 4203 14433 4215 14436
rect 4157 14427 4215 14433
rect 4246 14424 4252 14436
rect 4304 14424 4310 14476
rect 5442 14464 5448 14476
rect 5403 14436 5448 14464
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 5920 14473 5948 14504
rect 7926 14492 7932 14544
rect 7984 14532 7990 14544
rect 8128 14541 8156 14572
rect 9033 14569 9045 14572
rect 9079 14569 9091 14603
rect 9398 14600 9404 14612
rect 9359 14572 9404 14600
rect 9033 14563 9091 14569
rect 9398 14560 9404 14572
rect 9456 14560 9462 14612
rect 10781 14603 10839 14609
rect 10781 14569 10793 14603
rect 10827 14600 10839 14603
rect 11606 14600 11612 14612
rect 10827 14572 11612 14600
rect 10827 14569 10839 14572
rect 10781 14563 10839 14569
rect 11606 14560 11612 14572
rect 11664 14600 11670 14612
rect 12618 14600 12624 14612
rect 11664 14572 11836 14600
rect 12579 14572 12624 14600
rect 11664 14560 11670 14572
rect 8113 14535 8171 14541
rect 8113 14532 8125 14535
rect 7984 14504 8125 14532
rect 7984 14492 7990 14504
rect 8113 14501 8125 14504
rect 8159 14501 8171 14535
rect 8113 14495 8171 14501
rect 8205 14535 8263 14541
rect 8205 14501 8217 14535
rect 8251 14532 8263 14535
rect 8754 14532 8760 14544
rect 8251 14504 8760 14532
rect 8251 14501 8263 14504
rect 8205 14495 8263 14501
rect 8754 14492 8760 14504
rect 8812 14492 8818 14544
rect 5905 14467 5963 14473
rect 5905 14433 5917 14467
rect 5951 14464 5963 14467
rect 5994 14464 6000 14476
rect 5951 14436 6000 14464
rect 5951 14433 5963 14436
rect 5905 14427 5963 14433
rect 5994 14424 6000 14436
rect 6052 14424 6058 14476
rect 6178 14464 6184 14476
rect 6139 14436 6184 14464
rect 6178 14424 6184 14436
rect 6236 14424 6242 14476
rect 6546 14464 6552 14476
rect 6507 14436 6552 14464
rect 6546 14424 6552 14436
rect 6604 14424 6610 14476
rect 7282 14424 7288 14476
rect 7340 14464 7346 14476
rect 7653 14467 7711 14473
rect 7653 14464 7665 14467
rect 7340 14436 7665 14464
rect 7340 14424 7346 14436
rect 7653 14433 7665 14436
rect 7699 14433 7711 14467
rect 9416 14464 9444 14560
rect 10223 14535 10281 14541
rect 10223 14501 10235 14535
rect 10269 14532 10281 14535
rect 10410 14532 10416 14544
rect 10269 14504 10416 14532
rect 10269 14501 10281 14504
rect 10223 14495 10281 14501
rect 10410 14492 10416 14504
rect 10468 14532 10474 14544
rect 11330 14532 11336 14544
rect 10468 14504 11336 14532
rect 10468 14492 10474 14504
rect 11330 14492 11336 14504
rect 11388 14492 11394 14544
rect 11808 14541 11836 14572
rect 12618 14560 12624 14572
rect 12676 14560 12682 14612
rect 12986 14600 12992 14612
rect 12947 14572 12992 14600
rect 12986 14560 12992 14572
rect 13044 14560 13050 14612
rect 13170 14560 13176 14612
rect 13228 14600 13234 14612
rect 13228 14572 13308 14600
rect 13228 14560 13234 14572
rect 13280 14541 13308 14572
rect 13722 14560 13728 14612
rect 13780 14600 13786 14612
rect 14550 14600 14556 14612
rect 13780 14572 14556 14600
rect 13780 14560 13786 14572
rect 14550 14560 14556 14572
rect 14608 14560 14614 14612
rect 16206 14600 16212 14612
rect 16167 14572 16212 14600
rect 16206 14560 16212 14572
rect 16264 14560 16270 14612
rect 19518 14560 19524 14612
rect 19576 14600 19582 14612
rect 20254 14600 20260 14612
rect 19576 14572 20260 14600
rect 19576 14560 19582 14572
rect 20254 14560 20260 14572
rect 20312 14560 20318 14612
rect 11793 14535 11851 14541
rect 11793 14501 11805 14535
rect 11839 14501 11851 14535
rect 11793 14495 11851 14501
rect 13265 14535 13323 14541
rect 13265 14501 13277 14535
rect 13311 14501 13323 14535
rect 13265 14495 13323 14501
rect 13357 14535 13415 14541
rect 13357 14501 13369 14535
rect 13403 14532 13415 14535
rect 13630 14532 13636 14544
rect 13403 14504 13636 14532
rect 13403 14501 13415 14504
rect 13357 14495 13415 14501
rect 13630 14492 13636 14504
rect 13688 14492 13694 14544
rect 13906 14532 13912 14544
rect 13867 14504 13912 14532
rect 13906 14492 13912 14504
rect 13964 14492 13970 14544
rect 15470 14492 15476 14544
rect 15528 14532 15534 14544
rect 15610 14535 15668 14541
rect 15610 14532 15622 14535
rect 15528 14504 15622 14532
rect 15528 14492 15534 14504
rect 15610 14501 15622 14504
rect 15656 14501 15668 14535
rect 15610 14495 15668 14501
rect 9861 14467 9919 14473
rect 9861 14464 9873 14467
rect 9416 14436 9873 14464
rect 7653 14427 7711 14433
rect 9861 14433 9873 14436
rect 9907 14433 9919 14467
rect 9861 14427 9919 14433
rect 15289 14467 15347 14473
rect 15289 14433 15301 14467
rect 15335 14464 15347 14467
rect 15378 14464 15384 14476
rect 15335 14436 15384 14464
rect 15335 14433 15347 14436
rect 15289 14427 15347 14433
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 3786 14356 3792 14408
rect 3844 14396 3850 14408
rect 3881 14399 3939 14405
rect 3881 14396 3893 14399
rect 3844 14368 3893 14396
rect 3844 14356 3850 14368
rect 3881 14365 3893 14368
rect 3927 14396 3939 14399
rect 6564 14396 6592 14424
rect 3927 14368 6592 14396
rect 8757 14399 8815 14405
rect 3927 14365 3939 14368
rect 3881 14359 3939 14365
rect 8757 14365 8769 14399
rect 8803 14396 8815 14399
rect 11701 14399 11759 14405
rect 11701 14396 11713 14399
rect 8803 14368 11713 14396
rect 8803 14365 8815 14368
rect 8757 14359 8815 14365
rect 11701 14365 11713 14368
rect 11747 14365 11759 14399
rect 11701 14359 11759 14365
rect 4341 14331 4399 14337
rect 4341 14297 4353 14331
rect 4387 14328 4399 14331
rect 6546 14328 6552 14340
rect 4387 14300 6552 14328
rect 4387 14297 4399 14300
rect 4341 14291 4399 14297
rect 6546 14288 6552 14300
rect 6604 14288 6610 14340
rect 11716 14328 11744 14359
rect 11790 14356 11796 14408
rect 11848 14396 11854 14408
rect 12345 14399 12403 14405
rect 12345 14396 12357 14399
rect 11848 14368 12357 14396
rect 11848 14356 11854 14368
rect 12345 14365 12357 14368
rect 12391 14396 12403 14399
rect 18138 14396 18144 14408
rect 12391 14368 18144 14396
rect 12391 14365 12403 14368
rect 12345 14359 12403 14365
rect 18138 14356 18144 14368
rect 18196 14356 18202 14408
rect 11974 14328 11980 14340
rect 11716 14300 11980 14328
rect 11974 14288 11980 14300
rect 12032 14288 12038 14340
rect 14274 14260 14280 14272
rect 14235 14232 14280 14260
rect 14274 14220 14280 14232
rect 14332 14220 14338 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 3142 14016 3148 14068
rect 3200 14056 3206 14068
rect 3237 14059 3295 14065
rect 3237 14056 3249 14059
rect 3200 14028 3249 14056
rect 3200 14016 3206 14028
rect 3237 14025 3249 14028
rect 3283 14025 3295 14059
rect 3237 14019 3295 14025
rect 3881 14059 3939 14065
rect 3881 14025 3893 14059
rect 3927 14056 3939 14059
rect 5442 14056 5448 14068
rect 3927 14028 5448 14056
rect 3927 14025 3939 14028
rect 3881 14019 3939 14025
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13920 1639 13923
rect 1946 13920 1952 13932
rect 1627 13892 1952 13920
rect 1627 13889 1639 13892
rect 1581 13883 1639 13889
rect 1946 13880 1952 13892
rect 2004 13880 2010 13932
rect 2222 13920 2228 13932
rect 2183 13892 2228 13920
rect 2222 13880 2228 13892
rect 2280 13920 2286 13932
rect 2869 13923 2927 13929
rect 2869 13920 2881 13923
rect 2280 13892 2881 13920
rect 2280 13880 2286 13892
rect 2869 13889 2881 13892
rect 2915 13889 2927 13923
rect 2869 13883 2927 13889
rect 3050 13852 3056 13864
rect 3011 13824 3056 13852
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 4632 13861 4660 14028
rect 5442 14016 5448 14028
rect 5500 14056 5506 14068
rect 6181 14059 6239 14065
rect 6181 14056 6193 14059
rect 5500 14028 6193 14056
rect 5500 14016 5506 14028
rect 6181 14025 6193 14028
rect 6227 14025 6239 14059
rect 6181 14019 6239 14025
rect 6641 14059 6699 14065
rect 6641 14025 6653 14059
rect 6687 14056 6699 14059
rect 6730 14056 6736 14068
rect 6687 14028 6736 14056
rect 6687 14025 6699 14028
rect 6641 14019 6699 14025
rect 6730 14016 6736 14028
rect 6788 14016 6794 14068
rect 9950 14016 9956 14068
rect 10008 14056 10014 14068
rect 10410 14056 10416 14068
rect 10008 14028 10416 14056
rect 10008 14016 10014 14028
rect 10410 14016 10416 14028
rect 10468 14016 10474 14068
rect 10781 14059 10839 14065
rect 10781 14025 10793 14059
rect 10827 14056 10839 14059
rect 10962 14056 10968 14068
rect 10827 14028 10968 14056
rect 10827 14025 10839 14028
rect 10781 14019 10839 14025
rect 4982 13880 4988 13932
rect 5040 13920 5046 13932
rect 6748 13920 6776 14016
rect 9214 13948 9220 14000
rect 9272 13988 9278 14000
rect 9582 13988 9588 14000
rect 9272 13960 9588 13988
rect 9272 13948 9278 13960
rect 9582 13948 9588 13960
rect 9640 13988 9646 14000
rect 10045 13991 10103 13997
rect 10045 13988 10057 13991
rect 9640 13960 10057 13988
rect 9640 13948 9646 13960
rect 10045 13957 10057 13960
rect 10091 13957 10103 13991
rect 10045 13951 10103 13957
rect 10796 13920 10824 14019
rect 10962 14016 10968 14028
rect 11020 14016 11026 14068
rect 11793 14059 11851 14065
rect 11793 14025 11805 14059
rect 11839 14056 11851 14059
rect 11882 14056 11888 14068
rect 11839 14028 11888 14056
rect 11839 14025 11851 14028
rect 11793 14019 11851 14025
rect 11882 14016 11888 14028
rect 11940 14016 11946 14068
rect 13354 14056 13360 14068
rect 13315 14028 13360 14056
rect 13354 14016 13360 14028
rect 13412 14016 13418 14068
rect 14826 14016 14832 14068
rect 14884 14056 14890 14068
rect 15105 14059 15163 14065
rect 15105 14056 15117 14059
rect 14884 14028 15117 14056
rect 14884 14016 14890 14028
rect 15105 14025 15117 14028
rect 15151 14025 15163 14059
rect 15105 14019 15163 14025
rect 15378 14016 15384 14068
rect 15436 14056 15442 14068
rect 16945 14059 17003 14065
rect 16945 14056 16957 14059
rect 15436 14028 16957 14056
rect 15436 14016 15442 14028
rect 16945 14025 16957 14028
rect 16991 14025 17003 14059
rect 16945 14019 17003 14025
rect 11514 13948 11520 14000
rect 11572 13988 11578 14000
rect 13078 13988 13084 14000
rect 11572 13960 13084 13988
rect 11572 13948 11578 13960
rect 13078 13948 13084 13960
rect 13136 13948 13142 14000
rect 13446 13948 13452 14000
rect 13504 13988 13510 14000
rect 15749 13991 15807 13997
rect 15749 13988 15761 13991
rect 13504 13960 15761 13988
rect 13504 13948 13510 13960
rect 15749 13957 15761 13960
rect 15795 13957 15807 13991
rect 15749 13951 15807 13957
rect 5040 13892 5304 13920
rect 6748 13892 10824 13920
rect 12437 13923 12495 13929
rect 5040 13880 5046 13892
rect 4617 13855 4675 13861
rect 4617 13821 4629 13855
rect 4663 13821 4675 13855
rect 5166 13852 5172 13864
rect 5127 13824 5172 13852
rect 4617 13815 4675 13821
rect 5166 13812 5172 13824
rect 5224 13812 5230 13864
rect 5276 13861 5304 13892
rect 5261 13855 5319 13861
rect 5261 13821 5273 13855
rect 5307 13852 5319 13855
rect 5534 13852 5540 13864
rect 5307 13824 5540 13852
rect 5307 13821 5319 13824
rect 5261 13815 5319 13821
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 5813 13855 5871 13861
rect 5813 13821 5825 13855
rect 5859 13852 5871 13855
rect 6454 13852 6460 13864
rect 5859 13824 6460 13852
rect 5859 13821 5871 13824
rect 5813 13815 5871 13821
rect 6454 13812 6460 13824
rect 6512 13812 6518 13864
rect 7006 13852 7012 13864
rect 6967 13824 7012 13852
rect 7006 13812 7012 13824
rect 7064 13812 7070 13864
rect 7282 13852 7288 13864
rect 7243 13824 7288 13852
rect 7282 13812 7288 13824
rect 7340 13812 7346 13864
rect 7668 13861 7696 13892
rect 12437 13889 12449 13923
rect 12483 13920 12495 13923
rect 12618 13920 12624 13932
rect 12483 13892 12624 13920
rect 12483 13889 12495 13892
rect 12437 13883 12495 13889
rect 12618 13880 12624 13892
rect 12676 13880 12682 13932
rect 14093 13923 14151 13929
rect 14093 13920 14105 13923
rect 14003 13892 14105 13920
rect 14093 13889 14105 13892
rect 14139 13920 14151 13923
rect 14458 13920 14464 13932
rect 14139 13892 14464 13920
rect 14139 13889 14151 13892
rect 14093 13883 14151 13889
rect 7653 13855 7711 13861
rect 7653 13821 7665 13855
rect 7699 13821 7711 13855
rect 7653 13815 7711 13821
rect 8021 13855 8079 13861
rect 8021 13821 8033 13855
rect 8067 13852 8079 13855
rect 9122 13852 9128 13864
rect 8067 13824 8101 13852
rect 9083 13824 9128 13852
rect 8067 13821 8079 13824
rect 8021 13815 8079 13821
rect 1670 13784 1676 13796
rect 1583 13756 1676 13784
rect 1670 13744 1676 13756
rect 1728 13784 1734 13796
rect 2038 13784 2044 13796
rect 1728 13756 2044 13784
rect 1728 13744 1734 13756
rect 2038 13744 2044 13756
rect 2096 13744 2102 13796
rect 4246 13784 4252 13796
rect 4207 13756 4252 13784
rect 4246 13744 4252 13756
rect 4304 13744 4310 13796
rect 6822 13744 6828 13796
rect 6880 13784 6886 13796
rect 8036 13784 8064 13815
rect 9122 13812 9128 13824
rect 9180 13812 9186 13864
rect 11057 13855 11115 13861
rect 11057 13821 11069 13855
rect 11103 13852 11115 13855
rect 11882 13852 11888 13864
rect 11103 13824 11888 13852
rect 11103 13821 11115 13824
rect 11057 13815 11115 13821
rect 11882 13812 11888 13824
rect 11940 13812 11946 13864
rect 14108 13852 14136 13883
rect 14458 13880 14464 13892
rect 14516 13920 14522 13932
rect 15470 13920 15476 13932
rect 14516 13892 15476 13920
rect 14516 13880 14522 13892
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 15764 13920 15792 13951
rect 15838 13948 15844 14000
rect 15896 13988 15902 14000
rect 15896 13960 16436 13988
rect 15896 13948 15902 13960
rect 15764 13892 15976 13920
rect 13464 13824 14136 13852
rect 6880 13756 8064 13784
rect 6880 13744 6886 13756
rect 9306 13744 9312 13796
rect 9364 13784 9370 13796
rect 10873 13787 10931 13793
rect 9364 13756 10456 13784
rect 9364 13744 9370 13756
rect 2498 13716 2504 13728
rect 2459 13688 2504 13716
rect 2498 13676 2504 13688
rect 2556 13676 2562 13728
rect 4522 13716 4528 13728
rect 4483 13688 4528 13716
rect 4522 13676 4528 13688
rect 4580 13676 4586 13728
rect 6914 13716 6920 13728
rect 6875 13688 6920 13716
rect 6914 13676 6920 13688
rect 6972 13676 6978 13728
rect 8665 13719 8723 13725
rect 8665 13685 8677 13719
rect 8711 13716 8723 13719
rect 8754 13716 8760 13728
rect 8711 13688 8760 13716
rect 8711 13685 8723 13688
rect 8665 13679 8723 13685
rect 8754 13676 8760 13688
rect 8812 13676 8818 13728
rect 8846 13676 8852 13728
rect 8904 13716 8910 13728
rect 8941 13719 8999 13725
rect 8941 13716 8953 13719
rect 8904 13688 8953 13716
rect 8904 13676 8910 13688
rect 8941 13685 8953 13688
rect 8987 13716 8999 13719
rect 9493 13719 9551 13725
rect 9493 13716 9505 13719
rect 8987 13688 9505 13716
rect 8987 13685 8999 13688
rect 8941 13679 8999 13685
rect 9493 13685 9505 13688
rect 9539 13685 9551 13719
rect 10428 13716 10456 13756
rect 10873 13753 10885 13787
rect 10919 13784 10931 13787
rect 10962 13784 10968 13796
rect 10919 13756 10968 13784
rect 10919 13753 10931 13756
rect 10873 13747 10931 13753
rect 10962 13744 10968 13756
rect 11020 13744 11026 13796
rect 11330 13744 11336 13796
rect 11388 13784 11394 13796
rect 12253 13787 12311 13793
rect 12253 13784 12265 13787
rect 11388 13756 12265 13784
rect 11388 13744 11394 13756
rect 12253 13753 12265 13756
rect 12299 13784 12311 13787
rect 12526 13784 12532 13796
rect 12299 13756 12532 13784
rect 12299 13753 12311 13756
rect 12253 13747 12311 13753
rect 12526 13744 12532 13756
rect 12584 13784 12590 13796
rect 12799 13787 12857 13793
rect 12799 13784 12811 13787
rect 12584 13756 12811 13784
rect 12584 13744 12590 13756
rect 12799 13753 12811 13756
rect 12845 13784 12857 13787
rect 13464 13784 13492 13824
rect 13630 13784 13636 13796
rect 12845 13756 13492 13784
rect 13591 13756 13636 13784
rect 12845 13753 12857 13756
rect 12799 13747 12857 13753
rect 13630 13744 13636 13756
rect 13688 13744 13694 13796
rect 14108 13784 14136 13824
rect 14185 13855 14243 13861
rect 14185 13821 14197 13855
rect 14231 13852 14243 13855
rect 14274 13852 14280 13864
rect 14231 13824 14280 13852
rect 14231 13821 14243 13824
rect 14185 13815 14243 13821
rect 14274 13812 14280 13824
rect 14332 13852 14338 13864
rect 15948 13861 15976 13892
rect 16408 13861 16436 13960
rect 15933 13855 15991 13861
rect 14332 13824 15884 13852
rect 14332 13812 14338 13824
rect 14506 13787 14564 13793
rect 14506 13784 14518 13787
rect 14108 13756 14518 13784
rect 14506 13753 14518 13756
rect 14552 13753 14564 13787
rect 14506 13747 14564 13753
rect 11149 13719 11207 13725
rect 11149 13716 11161 13719
rect 10428 13688 11161 13716
rect 9493 13679 9551 13685
rect 11149 13685 11161 13688
rect 11195 13685 11207 13719
rect 15856 13716 15884 13824
rect 15933 13821 15945 13855
rect 15979 13821 15991 13855
rect 15933 13815 15991 13821
rect 16393 13855 16451 13861
rect 16393 13821 16405 13855
rect 16439 13821 16451 13855
rect 16393 13815 16451 13821
rect 16025 13719 16083 13725
rect 16025 13716 16037 13719
rect 15856 13688 16037 13716
rect 11149 13679 11207 13685
rect 16025 13685 16037 13688
rect 16071 13685 16083 13719
rect 16025 13679 16083 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1670 13512 1676 13524
rect 1631 13484 1676 13512
rect 1670 13472 1676 13484
rect 1728 13472 1734 13524
rect 2498 13512 2504 13524
rect 2459 13484 2504 13512
rect 2498 13472 2504 13484
rect 2556 13472 2562 13524
rect 3786 13512 3792 13524
rect 3747 13484 3792 13512
rect 3786 13472 3792 13484
rect 3844 13472 3850 13524
rect 5258 13512 5264 13524
rect 5219 13484 5264 13512
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 5350 13472 5356 13524
rect 5408 13512 5414 13524
rect 6086 13512 6092 13524
rect 5408 13484 6092 13512
rect 5408 13472 5414 13484
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 6178 13472 6184 13524
rect 6236 13512 6242 13524
rect 6917 13515 6975 13521
rect 6917 13512 6929 13515
rect 6236 13484 6929 13512
rect 6236 13472 6242 13484
rect 6917 13481 6929 13484
rect 6963 13481 6975 13515
rect 6917 13475 6975 13481
rect 7282 13472 7288 13524
rect 7340 13512 7346 13524
rect 7653 13515 7711 13521
rect 7653 13512 7665 13515
rect 7340 13484 7665 13512
rect 7340 13472 7346 13484
rect 7653 13481 7665 13484
rect 7699 13481 7711 13515
rect 7926 13512 7932 13524
rect 7887 13484 7932 13512
rect 7653 13475 7711 13481
rect 7926 13472 7932 13484
rect 7984 13472 7990 13524
rect 9122 13512 9128 13524
rect 9083 13484 9128 13512
rect 9122 13472 9128 13484
rect 9180 13512 9186 13524
rect 9769 13515 9827 13521
rect 9769 13512 9781 13515
rect 9180 13484 9781 13512
rect 9180 13472 9186 13484
rect 9769 13481 9781 13484
rect 9815 13481 9827 13515
rect 11606 13512 11612 13524
rect 11567 13484 11612 13512
rect 9769 13475 9827 13481
rect 11606 13472 11612 13484
rect 11664 13472 11670 13524
rect 11974 13512 11980 13524
rect 11935 13484 11980 13512
rect 11974 13472 11980 13484
rect 12032 13472 12038 13524
rect 12526 13512 12532 13524
rect 12487 13484 12532 13512
rect 12526 13472 12532 13484
rect 12584 13472 12590 13524
rect 13262 13472 13268 13524
rect 13320 13512 13326 13524
rect 13357 13515 13415 13521
rect 13357 13512 13369 13515
rect 13320 13484 13369 13512
rect 13320 13472 13326 13484
rect 13357 13481 13369 13484
rect 13403 13481 13415 13515
rect 15378 13512 15384 13524
rect 15339 13484 15384 13512
rect 13357 13475 13415 13481
rect 15378 13472 15384 13484
rect 15436 13472 15442 13524
rect 16942 13512 16948 13524
rect 16903 13484 16948 13512
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 5074 13404 5080 13456
rect 5132 13444 5138 13456
rect 8294 13444 8300 13456
rect 5132 13416 5672 13444
rect 5132 13404 5138 13416
rect 2869 13379 2927 13385
rect 2869 13345 2881 13379
rect 2915 13376 2927 13379
rect 2958 13376 2964 13388
rect 2915 13348 2964 13376
rect 2915 13345 2927 13348
rect 2869 13339 2927 13345
rect 2958 13336 2964 13348
rect 3016 13376 3022 13388
rect 3510 13376 3516 13388
rect 3016 13348 3516 13376
rect 3016 13336 3022 13348
rect 3510 13336 3516 13348
rect 3568 13336 3574 13388
rect 3970 13336 3976 13388
rect 4028 13376 4034 13388
rect 4100 13379 4158 13385
rect 4100 13376 4112 13379
rect 4028 13348 4112 13376
rect 4028 13336 4034 13348
rect 4100 13345 4112 13348
rect 4146 13345 4158 13379
rect 5442 13376 5448 13388
rect 5403 13348 5448 13376
rect 4100 13339 4158 13345
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 5644 13385 5672 13416
rect 8128 13416 8300 13444
rect 5629 13379 5687 13385
rect 5629 13345 5641 13379
rect 5675 13345 5687 13379
rect 5629 13339 5687 13345
rect 6181 13379 6239 13385
rect 6181 13345 6193 13379
rect 6227 13345 6239 13379
rect 6181 13339 6239 13345
rect 6549 13379 6607 13385
rect 6549 13345 6561 13379
rect 6595 13376 6607 13379
rect 6822 13376 6828 13388
rect 6595 13348 6828 13376
rect 6595 13345 6607 13348
rect 6549 13339 6607 13345
rect 2130 13268 2136 13320
rect 2188 13308 2194 13320
rect 3050 13308 3056 13320
rect 2188 13280 3056 13308
rect 2188 13268 2194 13280
rect 3050 13268 3056 13280
rect 3108 13308 3114 13320
rect 3237 13311 3295 13317
rect 3237 13308 3249 13311
rect 3108 13280 3249 13308
rect 3108 13268 3114 13280
rect 3237 13277 3249 13280
rect 3283 13277 3295 13311
rect 3237 13271 3295 13277
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13308 4675 13311
rect 5350 13308 5356 13320
rect 4663 13280 5356 13308
rect 4663 13277 4675 13280
rect 4617 13271 4675 13277
rect 5350 13268 5356 13280
rect 5408 13308 5414 13320
rect 5534 13308 5540 13320
rect 5408 13280 5540 13308
rect 5408 13268 5414 13280
rect 5534 13268 5540 13280
rect 5592 13308 5598 13320
rect 6196 13308 6224 13339
rect 6822 13336 6828 13348
rect 6880 13336 6886 13388
rect 7006 13336 7012 13388
rect 7064 13376 7070 13388
rect 7285 13379 7343 13385
rect 7285 13376 7297 13379
rect 7064 13348 7297 13376
rect 7064 13336 7070 13348
rect 7285 13345 7297 13348
rect 7331 13345 7343 13379
rect 7285 13339 7343 13345
rect 8018 13336 8024 13388
rect 8076 13376 8082 13388
rect 8128 13385 8156 13416
rect 8294 13404 8300 13416
rect 8352 13444 8358 13456
rect 10873 13447 10931 13453
rect 8352 13416 9674 13444
rect 8352 13404 8358 13416
rect 8113 13379 8171 13385
rect 8113 13376 8125 13379
rect 8076 13348 8125 13376
rect 8076 13336 8082 13348
rect 8113 13345 8125 13348
rect 8159 13345 8171 13379
rect 8386 13376 8392 13388
rect 8347 13348 8392 13376
rect 8113 13339 8171 13345
rect 8386 13336 8392 13348
rect 8444 13336 8450 13388
rect 9646 13376 9674 13416
rect 10873 13413 10885 13447
rect 10919 13444 10931 13447
rect 11330 13444 11336 13456
rect 10919 13416 11336 13444
rect 10919 13413 10931 13416
rect 10873 13407 10931 13413
rect 11330 13404 11336 13416
rect 11388 13444 11394 13456
rect 12342 13444 12348 13456
rect 11388 13416 12348 13444
rect 11388 13404 11394 13416
rect 12342 13404 12348 13416
rect 12400 13404 12406 13456
rect 13170 13404 13176 13456
rect 13228 13444 13234 13456
rect 13228 13416 16896 13444
rect 13228 13404 13234 13416
rect 16868 13388 16896 13416
rect 9858 13376 9864 13388
rect 9646 13348 9864 13376
rect 9858 13336 9864 13348
rect 9916 13336 9922 13388
rect 10134 13336 10140 13388
rect 10192 13376 10198 13388
rect 10229 13379 10287 13385
rect 10229 13376 10241 13379
rect 10192 13348 10241 13376
rect 10192 13336 10198 13348
rect 10229 13345 10241 13348
rect 10275 13376 10287 13379
rect 10686 13376 10692 13388
rect 10275 13348 10692 13376
rect 10275 13345 10287 13348
rect 10229 13339 10287 13345
rect 10686 13336 10692 13348
rect 10744 13376 10750 13388
rect 11698 13376 11704 13388
rect 10744 13348 11704 13376
rect 10744 13336 10750 13348
rect 11698 13336 11704 13348
rect 11756 13336 11762 13388
rect 13078 13376 13084 13388
rect 12991 13348 13084 13376
rect 13078 13336 13084 13348
rect 13136 13376 13142 13388
rect 13630 13376 13636 13388
rect 13136 13348 13636 13376
rect 13136 13336 13142 13348
rect 13630 13336 13636 13348
rect 13688 13336 13694 13388
rect 13976 13379 14034 13385
rect 13976 13345 13988 13379
rect 14022 13376 14034 13379
rect 14090 13376 14096 13388
rect 14022 13348 14096 13376
rect 14022 13345 14034 13348
rect 13976 13339 14034 13345
rect 14090 13336 14096 13348
rect 14148 13336 14154 13388
rect 15565 13379 15623 13385
rect 15565 13345 15577 13379
rect 15611 13345 15623 13379
rect 15746 13376 15752 13388
rect 15707 13348 15752 13376
rect 15565 13339 15623 13345
rect 11974 13308 11980 13320
rect 5592 13280 11980 13308
rect 5592 13268 5598 13280
rect 11974 13268 11980 13280
rect 12032 13268 12038 13320
rect 12158 13308 12164 13320
rect 12119 13280 12164 13308
rect 12158 13268 12164 13280
rect 12216 13268 12222 13320
rect 15580 13308 15608 13339
rect 15746 13336 15752 13348
rect 15804 13376 15810 13388
rect 16301 13379 16359 13385
rect 16301 13376 16313 13379
rect 15804 13348 16313 13376
rect 15804 13336 15810 13348
rect 16301 13345 16313 13348
rect 16347 13345 16359 13379
rect 16850 13376 16856 13388
rect 16763 13348 16856 13376
rect 16301 13339 16359 13345
rect 16850 13336 16856 13348
rect 16908 13336 16914 13388
rect 17310 13376 17316 13388
rect 17271 13348 17316 13376
rect 17310 13336 17316 13348
rect 17368 13336 17374 13388
rect 15838 13308 15844 13320
rect 15580 13280 15844 13308
rect 15838 13268 15844 13280
rect 15896 13268 15902 13320
rect 2038 13200 2044 13252
rect 2096 13240 2102 13252
rect 4203 13243 4261 13249
rect 4203 13240 4215 13243
rect 2096 13212 4215 13240
rect 2096 13200 2102 13212
rect 4203 13209 4215 13212
rect 4249 13209 4261 13243
rect 4203 13203 4261 13209
rect 8846 13200 8852 13252
rect 8904 13240 8910 13252
rect 9950 13240 9956 13252
rect 8904 13212 9956 13240
rect 8904 13200 8910 13212
rect 9950 13200 9956 13212
rect 10008 13200 10014 13252
rect 1946 13172 1952 13184
rect 1859 13144 1952 13172
rect 1946 13132 1952 13144
rect 2004 13172 2010 13184
rect 2406 13172 2412 13184
rect 2004 13144 2412 13172
rect 2004 13132 2010 13144
rect 2406 13132 2412 13144
rect 2464 13132 2470 13184
rect 5074 13172 5080 13184
rect 5035 13144 5080 13172
rect 5074 13132 5080 13144
rect 5132 13132 5138 13184
rect 13814 13132 13820 13184
rect 13872 13172 13878 13184
rect 14047 13175 14105 13181
rect 14047 13172 14059 13175
rect 13872 13144 14059 13172
rect 13872 13132 13878 13144
rect 14047 13141 14059 13144
rect 14093 13141 14105 13175
rect 14047 13135 14105 13141
rect 15105 13175 15163 13181
rect 15105 13141 15117 13175
rect 15151 13172 15163 13175
rect 15286 13172 15292 13184
rect 15151 13144 15292 13172
rect 15151 13141 15163 13144
rect 15105 13135 15163 13141
rect 15286 13132 15292 13144
rect 15344 13132 15350 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 2958 12968 2964 12980
rect 2919 12940 2964 12968
rect 2958 12928 2964 12940
rect 3016 12928 3022 12980
rect 3602 12968 3608 12980
rect 3563 12940 3608 12968
rect 3602 12928 3608 12940
rect 3660 12928 3666 12980
rect 3970 12928 3976 12980
rect 4028 12968 4034 12980
rect 4893 12971 4951 12977
rect 4893 12968 4905 12971
rect 4028 12940 4905 12968
rect 4028 12928 4034 12940
rect 4893 12937 4905 12940
rect 4939 12937 4951 12971
rect 5350 12968 5356 12980
rect 5311 12940 5356 12968
rect 4893 12931 4951 12937
rect 5350 12928 5356 12940
rect 5408 12928 5414 12980
rect 5442 12928 5448 12980
rect 5500 12968 5506 12980
rect 5905 12971 5963 12977
rect 5905 12968 5917 12971
rect 5500 12940 5917 12968
rect 5500 12928 5506 12940
rect 5905 12937 5917 12940
rect 5951 12937 5963 12971
rect 8018 12968 8024 12980
rect 7979 12940 8024 12968
rect 5905 12931 5963 12937
rect 8018 12928 8024 12940
rect 8076 12928 8082 12980
rect 9401 12971 9459 12977
rect 9401 12937 9413 12971
rect 9447 12968 9459 12971
rect 9582 12968 9588 12980
rect 9447 12940 9588 12968
rect 9447 12937 9459 12940
rect 9401 12931 9459 12937
rect 9582 12928 9588 12940
rect 9640 12928 9646 12980
rect 10134 12968 10140 12980
rect 10095 12940 10140 12968
rect 10134 12928 10140 12940
rect 10192 12928 10198 12980
rect 12253 12971 12311 12977
rect 12253 12937 12265 12971
rect 12299 12968 12311 12971
rect 12526 12968 12532 12980
rect 12299 12940 12532 12968
rect 12299 12937 12311 12940
rect 12253 12931 12311 12937
rect 12526 12928 12532 12940
rect 12584 12928 12590 12980
rect 14829 12971 14887 12977
rect 14829 12937 14841 12971
rect 14875 12968 14887 12971
rect 15746 12968 15752 12980
rect 14875 12940 15752 12968
rect 14875 12937 14887 12940
rect 14829 12931 14887 12937
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 16850 12968 16856 12980
rect 16811 12940 16856 12968
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 2038 12832 2044 12844
rect 1999 12804 2044 12832
rect 2038 12792 2044 12804
rect 2096 12792 2102 12844
rect 2498 12832 2504 12844
rect 2459 12804 2504 12832
rect 2498 12792 2504 12804
rect 2556 12792 2562 12844
rect 3697 12835 3755 12841
rect 3697 12801 3709 12835
rect 3743 12832 3755 12835
rect 3786 12832 3792 12844
rect 3743 12804 3792 12832
rect 3743 12801 3755 12804
rect 3697 12795 3755 12801
rect 3786 12792 3792 12804
rect 3844 12832 3850 12844
rect 4522 12832 4528 12844
rect 3844 12804 4528 12832
rect 3844 12792 3850 12804
rect 4522 12792 4528 12804
rect 4580 12792 4586 12844
rect 8036 12832 8064 12928
rect 9769 12903 9827 12909
rect 9769 12869 9781 12903
rect 9815 12900 9827 12903
rect 9858 12900 9864 12912
rect 9815 12872 9864 12900
rect 9815 12869 9827 12872
rect 9769 12863 9827 12869
rect 9858 12860 9864 12872
rect 9916 12900 9922 12912
rect 11698 12900 11704 12912
rect 9916 12872 11704 12900
rect 9916 12860 9922 12872
rect 11698 12860 11704 12872
rect 11756 12860 11762 12912
rect 14734 12860 14740 12912
rect 14792 12900 14798 12912
rect 15286 12900 15292 12912
rect 14792 12872 15292 12900
rect 14792 12860 14798 12872
rect 15286 12860 15292 12872
rect 15344 12900 15350 12912
rect 15764 12900 15792 12928
rect 17221 12903 17279 12909
rect 17221 12900 17233 12903
rect 15344 12872 15424 12900
rect 15764 12872 17233 12900
rect 15344 12860 15350 12872
rect 9950 12832 9956 12844
rect 7208 12804 8064 12832
rect 8582 12804 9956 12832
rect 3602 12724 3608 12776
rect 3660 12764 3666 12776
rect 3660 12736 4108 12764
rect 3660 12724 3666 12736
rect 1670 12656 1676 12708
rect 1728 12696 1734 12708
rect 4080 12705 4108 12736
rect 6546 12724 6552 12776
rect 6604 12764 6610 12776
rect 7208 12773 7236 12804
rect 6641 12767 6699 12773
rect 6641 12764 6653 12767
rect 6604 12736 6653 12764
rect 6604 12724 6610 12736
rect 6641 12733 6653 12736
rect 6687 12764 6699 12767
rect 7193 12767 7251 12773
rect 7193 12764 7205 12767
rect 6687 12736 7205 12764
rect 6687 12733 6699 12736
rect 6641 12727 6699 12733
rect 7193 12733 7205 12736
rect 7239 12733 7251 12767
rect 7193 12727 7251 12733
rect 7469 12767 7527 12773
rect 7469 12733 7481 12767
rect 7515 12733 7527 12767
rect 7469 12727 7527 12733
rect 7653 12767 7711 12773
rect 7653 12733 7665 12767
rect 7699 12764 7711 12767
rect 8478 12764 8484 12776
rect 7699 12736 8484 12764
rect 7699 12733 7711 12736
rect 7653 12727 7711 12733
rect 1857 12699 1915 12705
rect 1857 12696 1869 12699
rect 1728 12668 1869 12696
rect 1728 12656 1734 12668
rect 1857 12665 1869 12668
rect 1903 12696 1915 12699
rect 2133 12699 2191 12705
rect 2133 12696 2145 12699
rect 1903 12668 2145 12696
rect 1903 12665 1915 12668
rect 1857 12659 1915 12665
rect 2133 12665 2145 12668
rect 2179 12696 2191 12699
rect 4059 12699 4117 12705
rect 2179 12668 3693 12696
rect 2179 12665 2191 12668
rect 2133 12659 2191 12665
rect 3665 12628 3693 12668
rect 4059 12665 4071 12699
rect 4105 12696 4117 12699
rect 5350 12696 5356 12708
rect 4105 12668 5356 12696
rect 4105 12665 4117 12668
rect 4059 12659 4117 12665
rect 5350 12656 5356 12668
rect 5408 12656 5414 12708
rect 7006 12656 7012 12708
rect 7064 12696 7070 12708
rect 7484 12696 7512 12727
rect 8478 12724 8484 12736
rect 8536 12724 8542 12776
rect 8582 12696 8610 12804
rect 9950 12792 9956 12804
rect 10008 12832 10014 12844
rect 11238 12832 11244 12844
rect 10008 12804 11244 12832
rect 10008 12792 10014 12804
rect 11238 12792 11244 12804
rect 11296 12792 11302 12844
rect 11517 12835 11575 12841
rect 11517 12801 11529 12835
rect 11563 12832 11575 12835
rect 12158 12832 12164 12844
rect 11563 12804 12164 12832
rect 11563 12801 11575 12804
rect 11517 12795 11575 12801
rect 12158 12792 12164 12804
rect 12216 12832 12222 12844
rect 12621 12835 12679 12841
rect 12621 12832 12633 12835
rect 12216 12804 12633 12832
rect 12216 12792 12222 12804
rect 12621 12801 12633 12804
rect 12667 12801 12679 12835
rect 12621 12795 12679 12801
rect 13173 12835 13231 12841
rect 13173 12801 13185 12835
rect 13219 12832 13231 12835
rect 13814 12832 13820 12844
rect 13219 12804 13820 12832
rect 13219 12801 13231 12804
rect 13173 12795 13231 12801
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 15396 12841 15424 12872
rect 17221 12869 17233 12872
rect 17267 12900 17279 12903
rect 17310 12900 17316 12912
rect 17267 12872 17316 12900
rect 17267 12869 17279 12872
rect 17221 12863 17279 12869
rect 17310 12860 17316 12872
rect 17368 12860 17374 12912
rect 15381 12835 15439 12841
rect 15381 12801 15393 12835
rect 15427 12801 15439 12835
rect 15381 12795 15439 12801
rect 8846 12764 8852 12776
rect 8759 12736 8852 12764
rect 7064 12668 8610 12696
rect 7064 12656 7070 12668
rect 4617 12631 4675 12637
rect 4617 12628 4629 12631
rect 3665 12600 4629 12628
rect 4617 12597 4629 12600
rect 4663 12597 4675 12631
rect 5442 12628 5448 12640
rect 5403 12600 5448 12628
rect 4617 12591 4675 12597
rect 5442 12588 5448 12600
rect 5500 12588 5506 12640
rect 7834 12588 7840 12640
rect 7892 12628 7898 12640
rect 8297 12631 8355 12637
rect 8297 12628 8309 12631
rect 7892 12600 8309 12628
rect 7892 12588 7898 12600
rect 8297 12597 8309 12600
rect 8343 12628 8355 12631
rect 8772 12628 8800 12736
rect 8846 12724 8852 12736
rect 8904 12724 8910 12776
rect 10781 12767 10839 12773
rect 10781 12733 10793 12767
rect 10827 12733 10839 12767
rect 11330 12764 11336 12776
rect 11291 12736 11336 12764
rect 10781 12727 10839 12733
rect 8864 12637 8892 12724
rect 8343 12600 8800 12628
rect 8849 12631 8907 12637
rect 8343 12597 8355 12600
rect 8297 12591 8355 12597
rect 8849 12597 8861 12631
rect 8895 12597 8907 12631
rect 8849 12591 8907 12597
rect 10689 12631 10747 12637
rect 10689 12597 10701 12631
rect 10735 12628 10747 12631
rect 10796 12628 10824 12727
rect 11330 12724 11336 12736
rect 11388 12724 11394 12776
rect 13265 12699 13323 12705
rect 13265 12665 13277 12699
rect 13311 12696 13323 12699
rect 13354 12696 13360 12708
rect 13311 12668 13360 12696
rect 13311 12665 13323 12668
rect 13265 12659 13323 12665
rect 13354 12656 13360 12668
rect 13412 12656 13418 12708
rect 13814 12656 13820 12708
rect 13872 12696 13878 12708
rect 14182 12696 14188 12708
rect 13872 12668 14188 12696
rect 13872 12656 13878 12668
rect 14182 12656 14188 12668
rect 14240 12656 14246 12708
rect 15473 12699 15531 12705
rect 15473 12665 15485 12699
rect 15519 12665 15531 12699
rect 16022 12696 16028 12708
rect 15983 12668 16028 12696
rect 15473 12659 15531 12665
rect 11054 12628 11060 12640
rect 10735 12600 11060 12628
rect 10735 12597 10747 12600
rect 10689 12591 10747 12597
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 14090 12628 14096 12640
rect 14051 12600 14096 12628
rect 14090 12588 14096 12600
rect 14148 12588 14154 12640
rect 15194 12628 15200 12640
rect 15155 12600 15200 12628
rect 15194 12588 15200 12600
rect 15252 12588 15258 12640
rect 15488 12628 15516 12659
rect 16022 12656 16028 12668
rect 16080 12656 16086 12708
rect 15746 12628 15752 12640
rect 15488 12600 15752 12628
rect 15746 12588 15752 12600
rect 15804 12628 15810 12640
rect 16301 12631 16359 12637
rect 16301 12628 16313 12631
rect 15804 12600 16313 12628
rect 15804 12588 15810 12600
rect 16301 12597 16313 12600
rect 16347 12597 16359 12631
rect 16301 12591 16359 12597
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1397 12427 1455 12433
rect 1397 12393 1409 12427
rect 1443 12424 1455 12427
rect 1486 12424 1492 12436
rect 1443 12396 1492 12424
rect 1443 12393 1455 12396
rect 1397 12387 1455 12393
rect 1486 12384 1492 12396
rect 1544 12384 1550 12436
rect 1946 12424 1952 12436
rect 1859 12396 1952 12424
rect 1946 12384 1952 12396
rect 2004 12424 2010 12436
rect 3786 12424 3792 12436
rect 2004 12396 2728 12424
rect 3747 12396 3792 12424
rect 2004 12384 2010 12396
rect 2038 12316 2044 12368
rect 2096 12356 2102 12368
rect 2225 12359 2283 12365
rect 2225 12356 2237 12359
rect 2096 12328 2237 12356
rect 2096 12316 2102 12328
rect 2225 12325 2237 12328
rect 2271 12325 2283 12359
rect 2590 12356 2596 12368
rect 2551 12328 2596 12356
rect 2225 12319 2283 12325
rect 2590 12316 2596 12328
rect 2648 12316 2654 12368
rect 2700 12356 2728 12396
rect 3786 12384 3792 12396
rect 3844 12384 3850 12436
rect 4614 12424 4620 12436
rect 4575 12396 4620 12424
rect 4614 12384 4620 12396
rect 4672 12384 4678 12436
rect 5074 12424 5080 12436
rect 5035 12396 5080 12424
rect 5074 12384 5080 12396
rect 5132 12384 5138 12436
rect 7006 12424 7012 12436
rect 6967 12396 7012 12424
rect 7006 12384 7012 12396
rect 7064 12384 7070 12436
rect 7834 12384 7840 12436
rect 7892 12424 7898 12436
rect 7892 12396 8201 12424
rect 7892 12384 7898 12396
rect 4203 12359 4261 12365
rect 4203 12356 4215 12359
rect 2700 12328 4215 12356
rect 4203 12325 4215 12328
rect 4249 12325 4261 12359
rect 4203 12319 4261 12325
rect 5350 12316 5356 12368
rect 5408 12356 5414 12368
rect 8173 12365 8201 12396
rect 8478 12384 8484 12436
rect 8536 12424 8542 12436
rect 9033 12427 9091 12433
rect 9033 12424 9045 12427
rect 8536 12396 9045 12424
rect 8536 12384 8542 12396
rect 9033 12393 9045 12396
rect 9079 12393 9091 12427
rect 9033 12387 9091 12393
rect 12802 12384 12808 12436
rect 12860 12424 12866 12436
rect 13354 12424 13360 12436
rect 12860 12396 13360 12424
rect 12860 12384 12866 12396
rect 13354 12384 13360 12396
rect 13412 12384 13418 12436
rect 14826 12384 14832 12436
rect 14884 12424 14890 12436
rect 14921 12427 14979 12433
rect 14921 12424 14933 12427
rect 14884 12396 14933 12424
rect 14884 12384 14890 12396
rect 14921 12393 14933 12396
rect 14967 12424 14979 12427
rect 16942 12424 16948 12436
rect 14967 12396 16948 12424
rect 14967 12393 14979 12396
rect 14921 12387 14979 12393
rect 16942 12384 16948 12396
rect 17000 12384 17006 12436
rect 17126 12424 17132 12436
rect 17087 12396 17132 12424
rect 17126 12384 17132 12396
rect 17184 12384 17190 12436
rect 5490 12359 5548 12365
rect 5490 12356 5502 12359
rect 5408 12328 5502 12356
rect 5408 12316 5414 12328
rect 5490 12325 5502 12328
rect 5536 12325 5548 12359
rect 5490 12319 5548 12325
rect 8158 12359 8216 12365
rect 8158 12325 8170 12359
rect 8204 12325 8216 12359
rect 10778 12356 10784 12368
rect 10739 12328 10784 12356
rect 8158 12319 8216 12325
rect 10778 12316 10784 12328
rect 10836 12316 10842 12368
rect 11333 12359 11391 12365
rect 11333 12325 11345 12359
rect 11379 12356 11391 12359
rect 11422 12356 11428 12368
rect 11379 12328 11428 12356
rect 11379 12325 11391 12328
rect 11333 12319 11391 12325
rect 11422 12316 11428 12328
rect 11480 12356 11486 12368
rect 11790 12356 11796 12368
rect 11480 12328 11796 12356
rect 11480 12316 11486 12328
rect 11790 12316 11796 12328
rect 11848 12316 11854 12368
rect 11882 12316 11888 12368
rect 11940 12356 11946 12368
rect 13078 12356 13084 12368
rect 11940 12328 12388 12356
rect 13039 12328 13084 12356
rect 11940 12316 11946 12328
rect 4116 12291 4174 12297
rect 4116 12257 4128 12291
rect 4162 12288 4174 12291
rect 4430 12288 4436 12300
rect 4162 12260 4436 12288
rect 4162 12257 4174 12260
rect 4116 12251 4174 12257
rect 4430 12248 4436 12260
rect 4488 12248 4494 12300
rect 5169 12291 5227 12297
rect 5169 12257 5181 12291
rect 5215 12288 5227 12291
rect 5258 12288 5264 12300
rect 5215 12260 5264 12288
rect 5215 12257 5227 12260
rect 5169 12251 5227 12257
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 7837 12291 7895 12297
rect 7837 12257 7849 12291
rect 7883 12288 7895 12291
rect 7926 12288 7932 12300
rect 7883 12260 7932 12288
rect 7883 12257 7895 12260
rect 7837 12251 7895 12257
rect 7926 12248 7932 12260
rect 7984 12248 7990 12300
rect 8754 12288 8760 12300
rect 8715 12260 8760 12288
rect 8754 12248 8760 12260
rect 8812 12248 8818 12300
rect 11974 12248 11980 12300
rect 12032 12288 12038 12300
rect 12360 12297 12388 12328
rect 13078 12316 13084 12328
rect 13136 12316 13142 12368
rect 13538 12316 13544 12368
rect 13596 12356 13602 12368
rect 13817 12359 13875 12365
rect 13817 12356 13829 12359
rect 13596 12328 13829 12356
rect 13596 12316 13602 12328
rect 13817 12325 13829 12328
rect 13863 12325 13875 12359
rect 13817 12319 13875 12325
rect 14182 12316 14188 12368
rect 14240 12356 14246 12368
rect 14369 12359 14427 12365
rect 14369 12356 14381 12359
rect 14240 12328 14381 12356
rect 14240 12316 14246 12328
rect 14369 12325 14381 12328
rect 14415 12325 14427 12359
rect 14369 12319 14427 12325
rect 14642 12316 14648 12368
rect 14700 12356 14706 12368
rect 15651 12359 15709 12365
rect 14700 12328 15516 12356
rect 14700 12316 14706 12328
rect 15488 12300 15516 12328
rect 15651 12325 15663 12359
rect 15697 12325 15709 12359
rect 15651 12319 15709 12325
rect 12158 12291 12216 12297
rect 12158 12288 12170 12291
rect 12032 12260 12170 12288
rect 12032 12248 12038 12260
rect 12158 12257 12170 12260
rect 12204 12257 12216 12291
rect 12158 12251 12216 12257
rect 12345 12291 12403 12297
rect 12345 12257 12357 12291
rect 12391 12257 12403 12291
rect 12345 12251 12403 12257
rect 15289 12291 15347 12297
rect 15289 12257 15301 12291
rect 15335 12288 15347 12291
rect 15378 12288 15384 12300
rect 15335 12260 15384 12288
rect 15335 12257 15347 12260
rect 15289 12251 15347 12257
rect 15378 12248 15384 12260
rect 15436 12248 15442 12300
rect 15470 12248 15476 12300
rect 15528 12288 15534 12300
rect 15672 12288 15700 12319
rect 15930 12288 15936 12300
rect 15528 12260 15936 12288
rect 15528 12248 15534 12260
rect 15930 12248 15936 12260
rect 15988 12248 15994 12300
rect 17310 12288 17316 12300
rect 17271 12260 17316 12288
rect 17310 12248 17316 12260
rect 17368 12248 17374 12300
rect 17586 12288 17592 12300
rect 17547 12260 17592 12288
rect 17586 12248 17592 12260
rect 17644 12248 17650 12300
rect 2498 12220 2504 12232
rect 2459 12192 2504 12220
rect 2498 12180 2504 12192
rect 2556 12180 2562 12232
rect 3142 12220 3148 12232
rect 3103 12192 3148 12220
rect 3142 12180 3148 12192
rect 3200 12180 3206 12232
rect 10042 12180 10048 12232
rect 10100 12220 10106 12232
rect 10689 12223 10747 12229
rect 10689 12220 10701 12223
rect 10100 12192 10701 12220
rect 10100 12180 10106 12192
rect 10689 12189 10701 12192
rect 10735 12189 10747 12223
rect 10689 12183 10747 12189
rect 12713 12223 12771 12229
rect 12713 12189 12725 12223
rect 12759 12220 12771 12223
rect 13725 12223 13783 12229
rect 12759 12192 13400 12220
rect 12759 12189 12771 12192
rect 12713 12183 12771 12189
rect 13372 12152 13400 12192
rect 13725 12189 13737 12223
rect 13771 12220 13783 12223
rect 14182 12220 14188 12232
rect 13771 12192 14188 12220
rect 13771 12189 13783 12192
rect 13725 12183 13783 12189
rect 14182 12180 14188 12192
rect 14240 12180 14246 12232
rect 15194 12180 15200 12232
rect 15252 12220 15258 12232
rect 15838 12220 15844 12232
rect 15252 12192 15844 12220
rect 15252 12180 15258 12192
rect 15838 12180 15844 12192
rect 15896 12220 15902 12232
rect 17604 12220 17632 12248
rect 15896 12192 17632 12220
rect 15896 12180 15902 12192
rect 16850 12152 16856 12164
rect 13372 12124 16856 12152
rect 16850 12112 16856 12124
rect 16908 12112 16914 12164
rect 4706 12044 4712 12096
rect 4764 12084 4770 12096
rect 6089 12087 6147 12093
rect 6089 12084 6101 12087
rect 4764 12056 6101 12084
rect 4764 12044 4770 12056
rect 6089 12053 6101 12056
rect 6135 12053 6147 12087
rect 6089 12047 6147 12053
rect 7745 12087 7803 12093
rect 7745 12053 7757 12087
rect 7791 12084 7803 12087
rect 8386 12084 8392 12096
rect 7791 12056 8392 12084
rect 7791 12053 7803 12056
rect 7745 12047 7803 12053
rect 8386 12044 8392 12056
rect 8444 12084 8450 12096
rect 11054 12084 11060 12096
rect 8444 12056 11060 12084
rect 8444 12044 8450 12056
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 15470 12044 15476 12096
rect 15528 12084 15534 12096
rect 16209 12087 16267 12093
rect 16209 12084 16221 12087
rect 15528 12056 16221 12084
rect 15528 12044 15534 12056
rect 16209 12053 16221 12056
rect 16255 12053 16267 12087
rect 16209 12047 16267 12053
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 5077 11883 5135 11889
rect 5077 11849 5089 11883
rect 5123 11880 5135 11883
rect 5350 11880 5356 11892
rect 5123 11852 5356 11880
rect 5123 11849 5135 11852
rect 5077 11843 5135 11849
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 7926 11840 7932 11892
rect 7984 11880 7990 11892
rect 8205 11883 8263 11889
rect 8205 11880 8217 11883
rect 7984 11852 8217 11880
rect 7984 11840 7990 11852
rect 8205 11849 8217 11852
rect 8251 11849 8263 11883
rect 8205 11843 8263 11849
rect 10778 11840 10784 11892
rect 10836 11880 10842 11892
rect 11149 11883 11207 11889
rect 11149 11880 11161 11883
rect 10836 11852 11161 11880
rect 10836 11840 10842 11852
rect 11149 11849 11161 11852
rect 11195 11880 11207 11883
rect 11425 11883 11483 11889
rect 11425 11880 11437 11883
rect 11195 11852 11437 11880
rect 11195 11849 11207 11852
rect 11149 11843 11207 11849
rect 11425 11849 11437 11852
rect 11471 11849 11483 11883
rect 11425 11843 11483 11849
rect 11882 11840 11888 11892
rect 11940 11880 11946 11892
rect 12161 11883 12219 11889
rect 12161 11880 12173 11883
rect 11940 11852 12173 11880
rect 11940 11840 11946 11852
rect 12161 11849 12173 11852
rect 12207 11849 12219 11883
rect 12161 11843 12219 11849
rect 13538 11840 13544 11892
rect 13596 11880 13602 11892
rect 13633 11883 13691 11889
rect 13633 11880 13645 11883
rect 13596 11852 13645 11880
rect 13596 11840 13602 11852
rect 13633 11849 13645 11852
rect 13679 11849 13691 11883
rect 14642 11880 14648 11892
rect 14603 11852 14648 11880
rect 13633 11843 13691 11849
rect 14642 11840 14648 11852
rect 14700 11840 14706 11892
rect 15746 11880 15752 11892
rect 15707 11852 15752 11880
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 15930 11840 15936 11892
rect 15988 11880 15994 11892
rect 16025 11883 16083 11889
rect 16025 11880 16037 11883
rect 15988 11852 16037 11880
rect 15988 11840 15994 11852
rect 16025 11849 16037 11852
rect 16071 11849 16083 11883
rect 16025 11843 16083 11849
rect 16574 11840 16580 11892
rect 16632 11880 16638 11892
rect 16715 11883 16773 11889
rect 16715 11880 16727 11883
rect 16632 11852 16727 11880
rect 16632 11840 16638 11852
rect 16715 11849 16727 11852
rect 16761 11849 16773 11883
rect 16715 11843 16773 11849
rect 17310 11840 17316 11892
rect 17368 11880 17374 11892
rect 17405 11883 17463 11889
rect 17405 11880 17417 11883
rect 17368 11852 17417 11880
rect 17368 11840 17374 11852
rect 17405 11849 17417 11852
rect 17451 11849 17463 11883
rect 17405 11843 17463 11849
rect 4157 11815 4215 11821
rect 4157 11781 4169 11815
rect 4203 11812 4215 11815
rect 4430 11812 4436 11824
rect 4203 11784 4436 11812
rect 4203 11781 4215 11784
rect 4157 11775 4215 11781
rect 4430 11772 4436 11784
rect 4488 11812 4494 11824
rect 8018 11812 8024 11824
rect 4488 11784 8024 11812
rect 4488 11772 4494 11784
rect 8018 11772 8024 11784
rect 8076 11772 8082 11824
rect 11793 11815 11851 11821
rect 11793 11781 11805 11815
rect 11839 11812 11851 11815
rect 11974 11812 11980 11824
rect 11839 11784 11980 11812
rect 11839 11781 11851 11784
rect 11793 11775 11851 11781
rect 11974 11772 11980 11784
rect 12032 11772 12038 11824
rect 15378 11772 15384 11824
rect 15436 11812 15442 11824
rect 16393 11815 16451 11821
rect 16393 11812 16405 11815
rect 15436 11784 16405 11812
rect 15436 11772 15442 11784
rect 16393 11781 16405 11784
rect 16439 11781 16451 11815
rect 16393 11775 16451 11781
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11744 1639 11747
rect 1946 11744 1952 11756
rect 1627 11716 1952 11744
rect 1627 11713 1639 11716
rect 1581 11707 1639 11713
rect 1946 11704 1952 11716
rect 2004 11704 2010 11756
rect 2682 11704 2688 11756
rect 2740 11744 2746 11756
rect 3142 11744 3148 11756
rect 2740 11716 3148 11744
rect 2740 11704 2746 11716
rect 3142 11704 3148 11716
rect 3200 11744 3206 11756
rect 3421 11747 3479 11753
rect 3421 11744 3433 11747
rect 3200 11716 3433 11744
rect 3200 11704 3206 11716
rect 3421 11713 3433 11716
rect 3467 11713 3479 11747
rect 3421 11707 3479 11713
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11744 4767 11747
rect 5261 11747 5319 11753
rect 5261 11744 5273 11747
rect 4755 11716 5273 11744
rect 4755 11713 4767 11716
rect 4709 11707 4767 11713
rect 5261 11713 5273 11716
rect 5307 11744 5319 11747
rect 5442 11744 5448 11756
rect 5307 11716 5448 11744
rect 5307 11713 5319 11716
rect 5261 11707 5319 11713
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 5534 11704 5540 11756
rect 5592 11744 5598 11756
rect 5592 11716 5637 11744
rect 5592 11704 5598 11716
rect 8294 11704 8300 11756
rect 8352 11744 8358 11756
rect 9033 11747 9091 11753
rect 9033 11744 9045 11747
rect 8352 11716 9045 11744
rect 8352 11704 8358 11716
rect 9033 11713 9045 11716
rect 9079 11744 9091 11747
rect 9677 11747 9735 11753
rect 9677 11744 9689 11747
rect 9079 11716 9689 11744
rect 9079 11713 9091 11716
rect 9033 11707 9091 11713
rect 9677 11713 9689 11716
rect 9723 11744 9735 11747
rect 10042 11744 10048 11756
rect 9723 11716 10048 11744
rect 9723 11713 9735 11716
rect 9677 11707 9735 11713
rect 10042 11704 10048 11716
rect 10100 11704 10106 11756
rect 10134 11704 10140 11756
rect 10192 11744 10198 11756
rect 10229 11747 10287 11753
rect 10229 11744 10241 11747
rect 10192 11716 10241 11744
rect 10192 11704 10198 11716
rect 10229 11713 10241 11716
rect 10275 11744 10287 11747
rect 17126 11744 17132 11756
rect 10275 11716 17132 11744
rect 10275 11713 10287 11716
rect 10229 11707 10287 11713
rect 17126 11704 17132 11716
rect 17184 11704 17190 11756
rect 6641 11679 6699 11685
rect 6641 11645 6653 11679
rect 6687 11676 6699 11679
rect 6730 11676 6736 11688
rect 6687 11648 6736 11676
rect 6687 11645 6699 11648
rect 6641 11639 6699 11645
rect 6730 11636 6736 11648
rect 6788 11676 6794 11688
rect 6917 11679 6975 11685
rect 6917 11676 6929 11679
rect 6788 11648 6929 11676
rect 6788 11636 6794 11648
rect 6917 11645 6929 11648
rect 6963 11645 6975 11679
rect 14826 11676 14832 11688
rect 14787 11648 14832 11676
rect 6917 11639 6975 11645
rect 14826 11636 14832 11648
rect 14884 11636 14890 11688
rect 16644 11679 16702 11685
rect 16644 11645 16656 11679
rect 16690 11676 16702 11679
rect 17034 11676 17040 11688
rect 16690 11648 17040 11676
rect 16690 11645 16702 11648
rect 16644 11639 16702 11645
rect 17034 11636 17040 11648
rect 17092 11636 17098 11688
rect 1670 11608 1676 11620
rect 1631 11580 1676 11608
rect 1670 11568 1676 11580
rect 1728 11568 1734 11620
rect 2225 11611 2283 11617
rect 2225 11577 2237 11611
rect 2271 11608 2283 11611
rect 3142 11608 3148 11620
rect 2271 11580 3148 11608
rect 2271 11577 2283 11580
rect 2225 11571 2283 11577
rect 3142 11568 3148 11580
rect 3200 11568 3206 11620
rect 3234 11568 3240 11620
rect 3292 11608 3298 11620
rect 3292 11580 3337 11608
rect 3292 11568 3298 11580
rect 5074 11568 5080 11620
rect 5132 11608 5138 11620
rect 5330 11611 5388 11617
rect 5330 11608 5342 11611
rect 5132 11580 5342 11608
rect 5132 11568 5138 11580
rect 5330 11577 5342 11580
rect 5376 11577 5388 11611
rect 5330 11571 5388 11577
rect 5626 11568 5632 11620
rect 5684 11608 5690 11620
rect 6825 11611 6883 11617
rect 6825 11608 6837 11611
rect 5684 11580 6837 11608
rect 5684 11568 5690 11580
rect 6825 11577 6837 11580
rect 6871 11577 6883 11611
rect 6825 11571 6883 11577
rect 8757 11611 8815 11617
rect 8757 11577 8769 11611
rect 8803 11577 8815 11611
rect 8757 11571 8815 11577
rect 2590 11540 2596 11552
rect 2551 11512 2596 11540
rect 2590 11500 2596 11512
rect 2648 11500 2654 11552
rect 2961 11543 3019 11549
rect 2961 11509 2973 11543
rect 3007 11540 3019 11543
rect 3252 11540 3280 11568
rect 7834 11540 7840 11552
rect 3007 11512 3280 11540
rect 7795 11512 7840 11540
rect 3007 11509 3019 11512
rect 2961 11503 3019 11509
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 8772 11540 8800 11571
rect 8846 11568 8852 11620
rect 8904 11608 8910 11620
rect 9214 11608 9220 11620
rect 8904 11580 9220 11608
rect 8904 11568 8910 11580
rect 9214 11568 9220 11580
rect 9272 11568 9278 11620
rect 10137 11611 10195 11617
rect 10137 11577 10149 11611
rect 10183 11608 10195 11611
rect 10591 11611 10649 11617
rect 10591 11608 10603 11611
rect 10183 11580 10603 11608
rect 10183 11577 10195 11580
rect 10137 11571 10195 11577
rect 10591 11577 10603 11580
rect 10637 11608 10649 11611
rect 10778 11608 10784 11620
rect 10637 11580 10784 11608
rect 10637 11577 10649 11580
rect 10591 11571 10649 11577
rect 10778 11568 10784 11580
rect 10836 11608 10842 11620
rect 11882 11608 11888 11620
rect 10836 11580 11888 11608
rect 10836 11568 10842 11580
rect 11882 11568 11888 11580
rect 11940 11608 11946 11620
rect 12526 11608 12532 11620
rect 11940 11580 12532 11608
rect 11940 11568 11946 11580
rect 12526 11568 12532 11580
rect 12584 11568 12590 11620
rect 12710 11608 12716 11620
rect 12671 11580 12716 11608
rect 12710 11568 12716 11580
rect 12768 11568 12774 11620
rect 12805 11611 12863 11617
rect 12805 11577 12817 11611
rect 12851 11608 12863 11611
rect 13078 11608 13084 11620
rect 12851 11580 13084 11608
rect 12851 11577 12863 11580
rect 12805 11571 12863 11577
rect 13078 11568 13084 11580
rect 13136 11568 13142 11620
rect 13354 11608 13360 11620
rect 13315 11580 13360 11608
rect 13354 11568 13360 11580
rect 13412 11568 13418 11620
rect 14642 11568 14648 11620
rect 14700 11608 14706 11620
rect 15150 11611 15208 11617
rect 15150 11608 15162 11611
rect 14700 11580 15162 11608
rect 14700 11568 14706 11580
rect 15150 11577 15162 11580
rect 15196 11577 15208 11611
rect 15150 11571 15208 11577
rect 9122 11540 9128 11552
rect 8772 11512 9128 11540
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 14093 11543 14151 11549
rect 14093 11509 14105 11543
rect 14139 11540 14151 11543
rect 14274 11540 14280 11552
rect 14139 11512 14280 11540
rect 14139 11509 14151 11512
rect 14093 11503 14151 11509
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 16758 11500 16764 11552
rect 16816 11540 16822 11552
rect 17586 11540 17592 11552
rect 16816 11512 17592 11540
rect 16816 11500 16822 11512
rect 17586 11500 17592 11512
rect 17644 11540 17650 11552
rect 17773 11543 17831 11549
rect 17773 11540 17785 11543
rect 17644 11512 17785 11540
rect 17644 11500 17650 11512
rect 17773 11509 17785 11512
rect 17819 11509 17831 11543
rect 17773 11503 17831 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1670 11336 1676 11348
rect 1631 11308 1676 11336
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 3142 11296 3148 11348
rect 3200 11336 3206 11348
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 3200 11308 3433 11336
rect 3200 11296 3206 11308
rect 3421 11305 3433 11308
rect 3467 11305 3479 11339
rect 3421 11299 3479 11305
rect 5074 11296 5080 11348
rect 5132 11336 5138 11348
rect 5261 11339 5319 11345
rect 5261 11336 5273 11339
rect 5132 11308 5273 11336
rect 5132 11296 5138 11308
rect 5261 11305 5273 11308
rect 5307 11336 5319 11339
rect 5626 11336 5632 11348
rect 5307 11308 5632 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 6730 11336 6736 11348
rect 6691 11308 6736 11336
rect 6730 11296 6736 11308
rect 6788 11296 6794 11348
rect 7834 11296 7840 11348
rect 7892 11336 7898 11348
rect 7929 11339 7987 11345
rect 7929 11336 7941 11339
rect 7892 11308 7941 11336
rect 7892 11296 7898 11308
rect 7929 11305 7941 11308
rect 7975 11305 7987 11339
rect 7929 11299 7987 11305
rect 8202 11296 8208 11348
rect 8260 11336 8266 11348
rect 8846 11336 8852 11348
rect 8260 11308 8852 11336
rect 8260 11296 8266 11308
rect 8846 11296 8852 11308
rect 8904 11296 8910 11348
rect 10134 11296 10140 11348
rect 10192 11336 10198 11348
rect 10229 11339 10287 11345
rect 10229 11336 10241 11339
rect 10192 11308 10241 11336
rect 10192 11296 10198 11308
rect 10229 11305 10241 11308
rect 10275 11305 10287 11339
rect 10778 11336 10784 11348
rect 10739 11308 10784 11336
rect 10229 11299 10287 11305
rect 10778 11296 10784 11308
rect 10836 11296 10842 11348
rect 12529 11339 12587 11345
rect 12529 11305 12541 11339
rect 12575 11336 12587 11339
rect 12710 11336 12716 11348
rect 12575 11308 12716 11336
rect 12575 11305 12587 11308
rect 12529 11299 12587 11305
rect 12710 11296 12716 11308
rect 12768 11336 12774 11348
rect 12768 11308 13492 11336
rect 12768 11296 12774 11308
rect 2222 11268 2228 11280
rect 2183 11240 2228 11268
rect 2222 11228 2228 11240
rect 2280 11228 2286 11280
rect 2590 11228 2596 11280
rect 2648 11268 2654 11280
rect 4065 11271 4123 11277
rect 4065 11268 4077 11271
rect 2648 11240 4077 11268
rect 2648 11228 2654 11240
rect 4065 11237 4077 11240
rect 4111 11237 4123 11271
rect 4065 11231 4123 11237
rect 5350 11228 5356 11280
rect 5408 11268 5414 11280
rect 6178 11277 6184 11280
rect 6134 11271 6184 11277
rect 6134 11268 6146 11271
rect 5408 11240 6146 11268
rect 5408 11228 5414 11240
rect 6134 11237 6146 11240
rect 6180 11237 6184 11271
rect 6134 11231 6184 11237
rect 6178 11228 6184 11231
rect 6236 11228 6242 11280
rect 12802 11268 12808 11280
rect 12763 11240 12808 11268
rect 12802 11228 12808 11240
rect 12860 11228 12866 11280
rect 13464 11268 13492 11308
rect 13538 11296 13544 11348
rect 13596 11336 13602 11348
rect 14458 11336 14464 11348
rect 13596 11308 14464 11336
rect 13596 11296 13602 11308
rect 14458 11296 14464 11308
rect 14516 11336 14522 11348
rect 14645 11339 14703 11345
rect 14645 11336 14657 11339
rect 14516 11308 14657 11336
rect 14516 11296 14522 11308
rect 14645 11305 14657 11308
rect 14691 11305 14703 11339
rect 14645 11299 14703 11305
rect 14826 11268 14832 11280
rect 13464 11240 14832 11268
rect 14826 11228 14832 11240
rect 14884 11228 14890 11280
rect 15470 11268 15476 11280
rect 15431 11240 15476 11268
rect 15470 11228 15476 11240
rect 15528 11228 15534 11280
rect 16022 11268 16028 11280
rect 15983 11240 16028 11268
rect 16022 11228 16028 11240
rect 16080 11228 16086 11280
rect 3234 11160 3240 11212
rect 3292 11200 3298 11212
rect 4706 11200 4712 11212
rect 3292 11172 4712 11200
rect 3292 11160 3298 11172
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 5258 11160 5264 11212
rect 5316 11200 5322 11212
rect 5537 11203 5595 11209
rect 5537 11200 5549 11203
rect 5316 11172 5549 11200
rect 5316 11160 5322 11172
rect 5537 11169 5549 11172
rect 5583 11169 5595 11203
rect 5537 11163 5595 11169
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11200 5871 11203
rect 6914 11200 6920 11212
rect 5859 11172 6920 11200
rect 5859 11169 5871 11172
rect 5813 11163 5871 11169
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 7098 11160 7104 11212
rect 7156 11200 7162 11212
rect 7561 11203 7619 11209
rect 7561 11200 7573 11203
rect 7156 11172 7573 11200
rect 7156 11160 7162 11172
rect 7561 11169 7573 11172
rect 7607 11169 7619 11203
rect 7561 11163 7619 11169
rect 14252 11203 14310 11209
rect 14252 11169 14264 11203
rect 14298 11200 14310 11203
rect 14366 11200 14372 11212
rect 14298 11172 14372 11200
rect 14298 11169 14310 11172
rect 14252 11163 14310 11169
rect 14366 11160 14372 11172
rect 14424 11160 14430 11212
rect 2130 11132 2136 11144
rect 2091 11104 2136 11132
rect 2130 11092 2136 11104
rect 2188 11092 2194 11144
rect 2498 11092 2504 11144
rect 2556 11132 2562 11144
rect 2777 11135 2835 11141
rect 2777 11132 2789 11135
rect 2556 11104 2789 11132
rect 2556 11092 2562 11104
rect 2777 11101 2789 11104
rect 2823 11132 2835 11135
rect 3789 11135 3847 11141
rect 3789 11132 3801 11135
rect 2823 11104 3801 11132
rect 2823 11101 2835 11104
rect 2777 11095 2835 11101
rect 3789 11101 3801 11104
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 10413 11135 10471 11141
rect 10413 11101 10425 11135
rect 10459 11132 10471 11135
rect 11238 11132 11244 11144
rect 10459 11104 11244 11132
rect 10459 11101 10471 11104
rect 10413 11095 10471 11101
rect 11238 11092 11244 11104
rect 11296 11092 11302 11144
rect 12710 11132 12716 11144
rect 12671 11104 12716 11132
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 13354 11132 13360 11144
rect 13267 11104 13360 11132
rect 13354 11092 13360 11104
rect 13412 11132 13418 11144
rect 14734 11132 14740 11144
rect 13412 11104 14740 11132
rect 13412 11092 13418 11104
rect 14734 11092 14740 11104
rect 14792 11092 14798 11144
rect 15381 11135 15439 11141
rect 15381 11101 15393 11135
rect 15427 11101 15439 11135
rect 15381 11095 15439 11101
rect 13814 11024 13820 11076
rect 13872 11064 13878 11076
rect 15396 11064 15424 11095
rect 15562 11092 15568 11144
rect 15620 11132 15626 11144
rect 16853 11135 16911 11141
rect 16853 11132 16865 11135
rect 15620 11104 16865 11132
rect 15620 11092 15626 11104
rect 16853 11101 16865 11104
rect 16899 11101 16911 11135
rect 16853 11095 16911 11101
rect 15746 11064 15752 11076
rect 13872 11036 15752 11064
rect 13872 11024 13878 11036
rect 15746 11024 15752 11036
rect 15804 11024 15810 11076
rect 3050 10996 3056 11008
rect 3011 10968 3056 10996
rect 3050 10956 3056 10968
rect 3108 10956 3114 11008
rect 5350 10956 5356 11008
rect 5408 10996 5414 11008
rect 8481 10999 8539 11005
rect 8481 10996 8493 10999
rect 5408 10968 8493 10996
rect 5408 10956 5414 10968
rect 8481 10965 8493 10968
rect 8527 10965 8539 10999
rect 9122 10996 9128 11008
rect 9083 10968 9128 10996
rect 8481 10959 8539 10965
rect 9122 10956 9128 10968
rect 9180 10956 9186 11008
rect 11330 10996 11336 11008
rect 11291 10968 11336 10996
rect 11330 10956 11336 10968
rect 11388 10956 11394 11008
rect 11606 10996 11612 11008
rect 11567 10968 11612 10996
rect 11606 10956 11612 10968
rect 11664 10956 11670 11008
rect 13538 10956 13544 11008
rect 13596 10996 13602 11008
rect 14323 10999 14381 11005
rect 14323 10996 14335 10999
rect 13596 10968 14335 10996
rect 13596 10956 13602 10968
rect 14323 10965 14335 10968
rect 14369 10965 14381 10999
rect 14323 10959 14381 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 4706 10792 4712 10804
rect 4667 10764 4712 10792
rect 4706 10752 4712 10764
rect 4764 10752 4770 10804
rect 6178 10792 6184 10804
rect 6139 10764 6184 10792
rect 6178 10752 6184 10764
rect 6236 10752 6242 10804
rect 6641 10795 6699 10801
rect 6641 10761 6653 10795
rect 6687 10792 6699 10795
rect 6914 10792 6920 10804
rect 6687 10764 6920 10792
rect 6687 10761 6699 10764
rect 6641 10755 6699 10761
rect 6914 10752 6920 10764
rect 6972 10752 6978 10804
rect 7098 10792 7104 10804
rect 7059 10764 7104 10792
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 10505 10795 10563 10801
rect 10505 10761 10517 10795
rect 10551 10792 10563 10795
rect 10778 10792 10784 10804
rect 10551 10764 10784 10792
rect 10551 10761 10563 10764
rect 10505 10755 10563 10761
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 11330 10752 11336 10804
rect 11388 10792 11394 10804
rect 11793 10795 11851 10801
rect 11793 10792 11805 10795
rect 11388 10764 11805 10792
rect 11388 10752 11394 10764
rect 11793 10761 11805 10764
rect 11839 10761 11851 10795
rect 11793 10755 11851 10761
rect 14185 10795 14243 10801
rect 14185 10761 14197 10795
rect 14231 10792 14243 10795
rect 14366 10792 14372 10804
rect 14231 10764 14372 10792
rect 14231 10761 14243 10764
rect 14185 10755 14243 10761
rect 14366 10752 14372 10764
rect 14424 10752 14430 10804
rect 15381 10795 15439 10801
rect 15381 10761 15393 10795
rect 15427 10792 15439 10795
rect 15470 10792 15476 10804
rect 15427 10764 15476 10792
rect 15427 10761 15439 10764
rect 15381 10755 15439 10761
rect 15470 10752 15476 10764
rect 15528 10752 15534 10804
rect 15746 10792 15752 10804
rect 15707 10764 15752 10792
rect 15746 10752 15752 10764
rect 15804 10752 15810 10804
rect 3142 10724 3148 10736
rect 3103 10696 3148 10724
rect 3142 10684 3148 10696
rect 3200 10684 3206 10736
rect 6196 10724 6224 10752
rect 7469 10727 7527 10733
rect 7469 10724 7481 10727
rect 6196 10696 7481 10724
rect 7469 10693 7481 10696
rect 7515 10724 7527 10727
rect 7834 10724 7840 10736
rect 7515 10696 7840 10724
rect 7515 10693 7527 10696
rect 7469 10687 7527 10693
rect 7834 10684 7840 10696
rect 7892 10684 7898 10736
rect 8294 10724 8300 10736
rect 8255 10696 8300 10724
rect 8294 10684 8300 10696
rect 8352 10684 8358 10736
rect 11422 10724 11428 10736
rect 11383 10696 11428 10724
rect 11422 10684 11428 10696
rect 11480 10684 11486 10736
rect 12710 10684 12716 10736
rect 12768 10724 12774 10736
rect 15979 10727 16037 10733
rect 15979 10724 15991 10727
rect 12768 10696 15991 10724
rect 12768 10684 12774 10696
rect 15979 10693 15991 10696
rect 16025 10693 16037 10727
rect 15979 10687 16037 10693
rect 2590 10656 2596 10668
rect 2503 10628 2596 10656
rect 2590 10616 2596 10628
rect 2648 10656 2654 10668
rect 3050 10656 3056 10668
rect 2648 10628 3056 10656
rect 2648 10616 2654 10628
rect 3050 10616 3056 10628
rect 3108 10616 3114 10668
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10656 4215 10659
rect 9033 10659 9091 10665
rect 9033 10656 9045 10659
rect 4203 10628 9045 10656
rect 4203 10625 4215 10628
rect 4157 10619 4215 10625
rect 9033 10625 9045 10628
rect 9079 10656 9091 10659
rect 9309 10659 9367 10665
rect 9309 10656 9321 10659
rect 9079 10628 9321 10656
rect 9079 10625 9091 10628
rect 9033 10619 9091 10625
rect 9309 10625 9321 10628
rect 9355 10625 9367 10659
rect 9309 10619 9367 10625
rect 9398 10616 9404 10668
rect 9456 10656 9462 10668
rect 9953 10659 10011 10665
rect 9953 10656 9965 10659
rect 9456 10628 9965 10656
rect 9456 10616 9462 10628
rect 9953 10625 9965 10628
rect 9999 10656 10011 10659
rect 10873 10659 10931 10665
rect 10873 10656 10885 10659
rect 9999 10628 10885 10656
rect 9999 10625 10011 10628
rect 9953 10619 10011 10625
rect 10873 10625 10885 10628
rect 10919 10656 10931 10659
rect 11606 10656 11612 10668
rect 10919 10628 11612 10656
rect 10919 10625 10931 10628
rect 10873 10619 10931 10625
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 12805 10659 12863 10665
rect 12805 10625 12817 10659
rect 12851 10656 12863 10659
rect 13538 10656 13544 10668
rect 12851 10628 13544 10656
rect 12851 10625 12863 10628
rect 12805 10619 12863 10625
rect 13538 10616 13544 10628
rect 13596 10616 13602 10668
rect 13817 10659 13875 10665
rect 13817 10625 13829 10659
rect 13863 10656 13875 10659
rect 14369 10659 14427 10665
rect 14369 10656 14381 10659
rect 13863 10628 14381 10656
rect 13863 10625 13875 10628
rect 13817 10619 13875 10625
rect 14369 10625 14381 10628
rect 14415 10656 14427 10659
rect 15562 10656 15568 10668
rect 14415 10628 15568 10656
rect 14415 10625 14427 10628
rect 14369 10619 14427 10625
rect 15562 10616 15568 10628
rect 15620 10616 15626 10668
rect 15908 10591 15966 10597
rect 15908 10557 15920 10591
rect 15954 10557 15966 10591
rect 16850 10588 16856 10600
rect 16811 10560 16856 10588
rect 15908 10551 15966 10557
rect 1489 10523 1547 10529
rect 1489 10489 1501 10523
rect 1535 10520 1547 10523
rect 2130 10520 2136 10532
rect 1535 10492 2136 10520
rect 1535 10489 1547 10492
rect 1489 10483 1547 10489
rect 2130 10480 2136 10492
rect 2188 10480 2194 10532
rect 2685 10523 2743 10529
rect 2685 10489 2697 10523
rect 2731 10520 2743 10523
rect 2866 10520 2872 10532
rect 2731 10492 2872 10520
rect 2731 10489 2743 10492
rect 2685 10483 2743 10489
rect 2041 10455 2099 10461
rect 2041 10421 2053 10455
rect 2087 10452 2099 10455
rect 2222 10452 2228 10464
rect 2087 10424 2228 10452
rect 2087 10421 2099 10424
rect 2041 10415 2099 10421
rect 2222 10412 2228 10424
rect 2280 10452 2286 10464
rect 2700 10452 2728 10483
rect 2866 10480 2872 10492
rect 2924 10520 2930 10532
rect 3513 10523 3571 10529
rect 3513 10520 3525 10523
rect 2924 10492 3525 10520
rect 2924 10480 2930 10492
rect 3513 10489 3525 10492
rect 3559 10489 3571 10523
rect 5258 10520 5264 10532
rect 3513 10483 3571 10489
rect 4126 10492 5120 10520
rect 5219 10492 5264 10520
rect 2280 10424 2728 10452
rect 2280 10412 2286 10424
rect 3970 10412 3976 10464
rect 4028 10452 4034 10464
rect 4126 10452 4154 10492
rect 5092 10461 5120 10492
rect 5258 10480 5264 10492
rect 5316 10480 5322 10532
rect 5350 10480 5356 10532
rect 5408 10520 5414 10532
rect 5905 10523 5963 10529
rect 5408 10492 5453 10520
rect 5408 10480 5414 10492
rect 5905 10489 5917 10523
rect 5951 10520 5963 10523
rect 5994 10520 6000 10532
rect 5951 10492 6000 10520
rect 5951 10489 5963 10492
rect 5905 10483 5963 10489
rect 5994 10480 6000 10492
rect 6052 10480 6058 10532
rect 7742 10520 7748 10532
rect 7703 10492 7748 10520
rect 7742 10480 7748 10492
rect 7800 10480 7806 10532
rect 7834 10480 7840 10532
rect 7892 10520 7898 10532
rect 9401 10523 9459 10529
rect 9401 10520 9413 10523
rect 7892 10492 9413 10520
rect 7892 10480 7898 10492
rect 9401 10489 9413 10492
rect 9447 10520 9459 10523
rect 9582 10520 9588 10532
rect 9447 10492 9588 10520
rect 9447 10489 9459 10492
rect 9401 10483 9459 10489
rect 9582 10480 9588 10492
rect 9640 10480 9646 10532
rect 10965 10523 11023 10529
rect 10965 10489 10977 10523
rect 11011 10520 11023 10523
rect 11330 10520 11336 10532
rect 11011 10492 11336 10520
rect 11011 10489 11023 10492
rect 10965 10483 11023 10489
rect 11330 10480 11336 10492
rect 11388 10480 11394 10532
rect 12897 10523 12955 10529
rect 12897 10489 12909 10523
rect 12943 10520 12955 10523
rect 13078 10520 13084 10532
rect 12943 10492 13084 10520
rect 12943 10489 12955 10492
rect 12897 10483 12955 10489
rect 13078 10480 13084 10492
rect 13136 10480 13142 10532
rect 13449 10523 13507 10529
rect 13449 10489 13461 10523
rect 13495 10520 13507 10523
rect 13814 10520 13820 10532
rect 13495 10492 13820 10520
rect 13495 10489 13507 10492
rect 13449 10483 13507 10489
rect 13814 10480 13820 10492
rect 13872 10480 13878 10532
rect 14458 10520 14464 10532
rect 14419 10492 14464 10520
rect 14458 10480 14464 10492
rect 14516 10480 14522 10532
rect 14734 10480 14740 10532
rect 14792 10520 14798 10532
rect 15013 10523 15071 10529
rect 15013 10520 15025 10523
rect 14792 10492 15025 10520
rect 14792 10480 14798 10492
rect 15013 10489 15025 10492
rect 15059 10489 15071 10523
rect 15013 10483 15071 10489
rect 15746 10480 15752 10532
rect 15804 10520 15810 10532
rect 15923 10520 15951 10551
rect 16850 10548 16856 10560
rect 16908 10588 16914 10600
rect 17313 10591 17371 10597
rect 17313 10588 17325 10591
rect 16908 10560 17325 10588
rect 16908 10548 16914 10560
rect 17313 10557 17325 10560
rect 17359 10557 17371 10591
rect 17313 10551 17371 10557
rect 16301 10523 16359 10529
rect 16301 10520 16313 10523
rect 15804 10492 16313 10520
rect 15804 10480 15810 10492
rect 16301 10489 16313 10492
rect 16347 10489 16359 10523
rect 16301 10483 16359 10489
rect 4028 10424 4154 10452
rect 5077 10455 5135 10461
rect 4028 10412 4034 10424
rect 5077 10421 5089 10455
rect 5123 10452 5135 10455
rect 5368 10452 5396 10480
rect 5123 10424 5396 10452
rect 7760 10452 7788 10480
rect 8665 10455 8723 10461
rect 8665 10452 8677 10455
rect 7760 10424 8677 10452
rect 5123 10421 5135 10424
rect 5077 10415 5135 10421
rect 8665 10421 8677 10424
rect 8711 10421 8723 10455
rect 8665 10415 8723 10421
rect 11238 10412 11244 10464
rect 11296 10452 11302 10464
rect 12161 10455 12219 10461
rect 12161 10452 12173 10455
rect 11296 10424 12173 10452
rect 11296 10412 11302 10424
rect 12161 10421 12173 10424
rect 12207 10421 12219 10455
rect 12161 10415 12219 10421
rect 14182 10412 14188 10464
rect 14240 10452 14246 10464
rect 17037 10455 17095 10461
rect 17037 10452 17049 10455
rect 14240 10424 17049 10452
rect 14240 10412 14246 10424
rect 17037 10421 17049 10424
rect 17083 10421 17095 10455
rect 17037 10415 17095 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2041 10251 2099 10257
rect 2041 10217 2053 10251
rect 2087 10248 2099 10251
rect 2130 10248 2136 10260
rect 2087 10220 2136 10248
rect 2087 10217 2099 10220
rect 2041 10211 2099 10217
rect 2130 10208 2136 10220
rect 2188 10208 2194 10260
rect 5031 10251 5089 10257
rect 5031 10217 5043 10251
rect 5077 10248 5089 10251
rect 9122 10248 9128 10260
rect 5077 10220 9128 10248
rect 5077 10217 5089 10220
rect 5031 10211 5089 10217
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 9309 10251 9367 10257
rect 9309 10217 9321 10251
rect 9355 10248 9367 10251
rect 9582 10248 9588 10260
rect 9355 10220 9588 10248
rect 9355 10217 9367 10220
rect 9309 10211 9367 10217
rect 9582 10208 9588 10220
rect 9640 10208 9646 10260
rect 11238 10208 11244 10260
rect 11296 10248 11302 10260
rect 11333 10251 11391 10257
rect 11333 10248 11345 10251
rect 11296 10220 11345 10248
rect 11296 10208 11302 10220
rect 11333 10217 11345 10220
rect 11379 10217 11391 10251
rect 11333 10211 11391 10217
rect 12437 10251 12495 10257
rect 12437 10217 12449 10251
rect 12483 10248 12495 10251
rect 12710 10248 12716 10260
rect 12483 10220 12716 10248
rect 12483 10217 12495 10220
rect 12437 10211 12495 10217
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 12802 10208 12808 10260
rect 12860 10248 12866 10260
rect 13081 10251 13139 10257
rect 13081 10248 13093 10251
rect 12860 10220 13093 10248
rect 12860 10208 12866 10220
rect 13081 10217 13093 10220
rect 13127 10217 13139 10251
rect 13538 10248 13544 10260
rect 13499 10220 13544 10248
rect 13081 10211 13139 10217
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 13630 10208 13636 10260
rect 13688 10248 13694 10260
rect 13725 10251 13783 10257
rect 13725 10248 13737 10251
rect 13688 10220 13737 10248
rect 13688 10208 13694 10220
rect 13725 10217 13737 10220
rect 13771 10217 13783 10251
rect 13725 10211 13783 10217
rect 14826 10208 14832 10260
rect 14884 10248 14890 10260
rect 16439 10251 16497 10257
rect 16439 10248 16451 10251
rect 14884 10220 16451 10248
rect 14884 10208 14890 10220
rect 16439 10217 16451 10220
rect 16485 10217 16497 10251
rect 16439 10211 16497 10217
rect 2866 10180 2872 10192
rect 2827 10152 2872 10180
rect 2866 10140 2872 10152
rect 2924 10140 2930 10192
rect 5994 10180 6000 10192
rect 5955 10152 6000 10180
rect 5994 10140 6000 10152
rect 6052 10140 6058 10192
rect 6089 10183 6147 10189
rect 6089 10149 6101 10183
rect 6135 10180 6147 10183
rect 6270 10180 6276 10192
rect 6135 10152 6276 10180
rect 6135 10149 6147 10152
rect 6089 10143 6147 10149
rect 6270 10140 6276 10152
rect 6328 10180 6334 10192
rect 6730 10180 6736 10192
rect 6328 10152 6736 10180
rect 6328 10140 6334 10152
rect 6730 10140 6736 10152
rect 6788 10140 6794 10192
rect 7745 10183 7803 10189
rect 7745 10149 7757 10183
rect 7791 10180 7803 10183
rect 7834 10180 7840 10192
rect 7791 10152 7840 10180
rect 7791 10149 7803 10152
rect 7745 10143 7803 10149
rect 7834 10140 7840 10152
rect 7892 10140 7898 10192
rect 8202 10180 8208 10192
rect 8163 10152 8208 10180
rect 8202 10140 8208 10152
rect 8260 10140 8266 10192
rect 8757 10183 8815 10189
rect 8757 10149 8769 10183
rect 8803 10180 8815 10183
rect 8938 10180 8944 10192
rect 8803 10152 8944 10180
rect 8803 10149 8815 10152
rect 8757 10143 8815 10149
rect 8938 10140 8944 10152
rect 8996 10180 9002 10192
rect 9398 10180 9404 10192
rect 8996 10152 9404 10180
rect 8996 10140 9002 10152
rect 9398 10140 9404 10152
rect 9456 10140 9462 10192
rect 9858 10180 9864 10192
rect 9819 10152 9864 10180
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 14274 10140 14280 10192
rect 14332 10180 14338 10192
rect 15427 10183 15485 10189
rect 15427 10180 15439 10183
rect 14332 10152 15439 10180
rect 14332 10140 14338 10152
rect 15427 10149 15439 10152
rect 15473 10149 15485 10183
rect 15427 10143 15485 10149
rect 1670 10072 1676 10124
rect 1728 10112 1734 10124
rect 2130 10112 2136 10124
rect 1728 10084 2136 10112
rect 1728 10072 1734 10084
rect 2130 10072 2136 10084
rect 2188 10112 2194 10124
rect 2225 10115 2283 10121
rect 2225 10112 2237 10115
rect 2188 10084 2237 10112
rect 2188 10072 2194 10084
rect 2225 10081 2237 10084
rect 2271 10081 2283 10115
rect 11514 10112 11520 10124
rect 11475 10084 11520 10112
rect 2225 10075 2283 10081
rect 11514 10072 11520 10084
rect 11572 10072 11578 10124
rect 11793 10115 11851 10121
rect 11793 10081 11805 10115
rect 11839 10081 11851 10115
rect 11793 10075 11851 10081
rect 12805 10115 12863 10121
rect 12805 10081 12817 10115
rect 12851 10112 12863 10115
rect 13078 10112 13084 10124
rect 12851 10084 13084 10112
rect 12851 10081 12863 10084
rect 12805 10075 12863 10081
rect 5534 10004 5540 10056
rect 5592 10044 5598 10056
rect 6273 10047 6331 10053
rect 6273 10044 6285 10047
rect 5592 10016 6285 10044
rect 5592 10004 5598 10016
rect 6273 10013 6285 10016
rect 6319 10013 6331 10047
rect 6273 10007 6331 10013
rect 7558 10004 7564 10056
rect 7616 10044 7622 10056
rect 8113 10047 8171 10053
rect 8113 10044 8125 10047
rect 7616 10016 8125 10044
rect 7616 10004 7622 10016
rect 8113 10013 8125 10016
rect 8159 10013 8171 10047
rect 9766 10044 9772 10056
rect 9727 10016 9772 10044
rect 8113 10007 8171 10013
rect 9766 10004 9772 10016
rect 9824 10004 9830 10056
rect 10042 10044 10048 10056
rect 10003 10016 10048 10044
rect 10042 10004 10048 10016
rect 10100 10004 10106 10056
rect 11698 10004 11704 10056
rect 11756 10044 11762 10056
rect 11808 10044 11836 10075
rect 13078 10072 13084 10084
rect 13136 10072 13142 10124
rect 13538 10072 13544 10124
rect 13596 10112 13602 10124
rect 13633 10115 13691 10121
rect 13633 10112 13645 10115
rect 13596 10084 13645 10112
rect 13596 10072 13602 10084
rect 13633 10081 13645 10084
rect 13679 10081 13691 10115
rect 14090 10112 14096 10124
rect 14051 10084 14096 10112
rect 13633 10075 13691 10081
rect 14090 10072 14096 10084
rect 14148 10072 14154 10124
rect 15340 10115 15398 10121
rect 15340 10081 15352 10115
rect 15386 10112 15398 10115
rect 15562 10112 15568 10124
rect 15386 10084 15568 10112
rect 15386 10081 15398 10084
rect 15340 10075 15398 10081
rect 15562 10072 15568 10084
rect 15620 10072 15626 10124
rect 16368 10115 16426 10121
rect 16368 10081 16380 10115
rect 16414 10112 16426 10115
rect 16850 10112 16856 10124
rect 16414 10084 16856 10112
rect 16414 10081 16426 10084
rect 16368 10075 16426 10081
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 17218 10072 17224 10124
rect 17276 10112 17282 10124
rect 17313 10115 17371 10121
rect 17313 10112 17325 10115
rect 17276 10084 17325 10112
rect 17276 10072 17282 10084
rect 17313 10081 17325 10084
rect 17359 10081 17371 10115
rect 17313 10075 17371 10081
rect 11756 10016 13814 10044
rect 11756 10004 11762 10016
rect 4062 9936 4068 9988
rect 4120 9976 4126 9988
rect 5258 9976 5264 9988
rect 4120 9948 5264 9976
rect 4120 9936 4126 9948
rect 5258 9936 5264 9948
rect 5316 9976 5322 9988
rect 5353 9979 5411 9985
rect 5353 9976 5365 9979
rect 5316 9948 5365 9976
rect 5316 9936 5322 9948
rect 5353 9945 5365 9948
rect 5399 9945 5411 9979
rect 13786 9976 13814 10016
rect 17310 9976 17316 9988
rect 13786 9948 17316 9976
rect 5353 9939 5411 9945
rect 17310 9936 17316 9948
rect 17368 9936 17374 9988
rect 4338 9868 4344 9920
rect 4396 9908 4402 9920
rect 4801 9911 4859 9917
rect 4801 9908 4813 9911
rect 4396 9880 4813 9908
rect 4396 9868 4402 9880
rect 4801 9877 4813 9880
rect 4847 9908 4859 9911
rect 4890 9908 4896 9920
rect 4847 9880 4896 9908
rect 4847 9877 4859 9880
rect 4801 9871 4859 9877
rect 4890 9868 4896 9880
rect 4948 9868 4954 9920
rect 10134 9868 10140 9920
rect 10192 9908 10198 9920
rect 10781 9911 10839 9917
rect 10781 9908 10793 9911
rect 10192 9880 10793 9908
rect 10192 9868 10198 9880
rect 10781 9877 10793 9880
rect 10827 9877 10839 9911
rect 10781 9871 10839 9877
rect 13722 9868 13728 9920
rect 13780 9908 13786 9920
rect 14645 9911 14703 9917
rect 14645 9908 14657 9911
rect 13780 9880 14657 9908
rect 13780 9868 13786 9880
rect 14645 9877 14657 9880
rect 14691 9877 14703 9911
rect 17494 9908 17500 9920
rect 17455 9880 17500 9908
rect 14645 9871 14703 9877
rect 17494 9868 17500 9880
rect 17552 9868 17558 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 2130 9704 2136 9716
rect 2091 9676 2136 9704
rect 2130 9664 2136 9676
rect 2188 9664 2194 9716
rect 2363 9707 2421 9713
rect 2363 9673 2375 9707
rect 2409 9704 2421 9707
rect 2590 9704 2596 9716
rect 2409 9676 2596 9704
rect 2409 9673 2421 9676
rect 2363 9667 2421 9673
rect 2590 9664 2596 9676
rect 2648 9664 2654 9716
rect 3418 9664 3424 9716
rect 3476 9704 3482 9716
rect 3513 9707 3571 9713
rect 3513 9704 3525 9707
rect 3476 9676 3525 9704
rect 3476 9664 3482 9676
rect 3513 9673 3525 9676
rect 3559 9673 3571 9707
rect 6270 9704 6276 9716
rect 6231 9676 6276 9704
rect 3513 9667 3571 9673
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 7193 9707 7251 9713
rect 7193 9673 7205 9707
rect 7239 9704 7251 9707
rect 8202 9704 8208 9716
rect 7239 9676 8208 9704
rect 7239 9673 7251 9676
rect 7193 9667 7251 9673
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 10686 9704 10692 9716
rect 10647 9676 10692 9704
rect 10686 9664 10692 9676
rect 10744 9664 10750 9716
rect 11054 9664 11060 9716
rect 11112 9704 11118 9716
rect 13538 9704 13544 9716
rect 11112 9676 13544 9704
rect 11112 9664 11118 9676
rect 13538 9664 13544 9676
rect 13596 9704 13602 9716
rect 13633 9707 13691 9713
rect 13633 9704 13645 9707
rect 13596 9676 13645 9704
rect 13596 9664 13602 9676
rect 13633 9673 13645 9676
rect 13679 9673 13691 9707
rect 13633 9667 13691 9673
rect 17218 9664 17224 9716
rect 17276 9704 17282 9716
rect 17313 9707 17371 9713
rect 17313 9704 17325 9707
rect 17276 9676 17325 9704
rect 17276 9664 17282 9676
rect 17313 9673 17325 9676
rect 17359 9673 17371 9707
rect 17313 9667 17371 9673
rect 3789 9639 3847 9645
rect 3789 9605 3801 9639
rect 3835 9636 3847 9639
rect 5534 9636 5540 9648
rect 3835 9608 5540 9636
rect 3835 9605 3847 9608
rect 3789 9599 3847 9605
rect 2292 9503 2350 9509
rect 2292 9469 2304 9503
rect 2338 9500 2350 9503
rect 3304 9503 3362 9509
rect 2338 9472 2820 9500
rect 2338 9469 2350 9472
rect 2292 9463 2350 9469
rect 2792 9373 2820 9472
rect 3304 9469 3316 9503
rect 3350 9500 3362 9503
rect 3804 9500 3832 9599
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 5994 9596 6000 9648
rect 6052 9636 6058 9648
rect 6362 9636 6368 9648
rect 6052 9608 6368 9636
rect 6052 9596 6058 9608
rect 6362 9596 6368 9608
rect 6420 9636 6426 9648
rect 6549 9639 6607 9645
rect 6549 9636 6561 9639
rect 6420 9608 6561 9636
rect 6420 9596 6426 9608
rect 6549 9605 6561 9608
rect 6595 9605 6607 9639
rect 6549 9599 6607 9605
rect 7837 9639 7895 9645
rect 7837 9605 7849 9639
rect 7883 9636 7895 9639
rect 8018 9636 8024 9648
rect 7883 9608 8024 9636
rect 7883 9605 7895 9608
rect 7837 9599 7895 9605
rect 3350 9472 3832 9500
rect 3350 9469 3362 9472
rect 3304 9463 3362 9469
rect 3970 9460 3976 9512
rect 4028 9500 4034 9512
rect 4617 9503 4675 9509
rect 4617 9500 4629 9503
rect 4028 9472 4629 9500
rect 4028 9460 4034 9472
rect 4617 9469 4629 9472
rect 4663 9500 4675 9503
rect 5261 9503 5319 9509
rect 5261 9500 5273 9503
rect 4663 9472 5273 9500
rect 4663 9469 4675 9472
rect 4617 9463 4675 9469
rect 5261 9469 5273 9472
rect 5307 9469 5319 9503
rect 5261 9463 5319 9469
rect 7336 9503 7394 9509
rect 7336 9469 7348 9503
rect 7382 9500 7394 9503
rect 7852 9500 7880 9599
rect 8018 9596 8024 9608
rect 8076 9596 8082 9648
rect 8938 9636 8944 9648
rect 8899 9608 8944 9636
rect 8938 9596 8944 9608
rect 8996 9596 9002 9648
rect 11514 9596 11520 9648
rect 11572 9636 11578 9648
rect 11793 9639 11851 9645
rect 11793 9636 11805 9639
rect 11572 9608 11805 9636
rect 11572 9596 11578 9608
rect 11793 9605 11805 9608
rect 11839 9636 11851 9639
rect 12618 9636 12624 9648
rect 11839 9608 12624 9636
rect 11839 9605 11851 9608
rect 11793 9599 11851 9605
rect 12618 9596 12624 9608
rect 12676 9596 12682 9648
rect 7382 9472 7880 9500
rect 7382 9469 7394 9472
rect 7336 9463 7394 9469
rect 10686 9460 10692 9512
rect 10744 9500 10750 9512
rect 10781 9503 10839 9509
rect 10781 9500 10793 9503
rect 10744 9472 10793 9500
rect 10744 9460 10750 9472
rect 10781 9469 10793 9472
rect 10827 9469 10839 9503
rect 10781 9463 10839 9469
rect 11241 9503 11299 9509
rect 11241 9469 11253 9503
rect 11287 9469 11299 9503
rect 11241 9463 11299 9469
rect 5902 9432 5908 9444
rect 5863 9404 5908 9432
rect 5902 9392 5908 9404
rect 5960 9392 5966 9444
rect 7423 9435 7481 9441
rect 7423 9401 7435 9435
rect 7469 9432 7481 9435
rect 8202 9432 8208 9444
rect 7469 9404 8208 9432
rect 7469 9401 7481 9404
rect 7423 9395 7481 9401
rect 8202 9392 8208 9404
rect 8260 9392 8266 9444
rect 8386 9432 8392 9444
rect 8347 9404 8392 9432
rect 8386 9392 8392 9404
rect 8444 9392 8450 9444
rect 8481 9435 8539 9441
rect 8481 9401 8493 9435
rect 8527 9432 8539 9435
rect 8754 9432 8760 9444
rect 8527 9404 8760 9432
rect 8527 9401 8539 9404
rect 8481 9395 8539 9401
rect 2777 9367 2835 9373
rect 2777 9333 2789 9367
rect 2823 9364 2835 9367
rect 3142 9364 3148 9376
rect 2823 9336 3148 9364
rect 2823 9333 2835 9336
rect 2777 9327 2835 9333
rect 3142 9324 3148 9336
rect 3200 9324 3206 9376
rect 4890 9364 4896 9376
rect 4851 9336 4896 9364
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 8113 9367 8171 9373
rect 8113 9333 8125 9367
rect 8159 9364 8171 9367
rect 8496 9364 8524 9395
rect 8754 9392 8760 9404
rect 8812 9432 8818 9444
rect 9585 9435 9643 9441
rect 9585 9432 9597 9435
rect 8812 9404 9597 9432
rect 8812 9392 8818 9404
rect 9585 9401 9597 9404
rect 9631 9432 9643 9435
rect 9858 9432 9864 9444
rect 9631 9404 9864 9432
rect 9631 9401 9643 9404
rect 9585 9395 9643 9401
rect 9858 9392 9864 9404
rect 9916 9392 9922 9444
rect 11256 9432 11284 9463
rect 13722 9460 13728 9512
rect 13780 9500 13786 9512
rect 14369 9503 14427 9509
rect 14369 9500 14381 9503
rect 13780 9472 14381 9500
rect 13780 9460 13786 9472
rect 14369 9469 14381 9472
rect 14415 9469 14427 9503
rect 14369 9463 14427 9469
rect 15746 9460 15752 9512
rect 15804 9500 15810 9512
rect 16152 9503 16210 9509
rect 16152 9500 16164 9503
rect 15804 9472 16164 9500
rect 15804 9460 15810 9472
rect 16152 9469 16164 9472
rect 16198 9500 16210 9503
rect 16945 9503 17003 9509
rect 16945 9500 16957 9503
rect 16198 9472 16957 9500
rect 16198 9469 16210 9472
rect 16152 9463 16210 9469
rect 16945 9469 16957 9472
rect 16991 9469 17003 9503
rect 16945 9463 17003 9469
rect 17034 9460 17040 9512
rect 17092 9500 17098 9512
rect 18084 9503 18142 9509
rect 18084 9500 18096 9503
rect 17092 9472 18096 9500
rect 17092 9460 17098 9472
rect 18084 9469 18096 9472
rect 18130 9500 18142 9503
rect 18509 9503 18567 9509
rect 18509 9500 18521 9503
rect 18130 9472 18521 9500
rect 18130 9469 18142 9472
rect 18084 9463 18142 9469
rect 18509 9469 18521 9472
rect 18555 9469 18567 9503
rect 18509 9463 18567 9469
rect 11514 9432 11520 9444
rect 10152 9404 11284 9432
rect 11475 9404 11520 9432
rect 10152 9376 10180 9404
rect 11514 9392 11520 9404
rect 11572 9392 11578 9444
rect 12526 9432 12532 9444
rect 12487 9404 12532 9432
rect 12526 9392 12532 9404
rect 12584 9392 12590 9444
rect 12621 9435 12679 9441
rect 12621 9401 12633 9435
rect 12667 9401 12679 9435
rect 13170 9432 13176 9444
rect 13131 9404 13176 9432
rect 12621 9395 12679 9401
rect 8159 9336 8524 9364
rect 10045 9367 10103 9373
rect 8159 9333 8171 9336
rect 8113 9327 8171 9333
rect 10045 9333 10057 9367
rect 10091 9364 10103 9367
rect 10134 9364 10140 9376
rect 10091 9336 10140 9364
rect 10091 9333 10103 9336
rect 10045 9327 10103 9333
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 12253 9367 12311 9373
rect 12253 9333 12265 9367
rect 12299 9364 12311 9367
rect 12434 9364 12440 9376
rect 12299 9336 12440 9364
rect 12299 9333 12311 9336
rect 12253 9327 12311 9333
rect 12434 9324 12440 9336
rect 12492 9364 12498 9376
rect 12636 9364 12664 9395
rect 13170 9392 13176 9404
rect 13228 9392 13234 9444
rect 14690 9435 14748 9441
rect 14690 9432 14702 9435
rect 14292 9404 14702 9432
rect 14292 9376 14320 9404
rect 14690 9401 14702 9404
rect 14736 9401 14748 9435
rect 14690 9395 14748 9401
rect 14918 9392 14924 9444
rect 14976 9432 14982 9444
rect 16255 9435 16313 9441
rect 16255 9432 16267 9435
rect 14976 9404 16267 9432
rect 14976 9392 14982 9404
rect 16255 9401 16267 9404
rect 16301 9401 16313 9435
rect 16255 9395 16313 9401
rect 14274 9364 14280 9376
rect 12492 9336 12664 9364
rect 14235 9336 14280 9364
rect 12492 9324 12498 9336
rect 14274 9324 14280 9336
rect 14332 9324 14338 9376
rect 15289 9367 15347 9373
rect 15289 9333 15301 9367
rect 15335 9364 15347 9367
rect 15378 9364 15384 9376
rect 15335 9336 15384 9364
rect 15335 9333 15347 9336
rect 15289 9327 15347 9333
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 15562 9364 15568 9376
rect 15523 9336 15568 9364
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 16669 9367 16727 9373
rect 16669 9333 16681 9367
rect 16715 9364 16727 9367
rect 16850 9364 16856 9376
rect 16715 9336 16856 9364
rect 16715 9333 16727 9336
rect 16669 9327 16727 9333
rect 16850 9324 16856 9336
rect 16908 9324 16914 9376
rect 17034 9324 17040 9376
rect 17092 9364 17098 9376
rect 18187 9367 18245 9373
rect 18187 9364 18199 9367
rect 17092 9336 18199 9364
rect 17092 9324 17098 9336
rect 18187 9333 18199 9336
rect 18233 9333 18245 9367
rect 18187 9327 18245 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1811 9163 1869 9169
rect 1811 9129 1823 9163
rect 1857 9160 1869 9163
rect 2038 9160 2044 9172
rect 1857 9132 2044 9160
rect 1857 9129 1869 9132
rect 1811 9123 1869 9129
rect 2038 9120 2044 9132
rect 2096 9120 2102 9172
rect 2406 9120 2412 9172
rect 2464 9160 2470 9172
rect 2823 9163 2881 9169
rect 2823 9160 2835 9163
rect 2464 9132 2835 9160
rect 2464 9120 2470 9132
rect 2823 9129 2835 9132
rect 2869 9129 2881 9163
rect 2823 9123 2881 9129
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 5123 9163 5181 9169
rect 5123 9160 5135 9163
rect 4120 9132 5135 9160
rect 4120 9120 4126 9132
rect 5123 9129 5135 9132
rect 5169 9129 5181 9163
rect 7558 9160 7564 9172
rect 7519 9132 7564 9160
rect 5123 9123 5181 9129
rect 7558 9120 7564 9132
rect 7616 9120 7622 9172
rect 8110 9160 8116 9172
rect 8071 9132 8116 9160
rect 8110 9120 8116 9132
rect 8168 9120 8174 9172
rect 8202 9120 8208 9172
rect 8260 9160 8266 9172
rect 9401 9163 9459 9169
rect 9401 9160 9413 9163
rect 8260 9132 9413 9160
rect 8260 9120 8266 9132
rect 9401 9129 9413 9132
rect 9447 9160 9459 9163
rect 9766 9160 9772 9172
rect 9447 9132 9772 9160
rect 9447 9129 9459 9132
rect 9401 9123 9459 9129
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 11333 9163 11391 9169
rect 11333 9129 11345 9163
rect 11379 9160 11391 9163
rect 11698 9160 11704 9172
rect 11379 9132 11704 9160
rect 11379 9129 11391 9132
rect 11333 9123 11391 9129
rect 11698 9120 11704 9132
rect 11756 9120 11762 9172
rect 12526 9120 12532 9172
rect 12584 9160 12590 9172
rect 13081 9163 13139 9169
rect 13081 9160 13093 9163
rect 12584 9132 13093 9160
rect 12584 9120 12590 9132
rect 13081 9129 13093 9132
rect 13127 9129 13139 9163
rect 13722 9160 13728 9172
rect 13683 9132 13728 9160
rect 13081 9123 13139 9129
rect 1394 9052 1400 9104
rect 1452 9092 1458 9104
rect 1452 9064 2763 9092
rect 1452 9052 1458 9064
rect 1740 9027 1798 9033
rect 1740 8993 1752 9027
rect 1786 9024 1798 9027
rect 2590 9024 2596 9036
rect 1786 8996 2596 9024
rect 1786 8993 1798 8996
rect 1740 8987 1798 8993
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 2735 9033 2763 9064
rect 5902 9052 5908 9104
rect 5960 9092 5966 9104
rect 6181 9095 6239 9101
rect 6181 9092 6193 9095
rect 5960 9064 6193 9092
rect 5960 9052 5966 9064
rect 6181 9061 6193 9064
rect 6227 9092 6239 9095
rect 6546 9092 6552 9104
rect 6227 9064 6552 9092
rect 6227 9061 6239 9064
rect 6181 9055 6239 9061
rect 6546 9052 6552 9064
rect 6604 9052 6610 9104
rect 11054 9092 11060 9104
rect 8312 9064 11060 9092
rect 2720 9027 2778 9033
rect 2720 8993 2732 9027
rect 2766 9024 2778 9027
rect 2866 9024 2872 9036
rect 2766 8996 2872 9024
rect 2766 8993 2778 8996
rect 2720 8987 2778 8993
rect 2866 8984 2872 8996
rect 2924 8984 2930 9036
rect 5052 9027 5110 9033
rect 5052 8993 5064 9027
rect 5098 9024 5110 9027
rect 5166 9024 5172 9036
rect 5098 8996 5172 9024
rect 5098 8993 5110 8996
rect 5052 8987 5110 8993
rect 5166 8984 5172 8996
rect 5224 8984 5230 9036
rect 8312 9033 8340 9064
rect 8297 9027 8355 9033
rect 8297 8993 8309 9027
rect 8343 8993 8355 9027
rect 8297 8987 8355 8993
rect 8573 9027 8631 9033
rect 8573 8993 8585 9027
rect 8619 9024 8631 9027
rect 9490 9024 9496 9036
rect 8619 8996 9496 9024
rect 8619 8993 8631 8996
rect 8573 8987 8631 8993
rect 5534 8916 5540 8968
rect 5592 8956 5598 8968
rect 6089 8959 6147 8965
rect 6089 8956 6101 8959
rect 5592 8928 6101 8956
rect 5592 8916 5598 8928
rect 6089 8925 6101 8928
rect 6135 8925 6147 8959
rect 6362 8956 6368 8968
rect 6323 8928 6368 8956
rect 6089 8919 6147 8925
rect 6362 8916 6368 8928
rect 6420 8916 6426 8968
rect 6454 8916 6460 8968
rect 6512 8956 6518 8968
rect 7929 8959 7987 8965
rect 7929 8956 7941 8959
rect 6512 8928 7941 8956
rect 6512 8916 6518 8928
rect 7929 8925 7941 8928
rect 7975 8956 7987 8959
rect 8588 8956 8616 8987
rect 9490 8984 9496 8996
rect 9548 8984 9554 9036
rect 10060 9033 10088 9064
rect 11054 9052 11060 9064
rect 11112 9052 11118 9104
rect 11882 9101 11888 9104
rect 11879 9092 11888 9101
rect 11795 9064 11888 9092
rect 11879 9055 11888 9064
rect 11940 9092 11946 9104
rect 12250 9092 12256 9104
rect 11940 9064 12256 9092
rect 11882 9052 11888 9055
rect 11940 9052 11946 9064
rect 12250 9052 12256 9064
rect 12308 9052 12314 9104
rect 10045 9027 10103 9033
rect 10045 8993 10057 9027
rect 10091 8993 10103 9027
rect 10045 8987 10103 8993
rect 10134 8984 10140 9036
rect 10192 9024 10198 9036
rect 10413 9027 10471 9033
rect 10413 9024 10425 9027
rect 10192 8996 10425 9024
rect 10192 8984 10198 8996
rect 10413 8993 10425 8996
rect 10459 8993 10471 9027
rect 11514 9024 11520 9036
rect 11475 8996 11520 9024
rect 10413 8987 10471 8993
rect 11514 8984 11520 8996
rect 11572 8984 11578 9036
rect 10686 8956 10692 8968
rect 7975 8928 8616 8956
rect 10647 8928 10692 8956
rect 7975 8925 7987 8928
rect 7929 8919 7987 8925
rect 10686 8916 10692 8928
rect 10744 8916 10750 8968
rect 13096 8956 13124 9123
rect 13722 9120 13728 9132
rect 13780 9120 13786 9172
rect 15378 9052 15384 9104
rect 15436 9092 15442 9104
rect 15473 9095 15531 9101
rect 15473 9092 15485 9095
rect 15436 9064 15485 9092
rect 15436 9052 15442 9064
rect 15473 9061 15485 9064
rect 15519 9092 15531 9095
rect 15746 9092 15752 9104
rect 15519 9064 15752 9092
rect 15519 9061 15531 9064
rect 15473 9055 15531 9061
rect 15746 9052 15752 9064
rect 15804 9052 15810 9104
rect 13538 9024 13544 9036
rect 13499 8996 13544 9024
rect 13538 8984 13544 8996
rect 13596 8984 13602 9036
rect 14001 9027 14059 9033
rect 14001 8993 14013 9027
rect 14047 9024 14059 9027
rect 14090 9024 14096 9036
rect 14047 8996 14096 9024
rect 14047 8993 14059 8996
rect 14001 8987 14059 8993
rect 14090 8984 14096 8996
rect 14148 9024 14154 9036
rect 14550 9024 14556 9036
rect 14148 8996 14556 9024
rect 14148 8984 14154 8996
rect 14550 8984 14556 8996
rect 14608 8984 14614 9036
rect 16850 9024 16856 9036
rect 16811 8996 16856 9024
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 14918 8956 14924 8968
rect 13096 8928 14924 8956
rect 14918 8916 14924 8928
rect 14976 8916 14982 8968
rect 15105 8959 15163 8965
rect 15105 8925 15117 8959
rect 15151 8956 15163 8959
rect 15381 8959 15439 8965
rect 15381 8956 15393 8959
rect 15151 8928 15393 8956
rect 15151 8925 15163 8928
rect 15105 8919 15163 8925
rect 15381 8925 15393 8928
rect 15427 8956 15439 8959
rect 17034 8956 17040 8968
rect 15427 8928 17040 8956
rect 15427 8925 15439 8928
rect 15381 8919 15439 8925
rect 17034 8916 17040 8928
rect 17092 8916 17098 8968
rect 842 8848 848 8900
rect 900 8888 906 8900
rect 4430 8888 4436 8900
rect 900 8860 4436 8888
rect 900 8848 906 8860
rect 4430 8848 4436 8860
rect 4488 8848 4494 8900
rect 5994 8848 6000 8900
rect 6052 8888 6058 8900
rect 11146 8888 11152 8900
rect 6052 8860 11152 8888
rect 6052 8848 6058 8860
rect 11146 8848 11152 8860
rect 11204 8848 11210 8900
rect 12526 8848 12532 8900
rect 12584 8888 12590 8900
rect 12805 8891 12863 8897
rect 12805 8888 12817 8891
rect 12584 8860 12817 8888
rect 12584 8848 12590 8860
rect 12805 8857 12817 8860
rect 12851 8888 12863 8891
rect 15930 8888 15936 8900
rect 12851 8860 15148 8888
rect 15891 8860 15936 8888
rect 12851 8857 12863 8860
rect 12805 8851 12863 8857
rect 8386 8780 8392 8832
rect 8444 8820 8450 8832
rect 9033 8823 9091 8829
rect 9033 8820 9045 8823
rect 8444 8792 9045 8820
rect 8444 8780 8450 8792
rect 9033 8789 9045 8792
rect 9079 8789 9091 8823
rect 12434 8820 12440 8832
rect 12395 8792 12440 8820
rect 9033 8783 9091 8789
rect 12434 8780 12440 8792
rect 12492 8780 12498 8832
rect 14550 8820 14556 8832
rect 14511 8792 14556 8820
rect 14550 8780 14556 8792
rect 14608 8780 14614 8832
rect 15120 8820 15148 8860
rect 15930 8848 15936 8860
rect 15988 8848 15994 8900
rect 16991 8823 17049 8829
rect 16991 8820 17003 8823
rect 15120 8792 17003 8820
rect 16991 8789 17003 8792
rect 17037 8789 17049 8823
rect 16991 8783 17049 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1578 8576 1584 8628
rect 1636 8616 1642 8628
rect 1673 8619 1731 8625
rect 1673 8616 1685 8619
rect 1636 8588 1685 8616
rect 1636 8576 1642 8588
rect 1673 8585 1685 8588
rect 1719 8585 1731 8619
rect 1673 8579 1731 8585
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 2547 8619 2605 8625
rect 2547 8616 2559 8619
rect 2372 8588 2559 8616
rect 2372 8576 2378 8588
rect 2547 8585 2559 8588
rect 2593 8585 2605 8619
rect 2866 8616 2872 8628
rect 2827 8588 2872 8616
rect 2547 8579 2605 8585
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 3326 8616 3332 8628
rect 3287 8588 3332 8616
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 5077 8619 5135 8625
rect 5077 8585 5089 8619
rect 5123 8616 5135 8619
rect 5166 8616 5172 8628
rect 5123 8588 5172 8616
rect 5123 8585 5135 8588
rect 5077 8579 5135 8585
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 6546 8616 6552 8628
rect 6507 8588 6552 8616
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 7331 8619 7389 8625
rect 7331 8585 7343 8619
rect 7377 8616 7389 8619
rect 7742 8616 7748 8628
rect 7377 8588 7748 8616
rect 7377 8585 7389 8588
rect 7331 8579 7389 8585
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 7926 8576 7932 8628
rect 7984 8616 7990 8628
rect 8021 8619 8079 8625
rect 8021 8616 8033 8619
rect 7984 8588 8033 8616
rect 7984 8576 7990 8588
rect 8021 8585 8033 8588
rect 8067 8585 8079 8619
rect 8021 8579 8079 8585
rect 9493 8619 9551 8625
rect 9493 8585 9505 8619
rect 9539 8616 9551 8619
rect 11054 8616 11060 8628
rect 9539 8588 11060 8616
rect 9539 8585 9551 8588
rect 9493 8579 9551 8585
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 15654 8576 15660 8628
rect 15712 8616 15718 8628
rect 16255 8619 16313 8625
rect 16255 8616 16267 8619
rect 15712 8588 16267 8616
rect 15712 8576 15718 8588
rect 16255 8585 16267 8588
rect 16301 8585 16313 8619
rect 16255 8579 16313 8585
rect 5859 8551 5917 8557
rect 5859 8517 5871 8551
rect 5905 8548 5917 8551
rect 7558 8548 7564 8560
rect 5905 8520 7564 8548
rect 5905 8517 5917 8520
rect 5859 8511 5917 8517
rect 7558 8508 7564 8520
rect 7616 8508 7622 8560
rect 13449 8551 13507 8557
rect 13449 8548 13461 8551
rect 10612 8520 13461 8548
rect 10612 8492 10640 8520
rect 13449 8517 13461 8520
rect 13495 8548 13507 8551
rect 13538 8548 13544 8560
rect 13495 8520 13544 8548
rect 13495 8517 13507 8520
rect 13449 8511 13507 8517
rect 13538 8508 13544 8520
rect 13596 8508 13602 8560
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8480 2375 8483
rect 2682 8480 2688 8492
rect 2363 8452 2688 8480
rect 2363 8449 2375 8452
rect 2317 8443 2375 8449
rect 2682 8440 2688 8452
rect 2740 8440 2746 8492
rect 8110 8440 8116 8492
rect 8168 8480 8174 8492
rect 8205 8483 8263 8489
rect 8205 8480 8217 8483
rect 8168 8452 8217 8480
rect 8168 8440 8174 8452
rect 8205 8449 8217 8452
rect 8251 8449 8263 8483
rect 8205 8443 8263 8449
rect 9861 8483 9919 8489
rect 9861 8449 9873 8483
rect 9907 8480 9919 8483
rect 10594 8480 10600 8492
rect 9907 8452 10600 8480
rect 9907 8449 9919 8452
rect 9861 8443 9919 8449
rect 14 8372 20 8424
rect 72 8412 78 8424
rect 1432 8415 1490 8421
rect 1432 8412 1444 8415
rect 72 8384 1444 8412
rect 72 8372 78 8384
rect 1432 8381 1444 8384
rect 1478 8412 1490 8415
rect 1857 8415 1915 8421
rect 1857 8412 1869 8415
rect 1478 8384 1869 8412
rect 1478 8381 1490 8384
rect 1432 8375 1490 8381
rect 1857 8381 1869 8384
rect 1903 8412 1915 8415
rect 2222 8412 2228 8424
rect 1903 8384 2228 8412
rect 1903 8381 1915 8384
rect 1857 8375 1915 8381
rect 2222 8372 2228 8384
rect 2280 8372 2286 8424
rect 2476 8415 2534 8421
rect 2476 8381 2488 8415
rect 2522 8412 2534 8415
rect 3326 8412 3332 8424
rect 2522 8384 3332 8412
rect 2522 8381 2534 8384
rect 2476 8375 2534 8381
rect 3326 8372 3332 8384
rect 3384 8372 3390 8424
rect 5788 8415 5846 8421
rect 5788 8381 5800 8415
rect 5834 8412 5846 8415
rect 6178 8412 6184 8424
rect 5834 8384 6184 8412
rect 5834 8381 5846 8384
rect 5788 8375 5846 8381
rect 6178 8372 6184 8384
rect 6236 8372 6242 8424
rect 6822 8372 6828 8424
rect 6880 8412 6886 8424
rect 10244 8421 10272 8452
rect 10594 8440 10600 8452
rect 10652 8440 10658 8492
rect 11609 8483 11667 8489
rect 11609 8449 11621 8483
rect 11655 8480 11667 8483
rect 12250 8480 12256 8492
rect 11655 8452 12256 8480
rect 11655 8449 11667 8452
rect 11609 8443 11667 8449
rect 12250 8440 12256 8452
rect 12308 8440 12314 8492
rect 12526 8480 12532 8492
rect 12487 8452 12532 8480
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 13170 8480 13176 8492
rect 13131 8452 13176 8480
rect 13170 8440 13176 8452
rect 13228 8440 13234 8492
rect 13630 8440 13636 8492
rect 13688 8480 13694 8492
rect 13909 8483 13967 8489
rect 13688 8452 13814 8480
rect 13688 8440 13694 8452
rect 7228 8415 7286 8421
rect 7228 8412 7240 8415
rect 6880 8384 7240 8412
rect 6880 8372 6886 8384
rect 7228 8381 7240 8384
rect 7274 8412 7286 8415
rect 7653 8415 7711 8421
rect 7653 8412 7665 8415
rect 7274 8384 7665 8412
rect 7274 8381 7286 8384
rect 7228 8375 7286 8381
rect 7653 8381 7665 8384
rect 7699 8381 7711 8415
rect 7653 8375 7711 8381
rect 10229 8415 10287 8421
rect 10229 8381 10241 8415
rect 10275 8381 10287 8415
rect 10229 8375 10287 8381
rect 10413 8415 10471 8421
rect 10413 8381 10425 8415
rect 10459 8381 10471 8415
rect 13786 8412 13814 8452
rect 13909 8449 13921 8483
rect 13955 8480 13967 8483
rect 14550 8480 14556 8492
rect 13955 8452 14556 8480
rect 13955 8449 13967 8452
rect 13909 8443 13967 8449
rect 14550 8440 14556 8452
rect 14608 8440 14614 8492
rect 14366 8412 14372 8424
rect 13786 8384 14372 8412
rect 10413 8375 10471 8381
rect 1670 8304 1676 8356
rect 1728 8344 1734 8356
rect 5166 8344 5172 8356
rect 1728 8316 5172 8344
rect 1728 8304 1734 8316
rect 5166 8304 5172 8316
rect 5224 8304 5230 8356
rect 7926 8304 7932 8356
rect 7984 8344 7990 8356
rect 8526 8347 8584 8353
rect 8526 8344 8538 8347
rect 7984 8316 8538 8344
rect 7984 8304 7990 8316
rect 8526 8313 8538 8316
rect 8572 8313 8584 8347
rect 8526 8307 8584 8313
rect 9490 8304 9496 8356
rect 9548 8344 9554 8356
rect 10428 8344 10456 8375
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 16152 8415 16210 8421
rect 16152 8412 16164 8415
rect 15948 8384 16164 8412
rect 9548 8316 10456 8344
rect 12253 8347 12311 8353
rect 9548 8304 9554 8316
rect 12253 8313 12265 8347
rect 12299 8344 12311 8347
rect 12342 8344 12348 8356
rect 12299 8316 12348 8344
rect 12299 8313 12311 8316
rect 12253 8307 12311 8313
rect 12342 8304 12348 8316
rect 12400 8344 12406 8356
rect 12621 8347 12679 8353
rect 12621 8344 12633 8347
rect 12400 8316 12633 8344
rect 12400 8304 12406 8316
rect 12621 8313 12633 8316
rect 12667 8313 12679 8347
rect 12621 8307 12679 8313
rect 14690 8347 14748 8353
rect 14690 8313 14702 8347
rect 14736 8313 14748 8347
rect 14690 8307 14748 8313
rect 5534 8276 5540 8288
rect 5495 8248 5540 8276
rect 5534 8236 5540 8248
rect 5592 8236 5598 8288
rect 9122 8276 9128 8288
rect 9083 8248 9128 8276
rect 9122 8236 9128 8248
rect 9180 8236 9186 8288
rect 10042 8276 10048 8288
rect 10003 8248 10048 8276
rect 10042 8236 10048 8248
rect 10100 8236 10106 8288
rect 14274 8276 14280 8288
rect 14235 8248 14280 8276
rect 14274 8236 14280 8248
rect 14332 8276 14338 8288
rect 14705 8276 14733 8307
rect 14332 8248 14733 8276
rect 15289 8279 15347 8285
rect 14332 8236 14338 8248
rect 15289 8245 15301 8279
rect 15335 8276 15347 8279
rect 15470 8276 15476 8288
rect 15335 8248 15476 8276
rect 15335 8245 15347 8248
rect 15289 8239 15347 8245
rect 15470 8236 15476 8248
rect 15528 8236 15534 8288
rect 15657 8279 15715 8285
rect 15657 8245 15669 8279
rect 15703 8276 15715 8279
rect 15746 8276 15752 8288
rect 15703 8248 15752 8276
rect 15703 8245 15715 8248
rect 15657 8239 15715 8245
rect 15746 8236 15752 8248
rect 15804 8236 15810 8288
rect 15838 8236 15844 8288
rect 15896 8276 15902 8288
rect 15948 8285 15976 8384
rect 16152 8381 16164 8384
rect 16198 8381 16210 8415
rect 16152 8375 16210 8381
rect 15933 8279 15991 8285
rect 15933 8276 15945 8279
rect 15896 8248 15945 8276
rect 15896 8236 15902 8248
rect 15933 8245 15945 8248
rect 15979 8245 15991 8279
rect 16850 8276 16856 8288
rect 16811 8248 16856 8276
rect 15933 8239 15991 8245
rect 16850 8236 16856 8248
rect 16908 8236 16914 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 5997 8075 6055 8081
rect 5997 8041 6009 8075
rect 6043 8072 6055 8075
rect 6454 8072 6460 8084
rect 6043 8044 6460 8072
rect 6043 8041 6055 8044
rect 5997 8035 6055 8041
rect 6454 8032 6460 8044
rect 6512 8032 6518 8084
rect 6963 8075 7021 8081
rect 6963 8041 6975 8075
rect 7009 8072 7021 8075
rect 8386 8072 8392 8084
rect 7009 8044 8392 8072
rect 7009 8041 7021 8044
rect 6963 8035 7021 8041
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 9490 8072 9496 8084
rect 9451 8044 9496 8072
rect 9490 8032 9496 8044
rect 9548 8032 9554 8084
rect 11333 8075 11391 8081
rect 11333 8041 11345 8075
rect 11379 8072 11391 8075
rect 11514 8072 11520 8084
rect 11379 8044 11520 8072
rect 11379 8041 11391 8044
rect 11333 8035 11391 8041
rect 11514 8032 11520 8044
rect 11572 8032 11578 8084
rect 12342 8072 12348 8084
rect 12303 8044 12348 8072
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 12618 8072 12624 8084
rect 12579 8044 12624 8072
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 14366 8032 14372 8084
rect 14424 8072 14430 8084
rect 14829 8075 14887 8081
rect 14829 8072 14841 8075
rect 14424 8044 14841 8072
rect 14424 8032 14430 8044
rect 14829 8041 14841 8044
rect 14875 8041 14887 8075
rect 14829 8035 14887 8041
rect 7926 7964 7932 8016
rect 7984 8004 7990 8016
rect 8158 8007 8216 8013
rect 8158 8004 8170 8007
rect 7984 7976 8170 8004
rect 7984 7964 7990 7976
rect 8158 7973 8170 7976
rect 8204 7973 8216 8007
rect 10042 8004 10048 8016
rect 8158 7967 8216 7973
rect 8496 7976 10048 8004
rect 5813 7939 5871 7945
rect 5813 7905 5825 7939
rect 5859 7936 5871 7939
rect 5994 7936 6000 7948
rect 5859 7908 6000 7936
rect 5859 7905 5871 7908
rect 5813 7899 5871 7905
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 6892 7939 6950 7945
rect 6892 7905 6904 7939
rect 6938 7936 6950 7939
rect 7466 7936 7472 7948
rect 6938 7908 7472 7936
rect 6938 7905 6950 7908
rect 6892 7899 6950 7905
rect 7466 7896 7472 7908
rect 7524 7896 7530 7948
rect 7558 7896 7564 7948
rect 7616 7936 7622 7948
rect 7837 7939 7895 7945
rect 7837 7936 7849 7939
rect 7616 7908 7849 7936
rect 7616 7896 7622 7908
rect 7837 7905 7849 7908
rect 7883 7936 7895 7939
rect 8496 7936 8524 7976
rect 10042 7964 10048 7976
rect 10100 7964 10106 8016
rect 11787 8007 11845 8013
rect 11787 7973 11799 8007
rect 11833 8004 11845 8007
rect 12250 8004 12256 8016
rect 11833 7976 12256 8004
rect 11833 7973 11845 7976
rect 11787 7967 11845 7973
rect 12250 7964 12256 7976
rect 12308 7964 12314 8016
rect 15470 8004 15476 8016
rect 15431 7976 15476 8004
rect 15470 7964 15476 7976
rect 15528 7964 15534 8016
rect 15838 7964 15844 8016
rect 15896 8004 15902 8016
rect 15896 7976 16931 8004
rect 15896 7964 15902 7976
rect 9950 7936 9956 7948
rect 7883 7908 8524 7936
rect 9911 7908 9956 7936
rect 7883 7905 7895 7908
rect 7837 7899 7895 7905
rect 9950 7896 9956 7908
rect 10008 7896 10014 7948
rect 10318 7936 10324 7948
rect 10279 7908 10324 7936
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 10686 7896 10692 7948
rect 10744 7936 10750 7948
rect 11422 7936 11428 7948
rect 10744 7908 11428 7936
rect 10744 7896 10750 7908
rect 11422 7896 11428 7908
rect 11480 7896 11486 7948
rect 13262 7936 13268 7948
rect 13223 7908 13268 7936
rect 13262 7896 13268 7908
rect 13320 7896 13326 7948
rect 13633 7939 13691 7945
rect 13633 7905 13645 7939
rect 13679 7936 13691 7939
rect 14182 7936 14188 7948
rect 13679 7908 14188 7936
rect 13679 7905 13691 7908
rect 13633 7899 13691 7905
rect 8110 7828 8116 7880
rect 8168 7868 8174 7880
rect 9033 7871 9091 7877
rect 9033 7868 9045 7871
rect 8168 7840 9045 7868
rect 8168 7828 8174 7840
rect 9033 7837 9045 7840
rect 9079 7837 9091 7871
rect 9033 7831 9091 7837
rect 10597 7871 10655 7877
rect 10597 7837 10609 7871
rect 10643 7868 10655 7871
rect 11330 7868 11336 7880
rect 10643 7840 11336 7868
rect 10643 7837 10655 7840
rect 10597 7831 10655 7837
rect 11330 7828 11336 7840
rect 11388 7828 11394 7880
rect 13648 7868 13676 7899
rect 14182 7896 14188 7908
rect 14240 7896 14246 7948
rect 16903 7945 16931 7976
rect 16888 7939 16946 7945
rect 16888 7905 16900 7939
rect 16934 7936 16946 7939
rect 17126 7936 17132 7948
rect 16934 7908 17132 7936
rect 16934 7905 16946 7908
rect 16888 7899 16946 7905
rect 17126 7896 17132 7908
rect 17184 7896 17190 7948
rect 13004 7840 13676 7868
rect 10318 7760 10324 7812
rect 10376 7800 10382 7812
rect 13004 7809 13032 7840
rect 13814 7828 13820 7880
rect 13872 7868 13878 7880
rect 15378 7868 15384 7880
rect 13872 7840 13917 7868
rect 15291 7840 15384 7868
rect 13872 7828 13878 7840
rect 15378 7828 15384 7840
rect 15436 7868 15442 7880
rect 16991 7871 17049 7877
rect 16991 7868 17003 7871
rect 15436 7840 17003 7868
rect 15436 7828 15442 7840
rect 16991 7837 17003 7840
rect 17037 7837 17049 7871
rect 16991 7831 17049 7837
rect 12989 7803 13047 7809
rect 12989 7800 13001 7803
rect 10376 7772 13001 7800
rect 10376 7760 10382 7772
rect 12989 7769 13001 7772
rect 13035 7769 13047 7803
rect 15930 7800 15936 7812
rect 15843 7772 15936 7800
rect 12989 7763 13047 7769
rect 15930 7760 15936 7772
rect 15988 7760 15994 7812
rect 7282 7732 7288 7744
rect 7243 7704 7288 7732
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 7742 7732 7748 7744
rect 7703 7704 7748 7732
rect 7742 7692 7748 7704
rect 7800 7732 7806 7744
rect 8757 7735 8815 7741
rect 8757 7732 8769 7735
rect 7800 7704 8769 7732
rect 7800 7692 7806 7704
rect 8757 7701 8769 7704
rect 8803 7701 8815 7735
rect 14550 7732 14556 7744
rect 14511 7704 14556 7732
rect 8757 7695 8815 7701
rect 14550 7692 14556 7704
rect 14608 7692 14614 7744
rect 15948 7732 15976 7760
rect 16393 7735 16451 7741
rect 16393 7732 16405 7735
rect 15948 7704 16405 7732
rect 16393 7701 16405 7704
rect 16439 7732 16451 7735
rect 16482 7732 16488 7744
rect 16439 7704 16488 7732
rect 16439 7701 16451 7704
rect 16393 7695 16451 7701
rect 16482 7692 16488 7704
rect 16540 7692 16546 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 5905 7531 5963 7537
rect 5905 7497 5917 7531
rect 5951 7528 5963 7531
rect 5994 7528 6000 7540
rect 5951 7500 6000 7528
rect 5951 7497 5963 7500
rect 5905 7491 5963 7497
rect 5994 7488 6000 7500
rect 6052 7488 6058 7540
rect 7147 7531 7205 7537
rect 7147 7497 7159 7531
rect 7193 7528 7205 7531
rect 7282 7528 7288 7540
rect 7193 7500 7288 7528
rect 7193 7497 7205 7500
rect 7147 7491 7205 7497
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 9125 7531 9183 7537
rect 9125 7497 9137 7531
rect 9171 7528 9183 7531
rect 10318 7528 10324 7540
rect 9171 7500 10324 7528
rect 9171 7497 9183 7500
rect 9125 7491 9183 7497
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 13262 7488 13268 7540
rect 13320 7528 13326 7540
rect 13449 7531 13507 7537
rect 13449 7528 13461 7531
rect 13320 7500 13461 7528
rect 13320 7488 13326 7500
rect 13449 7497 13461 7500
rect 13495 7497 13507 7531
rect 13449 7491 13507 7497
rect 13909 7531 13967 7537
rect 13909 7497 13921 7531
rect 13955 7528 13967 7531
rect 14182 7528 14188 7540
rect 13955 7500 14188 7528
rect 13955 7497 13967 7500
rect 13909 7491 13967 7497
rect 14182 7488 14188 7500
rect 14240 7488 14246 7540
rect 17126 7528 17132 7540
rect 17087 7500 17132 7528
rect 17126 7488 17132 7500
rect 17184 7488 17190 7540
rect 7300 7392 7328 7488
rect 9950 7420 9956 7472
rect 10008 7460 10014 7472
rect 10597 7463 10655 7469
rect 10597 7460 10609 7463
rect 10008 7432 10609 7460
rect 10008 7420 10014 7432
rect 10597 7429 10609 7432
rect 10643 7460 10655 7463
rect 17034 7460 17040 7472
rect 10643 7432 17040 7460
rect 10643 7429 10655 7432
rect 10597 7423 10655 7429
rect 17034 7420 17040 7432
rect 17092 7420 17098 7472
rect 8113 7395 8171 7401
rect 8113 7392 8125 7395
rect 7300 7364 8125 7392
rect 8113 7361 8125 7364
rect 8159 7361 8171 7395
rect 8113 7355 8171 7361
rect 9490 7352 9496 7404
rect 9548 7392 9554 7404
rect 16117 7395 16175 7401
rect 9548 7364 10088 7392
rect 9548 7352 9554 7364
rect 6178 7284 6184 7336
rect 6236 7324 6242 7336
rect 10060 7333 10088 7364
rect 12636 7364 14412 7392
rect 12636 7336 12664 7364
rect 7044 7327 7102 7333
rect 7044 7324 7056 7327
rect 6236 7296 7056 7324
rect 6236 7284 6242 7296
rect 7044 7293 7056 7296
rect 7090 7324 7102 7327
rect 7837 7327 7895 7333
rect 7837 7324 7849 7327
rect 7090 7296 7849 7324
rect 7090 7293 7102 7296
rect 7044 7287 7102 7293
rect 7837 7293 7849 7296
rect 7883 7293 7895 7327
rect 7837 7287 7895 7293
rect 9861 7327 9919 7333
rect 9861 7293 9873 7327
rect 9907 7293 9919 7327
rect 9861 7287 9919 7293
rect 10045 7327 10103 7333
rect 10045 7293 10057 7327
rect 10091 7324 10103 7327
rect 10965 7327 11023 7333
rect 10965 7324 10977 7327
rect 10091 7296 10977 7324
rect 10091 7293 10103 7296
rect 10045 7287 10103 7293
rect 10965 7293 10977 7296
rect 11011 7293 11023 7327
rect 10965 7287 11023 7293
rect 7742 7216 7748 7268
rect 7800 7256 7806 7268
rect 8205 7259 8263 7265
rect 8205 7256 8217 7259
rect 7800 7228 8217 7256
rect 7800 7216 7806 7228
rect 8205 7225 8217 7228
rect 8251 7225 8263 7259
rect 8754 7256 8760 7268
rect 8715 7228 8760 7256
rect 8205 7219 8263 7225
rect 8754 7216 8760 7228
rect 8812 7216 8818 7268
rect 9493 7259 9551 7265
rect 9493 7225 9505 7259
rect 9539 7256 9551 7259
rect 9876 7256 9904 7287
rect 11238 7284 11244 7336
rect 11296 7324 11302 7336
rect 11368 7327 11426 7333
rect 11368 7324 11380 7327
rect 11296 7296 11380 7324
rect 11296 7284 11302 7296
rect 11368 7293 11380 7296
rect 11414 7324 11426 7327
rect 11793 7327 11851 7333
rect 11793 7324 11805 7327
rect 11414 7296 11805 7324
rect 11414 7293 11426 7296
rect 11368 7287 11426 7293
rect 11793 7293 11805 7296
rect 11839 7324 11851 7327
rect 11882 7324 11888 7336
rect 11839 7296 11888 7324
rect 11839 7293 11851 7296
rect 11793 7287 11851 7293
rect 11882 7284 11888 7296
rect 11940 7284 11946 7336
rect 12618 7324 12624 7336
rect 12579 7296 12624 7324
rect 12618 7284 12624 7296
rect 12676 7284 12682 7336
rect 12989 7327 13047 7333
rect 12989 7293 13001 7327
rect 13035 7324 13047 7327
rect 14182 7324 14188 7336
rect 13035 7296 14188 7324
rect 13035 7293 13047 7296
rect 12989 7287 13047 7293
rect 14182 7284 14188 7296
rect 14240 7284 14246 7336
rect 14384 7333 14412 7364
rect 16117 7361 16129 7395
rect 16163 7392 16175 7395
rect 16482 7392 16488 7404
rect 16163 7364 16488 7392
rect 16163 7361 16175 7364
rect 16117 7355 16175 7361
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 14369 7327 14427 7333
rect 14369 7293 14381 7327
rect 14415 7324 14427 7327
rect 14461 7327 14519 7333
rect 14461 7324 14473 7327
rect 14415 7296 14473 7324
rect 14415 7293 14427 7296
rect 14369 7287 14427 7293
rect 14461 7293 14473 7296
rect 14507 7293 14519 7327
rect 14461 7287 14519 7293
rect 14550 7284 14556 7336
rect 14608 7324 14614 7336
rect 15013 7327 15071 7333
rect 15013 7324 15025 7327
rect 14608 7296 15025 7324
rect 14608 7284 14614 7296
rect 15013 7293 15025 7296
rect 15059 7324 15071 7327
rect 15059 7296 15332 7324
rect 15059 7293 15071 7296
rect 15013 7287 15071 7293
rect 12636 7256 12664 7284
rect 15194 7256 15200 7268
rect 9539 7228 12664 7256
rect 15155 7228 15200 7256
rect 9539 7225 9551 7228
rect 9493 7219 9551 7225
rect 15194 7216 15200 7228
rect 15252 7216 15258 7268
rect 15304 7256 15332 7296
rect 16114 7256 16120 7268
rect 15304 7228 16120 7256
rect 16114 7216 16120 7228
rect 16172 7216 16178 7268
rect 16206 7216 16212 7268
rect 16264 7256 16270 7268
rect 16761 7259 16819 7265
rect 16264 7228 16309 7256
rect 16264 7216 16270 7228
rect 16761 7225 16773 7259
rect 16807 7256 16819 7259
rect 17770 7256 17776 7268
rect 16807 7228 17776 7256
rect 16807 7225 16819 7228
rect 16761 7219 16819 7225
rect 17770 7216 17776 7228
rect 17828 7216 17834 7268
rect 7466 7188 7472 7200
rect 7427 7160 7472 7188
rect 7466 7148 7472 7160
rect 7524 7148 7530 7200
rect 9674 7188 9680 7200
rect 9635 7160 9680 7188
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 11471 7191 11529 7197
rect 11471 7157 11483 7191
rect 11517 7188 11529 7191
rect 12066 7188 12072 7200
rect 11517 7160 12072 7188
rect 11517 7157 11529 7160
rect 11471 7151 11529 7157
rect 12066 7148 12072 7160
rect 12124 7148 12130 7200
rect 12250 7188 12256 7200
rect 12211 7160 12256 7188
rect 12250 7148 12256 7160
rect 12308 7148 12314 7200
rect 12526 7188 12532 7200
rect 12487 7160 12532 7188
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 15470 7188 15476 7200
rect 15431 7160 15476 7188
rect 15470 7148 15476 7160
rect 15528 7148 15534 7200
rect 15930 7188 15936 7200
rect 15891 7160 15936 7188
rect 15930 7148 15936 7160
rect 15988 7148 15994 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 7558 6984 7564 6996
rect 7519 6956 7564 6984
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 7926 6984 7932 6996
rect 7887 6956 7932 6984
rect 7926 6944 7932 6956
rect 7984 6984 7990 6996
rect 9490 6984 9496 6996
rect 7984 6956 9496 6984
rect 7984 6944 7990 6956
rect 9490 6944 9496 6956
rect 9548 6984 9554 6996
rect 11422 6984 11428 6996
rect 9548 6956 9674 6984
rect 11383 6956 11428 6984
rect 9548 6944 9554 6956
rect 8110 6876 8116 6928
rect 8168 6916 8174 6928
rect 8205 6919 8263 6925
rect 8205 6916 8217 6919
rect 8168 6888 8217 6916
rect 8168 6876 8174 6888
rect 8205 6885 8217 6888
rect 8251 6885 8263 6919
rect 8754 6916 8760 6928
rect 8715 6888 8760 6916
rect 8205 6879 8263 6885
rect 8754 6876 8760 6888
rect 8812 6916 8818 6928
rect 9033 6919 9091 6925
rect 9033 6916 9045 6919
rect 8812 6888 9045 6916
rect 8812 6876 8818 6888
rect 9033 6885 9045 6888
rect 9079 6885 9091 6919
rect 9646 6916 9674 6956
rect 11422 6944 11428 6956
rect 11480 6944 11486 6996
rect 12250 6944 12256 6996
rect 12308 6984 12314 6996
rect 12345 6987 12403 6993
rect 12345 6984 12357 6987
rect 12308 6956 12357 6984
rect 12308 6944 12314 6956
rect 12345 6953 12357 6956
rect 12391 6984 12403 6987
rect 14274 6984 14280 6996
rect 12391 6956 14280 6984
rect 12391 6953 12403 6956
rect 12345 6947 12403 6953
rect 14274 6944 14280 6956
rect 14332 6944 14338 6996
rect 15105 6987 15163 6993
rect 15105 6953 15117 6987
rect 15151 6984 15163 6987
rect 15378 6984 15384 6996
rect 15151 6956 15384 6984
rect 15151 6953 15163 6956
rect 15105 6947 15163 6953
rect 15378 6944 15384 6956
rect 15436 6944 15442 6996
rect 15654 6984 15660 6996
rect 15615 6956 15660 6984
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 15930 6944 15936 6996
rect 15988 6984 15994 6996
rect 16206 6984 16212 6996
rect 15988 6956 16212 6984
rect 15988 6944 15994 6956
rect 16206 6944 16212 6956
rect 16264 6944 16270 6996
rect 17129 6987 17187 6993
rect 17129 6984 17141 6987
rect 16316 6956 17141 6984
rect 9998 6919 10056 6925
rect 9998 6916 10010 6919
rect 9646 6888 10010 6916
rect 9033 6879 9091 6885
rect 9998 6885 10010 6888
rect 10044 6885 10056 6919
rect 9998 6879 10056 6885
rect 15838 6876 15844 6928
rect 15896 6916 15902 6928
rect 16316 6916 16344 6956
rect 17129 6953 17141 6956
rect 17175 6953 17187 6987
rect 17129 6947 17187 6953
rect 15896 6888 16344 6916
rect 15896 6876 15902 6888
rect 7060 6851 7118 6857
rect 7060 6817 7072 6851
rect 7106 6848 7118 6851
rect 7466 6848 7472 6860
rect 7106 6820 7472 6848
rect 7106 6817 7118 6820
rect 7060 6811 7118 6817
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6848 9551 6851
rect 9674 6848 9680 6860
rect 9539 6820 9680 6848
rect 9539 6817 9551 6820
rect 9493 6811 9551 6817
rect 9674 6808 9680 6820
rect 9732 6808 9738 6860
rect 11238 6808 11244 6860
rect 11296 6848 11302 6860
rect 11977 6851 12035 6857
rect 11977 6848 11989 6851
rect 11296 6820 11989 6848
rect 11296 6808 11302 6820
rect 11977 6817 11989 6820
rect 12023 6848 12035 6851
rect 12526 6848 12532 6860
rect 12023 6820 12532 6848
rect 12023 6817 12035 6820
rect 11977 6811 12035 6817
rect 12526 6808 12532 6820
rect 12584 6808 12590 6860
rect 15194 6808 15200 6860
rect 15252 6848 15258 6860
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 15252 6820 15301 6848
rect 15252 6808 15258 6820
rect 15289 6817 15301 6820
rect 15335 6817 15347 6851
rect 17034 6848 17040 6860
rect 16995 6820 17040 6848
rect 15289 6811 15347 6817
rect 17034 6808 17040 6820
rect 17092 6808 17098 6860
rect 17494 6848 17500 6860
rect 17455 6820 17500 6848
rect 17494 6808 17500 6820
rect 17552 6808 17558 6860
rect 6638 6740 6644 6792
rect 6696 6780 6702 6792
rect 7147 6783 7205 6789
rect 7147 6780 7159 6783
rect 6696 6752 7159 6780
rect 6696 6740 6702 6752
rect 7147 6749 7159 6752
rect 7193 6780 7205 6783
rect 8113 6783 8171 6789
rect 8113 6780 8125 6783
rect 7193 6752 8125 6780
rect 7193 6749 7205 6752
rect 7147 6743 7205 6749
rect 8113 6749 8125 6752
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 14185 6783 14243 6789
rect 14185 6749 14197 6783
rect 14231 6780 14243 6783
rect 15930 6780 15936 6792
rect 14231 6752 15936 6780
rect 14231 6749 14243 6752
rect 14185 6743 14243 6749
rect 15930 6740 15936 6752
rect 15988 6740 15994 6792
rect 16114 6740 16120 6792
rect 16172 6780 16178 6792
rect 17512 6780 17540 6808
rect 16172 6752 17540 6780
rect 16172 6740 16178 6752
rect 6362 6672 6368 6724
rect 6420 6712 6426 6724
rect 13262 6712 13268 6724
rect 6420 6684 13268 6712
rect 6420 6672 6426 6684
rect 13262 6672 13268 6684
rect 13320 6712 13326 6724
rect 18414 6712 18420 6724
rect 13320 6684 18420 6712
rect 13320 6672 13326 6684
rect 18414 6672 18420 6684
rect 18472 6672 18478 6724
rect 10594 6644 10600 6656
rect 10555 6616 10600 6644
rect 10594 6604 10600 6616
rect 10652 6604 10658 6656
rect 12894 6644 12900 6656
rect 12855 6616 12900 6644
rect 12894 6604 12900 6616
rect 12952 6604 12958 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 6638 6440 6644 6452
rect 6599 6412 6644 6440
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 9490 6440 9496 6452
rect 9451 6412 9496 6440
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 9766 6400 9772 6452
rect 9824 6440 9830 6452
rect 10594 6440 10600 6452
rect 9824 6412 10600 6440
rect 9824 6400 9830 6412
rect 10594 6400 10600 6412
rect 10652 6400 10658 6452
rect 11238 6440 11244 6452
rect 11199 6412 11244 6440
rect 11238 6400 11244 6412
rect 11296 6400 11302 6452
rect 12069 6443 12127 6449
rect 12069 6409 12081 6443
rect 12115 6440 12127 6443
rect 12250 6440 12256 6452
rect 12115 6412 12256 6440
rect 12115 6409 12127 6412
rect 12069 6403 12127 6409
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 15930 6440 15936 6452
rect 15891 6412 15936 6440
rect 15930 6400 15936 6412
rect 15988 6400 15994 6452
rect 17034 6400 17040 6452
rect 17092 6440 17098 6452
rect 17129 6443 17187 6449
rect 17129 6440 17141 6443
rect 17092 6412 17141 6440
rect 17092 6400 17098 6412
rect 17129 6409 17141 6412
rect 17175 6409 17187 6443
rect 17129 6403 17187 6409
rect 8110 6332 8116 6384
rect 8168 6372 8174 6384
rect 9033 6375 9091 6381
rect 9033 6372 9045 6375
rect 8168 6344 9045 6372
rect 8168 6332 8174 6344
rect 9033 6341 9045 6344
rect 9079 6372 9091 6375
rect 9122 6372 9128 6384
rect 9079 6344 9128 6372
rect 9079 6341 9091 6344
rect 9033 6335 9091 6341
rect 9122 6332 9128 6344
rect 9180 6332 9186 6384
rect 8754 6304 8760 6316
rect 8715 6276 8760 6304
rect 8754 6264 8760 6276
rect 8812 6304 8818 6316
rect 9677 6307 9735 6313
rect 9677 6304 9689 6307
rect 8812 6276 9689 6304
rect 8812 6264 8818 6276
rect 9677 6273 9689 6276
rect 9723 6273 9735 6307
rect 10134 6304 10140 6316
rect 10095 6276 10140 6304
rect 9677 6267 9735 6273
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 13170 6304 13176 6316
rect 13131 6276 13176 6304
rect 13170 6264 13176 6276
rect 13228 6264 13234 6316
rect 14369 6307 14427 6313
rect 14369 6273 14381 6307
rect 14415 6304 14427 6307
rect 14458 6304 14464 6316
rect 14415 6276 14464 6304
rect 14415 6273 14427 6276
rect 14369 6267 14427 6273
rect 14458 6264 14464 6276
rect 14516 6304 14522 6316
rect 15838 6304 15844 6316
rect 14516 6276 15844 6304
rect 14516 6264 14522 6276
rect 15838 6264 15844 6276
rect 15896 6264 15902 6316
rect 15948 6304 15976 6400
rect 16209 6307 16267 6313
rect 16209 6304 16221 6307
rect 15948 6276 16221 6304
rect 16209 6273 16221 6276
rect 16255 6273 16267 6307
rect 16482 6304 16488 6316
rect 16443 6276 16488 6304
rect 16209 6267 16267 6273
rect 16482 6264 16488 6276
rect 16540 6264 16546 6316
rect 15562 6236 15568 6248
rect 14746 6208 15568 6236
rect 7009 6171 7067 6177
rect 7009 6137 7021 6171
rect 7055 6168 7067 6171
rect 7837 6171 7895 6177
rect 7837 6168 7849 6171
rect 7055 6140 7849 6168
rect 7055 6137 7067 6140
rect 7009 6131 7067 6137
rect 7837 6137 7849 6140
rect 7883 6168 7895 6171
rect 8113 6171 8171 6177
rect 8113 6168 8125 6171
rect 7883 6140 8125 6168
rect 7883 6137 7895 6140
rect 7837 6131 7895 6137
rect 8113 6137 8125 6140
rect 8159 6137 8171 6171
rect 8113 6131 8171 6137
rect 8202 6128 8208 6180
rect 8260 6168 8266 6180
rect 8260 6140 8305 6168
rect 8260 6128 8266 6140
rect 9766 6128 9772 6180
rect 9824 6168 9830 6180
rect 11333 6171 11391 6177
rect 9824 6140 9869 6168
rect 9824 6128 9830 6140
rect 11333 6137 11345 6171
rect 11379 6168 11391 6171
rect 12526 6168 12532 6180
rect 11379 6140 12532 6168
rect 11379 6137 11391 6140
rect 11333 6131 11391 6137
rect 12526 6128 12532 6140
rect 12584 6128 12590 6180
rect 12618 6128 12624 6180
rect 12676 6168 12682 6180
rect 13449 6171 13507 6177
rect 13449 6168 13461 6171
rect 12676 6140 13461 6168
rect 12676 6128 12682 6140
rect 13449 6137 13461 6140
rect 13495 6137 13507 6171
rect 14274 6168 14280 6180
rect 14187 6140 14280 6168
rect 13449 6131 13507 6137
rect 14274 6128 14280 6140
rect 14332 6168 14338 6180
rect 14746 6177 14774 6208
rect 15562 6196 15568 6208
rect 15620 6196 15626 6248
rect 14731 6171 14789 6177
rect 14731 6168 14743 6171
rect 14332 6140 14743 6168
rect 14332 6128 14338 6140
rect 14731 6137 14743 6140
rect 14777 6137 14789 6171
rect 16301 6171 16359 6177
rect 16301 6168 16313 6171
rect 14731 6131 14789 6137
rect 15396 6140 16313 6168
rect 15396 6112 15424 6140
rect 16301 6137 16313 6140
rect 16347 6137 16359 6171
rect 16301 6131 16359 6137
rect 7466 6100 7472 6112
rect 7427 6072 7472 6100
rect 7466 6060 7472 6072
rect 7524 6060 7530 6112
rect 15289 6103 15347 6109
rect 15289 6069 15301 6103
rect 15335 6100 15347 6103
rect 15378 6100 15384 6112
rect 15335 6072 15384 6100
rect 15335 6069 15347 6072
rect 15289 6063 15347 6069
rect 15378 6060 15384 6072
rect 15436 6060 15442 6112
rect 15562 6100 15568 6112
rect 15523 6072 15568 6100
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 17494 6100 17500 6112
rect 17455 6072 17500 6100
rect 17494 6060 17500 6072
rect 17552 6060 17558 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 12526 5856 12532 5908
rect 12584 5896 12590 5908
rect 12621 5899 12679 5905
rect 12621 5896 12633 5899
rect 12584 5868 12633 5896
rect 12584 5856 12590 5868
rect 12621 5865 12633 5868
rect 12667 5865 12679 5899
rect 14458 5896 14464 5908
rect 14419 5868 14464 5896
rect 12621 5859 12679 5865
rect 14458 5856 14464 5868
rect 14516 5856 14522 5908
rect 15105 5899 15163 5905
rect 15105 5865 15117 5899
rect 15151 5896 15163 5899
rect 15286 5896 15292 5908
rect 15151 5868 15292 5896
rect 15151 5865 15163 5868
rect 15105 5859 15163 5865
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 16942 5896 16948 5908
rect 16903 5868 16948 5896
rect 16942 5856 16948 5868
rect 17000 5856 17006 5908
rect 18506 5896 18512 5908
rect 18467 5868 18512 5896
rect 18506 5856 18512 5868
rect 18564 5856 18570 5908
rect 7926 5788 7932 5840
rect 7984 5828 7990 5840
rect 8158 5831 8216 5837
rect 8158 5828 8170 5831
rect 7984 5800 8170 5828
rect 7984 5788 7990 5800
rect 8158 5797 8170 5800
rect 8204 5797 8216 5831
rect 9858 5828 9864 5840
rect 9819 5800 9864 5828
rect 8158 5791 8216 5797
rect 9858 5788 9864 5800
rect 9916 5788 9922 5840
rect 11787 5831 11845 5837
rect 11787 5797 11799 5831
rect 11833 5828 11845 5831
rect 12250 5828 12256 5840
rect 11833 5800 12256 5828
rect 11833 5797 11845 5800
rect 11787 5791 11845 5797
rect 12250 5788 12256 5800
rect 12308 5788 12314 5840
rect 12894 5788 12900 5840
rect 12952 5828 12958 5840
rect 13357 5831 13415 5837
rect 13357 5828 13369 5831
rect 12952 5800 13369 5828
rect 12952 5788 12958 5800
rect 13357 5797 13369 5800
rect 13403 5828 13415 5831
rect 13722 5828 13728 5840
rect 13403 5800 13728 5828
rect 13403 5797 13415 5800
rect 13357 5791 13415 5797
rect 13722 5788 13728 5800
rect 13780 5788 13786 5840
rect 14182 5788 14188 5840
rect 14240 5828 14246 5840
rect 17494 5828 17500 5840
rect 14240 5800 15792 5828
rect 17407 5800 17500 5828
rect 14240 5788 14246 5800
rect 6362 5760 6368 5772
rect 6323 5732 6368 5760
rect 6362 5720 6368 5732
rect 6420 5720 6426 5772
rect 6454 5720 6460 5772
rect 6512 5760 6518 5772
rect 6733 5763 6791 5769
rect 6733 5760 6745 5763
rect 6512 5732 6745 5760
rect 6512 5720 6518 5732
rect 6733 5729 6745 5732
rect 6779 5729 6791 5763
rect 6733 5723 6791 5729
rect 7009 5763 7067 5769
rect 7009 5729 7021 5763
rect 7055 5760 7067 5763
rect 9122 5760 9128 5772
rect 7055 5732 9128 5760
rect 7055 5729 7067 5732
rect 7009 5723 7067 5729
rect 9122 5720 9128 5732
rect 9180 5720 9186 5772
rect 11330 5720 11336 5772
rect 11388 5760 11394 5772
rect 11425 5763 11483 5769
rect 11425 5760 11437 5763
rect 11388 5732 11437 5760
rect 11388 5720 11394 5732
rect 11425 5729 11437 5732
rect 11471 5729 11483 5763
rect 11425 5723 11483 5729
rect 14642 5720 14648 5772
rect 14700 5760 14706 5772
rect 15764 5769 15792 5800
rect 15289 5763 15347 5769
rect 15289 5760 15301 5763
rect 14700 5732 15301 5760
rect 14700 5720 14706 5732
rect 15289 5729 15301 5732
rect 15335 5729 15347 5763
rect 15289 5723 15347 5729
rect 15749 5763 15807 5769
rect 15749 5729 15761 5763
rect 15795 5760 15807 5763
rect 16390 5760 16396 5772
rect 15795 5732 16396 5760
rect 15795 5729 15807 5732
rect 15749 5723 15807 5729
rect 16390 5720 16396 5732
rect 16448 5720 16454 5772
rect 16758 5720 16764 5772
rect 16816 5760 16822 5772
rect 16853 5763 16911 5769
rect 16853 5760 16865 5763
rect 16816 5732 16865 5760
rect 16816 5720 16822 5732
rect 16853 5729 16865 5732
rect 16899 5729 16911 5763
rect 16853 5723 16911 5729
rect 17034 5720 17040 5772
rect 17092 5760 17098 5772
rect 17420 5769 17448 5800
rect 17494 5788 17500 5800
rect 17552 5828 17558 5840
rect 17552 5800 18920 5828
rect 17552 5788 17558 5800
rect 18892 5772 18920 5800
rect 17405 5763 17463 5769
rect 17405 5760 17417 5763
rect 17092 5732 17417 5760
rect 17092 5720 17098 5732
rect 17405 5729 17417 5732
rect 17451 5729 17463 5763
rect 18414 5760 18420 5772
rect 18375 5732 18420 5760
rect 17405 5723 17463 5729
rect 18414 5720 18420 5732
rect 18472 5720 18478 5772
rect 18874 5760 18880 5772
rect 18835 5732 18880 5760
rect 18874 5720 18880 5732
rect 18932 5720 18938 5772
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5692 7435 5695
rect 7837 5695 7895 5701
rect 7837 5692 7849 5695
rect 7423 5664 7849 5692
rect 7423 5661 7435 5664
rect 7377 5655 7435 5661
rect 7837 5661 7849 5664
rect 7883 5692 7895 5695
rect 8018 5692 8024 5704
rect 7883 5664 8024 5692
rect 7883 5661 7895 5664
rect 7837 5655 7895 5661
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 9214 5652 9220 5704
rect 9272 5692 9278 5704
rect 9769 5695 9827 5701
rect 9769 5692 9781 5695
rect 9272 5664 9781 5692
rect 9272 5652 9278 5664
rect 9769 5661 9781 5664
rect 9815 5661 9827 5695
rect 10134 5692 10140 5704
rect 10095 5664 10140 5692
rect 9769 5655 9827 5661
rect 10134 5652 10140 5664
rect 10192 5692 10198 5704
rect 10962 5692 10968 5704
rect 10192 5664 10968 5692
rect 10192 5652 10198 5664
rect 10962 5652 10968 5664
rect 11020 5652 11026 5704
rect 13262 5692 13268 5704
rect 13223 5664 13268 5692
rect 13262 5652 13268 5664
rect 13320 5652 13326 5704
rect 13446 5652 13452 5704
rect 13504 5692 13510 5704
rect 15841 5695 15899 5701
rect 15841 5692 15853 5695
rect 13504 5664 15853 5692
rect 13504 5652 13510 5664
rect 15841 5661 15853 5664
rect 15887 5661 15899 5695
rect 15841 5655 15899 5661
rect 13078 5584 13084 5636
rect 13136 5624 13142 5636
rect 13817 5627 13875 5633
rect 13817 5624 13829 5627
rect 13136 5596 13829 5624
rect 13136 5584 13142 5596
rect 13817 5593 13829 5596
rect 13863 5624 13875 5627
rect 14274 5624 14280 5636
rect 13863 5596 14280 5624
rect 13863 5593 13875 5596
rect 13817 5587 13875 5593
rect 14274 5584 14280 5596
rect 14332 5584 14338 5636
rect 7558 5516 7564 5568
rect 7616 5556 7622 5568
rect 7653 5559 7711 5565
rect 7653 5556 7665 5559
rect 7616 5528 7665 5556
rect 7616 5516 7622 5528
rect 7653 5525 7665 5528
rect 7699 5556 7711 5559
rect 8202 5556 8208 5568
rect 7699 5528 8208 5556
rect 7699 5525 7711 5528
rect 7653 5519 7711 5525
rect 8202 5516 8208 5528
rect 8260 5556 8266 5568
rect 8757 5559 8815 5565
rect 8757 5556 8769 5559
rect 8260 5528 8769 5556
rect 8260 5516 8266 5528
rect 8757 5525 8769 5528
rect 8803 5525 8815 5559
rect 8757 5519 8815 5525
rect 11422 5516 11428 5568
rect 11480 5556 11486 5568
rect 12345 5559 12403 5565
rect 12345 5556 12357 5559
rect 11480 5528 12357 5556
rect 11480 5516 11486 5528
rect 12345 5525 12357 5528
rect 12391 5556 12403 5559
rect 12618 5556 12624 5568
rect 12391 5528 12624 5556
rect 12391 5525 12403 5528
rect 12345 5519 12403 5525
rect 12618 5516 12624 5528
rect 12676 5516 12682 5568
rect 12986 5556 12992 5568
rect 12947 5528 12992 5556
rect 12986 5516 12992 5528
rect 13044 5516 13050 5568
rect 15378 5516 15384 5568
rect 15436 5556 15442 5568
rect 16301 5559 16359 5565
rect 16301 5556 16313 5559
rect 15436 5528 16313 5556
rect 15436 5516 15442 5528
rect 16301 5525 16313 5528
rect 16347 5525 16359 5559
rect 16301 5519 16359 5525
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 6362 5352 6368 5364
rect 6323 5324 6368 5352
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 6454 5312 6460 5364
rect 6512 5352 6518 5364
rect 7009 5355 7067 5361
rect 7009 5352 7021 5355
rect 6512 5324 7021 5352
rect 6512 5312 6518 5324
rect 7009 5321 7021 5324
rect 7055 5321 7067 5355
rect 7009 5315 7067 5321
rect 7024 5284 7052 5315
rect 7926 5312 7932 5364
rect 7984 5352 7990 5364
rect 8573 5355 8631 5361
rect 8573 5352 8585 5355
rect 7984 5324 8585 5352
rect 7984 5312 7990 5324
rect 8573 5321 8585 5324
rect 8619 5352 8631 5355
rect 8941 5355 8999 5361
rect 8941 5352 8953 5355
rect 8619 5324 8953 5352
rect 8619 5321 8631 5324
rect 8573 5315 8631 5321
rect 8941 5321 8953 5324
rect 8987 5321 8999 5355
rect 8941 5315 8999 5321
rect 7650 5284 7656 5296
rect 7024 5256 7656 5284
rect 7650 5244 7656 5256
rect 7708 5284 7714 5296
rect 7708 5256 8064 5284
rect 7708 5244 7714 5256
rect 7834 5216 7840 5228
rect 7760 5188 7840 5216
rect 7760 5157 7788 5188
rect 7834 5176 7840 5188
rect 7892 5176 7898 5228
rect 8036 5157 8064 5256
rect 7469 5151 7527 5157
rect 7469 5117 7481 5151
rect 7515 5148 7527 5151
rect 7745 5151 7803 5157
rect 7745 5148 7757 5151
rect 7515 5120 7757 5148
rect 7515 5117 7527 5120
rect 7469 5111 7527 5117
rect 7745 5117 7757 5120
rect 7791 5117 7803 5151
rect 7745 5111 7803 5117
rect 8021 5151 8079 5157
rect 8021 5117 8033 5151
rect 8067 5117 8079 5151
rect 8956 5148 8984 5315
rect 9858 5312 9864 5364
rect 9916 5352 9922 5364
rect 10321 5355 10379 5361
rect 10321 5352 10333 5355
rect 9916 5324 10333 5352
rect 9916 5312 9922 5324
rect 10321 5321 10333 5324
rect 10367 5321 10379 5355
rect 10321 5315 10379 5321
rect 11330 5312 11336 5364
rect 11388 5352 11394 5364
rect 12069 5355 12127 5361
rect 12069 5352 12081 5355
rect 11388 5324 12081 5352
rect 11388 5312 11394 5324
rect 12069 5321 12081 5324
rect 12115 5321 12127 5355
rect 13722 5352 13728 5364
rect 13683 5324 13728 5352
rect 12069 5315 12127 5321
rect 13722 5312 13728 5324
rect 13780 5312 13786 5364
rect 16390 5352 16396 5364
rect 16351 5324 16396 5352
rect 16390 5312 16396 5324
rect 16448 5312 16454 5364
rect 17402 5352 17408 5364
rect 17363 5324 17408 5352
rect 17402 5312 17408 5324
rect 17460 5312 17466 5364
rect 17770 5352 17776 5364
rect 17731 5324 17776 5352
rect 17770 5312 17776 5324
rect 17828 5312 17834 5364
rect 18414 5312 18420 5364
rect 18472 5352 18478 5364
rect 18509 5355 18567 5361
rect 18509 5352 18521 5355
rect 18472 5324 18521 5352
rect 18472 5312 18478 5324
rect 18509 5321 18521 5324
rect 18555 5321 18567 5355
rect 18874 5352 18880 5364
rect 18835 5324 18880 5352
rect 18509 5315 18567 5321
rect 18874 5312 18880 5324
rect 18932 5312 18938 5364
rect 10870 5244 10876 5296
rect 10928 5284 10934 5296
rect 16574 5284 16580 5296
rect 10928 5256 16580 5284
rect 10928 5244 10934 5256
rect 16574 5244 16580 5256
rect 16632 5244 16638 5296
rect 9122 5216 9128 5228
rect 9083 5188 9128 5216
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 11238 5176 11244 5228
rect 11296 5216 11302 5228
rect 13078 5216 13084 5228
rect 11296 5188 13084 5216
rect 11296 5176 11302 5188
rect 13078 5176 13084 5188
rect 13136 5176 13142 5228
rect 14369 5219 14427 5225
rect 14369 5185 14381 5219
rect 14415 5216 14427 5219
rect 15197 5219 15255 5225
rect 15197 5216 15209 5219
rect 14415 5188 15209 5216
rect 14415 5185 14427 5188
rect 14369 5179 14427 5185
rect 15197 5185 15209 5188
rect 15243 5216 15255 5219
rect 18506 5216 18512 5228
rect 15243 5188 18512 5216
rect 15243 5185 15255 5188
rect 15197 5179 15255 5185
rect 18506 5176 18512 5188
rect 18564 5176 18570 5228
rect 8956 5120 9168 5148
rect 8021 5111 8079 5117
rect 8297 5083 8355 5089
rect 8297 5049 8309 5083
rect 8343 5080 8355 5083
rect 9030 5080 9036 5092
rect 8343 5052 9036 5080
rect 8343 5049 8355 5052
rect 8297 5043 8355 5049
rect 9030 5040 9036 5052
rect 9088 5040 9094 5092
rect 9140 5080 9168 5120
rect 9214 5108 9220 5160
rect 9272 5148 9278 5160
rect 10689 5151 10747 5157
rect 10689 5148 10701 5151
rect 9272 5120 10701 5148
rect 9272 5108 9278 5120
rect 10689 5117 10701 5120
rect 10735 5117 10747 5151
rect 10689 5111 10747 5117
rect 10940 5151 10998 5157
rect 10940 5117 10952 5151
rect 10986 5148 10998 5151
rect 17012 5151 17070 5157
rect 10986 5120 11468 5148
rect 10986 5117 10998 5120
rect 10940 5111 10998 5117
rect 9446 5083 9504 5089
rect 9446 5080 9458 5083
rect 9140 5052 9458 5080
rect 9446 5049 9458 5052
rect 9492 5080 9504 5083
rect 9766 5080 9772 5092
rect 9492 5052 9772 5080
rect 9492 5049 9504 5052
rect 9446 5043 9504 5049
rect 9766 5040 9772 5052
rect 9824 5040 9830 5092
rect 11440 5089 11468 5120
rect 17012 5117 17024 5151
rect 17058 5148 17070 5151
rect 17402 5148 17408 5160
rect 17058 5120 17408 5148
rect 17058 5117 17070 5120
rect 17012 5111 17070 5117
rect 17402 5108 17408 5120
rect 17460 5108 17466 5160
rect 17770 5108 17776 5160
rect 17828 5148 17834 5160
rect 18084 5151 18142 5157
rect 18084 5148 18096 5151
rect 17828 5120 18096 5148
rect 17828 5108 17834 5120
rect 18084 5117 18096 5120
rect 18130 5117 18142 5151
rect 18084 5111 18142 5117
rect 11425 5083 11483 5089
rect 11425 5049 11437 5083
rect 11471 5080 11483 5083
rect 12158 5080 12164 5092
rect 11471 5052 12164 5080
rect 11471 5049 11483 5052
rect 11425 5043 11483 5049
rect 12158 5040 12164 5052
rect 12216 5040 12222 5092
rect 12805 5083 12863 5089
rect 12805 5049 12817 5083
rect 12851 5049 12863 5083
rect 12805 5043 12863 5049
rect 12897 5083 12955 5089
rect 12897 5049 12909 5083
rect 12943 5080 12955 5083
rect 12986 5080 12992 5092
rect 12943 5052 12992 5080
rect 12943 5049 12955 5052
rect 12897 5043 12955 5049
rect 10042 5012 10048 5024
rect 10003 4984 10048 5012
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 10134 4972 10140 5024
rect 10192 5012 10198 5024
rect 11011 5015 11069 5021
rect 11011 5012 11023 5015
rect 10192 4984 11023 5012
rect 10192 4972 10198 4984
rect 11011 4981 11023 4984
rect 11057 4981 11069 5015
rect 11011 4975 11069 4981
rect 11793 5015 11851 5021
rect 11793 4981 11805 5015
rect 11839 5012 11851 5015
rect 12250 5012 12256 5024
rect 11839 4984 12256 5012
rect 11839 4981 11851 4984
rect 11793 4975 11851 4981
rect 12250 4972 12256 4984
rect 12308 4972 12314 5024
rect 12710 4972 12716 5024
rect 12768 5012 12774 5024
rect 12820 5012 12848 5043
rect 12986 5040 12992 5052
rect 13044 5040 13050 5092
rect 16758 5080 16764 5092
rect 14660 5052 16764 5080
rect 14660 5024 14688 5052
rect 16758 5040 16764 5052
rect 16816 5040 16822 5092
rect 14642 5012 14648 5024
rect 12768 4984 12848 5012
rect 14603 4984 14648 5012
rect 12768 4972 12774 4984
rect 14642 4972 14648 4984
rect 14700 4972 14706 5024
rect 14734 4972 14740 5024
rect 14792 5012 14798 5024
rect 15105 5015 15163 5021
rect 15105 5012 15117 5015
rect 14792 4984 15117 5012
rect 14792 4972 14798 4984
rect 15105 4981 15117 4984
rect 15151 5012 15163 5015
rect 15562 5012 15568 5024
rect 15151 4984 15568 5012
rect 15151 4981 15163 4984
rect 15105 4975 15163 4981
rect 15562 4972 15568 4984
rect 15620 4972 15626 5024
rect 16114 5012 16120 5024
rect 16075 4984 16120 5012
rect 16114 4972 16120 4984
rect 16172 4972 16178 5024
rect 16850 4972 16856 5024
rect 16908 5012 16914 5024
rect 17083 5015 17141 5021
rect 17083 5012 17095 5015
rect 16908 4984 17095 5012
rect 16908 4972 16914 4984
rect 17083 4981 17095 4984
rect 17129 4981 17141 5015
rect 17083 4975 17141 4981
rect 18187 5015 18245 5021
rect 18187 4981 18199 5015
rect 18233 5012 18245 5015
rect 18414 5012 18420 5024
rect 18233 4984 18420 5012
rect 18233 4981 18245 4984
rect 18187 4975 18245 4981
rect 18414 4972 18420 4984
rect 18472 4972 18478 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 7650 4808 7656 4820
rect 7611 4780 7656 4808
rect 7650 4768 7656 4780
rect 7708 4768 7714 4820
rect 8018 4808 8024 4820
rect 7979 4780 8024 4808
rect 8018 4768 8024 4780
rect 8076 4768 8082 4820
rect 9858 4768 9864 4820
rect 9916 4808 9922 4820
rect 10597 4811 10655 4817
rect 10597 4808 10609 4811
rect 9916 4780 10609 4808
rect 9916 4768 9922 4780
rect 10597 4777 10609 4780
rect 10643 4777 10655 4811
rect 10597 4771 10655 4777
rect 12250 4768 12256 4820
rect 12308 4808 12314 4820
rect 12345 4811 12403 4817
rect 12345 4808 12357 4811
rect 12308 4780 12357 4808
rect 12308 4768 12314 4780
rect 12345 4777 12357 4780
rect 12391 4777 12403 4811
rect 12345 4771 12403 4777
rect 12897 4811 12955 4817
rect 12897 4777 12909 4811
rect 12943 4808 12955 4811
rect 12986 4808 12992 4820
rect 12943 4780 12992 4808
rect 12943 4777 12955 4780
rect 12897 4771 12955 4777
rect 12986 4768 12992 4780
rect 13044 4768 13050 4820
rect 13262 4768 13268 4820
rect 13320 4808 13326 4820
rect 13541 4811 13599 4817
rect 13541 4808 13553 4811
rect 13320 4780 13553 4808
rect 13320 4768 13326 4780
rect 13541 4777 13553 4780
rect 13587 4777 13599 4811
rect 13541 4771 13599 4777
rect 15562 4768 15568 4820
rect 15620 4808 15626 4820
rect 15657 4811 15715 4817
rect 15657 4808 15669 4811
rect 15620 4780 15669 4808
rect 15620 4768 15626 4780
rect 15657 4777 15669 4780
rect 15703 4808 15715 4811
rect 16022 4808 16028 4820
rect 15703 4780 16028 4808
rect 15703 4777 15715 4780
rect 15657 4771 15715 4777
rect 16022 4768 16028 4780
rect 16080 4768 16086 4820
rect 16945 4811 17003 4817
rect 16945 4777 16957 4811
rect 16991 4808 17003 4811
rect 17034 4808 17040 4820
rect 16991 4780 17040 4808
rect 16991 4777 17003 4780
rect 16945 4771 17003 4777
rect 17034 4768 17040 4780
rect 17092 4768 17098 4820
rect 7668 4740 7696 4768
rect 7668 4712 8432 4740
rect 6822 4632 6828 4684
rect 6880 4672 6886 4684
rect 8404 4681 8432 4712
rect 9766 4700 9772 4752
rect 9824 4740 9830 4752
rect 9998 4743 10056 4749
rect 9998 4740 10010 4743
rect 9824 4712 10010 4740
rect 9824 4700 9830 4712
rect 9998 4709 10010 4712
rect 10044 4709 10056 4743
rect 9998 4703 10056 4709
rect 16114 4700 16120 4752
rect 16172 4740 16178 4752
rect 17221 4743 17279 4749
rect 17221 4740 17233 4743
rect 16172 4712 17233 4740
rect 16172 4700 16178 4712
rect 17221 4709 17233 4712
rect 17267 4740 17279 4743
rect 17494 4740 17500 4752
rect 17267 4712 17500 4740
rect 17267 4709 17279 4712
rect 17221 4703 17279 4709
rect 17494 4700 17500 4712
rect 17552 4700 17558 4752
rect 17770 4740 17776 4752
rect 17731 4712 17776 4740
rect 17770 4700 17776 4712
rect 17828 4700 17834 4752
rect 6952 4675 7010 4681
rect 6952 4672 6964 4675
rect 6880 4644 6964 4672
rect 6880 4632 6886 4644
rect 6952 4641 6964 4644
rect 6998 4641 7010 4675
rect 6952 4635 7010 4641
rect 8205 4675 8263 4681
rect 8205 4641 8217 4675
rect 8251 4641 8263 4675
rect 8205 4635 8263 4641
rect 8389 4675 8447 4681
rect 8389 4641 8401 4675
rect 8435 4672 8447 4675
rect 8754 4672 8760 4684
rect 8435 4644 8760 4672
rect 8435 4641 8447 4644
rect 8389 4635 8447 4641
rect 8220 4604 8248 4635
rect 8754 4632 8760 4644
rect 8812 4632 8818 4684
rect 9030 4632 9036 4684
rect 9088 4672 9094 4684
rect 9674 4672 9680 4684
rect 9088 4644 9680 4672
rect 9088 4632 9094 4644
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 10962 4632 10968 4684
rect 11020 4672 11026 4684
rect 13760 4675 13818 4681
rect 13760 4672 13772 4675
rect 11020 4644 13772 4672
rect 11020 4632 11026 4644
rect 13760 4641 13772 4644
rect 13806 4672 13818 4675
rect 13998 4672 14004 4684
rect 13806 4644 14004 4672
rect 13806 4641 13818 4644
rect 13760 4635 13818 4641
rect 13998 4632 14004 4644
rect 14056 4632 14062 4684
rect 14642 4632 14648 4684
rect 14700 4672 14706 4684
rect 15289 4675 15347 4681
rect 15289 4672 15301 4675
rect 14700 4644 15301 4672
rect 14700 4632 14706 4644
rect 15289 4641 15301 4644
rect 15335 4672 15347 4675
rect 16942 4672 16948 4684
rect 15335 4644 16948 4672
rect 15335 4641 15347 4644
rect 15289 4635 15347 4641
rect 16942 4632 16948 4644
rect 17000 4632 17006 4684
rect 8294 4604 8300 4616
rect 8207 4576 8300 4604
rect 8294 4564 8300 4576
rect 8352 4604 8358 4616
rect 9950 4604 9956 4616
rect 8352 4576 9956 4604
rect 8352 4564 8358 4576
rect 9950 4564 9956 4576
rect 10008 4564 10014 4616
rect 11977 4607 12035 4613
rect 11977 4573 11989 4607
rect 12023 4604 12035 4607
rect 13630 4604 13636 4616
rect 12023 4576 13636 4604
rect 12023 4573 12035 4576
rect 11977 4567 12035 4573
rect 13630 4564 13636 4576
rect 13688 4564 13694 4616
rect 17126 4604 17132 4616
rect 17087 4576 17132 4604
rect 17126 4564 17132 4576
rect 17184 4564 17190 4616
rect 11882 4496 11888 4548
rect 11940 4536 11946 4548
rect 11940 4508 17034 4536
rect 11940 4496 11946 4508
rect 6638 4428 6644 4480
rect 6696 4468 6702 4480
rect 7055 4471 7113 4477
rect 7055 4468 7067 4471
rect 6696 4440 7067 4468
rect 6696 4428 6702 4440
rect 7055 4437 7067 4440
rect 7101 4437 7113 4471
rect 7055 4431 7113 4437
rect 8846 4428 8852 4480
rect 8904 4468 8910 4480
rect 8941 4471 8999 4477
rect 8941 4468 8953 4471
rect 8904 4440 8953 4468
rect 8904 4428 8910 4440
rect 8941 4437 8953 4440
rect 8987 4437 8999 4471
rect 8941 4431 8999 4437
rect 9306 4428 9312 4480
rect 9364 4468 9370 4480
rect 10870 4468 10876 4480
rect 9364 4440 10876 4468
rect 9364 4428 9370 4440
rect 10870 4428 10876 4440
rect 10928 4428 10934 4480
rect 12710 4428 12716 4480
rect 12768 4468 12774 4480
rect 13173 4471 13231 4477
rect 13173 4468 13185 4471
rect 12768 4440 13185 4468
rect 12768 4428 12774 4440
rect 13173 4437 13185 4440
rect 13219 4437 13231 4471
rect 13173 4431 13231 4437
rect 13863 4471 13921 4477
rect 13863 4437 13875 4471
rect 13909 4468 13921 4471
rect 16022 4468 16028 4480
rect 13909 4440 16028 4468
rect 13909 4437 13921 4440
rect 13863 4431 13921 4437
rect 16022 4428 16028 4440
rect 16080 4428 16086 4480
rect 16206 4468 16212 4480
rect 16167 4440 16212 4468
rect 16206 4428 16212 4440
rect 16264 4428 16270 4480
rect 17006 4468 17034 4508
rect 17862 4468 17868 4480
rect 17006 4440 17868 4468
rect 17862 4428 17868 4440
rect 17920 4428 17926 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 6273 4267 6331 4273
rect 6273 4264 6285 4267
rect 6183 4236 6285 4264
rect 6273 4233 6285 4236
rect 6319 4264 6331 4267
rect 8754 4264 8760 4276
rect 6319 4236 8524 4264
rect 8715 4236 8760 4264
rect 6319 4233 6331 4236
rect 6273 4227 6331 4233
rect 5788 4063 5846 4069
rect 5788 4029 5800 4063
rect 5834 4060 5846 4063
rect 6288 4060 6316 4227
rect 6638 4196 6644 4208
rect 6599 4168 6644 4196
rect 6638 4156 6644 4168
rect 6696 4156 6702 4208
rect 8294 4156 8300 4208
rect 8352 4196 8358 4208
rect 8389 4199 8447 4205
rect 8389 4196 8401 4199
rect 8352 4168 8401 4196
rect 8352 4156 8358 4168
rect 8389 4165 8401 4168
rect 8435 4165 8447 4199
rect 8496 4196 8524 4236
rect 8754 4224 8760 4236
rect 8812 4224 8818 4276
rect 10042 4224 10048 4276
rect 10100 4264 10106 4276
rect 10321 4267 10379 4273
rect 10321 4264 10333 4267
rect 10100 4236 10333 4264
rect 10100 4224 10106 4236
rect 10321 4233 10333 4236
rect 10367 4233 10379 4267
rect 10321 4227 10379 4233
rect 13725 4267 13783 4273
rect 13725 4233 13737 4267
rect 13771 4264 13783 4267
rect 13814 4264 13820 4276
rect 13771 4236 13820 4264
rect 13771 4233 13783 4236
rect 13725 4227 13783 4233
rect 13814 4224 13820 4236
rect 13872 4224 13878 4276
rect 13998 4264 14004 4276
rect 13959 4236 14004 4264
rect 13998 4224 14004 4236
rect 14056 4224 14062 4276
rect 14642 4264 14648 4276
rect 14603 4236 14648 4264
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 16577 4267 16635 4273
rect 16577 4233 16589 4267
rect 16623 4264 16635 4267
rect 16850 4264 16856 4276
rect 16623 4236 16856 4264
rect 16623 4233 16635 4236
rect 16577 4227 16635 4233
rect 8938 4196 8944 4208
rect 8496 4168 8944 4196
rect 8389 4159 8447 4165
rect 8938 4156 8944 4168
rect 8996 4156 9002 4208
rect 10134 4196 10140 4208
rect 9048 4168 10140 4196
rect 6656 4128 6684 4156
rect 9048 4140 9076 4168
rect 10134 4156 10140 4168
rect 10192 4156 10198 4208
rect 7469 4131 7527 4137
rect 7469 4128 7481 4131
rect 6656 4100 7481 4128
rect 7469 4097 7481 4100
rect 7515 4097 7527 4131
rect 7469 4091 7527 4097
rect 7558 4088 7564 4140
rect 7616 4128 7622 4140
rect 8846 4128 8852 4140
rect 7616 4100 8852 4128
rect 7616 4088 7622 4100
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 9030 4088 9036 4140
rect 9088 4088 9094 4140
rect 9306 4128 9312 4140
rect 9267 4100 9312 4128
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 10597 4131 10655 4137
rect 10597 4097 10609 4131
rect 10643 4128 10655 4131
rect 10870 4128 10876 4140
rect 10643 4100 10876 4128
rect 10643 4097 10655 4100
rect 10597 4091 10655 4097
rect 10870 4088 10876 4100
rect 10928 4088 10934 4140
rect 10962 4088 10968 4140
rect 11020 4128 11026 4140
rect 15197 4131 15255 4137
rect 11020 4100 11065 4128
rect 11020 4088 11026 4100
rect 15197 4097 15209 4131
rect 15243 4128 15255 4131
rect 16592 4128 16620 4227
rect 16850 4224 16856 4236
rect 16908 4224 16914 4276
rect 19199 4267 19257 4273
rect 19199 4264 19211 4267
rect 16960 4236 19211 4264
rect 16666 4156 16672 4208
rect 16724 4196 16730 4208
rect 16960 4196 16988 4236
rect 19199 4233 19211 4236
rect 19245 4233 19257 4267
rect 19199 4227 19257 4233
rect 17494 4196 17500 4208
rect 16724 4168 16988 4196
rect 17455 4168 17500 4196
rect 16724 4156 16730 4168
rect 17494 4156 17500 4168
rect 17552 4156 17558 4208
rect 15243 4100 16620 4128
rect 17221 4131 17279 4137
rect 15243 4097 15255 4100
rect 15197 4091 15255 4097
rect 17221 4097 17233 4131
rect 17267 4128 17279 4131
rect 19334 4128 19340 4140
rect 17267 4100 19340 4128
rect 17267 4097 17279 4100
rect 17221 4091 17279 4097
rect 5834 4032 6316 4060
rect 12437 4063 12495 4069
rect 5834 4029 5846 4032
rect 5788 4023 5846 4029
rect 12437 4029 12449 4063
rect 12483 4060 12495 4063
rect 13446 4060 13452 4072
rect 12483 4032 13452 4060
rect 12483 4029 12495 4032
rect 12437 4023 12495 4029
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 16574 4020 16580 4072
rect 16632 4060 16638 4072
rect 16736 4063 16794 4069
rect 16736 4060 16748 4063
rect 16632 4032 16748 4060
rect 16632 4020 16638 4032
rect 16736 4029 16748 4032
rect 16782 4060 16794 4063
rect 17236 4060 17264 4091
rect 19334 4088 19340 4100
rect 19392 4088 19398 4140
rect 16782 4032 17264 4060
rect 16782 4029 16794 4032
rect 16736 4023 16794 4029
rect 17678 4020 17684 4072
rect 17736 4060 17742 4072
rect 18084 4063 18142 4069
rect 18084 4060 18096 4063
rect 17736 4032 18096 4060
rect 17736 4020 17742 4032
rect 18084 4029 18096 4032
rect 18130 4060 18142 4063
rect 18509 4063 18567 4069
rect 18509 4060 18521 4063
rect 18130 4032 18521 4060
rect 18130 4029 18142 4032
rect 18084 4023 18142 4029
rect 18509 4029 18521 4032
rect 18555 4029 18567 4063
rect 19096 4063 19154 4069
rect 19096 4060 19108 4063
rect 18509 4023 18567 4029
rect 18616 4032 19108 4060
rect 5997 3995 6055 4001
rect 5997 3961 6009 3995
rect 6043 3992 6055 3995
rect 7558 3992 7564 4004
rect 6043 3964 7190 3992
rect 7519 3964 7564 3992
rect 6043 3961 6055 3964
rect 5997 3955 6055 3961
rect 6822 3884 6828 3936
rect 6880 3924 6886 3936
rect 7009 3927 7067 3933
rect 7009 3924 7021 3927
rect 6880 3896 7021 3924
rect 6880 3884 6886 3896
rect 7009 3893 7021 3896
rect 7055 3893 7067 3927
rect 7162 3924 7190 3964
rect 7558 3952 7564 3964
rect 7616 3952 7622 4004
rect 7650 3952 7656 4004
rect 7708 3992 7714 4004
rect 8113 3995 8171 4001
rect 8113 3992 8125 3995
rect 7708 3964 8125 3992
rect 7708 3952 7714 3964
rect 8113 3961 8125 3964
rect 8159 3961 8171 3995
rect 9030 3992 9036 4004
rect 8991 3964 9036 3992
rect 8113 3955 8171 3961
rect 9030 3952 9036 3964
rect 9088 3952 9094 4004
rect 9125 3995 9183 4001
rect 9125 3961 9137 3995
rect 9171 3961 9183 3995
rect 9125 3955 9183 3961
rect 8754 3924 8760 3936
rect 7162 3896 8760 3924
rect 7009 3887 7067 3893
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 8846 3884 8852 3936
rect 8904 3924 8910 3936
rect 9140 3924 9168 3955
rect 10042 3952 10048 4004
rect 10100 3992 10106 4004
rect 10689 3995 10747 4001
rect 10689 3992 10701 3995
rect 10100 3964 10701 3992
rect 10100 3952 10106 3964
rect 10689 3961 10701 3964
rect 10735 3961 10747 3995
rect 10689 3955 10747 3961
rect 11885 3995 11943 4001
rect 11885 3961 11897 3995
rect 11931 3992 11943 3995
rect 12250 3992 12256 4004
rect 11931 3964 12256 3992
rect 11931 3961 11943 3964
rect 11885 3955 11943 3961
rect 8904 3896 9168 3924
rect 9953 3927 10011 3933
rect 8904 3884 8910 3896
rect 9953 3893 9965 3927
rect 9999 3924 10011 3927
rect 11900 3924 11928 3955
rect 12250 3952 12256 3964
rect 12308 3992 12314 4004
rect 12799 3995 12857 4001
rect 12799 3992 12811 3995
rect 12308 3964 12811 3992
rect 12308 3952 12314 3964
rect 12799 3961 12811 3964
rect 12845 3992 12857 3995
rect 14734 3992 14740 4004
rect 12845 3964 14740 3992
rect 12845 3961 12857 3964
rect 12799 3955 12857 3961
rect 14734 3952 14740 3964
rect 14792 3952 14798 4004
rect 15289 3995 15347 4001
rect 15289 3961 15301 3995
rect 15335 3992 15347 3995
rect 15378 3992 15384 4004
rect 15335 3964 15384 3992
rect 15335 3961 15347 3964
rect 15289 3955 15347 3961
rect 9999 3896 11928 3924
rect 9999 3893 10011 3896
rect 9953 3887 10011 3893
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 13357 3927 13415 3933
rect 13357 3924 13369 3927
rect 12492 3896 13369 3924
rect 12492 3884 12498 3896
rect 13357 3893 13369 3896
rect 13403 3893 13415 3927
rect 13357 3887 13415 3893
rect 15013 3927 15071 3933
rect 15013 3893 15025 3927
rect 15059 3924 15071 3927
rect 15304 3924 15332 3955
rect 15378 3952 15384 3964
rect 15436 3952 15442 4004
rect 15838 3992 15844 4004
rect 15799 3964 15844 3992
rect 15838 3952 15844 3964
rect 15896 3952 15902 4004
rect 16298 3952 16304 4004
rect 16356 3992 16362 4004
rect 18616 3992 18644 4032
rect 19096 4029 19108 4032
rect 19142 4060 19154 4063
rect 19521 4063 19579 4069
rect 19521 4060 19533 4063
rect 19142 4032 19533 4060
rect 19142 4029 19154 4032
rect 19096 4023 19154 4029
rect 19521 4029 19533 4032
rect 19567 4029 19579 4063
rect 19521 4023 19579 4029
rect 16356 3964 18644 3992
rect 16356 3952 16362 3964
rect 16114 3924 16120 3936
rect 15059 3896 15332 3924
rect 16075 3896 16120 3924
rect 15059 3893 15071 3896
rect 15013 3887 15071 3893
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 16574 3884 16580 3936
rect 16632 3924 16638 3936
rect 16807 3927 16865 3933
rect 16807 3924 16819 3927
rect 16632 3896 16819 3924
rect 16632 3884 16638 3896
rect 16807 3893 16819 3896
rect 16853 3893 16865 3927
rect 16807 3887 16865 3893
rect 17218 3884 17224 3936
rect 17276 3924 17282 3936
rect 18187 3927 18245 3933
rect 18187 3924 18199 3927
rect 17276 3896 18199 3924
rect 17276 3884 17282 3896
rect 18187 3893 18199 3896
rect 18233 3893 18245 3927
rect 18187 3887 18245 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 5721 3723 5779 3729
rect 5721 3720 5733 3723
rect 3936 3692 5733 3720
rect 3936 3680 3942 3692
rect 5721 3689 5733 3692
rect 5767 3720 5779 3723
rect 5994 3720 6000 3732
rect 5767 3692 6000 3720
rect 5767 3689 5779 3692
rect 5721 3683 5779 3689
rect 5994 3680 6000 3692
rect 6052 3680 6058 3732
rect 7558 3720 7564 3732
rect 7519 3692 7564 3720
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 9030 3720 9036 3732
rect 8991 3692 9036 3720
rect 9030 3680 9036 3692
rect 9088 3680 9094 3732
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 9861 3723 9919 3729
rect 9861 3720 9873 3723
rect 9732 3692 9873 3720
rect 9732 3680 9738 3692
rect 9861 3689 9873 3692
rect 9907 3689 9919 3723
rect 12434 3720 12440 3732
rect 9861 3683 9919 3689
rect 10704 3692 12440 3720
rect 8110 3612 8116 3664
rect 8168 3652 8174 3664
rect 8205 3655 8263 3661
rect 8205 3652 8217 3655
rect 8168 3624 8217 3652
rect 8168 3612 8174 3624
rect 8205 3621 8217 3624
rect 8251 3621 8263 3655
rect 8205 3615 8263 3621
rect 8754 3612 8760 3664
rect 8812 3652 8818 3664
rect 8812 3624 9812 3652
rect 8812 3612 8818 3624
rect 5052 3587 5110 3593
rect 5052 3553 5064 3587
rect 5098 3584 5110 3587
rect 5442 3584 5448 3596
rect 5098 3556 5448 3584
rect 5098 3553 5110 3556
rect 5052 3547 5110 3553
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 6064 3587 6122 3593
rect 6064 3553 6076 3587
rect 6110 3584 6122 3587
rect 6270 3584 6276 3596
rect 6110 3556 6276 3584
rect 6110 3553 6122 3556
rect 6064 3547 6122 3553
rect 6270 3544 6276 3556
rect 6328 3544 6334 3596
rect 6638 3544 6644 3596
rect 6696 3584 6702 3596
rect 7044 3587 7102 3593
rect 7044 3584 7056 3587
rect 6696 3556 7056 3584
rect 6696 3544 6702 3556
rect 7044 3553 7056 3556
rect 7090 3553 7102 3587
rect 7044 3547 7102 3553
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3485 8171 3519
rect 8113 3479 8171 3485
rect 8757 3519 8815 3525
rect 8757 3485 8769 3519
rect 8803 3516 8815 3519
rect 8846 3516 8852 3528
rect 8803 3488 8852 3516
rect 8803 3485 8815 3488
rect 8757 3479 8815 3485
rect 5123 3451 5181 3457
rect 5123 3417 5135 3451
rect 5169 3448 5181 3451
rect 5718 3448 5724 3460
rect 5169 3420 5724 3448
rect 5169 3417 5181 3420
rect 5123 3411 5181 3417
rect 5718 3408 5724 3420
rect 5776 3408 5782 3460
rect 7147 3451 7205 3457
rect 7147 3417 7159 3451
rect 7193 3448 7205 3451
rect 7837 3451 7895 3457
rect 7837 3448 7849 3451
rect 7193 3420 7849 3448
rect 7193 3417 7205 3420
rect 7147 3411 7205 3417
rect 7837 3417 7849 3420
rect 7883 3448 7895 3451
rect 8128 3448 8156 3479
rect 8846 3476 8852 3488
rect 8904 3516 8910 3528
rect 9306 3516 9312 3528
rect 8904 3488 9312 3516
rect 8904 3476 8910 3488
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 7883 3420 8156 3448
rect 9784 3448 9812 3624
rect 10318 3612 10324 3664
rect 10376 3652 10382 3664
rect 10704 3661 10732 3692
rect 12434 3680 12440 3692
rect 12492 3680 12498 3732
rect 13173 3723 13231 3729
rect 13173 3689 13185 3723
rect 13219 3720 13231 3723
rect 13446 3720 13452 3732
rect 13219 3692 13452 3720
rect 13219 3689 13231 3692
rect 13173 3683 13231 3689
rect 13446 3680 13452 3692
rect 13504 3680 13510 3732
rect 14090 3720 14096 3732
rect 13740 3692 14096 3720
rect 10689 3655 10747 3661
rect 10689 3652 10701 3655
rect 10376 3624 10701 3652
rect 10376 3612 10382 3624
rect 10689 3621 10701 3624
rect 10735 3621 10747 3655
rect 11238 3652 11244 3664
rect 11199 3624 11244 3652
rect 10689 3615 10747 3621
rect 11238 3612 11244 3624
rect 11296 3612 11302 3664
rect 11882 3612 11888 3664
rect 11940 3652 11946 3664
rect 12253 3655 12311 3661
rect 12253 3652 12265 3655
rect 11940 3624 12265 3652
rect 11940 3612 11946 3624
rect 12253 3621 12265 3624
rect 12299 3652 12311 3655
rect 12526 3652 12532 3664
rect 12299 3624 12532 3652
rect 12299 3621 12311 3624
rect 12253 3615 12311 3621
rect 12526 3612 12532 3624
rect 12584 3612 12590 3664
rect 13740 3661 13768 3692
rect 14090 3680 14096 3692
rect 14148 3720 14154 3732
rect 14148 3692 16068 3720
rect 14148 3680 14154 3692
rect 13725 3655 13783 3661
rect 13725 3621 13737 3655
rect 13771 3621 13783 3655
rect 13725 3615 13783 3621
rect 13814 3612 13820 3664
rect 13872 3652 13878 3664
rect 15470 3652 15476 3664
rect 13872 3624 13917 3652
rect 15431 3624 15476 3652
rect 13872 3612 13878 3624
rect 15470 3612 15476 3624
rect 15528 3612 15534 3664
rect 16040 3584 16068 3692
rect 16482 3680 16488 3732
rect 16540 3720 16546 3732
rect 16761 3723 16819 3729
rect 16761 3720 16773 3723
rect 16540 3692 16773 3720
rect 16540 3680 16546 3692
rect 16761 3689 16773 3692
rect 16807 3720 16819 3723
rect 17218 3720 17224 3732
rect 16807 3692 17224 3720
rect 16807 3689 16819 3692
rect 16761 3683 16819 3689
rect 17218 3680 17224 3692
rect 17276 3680 17282 3732
rect 16206 3612 16212 3664
rect 16264 3652 16270 3664
rect 17037 3655 17095 3661
rect 17037 3652 17049 3655
rect 16264 3624 17049 3652
rect 16264 3612 16270 3624
rect 17037 3621 17049 3624
rect 17083 3652 17095 3655
rect 17402 3652 17408 3664
rect 17083 3624 17408 3652
rect 17083 3621 17095 3624
rect 17037 3615 17095 3621
rect 17402 3612 17408 3624
rect 17460 3612 17466 3664
rect 17589 3655 17647 3661
rect 17589 3621 17601 3655
rect 17635 3652 17647 3655
rect 17770 3652 17776 3664
rect 17635 3624 17776 3652
rect 17635 3621 17647 3624
rect 17589 3615 17647 3621
rect 17770 3612 17776 3624
rect 17828 3612 17834 3664
rect 18598 3652 18604 3664
rect 18559 3624 18604 3652
rect 18598 3612 18604 3624
rect 18656 3612 18662 3664
rect 16666 3584 16672 3596
rect 16040 3556 16672 3584
rect 16666 3544 16672 3556
rect 16724 3544 16730 3596
rect 10413 3519 10471 3525
rect 10413 3485 10425 3519
rect 10459 3516 10471 3519
rect 10597 3519 10655 3525
rect 10597 3516 10609 3519
rect 10459 3488 10609 3516
rect 10459 3485 10471 3488
rect 10413 3479 10471 3485
rect 10597 3485 10609 3488
rect 10643 3516 10655 3519
rect 11238 3516 11244 3528
rect 10643 3488 11244 3516
rect 10643 3485 10655 3488
rect 10597 3479 10655 3485
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 12161 3519 12219 3525
rect 12161 3485 12173 3519
rect 12207 3485 12219 3519
rect 13998 3516 14004 3528
rect 13959 3488 14004 3516
rect 12161 3479 12219 3485
rect 11974 3448 11980 3460
rect 9784 3420 11980 3448
rect 7883 3417 7895 3420
rect 7837 3411 7895 3417
rect 11974 3408 11980 3420
rect 12032 3448 12038 3460
rect 12176 3448 12204 3479
rect 13998 3476 14004 3488
rect 14056 3476 14062 3528
rect 15381 3519 15439 3525
rect 15381 3485 15393 3519
rect 15427 3485 15439 3519
rect 15838 3516 15844 3528
rect 15799 3488 15844 3516
rect 15381 3479 15439 3485
rect 12710 3448 12716 3460
rect 12032 3420 12204 3448
rect 12671 3420 12716 3448
rect 12032 3408 12038 3420
rect 12710 3408 12716 3420
rect 12768 3408 12774 3460
rect 15396 3448 15424 3479
rect 15838 3476 15844 3488
rect 15896 3516 15902 3528
rect 16758 3516 16764 3528
rect 15896 3488 16764 3516
rect 15896 3476 15902 3488
rect 16758 3476 16764 3488
rect 16816 3516 16822 3528
rect 16945 3519 17003 3525
rect 16945 3516 16957 3519
rect 16816 3488 16957 3516
rect 16816 3476 16822 3488
rect 16945 3485 16957 3488
rect 16991 3485 17003 3519
rect 18506 3516 18512 3528
rect 18467 3488 18512 3516
rect 16945 3479 17003 3485
rect 18506 3476 18512 3488
rect 18564 3476 18570 3528
rect 18785 3519 18843 3525
rect 18785 3516 18797 3519
rect 18616 3488 18797 3516
rect 15396 3420 16436 3448
rect 16408 3392 16436 3420
rect 17126 3408 17132 3460
rect 17184 3448 17190 3460
rect 17957 3451 18015 3457
rect 17957 3448 17969 3451
rect 17184 3420 17969 3448
rect 17184 3408 17190 3420
rect 17957 3417 17969 3420
rect 18003 3448 18015 3451
rect 18616 3448 18644 3488
rect 18785 3485 18797 3488
rect 18831 3485 18843 3519
rect 18785 3479 18843 3485
rect 18003 3420 18644 3448
rect 18003 3417 18015 3420
rect 17957 3411 18015 3417
rect 6135 3383 6193 3389
rect 6135 3349 6147 3383
rect 6181 3380 6193 3383
rect 6825 3383 6883 3389
rect 6825 3380 6837 3383
rect 6181 3352 6837 3380
rect 6181 3349 6193 3352
rect 6135 3343 6193 3349
rect 6825 3349 6837 3352
rect 6871 3380 6883 3383
rect 6914 3380 6920 3392
rect 6871 3352 6920 3380
rect 6871 3349 6883 3352
rect 6825 3343 6883 3349
rect 6914 3340 6920 3352
rect 6972 3340 6978 3392
rect 8570 3340 8576 3392
rect 8628 3380 8634 3392
rect 9401 3383 9459 3389
rect 9401 3380 9413 3383
rect 8628 3352 9413 3380
rect 8628 3340 8634 3352
rect 9401 3349 9413 3352
rect 9447 3349 9459 3383
rect 9401 3343 9459 3349
rect 14550 3340 14556 3392
rect 14608 3380 14614 3392
rect 14829 3383 14887 3389
rect 14829 3380 14841 3383
rect 14608 3352 14841 3380
rect 14608 3340 14614 3352
rect 14829 3349 14841 3352
rect 14875 3349 14887 3383
rect 16390 3380 16396 3392
rect 16351 3352 16396 3380
rect 14829 3343 14887 3349
rect 16390 3340 16396 3352
rect 16448 3340 16454 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 4246 3176 4252 3188
rect 4207 3148 4252 3176
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 4847 3179 4905 3185
rect 4847 3145 4859 3179
rect 4893 3176 4905 3179
rect 7745 3179 7803 3185
rect 7745 3176 7757 3179
rect 4893 3148 7757 3176
rect 4893 3145 4905 3148
rect 4847 3139 4905 3145
rect 7745 3145 7757 3148
rect 7791 3145 7803 3179
rect 7745 3139 7803 3145
rect 8021 3179 8079 3185
rect 8021 3145 8033 3179
rect 8067 3176 8079 3179
rect 8110 3176 8116 3188
rect 8067 3148 8116 3176
rect 8067 3145 8079 3148
rect 8021 3139 8079 3145
rect 8110 3136 8116 3148
rect 8168 3176 8174 3188
rect 8297 3179 8355 3185
rect 8297 3176 8309 3179
rect 8168 3148 8309 3176
rect 8168 3136 8174 3148
rect 8297 3145 8309 3148
rect 8343 3145 8355 3179
rect 10318 3176 10324 3188
rect 10279 3148 10324 3176
rect 8297 3139 8355 3145
rect 10318 3136 10324 3148
rect 10376 3136 10382 3188
rect 11882 3176 11888 3188
rect 11843 3148 11888 3176
rect 11882 3136 11888 3148
rect 11940 3136 11946 3188
rect 12253 3179 12311 3185
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 12342 3176 12348 3188
rect 12299 3148 12348 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 12342 3136 12348 3148
rect 12400 3136 12406 3188
rect 12526 3136 12532 3188
rect 12584 3176 12590 3188
rect 13633 3179 13691 3185
rect 13633 3176 13645 3179
rect 12584 3148 13645 3176
rect 12584 3136 12590 3148
rect 13633 3145 13645 3148
rect 13679 3176 13691 3179
rect 13814 3176 13820 3188
rect 13679 3148 13820 3176
rect 13679 3145 13691 3148
rect 13633 3139 13691 3145
rect 13814 3136 13820 3148
rect 13872 3136 13878 3188
rect 15470 3136 15476 3188
rect 15528 3176 15534 3188
rect 15654 3176 15660 3188
rect 15528 3148 15660 3176
rect 15528 3136 15534 3148
rect 15654 3136 15660 3148
rect 15712 3176 15718 3188
rect 15841 3179 15899 3185
rect 15841 3176 15853 3179
rect 15712 3148 15853 3176
rect 15712 3136 15718 3148
rect 15841 3145 15853 3148
rect 15887 3145 15899 3179
rect 17402 3176 17408 3188
rect 17363 3148 17408 3176
rect 15841 3139 15899 3145
rect 17402 3136 17408 3148
rect 17460 3136 17466 3188
rect 17865 3179 17923 3185
rect 17865 3145 17877 3179
rect 17911 3176 17923 3179
rect 18187 3179 18245 3185
rect 18187 3176 18199 3179
rect 17911 3148 18199 3176
rect 17911 3145 17923 3148
rect 17865 3139 17923 3145
rect 18187 3145 18199 3148
rect 18233 3176 18245 3179
rect 18506 3176 18512 3188
rect 18233 3148 18512 3176
rect 18233 3145 18245 3148
rect 18187 3139 18245 3145
rect 18506 3136 18512 3148
rect 18564 3136 18570 3188
rect 5859 3111 5917 3117
rect 5859 3077 5871 3111
rect 5905 3108 5917 3111
rect 7926 3108 7932 3120
rect 5905 3080 7932 3108
rect 5905 3077 5917 3080
rect 5859 3071 5917 3077
rect 7926 3068 7932 3080
rect 7984 3068 7990 3120
rect 8386 3068 8392 3120
rect 8444 3108 8450 3120
rect 8444 3080 9674 3108
rect 8444 3068 8450 3080
rect 6270 3040 6276 3052
rect 6231 3012 6276 3040
rect 6270 3000 6276 3012
rect 6328 3000 6334 3052
rect 7006 3040 7012 3052
rect 6967 3012 7012 3040
rect 7006 3000 7012 3012
rect 7064 3000 7070 3052
rect 7650 3040 7656 3052
rect 7611 3012 7656 3040
rect 7650 3000 7656 3012
rect 7708 3040 7714 3052
rect 8849 3043 8907 3049
rect 8849 3040 8861 3043
rect 7708 3012 8861 3040
rect 7708 3000 7714 3012
rect 8849 3009 8861 3012
rect 8895 3040 8907 3043
rect 9214 3040 9220 3052
rect 8895 3012 9220 3040
rect 8895 3009 8907 3012
rect 8849 3003 8907 3009
rect 9214 3000 9220 3012
rect 9272 3000 9278 3052
rect 3748 2975 3806 2981
rect 3748 2941 3760 2975
rect 3794 2972 3806 2975
rect 4062 2972 4068 2984
rect 3794 2944 4068 2972
rect 3794 2941 3806 2944
rect 3748 2935 3806 2941
rect 4062 2932 4068 2944
rect 4120 2972 4126 2984
rect 4246 2972 4252 2984
rect 4120 2944 4252 2972
rect 4120 2932 4126 2944
rect 4246 2932 4252 2944
rect 4304 2932 4310 2984
rect 4776 2975 4834 2981
rect 4776 2941 4788 2975
rect 4822 2972 4834 2975
rect 5788 2975 5846 2981
rect 4822 2944 5304 2972
rect 4822 2941 4834 2944
rect 4776 2935 4834 2941
rect 3835 2907 3893 2913
rect 3835 2873 3847 2907
rect 3881 2904 3893 2907
rect 5166 2904 5172 2916
rect 3881 2876 5172 2904
rect 3881 2873 3893 2876
rect 3835 2867 3893 2873
rect 5166 2864 5172 2876
rect 5224 2864 5230 2916
rect 5276 2848 5304 2944
rect 5788 2941 5800 2975
rect 5834 2972 5846 2975
rect 5994 2972 6000 2984
rect 5834 2944 6000 2972
rect 5834 2941 5846 2944
rect 5788 2935 5846 2941
rect 5994 2932 6000 2944
rect 6052 2932 6058 2984
rect 7745 2975 7803 2981
rect 7745 2941 7757 2975
rect 7791 2972 7803 2975
rect 8386 2972 8392 2984
rect 7791 2944 8392 2972
rect 7791 2941 7803 2944
rect 7745 2935 7803 2941
rect 8386 2932 8392 2944
rect 8444 2932 8450 2984
rect 7101 2907 7159 2913
rect 7101 2873 7113 2907
rect 7147 2873 7159 2907
rect 8570 2904 8576 2916
rect 8531 2876 8576 2904
rect 7101 2867 7159 2873
rect 5258 2836 5264 2848
rect 5219 2808 5264 2836
rect 5258 2796 5264 2808
rect 5316 2796 5322 2848
rect 5442 2796 5448 2848
rect 5500 2836 5506 2848
rect 5629 2839 5687 2845
rect 5629 2836 5641 2839
rect 5500 2808 5641 2836
rect 5500 2796 5506 2808
rect 5629 2805 5641 2808
rect 5675 2836 5687 2839
rect 5994 2836 6000 2848
rect 5675 2808 6000 2836
rect 5675 2805 5687 2808
rect 5629 2799 5687 2805
rect 5994 2796 6000 2808
rect 6052 2796 6058 2848
rect 6638 2836 6644 2848
rect 6599 2808 6644 2836
rect 6638 2796 6644 2808
rect 6696 2796 6702 2848
rect 7116 2836 7144 2867
rect 8570 2864 8576 2876
rect 8628 2864 8634 2916
rect 8674 2907 8732 2913
rect 8674 2873 8686 2907
rect 8720 2873 8732 2907
rect 9646 2904 9674 3080
rect 12066 3068 12072 3120
rect 12124 3108 12130 3120
rect 14001 3111 14059 3117
rect 14001 3108 14013 3111
rect 12124 3080 14013 3108
rect 12124 3068 12130 3080
rect 14001 3077 14013 3080
rect 14047 3077 14059 3111
rect 14001 3071 14059 3077
rect 15746 3068 15752 3120
rect 15804 3108 15810 3120
rect 16209 3111 16267 3117
rect 16209 3108 16221 3111
rect 15804 3080 16221 3108
rect 15804 3068 15810 3080
rect 16209 3077 16221 3080
rect 16255 3077 16267 3111
rect 16209 3071 16267 3077
rect 11517 3043 11575 3049
rect 11517 3009 11529 3043
rect 11563 3040 11575 3043
rect 12710 3040 12716 3052
rect 11563 3012 12716 3040
rect 11563 3009 11575 3012
rect 11517 3003 11575 3009
rect 12710 3000 12716 3012
rect 12768 3040 12774 3052
rect 12805 3043 12863 3049
rect 12805 3040 12817 3043
rect 12768 3012 12817 3040
rect 12768 3000 12774 3012
rect 12805 3009 12817 3012
rect 12851 3009 12863 3043
rect 12805 3003 12863 3009
rect 9861 2907 9919 2913
rect 9861 2904 9873 2907
rect 9646 2876 9873 2904
rect 8674 2867 8732 2873
rect 9861 2873 9873 2876
rect 9907 2904 9919 2907
rect 10873 2907 10931 2913
rect 10873 2904 10885 2907
rect 9907 2876 10885 2904
rect 9907 2873 9919 2876
rect 9861 2867 9919 2873
rect 10873 2873 10885 2876
rect 10919 2873 10931 2907
rect 10873 2867 10931 2873
rect 10965 2907 11023 2913
rect 10965 2873 10977 2907
rect 11011 2904 11023 2907
rect 11330 2904 11336 2916
rect 11011 2876 11336 2904
rect 11011 2873 11023 2876
rect 10965 2867 11023 2873
rect 8110 2836 8116 2848
rect 7116 2808 8116 2836
rect 8110 2796 8116 2808
rect 8168 2796 8174 2848
rect 8680 2836 8708 2867
rect 8754 2836 8760 2848
rect 8680 2808 8760 2836
rect 8754 2796 8760 2808
rect 8812 2836 8818 2848
rect 9493 2839 9551 2845
rect 9493 2836 9505 2839
rect 8812 2808 9505 2836
rect 8812 2796 8818 2808
rect 9493 2805 9505 2808
rect 9539 2805 9551 2839
rect 9493 2799 9551 2805
rect 10689 2839 10747 2845
rect 10689 2805 10701 2839
rect 10735 2836 10747 2839
rect 10778 2836 10784 2848
rect 10735 2808 10784 2836
rect 10735 2805 10747 2808
rect 10689 2799 10747 2805
rect 10778 2796 10784 2808
rect 10836 2836 10842 2848
rect 10980 2836 11008 2867
rect 11330 2864 11336 2876
rect 11388 2864 11394 2916
rect 12066 2864 12072 2916
rect 12124 2904 12130 2916
rect 12529 2907 12587 2913
rect 12529 2904 12541 2907
rect 12124 2876 12541 2904
rect 12124 2864 12130 2876
rect 12529 2873 12541 2876
rect 12575 2873 12587 2907
rect 12529 2867 12587 2873
rect 12618 2864 12624 2916
rect 12676 2904 12682 2916
rect 12676 2876 12721 2904
rect 12676 2864 12682 2876
rect 14550 2864 14556 2916
rect 14608 2904 14614 2916
rect 14921 2907 14979 2913
rect 14921 2904 14933 2907
rect 14608 2876 14933 2904
rect 14608 2864 14614 2876
rect 14921 2873 14933 2876
rect 14967 2873 14979 2907
rect 14921 2867 14979 2873
rect 15013 2907 15071 2913
rect 15013 2873 15025 2907
rect 15059 2904 15071 2907
rect 15378 2904 15384 2916
rect 15059 2876 15384 2904
rect 15059 2873 15071 2876
rect 15013 2867 15071 2873
rect 10836 2808 11008 2836
rect 14737 2839 14795 2845
rect 10836 2796 10842 2808
rect 14737 2805 14749 2839
rect 14783 2836 14795 2839
rect 15028 2836 15056 2867
rect 15378 2864 15384 2876
rect 15436 2864 15442 2916
rect 15565 2907 15623 2913
rect 15565 2873 15577 2907
rect 15611 2904 15623 2907
rect 16114 2904 16120 2916
rect 15611 2876 16120 2904
rect 15611 2873 15623 2876
rect 15565 2867 15623 2873
rect 16114 2864 16120 2876
rect 16172 2864 16178 2916
rect 16224 2904 16252 3071
rect 16390 3068 16396 3120
rect 16448 3108 16454 3120
rect 19199 3111 19257 3117
rect 19199 3108 19211 3111
rect 16448 3080 19211 3108
rect 16448 3068 16454 3080
rect 19199 3077 19211 3080
rect 19245 3077 19257 3111
rect 19199 3071 19257 3077
rect 20625 3111 20683 3117
rect 20625 3077 20637 3111
rect 20671 3108 20683 3111
rect 22094 3108 22100 3120
rect 20671 3080 22100 3108
rect 20671 3077 20683 3080
rect 20625 3071 20683 3077
rect 22094 3068 22100 3080
rect 22152 3068 22158 3120
rect 16482 3040 16488 3052
rect 16443 3012 16488 3040
rect 16482 3000 16488 3012
rect 16540 3000 16546 3052
rect 16758 3040 16764 3052
rect 16719 3012 16764 3040
rect 16758 3000 16764 3012
rect 16816 3000 16822 3052
rect 18601 3043 18659 3049
rect 18601 3009 18613 3043
rect 18647 3040 18659 3043
rect 18647 3012 23474 3040
rect 18647 3009 18659 3012
rect 18601 3003 18659 3009
rect 17954 2932 17960 2984
rect 18012 2972 18018 2984
rect 18116 2975 18174 2981
rect 18116 2972 18128 2975
rect 18012 2944 18128 2972
rect 18012 2932 18018 2944
rect 18116 2941 18128 2944
rect 18162 2972 18174 2975
rect 18616 2972 18644 3003
rect 18162 2944 18644 2972
rect 19128 2975 19186 2981
rect 18162 2941 18174 2944
rect 18116 2935 18174 2941
rect 19128 2941 19140 2975
rect 19174 2972 19186 2975
rect 19518 2972 19524 2984
rect 19174 2944 19524 2972
rect 19174 2941 19186 2944
rect 19128 2935 19186 2941
rect 19518 2932 19524 2944
rect 19576 2932 19582 2984
rect 20438 2972 20444 2984
rect 20399 2944 20444 2972
rect 20438 2932 20444 2944
rect 20496 2972 20502 2984
rect 20993 2975 21051 2981
rect 20993 2972 21005 2975
rect 20496 2944 21005 2972
rect 20496 2932 20502 2944
rect 20993 2941 21005 2944
rect 21039 2941 21051 2975
rect 23446 2972 23474 3012
rect 23661 2975 23719 2981
rect 23661 2972 23673 2975
rect 23446 2944 23673 2972
rect 20993 2935 21051 2941
rect 23661 2941 23673 2944
rect 23707 2972 23719 2975
rect 24213 2975 24271 2981
rect 24213 2972 24225 2975
rect 23707 2944 24225 2972
rect 23707 2941 23719 2944
rect 23661 2935 23719 2941
rect 24213 2941 24225 2944
rect 24259 2941 24271 2975
rect 24213 2935 24271 2941
rect 16577 2907 16635 2913
rect 16577 2904 16589 2907
rect 16224 2876 16589 2904
rect 16577 2873 16589 2876
rect 16623 2904 16635 2907
rect 18598 2904 18604 2916
rect 16623 2876 18604 2904
rect 16623 2873 16635 2876
rect 16577 2867 16635 2873
rect 18598 2864 18604 2876
rect 18656 2904 18662 2916
rect 18877 2907 18935 2913
rect 18877 2904 18889 2907
rect 18656 2876 18889 2904
rect 18656 2864 18662 2876
rect 18877 2873 18889 2876
rect 18923 2873 18935 2907
rect 18877 2867 18935 2873
rect 14783 2808 15056 2836
rect 14783 2805 14795 2808
rect 14737 2799 14795 2805
rect 16206 2796 16212 2848
rect 16264 2836 16270 2848
rect 18138 2836 18144 2848
rect 16264 2808 18144 2836
rect 16264 2796 16270 2808
rect 18138 2796 18144 2808
rect 18196 2796 18202 2848
rect 23845 2839 23903 2845
rect 23845 2805 23857 2839
rect 23891 2836 23903 2839
rect 25498 2836 25504 2848
rect 23891 2808 25504 2836
rect 23891 2805 23903 2808
rect 23845 2799 23903 2805
rect 25498 2796 25504 2808
rect 25556 2796 25562 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 3099 2635 3157 2641
rect 3099 2601 3111 2635
rect 3145 2632 3157 2635
rect 5534 2632 5540 2644
rect 3145 2604 5540 2632
rect 3145 2601 3157 2604
rect 3099 2595 3157 2601
rect 5534 2592 5540 2604
rect 5592 2592 5598 2644
rect 5951 2635 6009 2641
rect 5951 2601 5963 2635
rect 5997 2632 6009 2635
rect 7098 2632 7104 2644
rect 5997 2604 7104 2632
rect 5997 2601 6009 2604
rect 5951 2595 6009 2601
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 7377 2635 7435 2641
rect 7377 2632 7389 2635
rect 7248 2604 7389 2632
rect 7248 2592 7254 2604
rect 7377 2601 7389 2604
rect 7423 2601 7435 2635
rect 9030 2632 9036 2644
rect 7377 2595 7435 2601
rect 7576 2604 9036 2632
rect 6365 2567 6423 2573
rect 6365 2564 6377 2567
rect 5895 2536 6377 2564
rect 3028 2499 3086 2505
rect 3028 2465 3040 2499
rect 3074 2496 3086 2499
rect 4868 2499 4926 2505
rect 3074 2468 3556 2496
rect 3074 2465 3086 2468
rect 3028 2459 3086 2465
rect 3528 2369 3556 2468
rect 4868 2465 4880 2499
rect 4914 2496 4926 2499
rect 5442 2496 5448 2508
rect 4914 2468 5448 2496
rect 4914 2465 4926 2468
rect 4868 2459 4926 2465
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 5895 2505 5923 2536
rect 6365 2533 6377 2536
rect 6411 2564 6423 2567
rect 7576 2564 7604 2604
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 10778 2632 10784 2644
rect 10739 2604 10784 2632
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 11974 2632 11980 2644
rect 11935 2604 11980 2632
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 12342 2632 12348 2644
rect 12303 2604 12348 2632
rect 12342 2592 12348 2604
rect 12400 2592 12406 2644
rect 14090 2632 14096 2644
rect 14051 2604 14096 2632
rect 14090 2592 14096 2604
rect 14148 2592 14154 2644
rect 14507 2635 14565 2641
rect 14507 2601 14519 2635
rect 14553 2632 14565 2635
rect 18601 2635 18659 2641
rect 14553 2604 17172 2632
rect 14553 2601 14565 2604
rect 14507 2595 14565 2601
rect 6411 2536 7604 2564
rect 6411 2533 6423 2536
rect 6365 2527 6423 2533
rect 7742 2524 7748 2576
rect 7800 2564 7806 2576
rect 8018 2564 8024 2576
rect 7800 2536 8024 2564
rect 7800 2524 7806 2536
rect 8018 2524 8024 2536
rect 8076 2524 8082 2576
rect 8294 2564 8300 2576
rect 8255 2536 8300 2564
rect 8294 2524 8300 2536
rect 8352 2564 8358 2576
rect 8662 2564 8668 2576
rect 8352 2536 8668 2564
rect 8352 2524 8358 2536
rect 8662 2524 8668 2536
rect 8720 2524 8726 2576
rect 8846 2564 8852 2576
rect 8807 2536 8852 2564
rect 8846 2524 8852 2536
rect 8904 2524 8910 2576
rect 9490 2564 9496 2576
rect 9451 2536 9496 2564
rect 9490 2524 9496 2536
rect 9548 2524 9554 2576
rect 10796 2564 10824 2592
rect 11149 2567 11207 2573
rect 11149 2564 11161 2567
rect 10796 2536 11161 2564
rect 11149 2533 11161 2536
rect 11195 2533 11207 2567
rect 11149 2527 11207 2533
rect 12250 2524 12256 2576
rect 12308 2564 12314 2576
rect 12710 2564 12716 2576
rect 12308 2536 12716 2564
rect 12308 2524 12314 2536
rect 12710 2524 12716 2536
rect 12768 2524 12774 2576
rect 12802 2524 12808 2576
rect 12860 2564 12866 2576
rect 15289 2567 15347 2573
rect 12860 2536 12905 2564
rect 12860 2524 12866 2536
rect 15289 2533 15301 2567
rect 15335 2564 15347 2567
rect 15654 2564 15660 2576
rect 15335 2536 15660 2564
rect 15335 2533 15347 2536
rect 15289 2527 15347 2533
rect 15654 2524 15660 2536
rect 15712 2524 15718 2576
rect 16574 2564 16580 2576
rect 16535 2536 16580 2564
rect 16574 2524 16580 2536
rect 16632 2524 16638 2576
rect 16758 2524 16764 2576
rect 16816 2564 16822 2576
rect 16853 2567 16911 2573
rect 16853 2564 16865 2567
rect 16816 2536 16865 2564
rect 16816 2524 16822 2536
rect 16853 2533 16865 2536
rect 16899 2533 16911 2567
rect 16853 2527 16911 2533
rect 5880 2499 5938 2505
rect 5880 2465 5892 2499
rect 5926 2465 5938 2499
rect 5880 2459 5938 2465
rect 7168 2499 7226 2505
rect 7168 2465 7180 2499
rect 7214 2496 7226 2499
rect 7214 2468 7696 2496
rect 7214 2465 7226 2468
rect 7168 2459 7226 2465
rect 3513 2363 3571 2369
rect 3513 2329 3525 2363
rect 3559 2360 3571 2363
rect 7190 2360 7196 2372
rect 3559 2332 7196 2360
rect 3559 2329 3571 2332
rect 3513 2323 3571 2329
rect 7190 2320 7196 2332
rect 7248 2320 7254 2372
rect 7668 2369 7696 2468
rect 7926 2388 7932 2440
rect 7984 2428 7990 2440
rect 8205 2431 8263 2437
rect 8205 2428 8217 2431
rect 7984 2400 8217 2428
rect 7984 2388 7990 2400
rect 8205 2397 8217 2400
rect 8251 2428 8263 2431
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8251 2400 9137 2428
rect 8251 2397 8263 2400
rect 8205 2391 8263 2397
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9508 2428 9536 2524
rect 9582 2456 9588 2508
rect 9640 2496 9646 2508
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 9640 2468 9781 2496
rect 9640 2456 9646 2468
rect 9769 2465 9781 2468
rect 9815 2496 9827 2499
rect 10321 2499 10379 2505
rect 10321 2496 10333 2499
rect 9815 2468 10333 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 10321 2465 10333 2468
rect 10367 2465 10379 2499
rect 10321 2459 10379 2465
rect 14274 2456 14280 2508
rect 14332 2496 14338 2508
rect 14404 2499 14462 2505
rect 14404 2496 14416 2499
rect 14332 2468 14416 2496
rect 14332 2456 14338 2468
rect 14404 2465 14416 2468
rect 14450 2496 14462 2499
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 14450 2468 14841 2496
rect 14450 2465 14462 2468
rect 14404 2459 14462 2465
rect 14829 2465 14841 2468
rect 14875 2465 14887 2499
rect 14829 2459 14887 2465
rect 11057 2431 11115 2437
rect 11057 2428 11069 2431
rect 9508 2400 11069 2428
rect 9125 2391 9183 2397
rect 11057 2397 11069 2400
rect 11103 2397 11115 2431
rect 11057 2391 11115 2397
rect 11238 2388 11244 2440
rect 11296 2428 11302 2440
rect 11333 2431 11391 2437
rect 11333 2428 11345 2431
rect 11296 2400 11345 2428
rect 11296 2388 11302 2400
rect 11333 2397 11345 2400
rect 11379 2428 11391 2431
rect 12989 2431 13047 2437
rect 11379 2400 11928 2428
rect 11379 2397 11391 2400
rect 11333 2391 11391 2397
rect 7653 2363 7711 2369
rect 7653 2329 7665 2363
rect 7699 2360 7711 2363
rect 8110 2360 8116 2372
rect 7699 2332 8116 2360
rect 7699 2329 7711 2332
rect 7653 2323 7711 2329
rect 8110 2320 8116 2332
rect 8168 2320 8174 2372
rect 9953 2363 10011 2369
rect 9953 2329 9965 2363
rect 9999 2360 10011 2363
rect 11514 2360 11520 2372
rect 9999 2332 11520 2360
rect 9999 2329 10011 2332
rect 9953 2323 10011 2329
rect 11514 2320 11520 2332
rect 11572 2320 11578 2372
rect 11900 2360 11928 2400
rect 12989 2397 13001 2431
rect 13035 2428 13047 2431
rect 13998 2428 14004 2440
rect 13035 2400 14004 2428
rect 13035 2397 13047 2400
rect 12989 2391 13047 2397
rect 13004 2360 13032 2391
rect 13998 2388 14004 2400
rect 14056 2388 14062 2440
rect 15565 2431 15623 2437
rect 15565 2397 15577 2431
rect 15611 2428 15623 2431
rect 16592 2428 16620 2524
rect 17144 2505 17172 2604
rect 18601 2601 18613 2635
rect 18647 2632 18659 2635
rect 20530 2632 20536 2644
rect 18647 2604 20536 2632
rect 18647 2601 18659 2604
rect 18601 2595 18659 2601
rect 20530 2592 20536 2604
rect 20588 2592 20594 2644
rect 21453 2635 21511 2641
rect 21453 2601 21465 2635
rect 21499 2632 21511 2635
rect 23474 2632 23480 2644
rect 21499 2604 23480 2632
rect 21499 2601 21511 2604
rect 21453 2595 21511 2601
rect 23474 2592 23480 2604
rect 23532 2592 23538 2644
rect 18506 2524 18512 2576
rect 18564 2564 18570 2576
rect 21821 2567 21879 2573
rect 21821 2564 21833 2567
rect 18564 2536 21833 2564
rect 18564 2524 18570 2536
rect 17129 2499 17187 2505
rect 17129 2465 17141 2499
rect 17175 2496 17187 2499
rect 17681 2499 17739 2505
rect 17681 2496 17693 2499
rect 17175 2468 17693 2496
rect 17175 2465 17187 2468
rect 17129 2459 17187 2465
rect 17681 2465 17693 2468
rect 17727 2465 17739 2499
rect 17681 2459 17739 2465
rect 17862 2456 17868 2508
rect 17920 2496 17926 2508
rect 18417 2499 18475 2505
rect 18417 2496 18429 2499
rect 17920 2468 18429 2496
rect 17920 2456 17926 2468
rect 18417 2465 18429 2468
rect 18463 2496 18475 2499
rect 18969 2499 19027 2505
rect 18969 2496 18981 2499
rect 18463 2468 18981 2496
rect 18463 2465 18475 2468
rect 18417 2459 18475 2465
rect 18969 2465 18981 2468
rect 19015 2465 19027 2499
rect 18969 2459 19027 2465
rect 19334 2456 19340 2508
rect 19392 2496 19398 2508
rect 21284 2505 21312 2536
rect 21821 2533 21833 2536
rect 21867 2533 21879 2567
rect 21821 2527 21879 2533
rect 19521 2499 19579 2505
rect 19521 2496 19533 2499
rect 19392 2468 19533 2496
rect 19392 2456 19398 2468
rect 19521 2465 19533 2468
rect 19567 2496 19579 2499
rect 20073 2499 20131 2505
rect 20073 2496 20085 2499
rect 19567 2468 20085 2496
rect 19567 2465 19579 2468
rect 19521 2459 19579 2465
rect 20073 2465 20085 2468
rect 20119 2465 20131 2499
rect 20073 2459 20131 2465
rect 21269 2499 21327 2505
rect 21269 2465 21281 2499
rect 21315 2465 21327 2499
rect 22370 2496 22376 2508
rect 22331 2468 22376 2496
rect 21269 2459 21327 2465
rect 22370 2456 22376 2468
rect 22428 2496 22434 2508
rect 22925 2499 22983 2505
rect 22925 2496 22937 2499
rect 22428 2468 22937 2496
rect 22428 2456 22434 2468
rect 22925 2465 22937 2468
rect 22971 2465 22983 2499
rect 22925 2459 22983 2465
rect 24210 2456 24216 2508
rect 24268 2496 24274 2508
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 24268 2468 24593 2496
rect 24268 2456 24274 2468
rect 24581 2465 24593 2468
rect 24627 2496 24639 2499
rect 25133 2499 25191 2505
rect 25133 2496 25145 2499
rect 24627 2468 25145 2496
rect 24627 2465 24639 2468
rect 24581 2459 24639 2465
rect 25133 2465 25145 2468
rect 25179 2465 25191 2499
rect 25133 2459 25191 2465
rect 15611 2400 16620 2428
rect 15611 2397 15623 2400
rect 15565 2391 15623 2397
rect 16114 2360 16120 2372
rect 11900 2332 13032 2360
rect 16027 2332 16120 2360
rect 16114 2320 16120 2332
rect 16172 2360 16178 2372
rect 17126 2360 17132 2372
rect 16172 2332 17132 2360
rect 16172 2320 16178 2332
rect 17126 2320 17132 2332
rect 17184 2320 17190 2372
rect 17313 2363 17371 2369
rect 17313 2329 17325 2363
rect 17359 2360 17371 2363
rect 19150 2360 19156 2372
rect 17359 2332 19156 2360
rect 17359 2329 17371 2332
rect 17313 2323 17371 2329
rect 19150 2320 19156 2332
rect 19208 2320 19214 2372
rect 19705 2363 19763 2369
rect 19705 2329 19717 2363
rect 19751 2360 19763 2363
rect 21174 2360 21180 2372
rect 19751 2332 21180 2360
rect 19751 2329 19763 2332
rect 19705 2323 19763 2329
rect 21174 2320 21180 2332
rect 21232 2320 21238 2372
rect 22557 2363 22615 2369
rect 22557 2329 22569 2363
rect 22603 2360 22615 2363
rect 24118 2360 24124 2372
rect 22603 2332 24124 2360
rect 22603 2329 22615 2332
rect 22557 2323 22615 2329
rect 24118 2320 24124 2332
rect 24176 2320 24182 2372
rect 24765 2363 24823 2369
rect 24765 2329 24777 2363
rect 24811 2360 24823 2363
rect 27522 2360 27528 2372
rect 24811 2332 27528 2360
rect 24811 2329 24823 2332
rect 24765 2323 24823 2329
rect 27522 2320 27528 2332
rect 27580 2320 27586 2372
rect 4939 2295 4997 2301
rect 4939 2261 4951 2295
rect 4985 2292 4997 2295
rect 5166 2292 5172 2304
rect 4985 2264 5172 2292
rect 4985 2261 4997 2264
rect 4939 2255 4997 2261
rect 5166 2252 5172 2264
rect 5224 2252 5230 2304
rect 5353 2295 5411 2301
rect 5353 2261 5365 2295
rect 5399 2292 5411 2295
rect 5442 2292 5448 2304
rect 5399 2264 5448 2292
rect 5399 2261 5411 2264
rect 5353 2255 5411 2261
rect 5442 2252 5448 2264
rect 5500 2252 5506 2304
rect 6086 2252 6092 2304
rect 6144 2292 6150 2304
rect 9582 2292 9588 2304
rect 6144 2264 9588 2292
rect 6144 2252 6150 2264
rect 9582 2252 9588 2264
rect 9640 2252 9646 2304
rect 12710 2252 12716 2304
rect 12768 2292 12774 2304
rect 13633 2295 13691 2301
rect 13633 2292 13645 2295
rect 12768 2264 13645 2292
rect 12768 2252 12774 2264
rect 13633 2261 13645 2264
rect 13679 2261 13691 2295
rect 13633 2255 13691 2261
rect 14734 2252 14740 2304
rect 14792 2292 14798 2304
rect 19518 2292 19524 2304
rect 14792 2264 19524 2292
rect 14792 2252 14798 2264
rect 19518 2252 19524 2264
rect 19576 2252 19582 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 5442 2048 5448 2100
rect 5500 2088 5506 2100
rect 11054 2088 11060 2100
rect 5500 2060 11060 2088
rect 5500 2048 5506 2060
rect 11054 2048 11060 2060
rect 11112 2048 11118 2100
rect 5994 1980 6000 2032
rect 6052 2020 6058 2032
rect 13078 2020 13084 2032
rect 6052 1992 13084 2020
rect 6052 1980 6058 1992
rect 13078 1980 13084 1992
rect 13136 1980 13142 2032
rect 5258 1912 5264 1964
rect 5316 1952 5322 1964
rect 10134 1952 10140 1964
rect 5316 1924 10140 1952
rect 5316 1912 5322 1924
rect 10134 1912 10140 1924
rect 10192 1912 10198 1964
rect 2682 824 2688 876
rect 2740 864 2746 876
rect 4798 864 4804 876
rect 2740 836 4804 864
rect 2740 824 2746 836
rect 4798 824 4804 836
rect 4856 824 4862 876
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 4528 25440 4580 25492
rect 5908 25440 5960 25492
rect 2780 25304 2832 25356
rect 6000 25304 6052 25356
rect 6736 25304 6788 25356
rect 7380 25347 7432 25356
rect 7380 25313 7389 25347
rect 7389 25313 7423 25347
rect 7423 25313 7432 25347
rect 7380 25304 7432 25313
rect 8208 25304 8260 25356
rect 9128 25304 9180 25356
rect 11704 25304 11756 25356
rect 13360 25304 13412 25356
rect 10140 25236 10192 25288
rect 7012 25168 7064 25220
rect 1216 25100 1268 25152
rect 2872 25143 2924 25152
rect 2872 25109 2881 25143
rect 2881 25109 2915 25143
rect 2915 25109 2924 25143
rect 2872 25100 2924 25109
rect 3792 25100 3844 25152
rect 4712 25100 4764 25152
rect 6920 25100 6972 25152
rect 7196 25143 7248 25152
rect 7196 25109 7205 25143
rect 7205 25109 7239 25143
rect 7239 25109 7248 25143
rect 7196 25100 7248 25109
rect 8024 25100 8076 25152
rect 13176 25100 13228 25152
rect 13544 25100 13596 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 2780 24896 2832 24948
rect 4528 24939 4580 24948
rect 4528 24905 4537 24939
rect 4537 24905 4571 24939
rect 4571 24905 4580 24939
rect 4528 24896 4580 24905
rect 6000 24896 6052 24948
rect 11704 24896 11756 24948
rect 8024 24828 8076 24880
rect 10692 24828 10744 24880
rect 13360 24828 13412 24880
rect 4712 24803 4764 24812
rect 4712 24769 4721 24803
rect 4721 24769 4755 24803
rect 4755 24769 4764 24803
rect 4712 24760 4764 24769
rect 4988 24803 5040 24812
rect 4988 24769 4997 24803
rect 4997 24769 5031 24803
rect 5031 24769 5040 24803
rect 4988 24760 5040 24769
rect 7012 24760 7064 24812
rect 7564 24803 7616 24812
rect 7564 24769 7573 24803
rect 7573 24769 7607 24803
rect 7607 24769 7616 24803
rect 7564 24760 7616 24769
rect 4528 24692 4580 24744
rect 8576 24735 8628 24744
rect 8576 24701 8585 24735
rect 8585 24701 8619 24735
rect 8619 24701 8628 24735
rect 8576 24692 8628 24701
rect 8852 24692 8904 24744
rect 11796 24692 11848 24744
rect 2872 24624 2924 24676
rect 1584 24599 1636 24608
rect 1584 24565 1593 24599
rect 1593 24565 1627 24599
rect 1627 24565 1636 24599
rect 1584 24556 1636 24565
rect 2412 24556 2464 24608
rect 4804 24667 4856 24676
rect 4804 24633 4813 24667
rect 4813 24633 4847 24667
rect 4847 24633 4856 24667
rect 4804 24624 4856 24633
rect 4344 24556 4396 24608
rect 5356 24556 5408 24608
rect 7380 24624 7432 24676
rect 7932 24624 7984 24676
rect 11980 24624 12032 24676
rect 8208 24599 8260 24608
rect 8208 24565 8217 24599
rect 8217 24565 8251 24599
rect 8251 24565 8260 24599
rect 8208 24556 8260 24565
rect 10692 24556 10744 24608
rect 12256 24556 12308 24608
rect 13728 24599 13780 24608
rect 13728 24565 13737 24599
rect 13737 24565 13771 24599
rect 13771 24565 13780 24599
rect 13728 24556 13780 24565
rect 14096 24599 14148 24608
rect 14096 24565 14105 24599
rect 14105 24565 14139 24599
rect 14139 24565 14148 24599
rect 14096 24556 14148 24565
rect 14464 24556 14516 24608
rect 17960 24556 18012 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1492 24352 1544 24404
rect 14280 24395 14332 24404
rect 14280 24361 14289 24395
rect 14289 24361 14323 24395
rect 14323 24361 14332 24395
rect 14280 24352 14332 24361
rect 18696 24352 18748 24404
rect 23480 24352 23532 24404
rect 4712 24327 4764 24336
rect 4712 24293 4721 24327
rect 4721 24293 4755 24327
rect 4755 24293 4764 24327
rect 4712 24284 4764 24293
rect 6920 24327 6972 24336
rect 6920 24293 6929 24327
rect 6929 24293 6963 24327
rect 6963 24293 6972 24327
rect 6920 24284 6972 24293
rect 7196 24284 7248 24336
rect 7564 24327 7616 24336
rect 7564 24293 7573 24327
rect 7573 24293 7607 24327
rect 7607 24293 7616 24327
rect 7564 24284 7616 24293
rect 8208 24284 8260 24336
rect 10600 24284 10652 24336
rect 1676 24216 1728 24268
rect 2964 24216 3016 24268
rect 10692 24259 10744 24268
rect 10692 24225 10701 24259
rect 10701 24225 10735 24259
rect 10735 24225 10744 24259
rect 10692 24216 10744 24225
rect 11704 24259 11756 24268
rect 11704 24225 11722 24259
rect 11722 24225 11756 24259
rect 11704 24216 11756 24225
rect 12348 24216 12400 24268
rect 13636 24259 13688 24268
rect 13636 24225 13645 24259
rect 13645 24225 13679 24259
rect 13679 24225 13688 24259
rect 13636 24216 13688 24225
rect 14740 24216 14792 24268
rect 20720 24216 20772 24268
rect 4988 24148 5040 24200
rect 7656 24148 7708 24200
rect 10048 24191 10100 24200
rect 10048 24157 10057 24191
rect 10057 24157 10091 24191
rect 10091 24157 10100 24191
rect 10048 24148 10100 24157
rect 14188 24148 14240 24200
rect 4528 24080 4580 24132
rect 1676 24012 1728 24064
rect 10232 24012 10284 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1676 23851 1728 23860
rect 1676 23817 1685 23851
rect 1685 23817 1719 23851
rect 1719 23817 1728 23851
rect 1676 23808 1728 23817
rect 2412 23808 2464 23860
rect 2504 23851 2556 23860
rect 2504 23817 2513 23851
rect 2513 23817 2547 23851
rect 2547 23817 2556 23851
rect 2504 23808 2556 23817
rect 4712 23808 4764 23860
rect 5448 23808 5500 23860
rect 6920 23808 6972 23860
rect 7196 23808 7248 23860
rect 9680 23851 9732 23860
rect 9680 23817 9689 23851
rect 9689 23817 9723 23851
rect 9723 23817 9732 23851
rect 9680 23808 9732 23817
rect 10048 23851 10100 23860
rect 10048 23817 10057 23851
rect 10057 23817 10091 23851
rect 10091 23817 10100 23851
rect 10048 23808 10100 23817
rect 10692 23808 10744 23860
rect 11704 23851 11756 23860
rect 11704 23817 11713 23851
rect 11713 23817 11747 23851
rect 11747 23817 11756 23851
rect 11704 23808 11756 23817
rect 13636 23851 13688 23860
rect 13636 23817 13645 23851
rect 13645 23817 13679 23851
rect 13679 23817 13688 23851
rect 13636 23808 13688 23817
rect 14464 23808 14516 23860
rect 21088 23808 21140 23860
rect 22744 23808 22796 23860
rect 27528 23808 27580 23860
rect 2964 23783 3016 23792
rect 2964 23749 2973 23783
rect 2973 23749 3007 23783
rect 3007 23749 3016 23783
rect 2964 23740 3016 23749
rect 4436 23740 4488 23792
rect 4528 23740 4580 23792
rect 4988 23740 5040 23792
rect 9772 23740 9824 23792
rect 10140 23740 10192 23792
rect 14280 23783 14332 23792
rect 7656 23715 7708 23724
rect 7656 23681 7665 23715
rect 7665 23681 7699 23715
rect 7699 23681 7708 23715
rect 7656 23672 7708 23681
rect 10692 23715 10744 23724
rect 10692 23681 10701 23715
rect 10701 23681 10735 23715
rect 10735 23681 10744 23715
rect 10692 23672 10744 23681
rect 9680 23604 9732 23656
rect 12348 23604 12400 23656
rect 14280 23749 14289 23783
rect 14289 23749 14323 23783
rect 14323 23749 14332 23783
rect 14280 23740 14332 23749
rect 21640 23740 21692 23792
rect 13912 23672 13964 23724
rect 14188 23647 14240 23656
rect 14188 23613 14197 23647
rect 14197 23613 14231 23647
rect 14231 23613 14240 23647
rect 14188 23604 14240 23613
rect 14464 23647 14516 23656
rect 14464 23613 14473 23647
rect 14473 23613 14507 23647
rect 14507 23613 14516 23647
rect 14464 23604 14516 23613
rect 20720 23672 20772 23724
rect 18420 23604 18472 23656
rect 20260 23647 20312 23656
rect 20260 23613 20269 23647
rect 20269 23613 20303 23647
rect 20303 23613 20312 23647
rect 20260 23604 20312 23613
rect 21364 23647 21416 23656
rect 21364 23613 21373 23647
rect 21373 23613 21407 23647
rect 21407 23613 21416 23647
rect 21364 23604 21416 23613
rect 23480 23604 23532 23656
rect 3976 23468 4028 23520
rect 7932 23536 7984 23588
rect 4436 23468 4488 23520
rect 8024 23468 8076 23520
rect 9404 23468 9456 23520
rect 10048 23468 10100 23520
rect 12716 23468 12768 23520
rect 12992 23468 13044 23520
rect 14556 23536 14608 23588
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 2504 23128 2556 23180
rect 5448 23264 5500 23316
rect 9680 23264 9732 23316
rect 12624 23264 12676 23316
rect 14188 23264 14240 23316
rect 3976 23196 4028 23248
rect 4528 23196 4580 23248
rect 8116 23196 8168 23248
rect 8576 23196 8628 23248
rect 10784 23196 10836 23248
rect 11520 23196 11572 23248
rect 6276 23128 6328 23180
rect 7288 23128 7340 23180
rect 14464 23128 14516 23180
rect 15292 23128 15344 23180
rect 1492 23060 1544 23112
rect 4712 23103 4764 23112
rect 4712 23069 4721 23103
rect 4721 23069 4755 23103
rect 4755 23069 4764 23103
rect 4712 23060 4764 23069
rect 4988 23103 5040 23112
rect 4988 23069 4997 23103
rect 4997 23069 5031 23103
rect 5031 23069 5040 23103
rect 4988 23060 5040 23069
rect 7472 23060 7524 23112
rect 8024 23103 8076 23112
rect 8024 23069 8033 23103
rect 8033 23069 8067 23103
rect 8067 23069 8076 23103
rect 8024 23060 8076 23069
rect 10416 23103 10468 23112
rect 10416 23069 10425 23103
rect 10425 23069 10459 23103
rect 10459 23069 10468 23103
rect 10416 23060 10468 23069
rect 10692 23103 10744 23112
rect 10692 23069 10701 23103
rect 10701 23069 10735 23103
rect 10735 23069 10744 23103
rect 10692 23060 10744 23069
rect 12256 23103 12308 23112
rect 12256 23069 12265 23103
rect 12265 23069 12299 23103
rect 12299 23069 12308 23103
rect 12256 23060 12308 23069
rect 12900 23060 12952 23112
rect 12072 22992 12124 23044
rect 4528 22967 4580 22976
rect 4528 22933 4537 22967
rect 4537 22933 4571 22967
rect 4571 22933 4580 22967
rect 4528 22924 4580 22933
rect 7932 22924 7984 22976
rect 8576 22924 8628 22976
rect 12992 22924 13044 22976
rect 14188 22924 14240 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 2504 22763 2556 22772
rect 2504 22729 2513 22763
rect 2513 22729 2547 22763
rect 2547 22729 2556 22763
rect 2504 22720 2556 22729
rect 4712 22720 4764 22772
rect 6276 22763 6328 22772
rect 6276 22729 6285 22763
rect 6285 22729 6319 22763
rect 6319 22729 6328 22763
rect 6276 22720 6328 22729
rect 7380 22720 7432 22772
rect 8116 22763 8168 22772
rect 8116 22729 8125 22763
rect 8125 22729 8159 22763
rect 8159 22729 8168 22763
rect 8116 22720 8168 22729
rect 10784 22720 10836 22772
rect 11520 22763 11572 22772
rect 11520 22729 11529 22763
rect 11529 22729 11563 22763
rect 11563 22729 11572 22763
rect 11520 22720 11572 22729
rect 12348 22720 12400 22772
rect 4528 22652 4580 22704
rect 14464 22720 14516 22772
rect 23940 22720 23992 22772
rect 12808 22652 12860 22704
rect 14280 22652 14332 22704
rect 14740 22652 14792 22704
rect 1124 22584 1176 22636
rect 1400 22559 1452 22568
rect 1400 22525 1409 22559
rect 1409 22525 1443 22559
rect 1443 22525 1452 22559
rect 1400 22516 1452 22525
rect 3424 22516 3476 22568
rect 10416 22584 10468 22636
rect 12256 22584 12308 22636
rect 13452 22584 13504 22636
rect 4252 22516 4304 22568
rect 4712 22559 4764 22568
rect 4712 22525 4721 22559
rect 4721 22525 4755 22559
rect 4755 22525 4764 22559
rect 4712 22516 4764 22525
rect 6920 22516 6972 22568
rect 9312 22559 9364 22568
rect 9312 22525 9321 22559
rect 9321 22525 9355 22559
rect 9355 22525 9364 22559
rect 9312 22516 9364 22525
rect 12624 22559 12676 22568
rect 12624 22525 12633 22559
rect 12633 22525 12667 22559
rect 12667 22525 12676 22559
rect 12624 22516 12676 22525
rect 12900 22559 12952 22568
rect 12900 22525 12909 22559
rect 12909 22525 12943 22559
rect 12943 22525 12952 22559
rect 12900 22516 12952 22525
rect 14188 22559 14240 22568
rect 14188 22525 14197 22559
rect 14197 22525 14231 22559
rect 14231 22525 14240 22559
rect 14188 22516 14240 22525
rect 14280 22559 14332 22568
rect 14280 22525 14289 22559
rect 14289 22525 14323 22559
rect 14323 22525 14332 22559
rect 14464 22559 14516 22568
rect 14280 22516 14332 22525
rect 14464 22525 14473 22559
rect 14473 22525 14507 22559
rect 14507 22525 14516 22559
rect 14464 22516 14516 22525
rect 112 22380 164 22432
rect 4344 22448 4396 22500
rect 4436 22448 4488 22500
rect 8024 22448 8076 22500
rect 3424 22380 3476 22432
rect 4252 22423 4304 22432
rect 4252 22389 4261 22423
rect 4261 22389 4295 22423
rect 4295 22389 4304 22423
rect 4252 22380 4304 22389
rect 6092 22380 6144 22432
rect 10140 22448 10192 22500
rect 16396 22516 16448 22568
rect 22284 22559 22336 22568
rect 22284 22525 22293 22559
rect 22293 22525 22327 22559
rect 22327 22525 22336 22559
rect 22284 22516 22336 22525
rect 15292 22423 15344 22432
rect 15292 22389 15301 22423
rect 15301 22389 15335 22423
rect 15335 22389 15344 22423
rect 15292 22380 15344 22389
rect 16028 22380 16080 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 1584 22219 1636 22228
rect 1584 22185 1593 22219
rect 1593 22185 1627 22219
rect 1627 22185 1636 22219
rect 1584 22176 1636 22185
rect 5448 22219 5500 22228
rect 5448 22185 5457 22219
rect 5457 22185 5491 22219
rect 5491 22185 5500 22219
rect 5448 22176 5500 22185
rect 7012 22176 7064 22228
rect 7472 22219 7524 22228
rect 7472 22185 7481 22219
rect 7481 22185 7515 22219
rect 7515 22185 7524 22219
rect 7472 22176 7524 22185
rect 8116 22176 8168 22228
rect 9956 22176 10008 22228
rect 10140 22176 10192 22228
rect 12164 22176 12216 22228
rect 14280 22176 14332 22228
rect 22284 22176 22336 22228
rect 4436 22108 4488 22160
rect 8024 22108 8076 22160
rect 12072 22151 12124 22160
rect 12072 22117 12081 22151
rect 12081 22117 12115 22151
rect 12115 22117 12124 22151
rect 12072 22108 12124 22117
rect 15200 22108 15252 22160
rect 2044 22040 2096 22092
rect 2320 22040 2372 22092
rect 6552 22083 6604 22092
rect 6552 22049 6561 22083
rect 6561 22049 6595 22083
rect 6595 22049 6604 22083
rect 6552 22040 6604 22049
rect 11244 22040 11296 22092
rect 12624 22083 12676 22092
rect 12624 22049 12633 22083
rect 12633 22049 12667 22083
rect 12667 22049 12676 22083
rect 12624 22040 12676 22049
rect 12716 22083 12768 22092
rect 12716 22049 12725 22083
rect 12725 22049 12759 22083
rect 12759 22049 12768 22083
rect 12900 22083 12952 22092
rect 12716 22040 12768 22049
rect 12900 22049 12909 22083
rect 12909 22049 12943 22083
rect 12943 22049 12952 22083
rect 12900 22040 12952 22049
rect 13084 22040 13136 22092
rect 14648 22040 14700 22092
rect 2504 22015 2556 22024
rect 2504 21981 2513 22015
rect 2513 21981 2547 22015
rect 2547 21981 2556 22015
rect 2504 21972 2556 21981
rect 4620 21972 4672 22024
rect 7288 21972 7340 22024
rect 11152 21972 11204 22024
rect 13360 22015 13412 22024
rect 13360 21981 13369 22015
rect 13369 21981 13403 22015
rect 13403 21981 13412 22015
rect 13360 21972 13412 21981
rect 13820 21972 13872 22024
rect 14464 21972 14516 22024
rect 15384 22015 15436 22024
rect 15384 21981 15393 22015
rect 15393 21981 15427 22015
rect 15427 21981 15436 22015
rect 15384 21972 15436 21981
rect 15844 22015 15896 22024
rect 15844 21981 15853 22015
rect 15853 21981 15887 22015
rect 15887 21981 15896 22015
rect 15844 21972 15896 21981
rect 9312 21904 9364 21956
rect 11520 21904 11572 21956
rect 2044 21879 2096 21888
rect 2044 21845 2053 21879
rect 2053 21845 2087 21879
rect 2087 21845 2096 21879
rect 2044 21836 2096 21845
rect 3240 21879 3292 21888
rect 3240 21845 3249 21879
rect 3249 21845 3283 21879
rect 3283 21845 3292 21879
rect 3240 21836 3292 21845
rect 4712 21836 4764 21888
rect 6276 21836 6328 21888
rect 6920 21836 6972 21888
rect 9772 21836 9824 21888
rect 11704 21879 11756 21888
rect 11704 21845 11713 21879
rect 11713 21845 11747 21879
rect 11747 21845 11756 21879
rect 11704 21836 11756 21845
rect 13728 21836 13780 21888
rect 16856 21836 16908 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 2504 21675 2556 21684
rect 2504 21641 2513 21675
rect 2513 21641 2547 21675
rect 2547 21641 2556 21675
rect 2504 21632 2556 21641
rect 4436 21632 4488 21684
rect 4804 21632 4856 21684
rect 8576 21632 8628 21684
rect 10784 21632 10836 21684
rect 14464 21632 14516 21684
rect 14648 21675 14700 21684
rect 14648 21641 14657 21675
rect 14657 21641 14691 21675
rect 14691 21641 14700 21675
rect 14648 21632 14700 21641
rect 14832 21632 14884 21684
rect 15292 21632 15344 21684
rect 15384 21632 15436 21684
rect 25872 21632 25924 21684
rect 4528 21428 4580 21480
rect 9956 21564 10008 21616
rect 12624 21564 12676 21616
rect 13360 21564 13412 21616
rect 8484 21496 8536 21548
rect 9496 21428 9548 21480
rect 9772 21428 9824 21480
rect 11796 21471 11848 21480
rect 11796 21437 11805 21471
rect 11805 21437 11839 21471
rect 11839 21437 11848 21471
rect 11796 21428 11848 21437
rect 13728 21539 13780 21548
rect 13728 21505 13737 21539
rect 13737 21505 13771 21539
rect 13771 21505 13780 21539
rect 13728 21496 13780 21505
rect 16580 21539 16632 21548
rect 16580 21505 16589 21539
rect 16589 21505 16623 21539
rect 16623 21505 16632 21539
rect 16580 21496 16632 21505
rect 23940 21471 23992 21480
rect 23940 21437 23949 21471
rect 23949 21437 23983 21471
rect 23983 21437 23992 21471
rect 23940 21428 23992 21437
rect 1584 21403 1636 21412
rect 1584 21369 1593 21403
rect 1593 21369 1627 21403
rect 1627 21369 1636 21403
rect 1584 21360 1636 21369
rect 2964 21360 3016 21412
rect 3240 21403 3292 21412
rect 3240 21369 3249 21403
rect 3249 21369 3283 21403
rect 3283 21369 3292 21403
rect 3240 21360 3292 21369
rect 3332 21403 3384 21412
rect 3332 21369 3341 21403
rect 3341 21369 3375 21403
rect 3375 21369 3384 21403
rect 3332 21360 3384 21369
rect 4252 21360 4304 21412
rect 4620 21360 4672 21412
rect 6644 21360 6696 21412
rect 8024 21360 8076 21412
rect 11244 21360 11296 21412
rect 13820 21403 13872 21412
rect 13820 21369 13829 21403
rect 13829 21369 13863 21403
rect 13863 21369 13872 21403
rect 14372 21403 14424 21412
rect 13820 21360 13872 21369
rect 14372 21369 14381 21403
rect 14381 21369 14415 21403
rect 14415 21369 14424 21403
rect 14372 21360 14424 21369
rect 15384 21403 15436 21412
rect 15384 21369 15393 21403
rect 15393 21369 15427 21403
rect 15427 21369 15436 21403
rect 15384 21360 15436 21369
rect 15660 21360 15712 21412
rect 16856 21360 16908 21412
rect 3516 21292 3568 21344
rect 4436 21292 4488 21344
rect 6552 21335 6604 21344
rect 6552 21301 6561 21335
rect 6561 21301 6595 21335
rect 6595 21301 6604 21335
rect 6552 21292 6604 21301
rect 7288 21292 7340 21344
rect 7472 21335 7524 21344
rect 7472 21301 7481 21335
rect 7481 21301 7515 21335
rect 7515 21301 7524 21335
rect 7472 21292 7524 21301
rect 7748 21335 7800 21344
rect 7748 21301 7757 21335
rect 7757 21301 7791 21335
rect 7791 21301 7800 21335
rect 7748 21292 7800 21301
rect 9128 21292 9180 21344
rect 9956 21335 10008 21344
rect 9956 21301 9965 21335
rect 9965 21301 9999 21335
rect 9999 21301 10008 21335
rect 9956 21292 10008 21301
rect 11152 21335 11204 21344
rect 11152 21301 11161 21335
rect 11161 21301 11195 21335
rect 11195 21301 11204 21335
rect 11152 21292 11204 21301
rect 11520 21335 11572 21344
rect 11520 21301 11529 21335
rect 11529 21301 11563 21335
rect 11563 21301 11572 21335
rect 11520 21292 11572 21301
rect 14648 21292 14700 21344
rect 16948 21335 17000 21344
rect 16948 21301 16957 21335
rect 16957 21301 16991 21335
rect 16991 21301 17000 21335
rect 16948 21292 17000 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 3792 21131 3844 21140
rect 3792 21097 3801 21131
rect 3801 21097 3835 21131
rect 3835 21097 3844 21131
rect 3792 21088 3844 21097
rect 4344 21088 4396 21140
rect 6920 21131 6972 21140
rect 2412 21063 2464 21072
rect 2412 21029 2421 21063
rect 2421 21029 2455 21063
rect 2455 21029 2464 21063
rect 2412 21020 2464 21029
rect 2964 21063 3016 21072
rect 2964 21029 2973 21063
rect 2973 21029 3007 21063
rect 3007 21029 3016 21063
rect 2964 21020 3016 21029
rect 4160 21020 4212 21072
rect 6920 21097 6929 21131
rect 6929 21097 6963 21131
rect 6963 21097 6972 21131
rect 6920 21088 6972 21097
rect 9772 21131 9824 21140
rect 9772 21097 9781 21131
rect 9781 21097 9815 21131
rect 9815 21097 9824 21131
rect 9772 21088 9824 21097
rect 12900 21088 12952 21140
rect 16580 21088 16632 21140
rect 7012 20952 7064 21004
rect 7472 20952 7524 21004
rect 7656 20995 7708 21004
rect 7656 20961 7665 20995
rect 7665 20961 7699 20995
rect 7699 20961 7708 20995
rect 7656 20952 7708 20961
rect 9128 21020 9180 21072
rect 9220 21020 9272 21072
rect 12716 21020 12768 21072
rect 14188 21020 14240 21072
rect 15936 21063 15988 21072
rect 15936 21029 15945 21063
rect 15945 21029 15979 21063
rect 15979 21029 15988 21063
rect 15936 21020 15988 21029
rect 9036 20952 9088 21004
rect 10324 20995 10376 21004
rect 3792 20884 3844 20936
rect 4252 20884 4304 20936
rect 8484 20884 8536 20936
rect 10324 20961 10333 20995
rect 10333 20961 10367 20995
rect 10367 20961 10376 20995
rect 10324 20952 10376 20961
rect 10508 20995 10560 21004
rect 10508 20961 10517 20995
rect 10517 20961 10551 20995
rect 10551 20961 10560 20995
rect 10508 20952 10560 20961
rect 10784 20952 10836 21004
rect 11520 20952 11572 21004
rect 12072 20995 12124 21004
rect 12072 20961 12081 20995
rect 12081 20961 12115 20995
rect 12115 20961 12124 20995
rect 12072 20952 12124 20961
rect 17500 20952 17552 21004
rect 11612 20884 11664 20936
rect 13544 20884 13596 20936
rect 14372 20927 14424 20936
rect 14372 20893 14381 20927
rect 14381 20893 14415 20927
rect 14415 20893 14424 20927
rect 15844 20927 15896 20936
rect 14372 20884 14424 20893
rect 15844 20893 15853 20927
rect 15853 20893 15887 20927
rect 15887 20893 15896 20927
rect 15844 20884 15896 20893
rect 16488 20884 16540 20936
rect 11704 20816 11756 20868
rect 1584 20791 1636 20800
rect 1584 20757 1593 20791
rect 1593 20757 1627 20791
rect 1627 20757 1636 20791
rect 1584 20748 1636 20757
rect 1676 20748 1728 20800
rect 2780 20748 2832 20800
rect 6828 20748 6880 20800
rect 9036 20791 9088 20800
rect 9036 20757 9045 20791
rect 9045 20757 9079 20791
rect 9079 20757 9088 20791
rect 9036 20748 9088 20757
rect 16856 20816 16908 20868
rect 14004 20748 14056 20800
rect 14372 20748 14424 20800
rect 15384 20748 15436 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1400 20544 1452 20596
rect 10416 20544 10468 20596
rect 2228 20476 2280 20528
rect 2412 20476 2464 20528
rect 7748 20476 7800 20528
rect 10508 20476 10560 20528
rect 13544 20544 13596 20596
rect 15292 20544 15344 20596
rect 15936 20544 15988 20596
rect 16488 20587 16540 20596
rect 16488 20553 16497 20587
rect 16497 20553 16531 20587
rect 16531 20553 16540 20587
rect 16488 20544 16540 20553
rect 1676 20340 1728 20392
rect 2596 20340 2648 20392
rect 4344 20340 4396 20392
rect 4896 20383 4948 20392
rect 4896 20349 4905 20383
rect 4905 20349 4939 20383
rect 4939 20349 4948 20383
rect 4896 20340 4948 20349
rect 5448 20383 5500 20392
rect 5448 20349 5457 20383
rect 5457 20349 5491 20383
rect 5491 20349 5500 20383
rect 5448 20340 5500 20349
rect 2872 20272 2924 20324
rect 3516 20272 3568 20324
rect 4528 20247 4580 20256
rect 4528 20213 4537 20247
rect 4537 20213 4571 20247
rect 4571 20213 4580 20247
rect 4528 20204 4580 20213
rect 5264 20204 5316 20256
rect 7012 20340 7064 20392
rect 7472 20340 7524 20392
rect 8208 20383 8260 20392
rect 8208 20349 8217 20383
rect 8217 20349 8251 20383
rect 8251 20349 8260 20383
rect 8208 20340 8260 20349
rect 9036 20408 9088 20460
rect 7656 20272 7708 20324
rect 6736 20204 6788 20256
rect 7288 20204 7340 20256
rect 10416 20383 10468 20392
rect 10416 20349 10425 20383
rect 10425 20349 10459 20383
rect 10459 20349 10468 20383
rect 10416 20340 10468 20349
rect 11152 20451 11204 20460
rect 11152 20417 11161 20451
rect 11161 20417 11195 20451
rect 11195 20417 11204 20451
rect 11152 20408 11204 20417
rect 15660 20408 15712 20460
rect 10968 20340 11020 20392
rect 11336 20340 11388 20392
rect 15384 20340 15436 20392
rect 15936 20340 15988 20392
rect 21364 20408 21416 20460
rect 18512 20340 18564 20392
rect 13452 20315 13504 20324
rect 13452 20281 13461 20315
rect 13461 20281 13495 20315
rect 13495 20281 13504 20315
rect 13452 20272 13504 20281
rect 9864 20204 9916 20256
rect 12072 20247 12124 20256
rect 12072 20213 12081 20247
rect 12081 20213 12115 20247
rect 12115 20213 12124 20247
rect 12072 20204 12124 20213
rect 14832 20272 14884 20324
rect 23940 20340 23992 20392
rect 14372 20247 14424 20256
rect 14372 20213 14381 20247
rect 14381 20213 14415 20247
rect 14415 20213 14424 20247
rect 14372 20204 14424 20213
rect 15286 20247 15338 20256
rect 15286 20213 15295 20247
rect 15295 20213 15329 20247
rect 15329 20213 15338 20247
rect 15286 20204 15338 20213
rect 16580 20204 16632 20256
rect 17500 20247 17552 20256
rect 17500 20213 17509 20247
rect 17509 20213 17543 20247
rect 17543 20213 17552 20247
rect 17500 20204 17552 20213
rect 18512 20247 18564 20256
rect 18512 20213 18521 20247
rect 18521 20213 18555 20247
rect 18555 20213 18564 20247
rect 18512 20204 18564 20213
rect 18604 20204 18656 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 3424 20000 3476 20052
rect 6276 20043 6328 20052
rect 1584 19975 1636 19984
rect 1584 19941 1593 19975
rect 1593 19941 1627 19975
rect 1627 19941 1636 19975
rect 1584 19932 1636 19941
rect 3332 19932 3384 19984
rect 2228 19907 2280 19916
rect 2228 19873 2237 19907
rect 2237 19873 2271 19907
rect 2271 19873 2280 19907
rect 2228 19864 2280 19873
rect 4160 19907 4212 19916
rect 4160 19873 4169 19907
rect 4169 19873 4203 19907
rect 4203 19873 4212 19907
rect 6276 20009 6285 20043
rect 6285 20009 6319 20043
rect 6319 20009 6328 20043
rect 6276 20000 6328 20009
rect 7012 20000 7064 20052
rect 9036 20000 9088 20052
rect 11796 20043 11848 20052
rect 11796 20009 11805 20043
rect 11805 20009 11839 20043
rect 11839 20009 11848 20043
rect 11796 20000 11848 20009
rect 12440 20000 12492 20052
rect 13452 20000 13504 20052
rect 16580 20000 16632 20052
rect 6736 19932 6788 19984
rect 4160 19864 4212 19873
rect 6460 19907 6512 19916
rect 6460 19873 6469 19907
rect 6469 19873 6503 19907
rect 6503 19873 6512 19907
rect 6460 19864 6512 19873
rect 6828 19907 6880 19916
rect 6828 19873 6837 19907
rect 6837 19873 6871 19907
rect 6871 19873 6880 19907
rect 6828 19864 6880 19873
rect 9128 19932 9180 19984
rect 9496 19932 9548 19984
rect 8576 19907 8628 19916
rect 8576 19873 8585 19907
rect 8585 19873 8619 19907
rect 8619 19873 8628 19907
rect 8576 19864 8628 19873
rect 9864 19864 9916 19916
rect 10140 19864 10192 19916
rect 12072 19932 12124 19984
rect 16396 19975 16448 19984
rect 11796 19864 11848 19916
rect 13268 19864 13320 19916
rect 16396 19941 16405 19975
rect 16405 19941 16439 19975
rect 16439 19941 16448 19975
rect 16396 19932 16448 19941
rect 14004 19864 14056 19916
rect 16120 19864 16172 19916
rect 17776 19907 17828 19916
rect 17776 19873 17785 19907
rect 17785 19873 17819 19907
rect 17819 19873 17828 19907
rect 17776 19864 17828 19873
rect 18788 19907 18840 19916
rect 18788 19873 18797 19907
rect 18797 19873 18831 19907
rect 18831 19873 18840 19907
rect 18788 19864 18840 19873
rect 2688 19703 2740 19712
rect 2688 19669 2697 19703
rect 2697 19669 2731 19703
rect 2731 19669 2740 19703
rect 2688 19660 2740 19669
rect 2964 19703 3016 19712
rect 2964 19669 2973 19703
rect 2973 19669 3007 19703
rect 3007 19669 3016 19703
rect 2964 19660 3016 19669
rect 3608 19660 3660 19712
rect 5264 19660 5316 19712
rect 5540 19660 5592 19712
rect 7288 19796 7340 19848
rect 9220 19796 9272 19848
rect 10692 19839 10744 19848
rect 10692 19805 10701 19839
rect 10701 19805 10735 19839
rect 10735 19805 10744 19839
rect 10692 19796 10744 19805
rect 13728 19839 13780 19848
rect 13728 19805 13737 19839
rect 13737 19805 13771 19839
rect 13771 19805 13780 19839
rect 13728 19796 13780 19805
rect 15660 19796 15712 19848
rect 16028 19796 16080 19848
rect 9956 19728 10008 19780
rect 12532 19728 12584 19780
rect 18512 19796 18564 19848
rect 16856 19771 16908 19780
rect 7656 19660 7708 19712
rect 8208 19660 8260 19712
rect 8668 19660 8720 19712
rect 9128 19660 9180 19712
rect 9772 19660 9824 19712
rect 10968 19703 11020 19712
rect 10968 19669 10977 19703
rect 10977 19669 11011 19703
rect 11011 19669 11020 19703
rect 10968 19660 11020 19669
rect 11428 19703 11480 19712
rect 11428 19669 11437 19703
rect 11437 19669 11471 19703
rect 11471 19669 11480 19703
rect 16856 19737 16865 19771
rect 16865 19737 16899 19771
rect 16899 19737 16908 19771
rect 16856 19728 16908 19737
rect 11428 19660 11480 19669
rect 15384 19660 15436 19712
rect 15568 19703 15620 19712
rect 15568 19669 15577 19703
rect 15577 19669 15611 19703
rect 15611 19669 15620 19703
rect 15568 19660 15620 19669
rect 15844 19660 15896 19712
rect 18972 19703 19024 19712
rect 18972 19669 18981 19703
rect 18981 19669 19015 19703
rect 19015 19669 19024 19703
rect 18972 19660 19024 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 2228 19456 2280 19508
rect 2872 19499 2924 19508
rect 2872 19465 2881 19499
rect 2881 19465 2915 19499
rect 2915 19465 2924 19499
rect 2872 19456 2924 19465
rect 4160 19456 4212 19508
rect 6828 19456 6880 19508
rect 7472 19456 7524 19508
rect 9864 19456 9916 19508
rect 10784 19456 10836 19508
rect 11796 19499 11848 19508
rect 11796 19465 11805 19499
rect 11805 19465 11839 19499
rect 11839 19465 11848 19499
rect 11796 19456 11848 19465
rect 13268 19456 13320 19508
rect 15476 19456 15528 19508
rect 16396 19499 16448 19508
rect 16396 19465 16405 19499
rect 16405 19465 16439 19499
rect 16439 19465 16448 19499
rect 16396 19456 16448 19465
rect 10876 19431 10928 19440
rect 3148 19320 3200 19372
rect 4528 19320 4580 19372
rect 6460 19320 6512 19372
rect 2228 19252 2280 19304
rect 2964 19252 3016 19304
rect 2872 19184 2924 19236
rect 6736 19252 6788 19304
rect 7564 19320 7616 19372
rect 7380 19295 7432 19304
rect 7380 19261 7389 19295
rect 7389 19261 7423 19295
rect 7423 19261 7432 19295
rect 7380 19252 7432 19261
rect 7288 19184 7340 19236
rect 7748 19252 7800 19304
rect 10876 19397 10885 19431
rect 10885 19397 10919 19431
rect 10919 19397 10928 19431
rect 10876 19388 10928 19397
rect 11428 19388 11480 19440
rect 16028 19388 16080 19440
rect 9956 19363 10008 19372
rect 9956 19329 9965 19363
rect 9965 19329 9999 19363
rect 9999 19329 10008 19363
rect 9956 19320 10008 19329
rect 1676 19159 1728 19168
rect 1676 19125 1685 19159
rect 1685 19125 1719 19159
rect 1719 19125 1728 19159
rect 1676 19116 1728 19125
rect 4620 19159 4672 19168
rect 4620 19125 4629 19159
rect 4629 19125 4663 19159
rect 4663 19125 4672 19159
rect 4620 19116 4672 19125
rect 4988 19159 5040 19168
rect 4988 19125 4997 19159
rect 4997 19125 5031 19159
rect 5031 19125 5040 19159
rect 4988 19116 5040 19125
rect 5540 19159 5592 19168
rect 5540 19125 5549 19159
rect 5549 19125 5583 19159
rect 5583 19125 5592 19159
rect 5540 19116 5592 19125
rect 6644 19116 6696 19168
rect 7196 19116 7248 19168
rect 10968 19252 11020 19304
rect 11060 19295 11112 19304
rect 11060 19261 11069 19295
rect 11069 19261 11103 19295
rect 11103 19261 11112 19295
rect 11060 19252 11112 19261
rect 9864 19184 9916 19236
rect 12072 19252 12124 19304
rect 12440 19295 12492 19304
rect 12440 19261 12449 19295
rect 12449 19261 12483 19295
rect 12483 19261 12492 19295
rect 12440 19252 12492 19261
rect 12532 19295 12584 19304
rect 12532 19261 12541 19295
rect 12541 19261 12575 19295
rect 12575 19261 12584 19295
rect 13728 19320 13780 19372
rect 17776 19456 17828 19508
rect 17776 19320 17828 19372
rect 12532 19252 12584 19261
rect 15568 19252 15620 19304
rect 7840 19116 7892 19168
rect 8576 19159 8628 19168
rect 8576 19125 8585 19159
rect 8585 19125 8619 19159
rect 8619 19125 8628 19159
rect 8576 19116 8628 19125
rect 10140 19116 10192 19168
rect 12256 19184 12308 19236
rect 14464 19184 14516 19236
rect 14004 19116 14056 19168
rect 14188 19159 14240 19168
rect 14188 19125 14197 19159
rect 14197 19125 14231 19159
rect 14231 19125 14240 19159
rect 14188 19116 14240 19125
rect 15292 19159 15344 19168
rect 15292 19125 15301 19159
rect 15301 19125 15335 19159
rect 15335 19125 15344 19159
rect 15292 19116 15344 19125
rect 15660 19184 15712 19236
rect 16764 19116 16816 19168
rect 17776 19159 17828 19168
rect 17776 19125 17785 19159
rect 17785 19125 17819 19159
rect 17819 19125 17828 19159
rect 17776 19116 17828 19125
rect 18144 19252 18196 19304
rect 18788 19252 18840 19304
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1492 18912 1544 18964
rect 3148 18955 3200 18964
rect 3148 18921 3157 18955
rect 3157 18921 3191 18955
rect 3191 18921 3200 18955
rect 3148 18912 3200 18921
rect 4620 18912 4672 18964
rect 5172 18955 5224 18964
rect 5172 18921 5181 18955
rect 5181 18921 5215 18955
rect 5215 18921 5224 18955
rect 5172 18912 5224 18921
rect 7104 18912 7156 18964
rect 7748 18912 7800 18964
rect 2228 18887 2280 18896
rect 2228 18853 2237 18887
rect 2237 18853 2271 18887
rect 2271 18853 2280 18887
rect 2228 18844 2280 18853
rect 2780 18887 2832 18896
rect 2780 18853 2789 18887
rect 2789 18853 2823 18887
rect 2823 18853 2832 18887
rect 2780 18844 2832 18853
rect 4344 18844 4396 18896
rect 7472 18844 7524 18896
rect 10876 18912 10928 18964
rect 15384 18912 15436 18964
rect 18144 18955 18196 18964
rect 18144 18921 18153 18955
rect 18153 18921 18187 18955
rect 18187 18921 18196 18955
rect 18144 18912 18196 18921
rect 10416 18844 10468 18896
rect 14648 18844 14700 18896
rect 16028 18887 16080 18896
rect 16028 18853 16037 18887
rect 16037 18853 16071 18887
rect 16071 18853 16080 18887
rect 16028 18844 16080 18853
rect 3608 18708 3660 18760
rect 6000 18819 6052 18828
rect 4896 18708 4948 18760
rect 6000 18785 6009 18819
rect 6009 18785 6043 18819
rect 6043 18785 6052 18819
rect 6000 18776 6052 18785
rect 6368 18819 6420 18828
rect 6368 18785 6377 18819
rect 6377 18785 6411 18819
rect 6411 18785 6420 18819
rect 6368 18776 6420 18785
rect 8208 18819 8260 18828
rect 8208 18785 8217 18819
rect 8217 18785 8251 18819
rect 8251 18785 8260 18819
rect 8208 18776 8260 18785
rect 9772 18819 9824 18828
rect 9772 18785 9781 18819
rect 9781 18785 9815 18819
rect 9815 18785 9824 18819
rect 9772 18776 9824 18785
rect 9956 18776 10008 18828
rect 10140 18776 10192 18828
rect 11244 18776 11296 18828
rect 11336 18819 11388 18828
rect 11336 18785 11345 18819
rect 11345 18785 11379 18819
rect 11379 18785 11388 18819
rect 11612 18819 11664 18828
rect 11336 18776 11388 18785
rect 11612 18785 11621 18819
rect 11621 18785 11655 18819
rect 11655 18785 11664 18819
rect 11612 18776 11664 18785
rect 13268 18819 13320 18828
rect 13268 18785 13277 18819
rect 13277 18785 13311 18819
rect 13311 18785 13320 18819
rect 13268 18776 13320 18785
rect 9312 18708 9364 18760
rect 9496 18751 9548 18760
rect 9496 18717 9505 18751
rect 9505 18717 9539 18751
rect 9539 18717 9548 18751
rect 11796 18751 11848 18760
rect 9496 18708 9548 18717
rect 9036 18640 9088 18692
rect 2964 18572 3016 18624
rect 3884 18615 3936 18624
rect 3884 18581 3893 18615
rect 3893 18581 3927 18615
rect 3927 18581 3936 18615
rect 3884 18572 3936 18581
rect 7564 18572 7616 18624
rect 8024 18572 8076 18624
rect 9128 18615 9180 18624
rect 9128 18581 9137 18615
rect 9137 18581 9171 18615
rect 9171 18581 9180 18615
rect 9128 18572 9180 18581
rect 11796 18717 11805 18751
rect 11805 18717 11839 18751
rect 11839 18717 11848 18751
rect 11796 18708 11848 18717
rect 13728 18776 13780 18828
rect 17224 18776 17276 18828
rect 17408 18819 17460 18828
rect 17408 18785 17417 18819
rect 17417 18785 17451 18819
rect 17451 18785 17460 18819
rect 17408 18776 17460 18785
rect 18328 18776 18380 18828
rect 13912 18751 13964 18760
rect 13912 18717 13921 18751
rect 13921 18717 13955 18751
rect 13955 18717 13964 18751
rect 13912 18708 13964 18717
rect 15384 18751 15436 18760
rect 15384 18717 15393 18751
rect 15393 18717 15427 18751
rect 15427 18717 15436 18751
rect 15384 18708 15436 18717
rect 9864 18640 9916 18692
rect 11336 18640 11388 18692
rect 12532 18640 12584 18692
rect 14464 18640 14516 18692
rect 9956 18572 10008 18624
rect 11060 18572 11112 18624
rect 16304 18572 16356 18624
rect 16488 18615 16540 18624
rect 16488 18581 16497 18615
rect 16497 18581 16531 18615
rect 16531 18581 16540 18615
rect 16488 18572 16540 18581
rect 18604 18615 18656 18624
rect 18604 18581 18613 18615
rect 18613 18581 18647 18615
rect 18647 18581 18656 18615
rect 18604 18572 18656 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 2228 18368 2280 18420
rect 2872 18368 2924 18420
rect 1492 18275 1544 18284
rect 1492 18241 1501 18275
rect 1501 18241 1535 18275
rect 1535 18241 1544 18275
rect 1492 18232 1544 18241
rect 2780 18232 2832 18284
rect 4896 18368 4948 18420
rect 6000 18368 6052 18420
rect 8208 18411 8260 18420
rect 8208 18377 8217 18411
rect 8217 18377 8251 18411
rect 8251 18377 8260 18411
rect 8208 18368 8260 18377
rect 8852 18368 8904 18420
rect 10140 18368 10192 18420
rect 11336 18411 11388 18420
rect 11336 18377 11345 18411
rect 11345 18377 11379 18411
rect 11379 18377 11388 18411
rect 11336 18368 11388 18377
rect 11428 18368 11480 18420
rect 18328 18368 18380 18420
rect 6276 18343 6328 18352
rect 3332 18207 3384 18216
rect 3332 18173 3341 18207
rect 3341 18173 3375 18207
rect 3375 18173 3384 18207
rect 3332 18164 3384 18173
rect 1676 18096 1728 18148
rect 4988 18232 5040 18284
rect 5448 18164 5500 18216
rect 6276 18309 6285 18343
rect 6285 18309 6319 18343
rect 6319 18309 6328 18343
rect 6276 18300 6328 18309
rect 8484 18343 8536 18352
rect 8484 18309 8493 18343
rect 8493 18309 8527 18343
rect 8527 18309 8536 18343
rect 8484 18300 8536 18309
rect 10324 18300 10376 18352
rect 14648 18300 14700 18352
rect 15568 18300 15620 18352
rect 6460 18232 6512 18284
rect 7840 18275 7892 18284
rect 7104 18207 7156 18216
rect 7104 18173 7113 18207
rect 7113 18173 7147 18207
rect 7147 18173 7156 18207
rect 7104 18164 7156 18173
rect 7196 18207 7248 18216
rect 7196 18173 7205 18207
rect 7205 18173 7239 18207
rect 7239 18173 7248 18207
rect 7840 18241 7849 18275
rect 7849 18241 7883 18275
rect 7883 18241 7892 18275
rect 7840 18232 7892 18241
rect 9128 18232 9180 18284
rect 10048 18232 10100 18284
rect 7196 18164 7248 18173
rect 4344 18028 4396 18080
rect 8852 18139 8904 18148
rect 8852 18105 8861 18139
rect 8861 18105 8895 18139
rect 8895 18105 8904 18139
rect 8852 18096 8904 18105
rect 9036 18096 9088 18148
rect 13912 18275 13964 18284
rect 13912 18241 13921 18275
rect 13921 18241 13955 18275
rect 13955 18241 13964 18275
rect 13912 18232 13964 18241
rect 16488 18275 16540 18284
rect 16488 18241 16497 18275
rect 16497 18241 16531 18275
rect 16531 18241 16540 18275
rect 16488 18232 16540 18241
rect 16856 18275 16908 18284
rect 16856 18241 16865 18275
rect 16865 18241 16899 18275
rect 16899 18241 16908 18275
rect 16856 18232 16908 18241
rect 12624 18207 12676 18216
rect 12624 18173 12633 18207
rect 12633 18173 12667 18207
rect 12667 18173 12676 18207
rect 12624 18164 12676 18173
rect 10324 18139 10376 18148
rect 10324 18105 10333 18139
rect 10333 18105 10367 18139
rect 10367 18105 10376 18139
rect 10324 18096 10376 18105
rect 10416 18139 10468 18148
rect 10416 18105 10425 18139
rect 10425 18105 10459 18139
rect 10459 18105 10468 18139
rect 10416 18096 10468 18105
rect 11612 18096 11664 18148
rect 11520 18028 11572 18080
rect 12900 18096 12952 18148
rect 16120 18164 16172 18216
rect 14004 18028 14056 18080
rect 15384 18028 15436 18080
rect 16212 18028 16264 18080
rect 16672 18028 16724 18080
rect 17316 18028 17368 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1676 17867 1728 17876
rect 1676 17833 1685 17867
rect 1685 17833 1719 17867
rect 1719 17833 1728 17867
rect 1676 17824 1728 17833
rect 2228 17824 2280 17876
rect 3332 17824 3384 17876
rect 4252 17867 4304 17876
rect 2872 17756 2924 17808
rect 4252 17833 4261 17867
rect 4261 17833 4295 17867
rect 4295 17833 4304 17867
rect 4252 17824 4304 17833
rect 7196 17867 7248 17876
rect 7196 17833 7205 17867
rect 7205 17833 7239 17867
rect 7239 17833 7248 17867
rect 7196 17824 7248 17833
rect 8852 17824 8904 17876
rect 9496 17867 9548 17876
rect 9496 17833 9505 17867
rect 9505 17833 9539 17867
rect 9539 17833 9548 17867
rect 9496 17824 9548 17833
rect 9772 17824 9824 17876
rect 11612 17824 11664 17876
rect 5172 17756 5224 17808
rect 5540 17756 5592 17808
rect 2780 17620 2832 17672
rect 2136 17484 2188 17536
rect 3332 17484 3384 17536
rect 5632 17731 5684 17740
rect 4712 17620 4764 17672
rect 5632 17697 5641 17731
rect 5641 17697 5675 17731
rect 5675 17697 5684 17731
rect 5632 17688 5684 17697
rect 7472 17756 7524 17808
rect 6552 17731 6604 17740
rect 6552 17697 6561 17731
rect 6561 17697 6595 17731
rect 6595 17697 6604 17731
rect 6552 17688 6604 17697
rect 8208 17688 8260 17740
rect 9312 17688 9364 17740
rect 10140 17688 10192 17740
rect 11520 17688 11572 17740
rect 11704 17688 11756 17740
rect 14188 17824 14240 17876
rect 16672 17867 16724 17876
rect 16672 17833 16681 17867
rect 16681 17833 16715 17867
rect 16715 17833 16724 17867
rect 16672 17824 16724 17833
rect 17408 17824 17460 17876
rect 12716 17756 12768 17808
rect 15476 17756 15528 17808
rect 16212 17756 16264 17808
rect 13268 17731 13320 17740
rect 13268 17697 13277 17731
rect 13277 17697 13311 17731
rect 13311 17697 13320 17731
rect 13268 17688 13320 17697
rect 13636 17731 13688 17740
rect 13636 17697 13645 17731
rect 13645 17697 13679 17731
rect 13679 17697 13688 17731
rect 13636 17688 13688 17697
rect 13728 17688 13780 17740
rect 5264 17552 5316 17604
rect 6552 17552 6604 17604
rect 8300 17620 8352 17672
rect 12808 17663 12860 17672
rect 12808 17629 12817 17663
rect 12817 17629 12851 17663
rect 12851 17629 12860 17663
rect 12808 17620 12860 17629
rect 17408 17688 17460 17740
rect 17040 17620 17092 17672
rect 18328 17620 18380 17672
rect 15292 17552 15344 17604
rect 4896 17484 4948 17536
rect 5540 17484 5592 17536
rect 6828 17484 6880 17536
rect 10784 17484 10836 17536
rect 13268 17484 13320 17536
rect 15844 17484 15896 17536
rect 18696 17527 18748 17536
rect 18696 17493 18705 17527
rect 18705 17493 18739 17527
rect 18739 17493 18748 17527
rect 18696 17484 18748 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2688 17280 2740 17332
rect 2872 17280 2924 17332
rect 10140 17323 10192 17332
rect 10140 17289 10149 17323
rect 10149 17289 10183 17323
rect 10183 17289 10192 17323
rect 10140 17280 10192 17289
rect 13084 17280 13136 17332
rect 13636 17280 13688 17332
rect 13820 17280 13872 17332
rect 17040 17323 17092 17332
rect 4620 17212 4672 17264
rect 5540 17212 5592 17264
rect 14832 17255 14884 17264
rect 14832 17221 14841 17255
rect 14841 17221 14875 17255
rect 14875 17221 14884 17255
rect 14832 17212 14884 17221
rect 15292 17212 15344 17264
rect 16488 17212 16540 17264
rect 17040 17289 17049 17323
rect 17049 17289 17083 17323
rect 17083 17289 17092 17323
rect 17040 17280 17092 17289
rect 18328 17280 18380 17332
rect 2136 17076 2188 17128
rect 4712 17119 4764 17128
rect 4712 17085 4721 17119
rect 4721 17085 4755 17119
rect 4755 17085 4764 17119
rect 4712 17076 4764 17085
rect 4896 17119 4948 17128
rect 4896 17085 4905 17119
rect 4905 17085 4939 17119
rect 4939 17085 4948 17119
rect 4896 17076 4948 17085
rect 5264 17119 5316 17128
rect 5264 17085 5273 17119
rect 5273 17085 5307 17119
rect 5307 17085 5316 17119
rect 5264 17076 5316 17085
rect 5540 17076 5592 17128
rect 6828 17119 6880 17128
rect 2964 17051 3016 17060
rect 2964 17017 2973 17051
rect 2973 17017 3007 17051
rect 3007 17017 3016 17051
rect 2964 17008 3016 17017
rect 3608 17051 3660 17060
rect 112 16940 164 16992
rect 3608 17017 3617 17051
rect 3617 17017 3651 17051
rect 3651 17017 3660 17051
rect 3608 17008 3660 17017
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 7288 17119 7340 17128
rect 7288 17085 7297 17119
rect 7297 17085 7331 17119
rect 7331 17085 7340 17119
rect 7288 17076 7340 17085
rect 7656 17076 7708 17128
rect 8208 17119 8260 17128
rect 6368 17008 6420 17060
rect 8208 17085 8217 17119
rect 8217 17085 8251 17119
rect 8251 17085 8260 17119
rect 8208 17076 8260 17085
rect 8300 17051 8352 17060
rect 8300 17017 8309 17051
rect 8309 17017 8343 17051
rect 8343 17017 8352 17051
rect 8300 17008 8352 17017
rect 9220 17051 9272 17060
rect 9220 17017 9229 17051
rect 9229 17017 9263 17051
rect 9263 17017 9272 17051
rect 9220 17008 9272 17017
rect 3516 16940 3568 16992
rect 4528 16983 4580 16992
rect 4528 16949 4537 16983
rect 4537 16949 4571 16983
rect 4571 16949 4580 16983
rect 4528 16940 4580 16949
rect 7472 16940 7524 16992
rect 9404 17008 9456 17060
rect 10048 17008 10100 17060
rect 10784 17119 10836 17128
rect 10784 17085 10793 17119
rect 10793 17085 10827 17119
rect 10827 17085 10836 17119
rect 11888 17144 11940 17196
rect 10784 17076 10836 17085
rect 12532 17076 12584 17128
rect 13728 17144 13780 17196
rect 14004 17144 14056 17196
rect 12900 17076 12952 17128
rect 13912 17119 13964 17128
rect 13912 17085 13921 17119
rect 13921 17085 13955 17119
rect 13955 17085 13964 17119
rect 13912 17076 13964 17085
rect 11060 17008 11112 17060
rect 12440 17051 12492 17060
rect 12440 17017 12449 17051
rect 12449 17017 12483 17051
rect 12483 17017 12492 17051
rect 12440 17008 12492 17017
rect 14004 17008 14056 17060
rect 16856 17144 16908 17196
rect 18512 17212 18564 17264
rect 11152 16983 11204 16992
rect 11152 16949 11161 16983
rect 11161 16949 11195 16983
rect 11195 16949 11204 16983
rect 11152 16940 11204 16949
rect 11704 16940 11756 16992
rect 15568 17008 15620 17060
rect 14464 16940 14516 16992
rect 15476 16983 15528 16992
rect 15476 16949 15485 16983
rect 15485 16949 15519 16983
rect 15519 16949 15528 16983
rect 15476 16940 15528 16949
rect 17408 16940 17460 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 2780 16779 2832 16788
rect 2780 16745 2789 16779
rect 2789 16745 2823 16779
rect 2823 16745 2832 16779
rect 2780 16736 2832 16745
rect 4528 16736 4580 16788
rect 4896 16736 4948 16788
rect 3884 16668 3936 16720
rect 4344 16668 4396 16720
rect 8300 16736 8352 16788
rect 13728 16736 13780 16788
rect 15568 16736 15620 16788
rect 16856 16779 16908 16788
rect 16856 16745 16865 16779
rect 16865 16745 16899 16779
rect 16899 16745 16908 16779
rect 16856 16736 16908 16745
rect 2044 16643 2096 16652
rect 2044 16609 2053 16643
rect 2053 16609 2087 16643
rect 2087 16609 2096 16643
rect 2044 16600 2096 16609
rect 2872 16600 2924 16652
rect 5540 16600 5592 16652
rect 6184 16600 6236 16652
rect 6828 16600 6880 16652
rect 7288 16668 7340 16720
rect 9864 16711 9916 16720
rect 9864 16677 9873 16711
rect 9873 16677 9907 16711
rect 9907 16677 9916 16711
rect 9864 16668 9916 16677
rect 11060 16668 11112 16720
rect 14372 16668 14424 16720
rect 15844 16668 15896 16720
rect 16488 16668 16540 16720
rect 7656 16643 7708 16652
rect 7656 16609 7665 16643
rect 7665 16609 7699 16643
rect 7699 16609 7708 16643
rect 7656 16600 7708 16609
rect 8116 16600 8168 16652
rect 11704 16600 11756 16652
rect 12348 16643 12400 16652
rect 12348 16609 12357 16643
rect 12357 16609 12391 16643
rect 12391 16609 12400 16643
rect 12348 16600 12400 16609
rect 12440 16600 12492 16652
rect 3608 16532 3660 16584
rect 7196 16532 7248 16584
rect 9220 16532 9272 16584
rect 9772 16575 9824 16584
rect 9772 16541 9781 16575
rect 9781 16541 9815 16575
rect 9815 16541 9824 16575
rect 9772 16532 9824 16541
rect 10048 16575 10100 16584
rect 10048 16541 10057 16575
rect 10057 16541 10091 16575
rect 10091 16541 10100 16575
rect 10048 16532 10100 16541
rect 12624 16575 12676 16584
rect 12624 16541 12633 16575
rect 12633 16541 12667 16575
rect 12667 16541 12676 16575
rect 12624 16532 12676 16541
rect 12808 16600 12860 16652
rect 13452 16643 13504 16652
rect 13452 16609 13461 16643
rect 13461 16609 13495 16643
rect 13495 16609 13504 16643
rect 13452 16600 13504 16609
rect 16120 16600 16172 16652
rect 18604 16600 18656 16652
rect 14740 16532 14792 16584
rect 16580 16532 16632 16584
rect 1492 16464 1544 16516
rect 4712 16464 4764 16516
rect 8024 16507 8076 16516
rect 8024 16473 8033 16507
rect 8033 16473 8067 16507
rect 8067 16473 8076 16507
rect 8024 16464 8076 16473
rect 10784 16464 10836 16516
rect 13820 16464 13872 16516
rect 13912 16464 13964 16516
rect 16028 16464 16080 16516
rect 1676 16439 1728 16448
rect 1676 16405 1685 16439
rect 1685 16405 1719 16439
rect 1719 16405 1728 16439
rect 1676 16396 1728 16405
rect 3424 16439 3476 16448
rect 3424 16405 3433 16439
rect 3433 16405 3467 16439
rect 3467 16405 3476 16439
rect 3424 16396 3476 16405
rect 5172 16439 5224 16448
rect 5172 16405 5181 16439
rect 5181 16405 5215 16439
rect 5215 16405 5224 16439
rect 5172 16396 5224 16405
rect 6000 16396 6052 16448
rect 6184 16439 6236 16448
rect 6184 16405 6193 16439
rect 6193 16405 6227 16439
rect 6227 16405 6236 16439
rect 6184 16396 6236 16405
rect 7288 16396 7340 16448
rect 8392 16439 8444 16448
rect 8392 16405 8401 16439
rect 8401 16405 8435 16439
rect 8435 16405 8444 16439
rect 8392 16396 8444 16405
rect 14372 16439 14424 16448
rect 14372 16405 14381 16439
rect 14381 16405 14415 16439
rect 14415 16405 14424 16439
rect 14372 16396 14424 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 4344 16192 4396 16244
rect 6000 16192 6052 16244
rect 9772 16192 9824 16244
rect 11888 16235 11940 16244
rect 11888 16201 11897 16235
rect 11897 16201 11931 16235
rect 11931 16201 11940 16235
rect 11888 16192 11940 16201
rect 12716 16235 12768 16244
rect 12716 16201 12725 16235
rect 12725 16201 12759 16235
rect 12759 16201 12768 16235
rect 12716 16192 12768 16201
rect 13728 16192 13780 16244
rect 14372 16192 14424 16244
rect 14832 16192 14884 16244
rect 15384 16192 15436 16244
rect 16304 16192 16356 16244
rect 18604 16235 18656 16244
rect 18604 16201 18613 16235
rect 18613 16201 18647 16235
rect 18647 16201 18656 16235
rect 18604 16192 18656 16201
rect 19524 16192 19576 16244
rect 2872 16167 2924 16176
rect 2872 16133 2881 16167
rect 2881 16133 2915 16167
rect 2915 16133 2924 16167
rect 2872 16124 2924 16133
rect 3884 16124 3936 16176
rect 5080 16124 5132 16176
rect 6552 16167 6604 16176
rect 6552 16133 6561 16167
rect 6561 16133 6595 16167
rect 6595 16133 6604 16167
rect 6552 16124 6604 16133
rect 7564 16124 7616 16176
rect 3424 16056 3476 16108
rect 3516 16056 3568 16108
rect 8024 16056 8076 16108
rect 9404 16099 9456 16108
rect 9404 16065 9413 16099
rect 9413 16065 9447 16099
rect 9447 16065 9456 16099
rect 9404 16056 9456 16065
rect 11060 16056 11112 16108
rect 15844 16167 15896 16176
rect 15844 16133 15853 16167
rect 15853 16133 15887 16167
rect 15887 16133 15896 16167
rect 15844 16124 15896 16133
rect 19984 16124 20036 16176
rect 13912 16099 13964 16108
rect 4344 15988 4396 16040
rect 9864 15988 9916 16040
rect 11888 15988 11940 16040
rect 13268 15988 13320 16040
rect 13912 16065 13921 16099
rect 13921 16065 13955 16099
rect 13955 16065 13964 16099
rect 13912 16056 13964 16065
rect 14280 15988 14332 16040
rect 1492 15963 1544 15972
rect 1492 15929 1501 15963
rect 1501 15929 1535 15963
rect 1535 15929 1544 15963
rect 1492 15920 1544 15929
rect 1676 15920 1728 15972
rect 2228 15920 2280 15972
rect 3516 15920 3568 15972
rect 3700 15963 3752 15972
rect 3700 15929 3709 15963
rect 3709 15929 3743 15963
rect 3743 15929 3752 15963
rect 3700 15920 3752 15929
rect 4804 15920 4856 15972
rect 6184 15920 6236 15972
rect 7104 15920 7156 15972
rect 7472 15963 7524 15972
rect 7472 15929 7481 15963
rect 7481 15929 7515 15963
rect 7515 15929 7524 15963
rect 7472 15920 7524 15929
rect 11520 15963 11572 15972
rect 5264 15852 5316 15904
rect 5724 15895 5776 15904
rect 5724 15861 5733 15895
rect 5733 15861 5767 15895
rect 5767 15861 5776 15895
rect 5724 15852 5776 15861
rect 5908 15852 5960 15904
rect 9128 15852 9180 15904
rect 11520 15929 11529 15963
rect 11529 15929 11563 15963
rect 11563 15929 11572 15963
rect 11520 15920 11572 15929
rect 13544 15920 13596 15972
rect 16764 16031 16816 16040
rect 16764 15997 16773 16031
rect 16773 15997 16807 16031
rect 16807 15997 16816 16031
rect 16764 15988 16816 15997
rect 11704 15852 11756 15904
rect 15384 15963 15436 15972
rect 15384 15929 15393 15963
rect 15393 15929 15427 15963
rect 15427 15929 15436 15963
rect 15384 15920 15436 15929
rect 15568 15852 15620 15904
rect 16580 15895 16632 15904
rect 16580 15861 16589 15895
rect 16589 15861 16623 15895
rect 16623 15861 16632 15895
rect 16580 15852 16632 15861
rect 18236 15895 18288 15904
rect 18236 15861 18245 15895
rect 18245 15861 18279 15895
rect 18279 15861 18288 15895
rect 18236 15852 18288 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2044 15648 2096 15700
rect 4344 15648 4396 15700
rect 4620 15691 4672 15700
rect 4620 15657 4629 15691
rect 4629 15657 4663 15691
rect 4663 15657 4672 15691
rect 4620 15648 4672 15657
rect 5264 15691 5316 15700
rect 5264 15657 5273 15691
rect 5273 15657 5307 15691
rect 5307 15657 5316 15691
rect 5264 15648 5316 15657
rect 6552 15648 6604 15700
rect 7288 15691 7340 15700
rect 7288 15657 7297 15691
rect 7297 15657 7331 15691
rect 7331 15657 7340 15691
rect 7288 15648 7340 15657
rect 8024 15648 8076 15700
rect 9956 15648 10008 15700
rect 11244 15648 11296 15700
rect 13360 15648 13412 15700
rect 13452 15648 13504 15700
rect 14280 15691 14332 15700
rect 14280 15657 14289 15691
rect 14289 15657 14323 15691
rect 14323 15657 14332 15691
rect 14280 15648 14332 15657
rect 15384 15691 15436 15700
rect 15384 15657 15393 15691
rect 15393 15657 15427 15691
rect 15427 15657 15436 15691
rect 15384 15648 15436 15657
rect 1676 15623 1728 15632
rect 1676 15589 1685 15623
rect 1685 15589 1719 15623
rect 1719 15589 1728 15623
rect 1676 15580 1728 15589
rect 2320 15580 2372 15632
rect 3424 15580 3476 15632
rect 4252 15580 4304 15632
rect 8760 15580 8812 15632
rect 9588 15580 9640 15632
rect 12716 15623 12768 15632
rect 12716 15589 12725 15623
rect 12725 15589 12759 15623
rect 12759 15589 12768 15623
rect 12716 15580 12768 15589
rect 18420 15623 18472 15632
rect 18420 15589 18429 15623
rect 18429 15589 18463 15623
rect 18463 15589 18472 15623
rect 18420 15580 18472 15589
rect 5448 15555 5500 15564
rect 5448 15521 5457 15555
rect 5457 15521 5491 15555
rect 5491 15521 5500 15555
rect 5448 15512 5500 15521
rect 5908 15555 5960 15564
rect 5908 15521 5917 15555
rect 5917 15521 5951 15555
rect 5951 15521 5960 15555
rect 5908 15512 5960 15521
rect 6184 15555 6236 15564
rect 6184 15521 6193 15555
rect 6193 15521 6227 15555
rect 6227 15521 6236 15555
rect 6184 15512 6236 15521
rect 6368 15555 6420 15564
rect 6368 15521 6377 15555
rect 6377 15521 6411 15555
rect 6411 15521 6420 15555
rect 6368 15512 6420 15521
rect 8300 15555 8352 15564
rect 8300 15521 8309 15555
rect 8309 15521 8343 15555
rect 8343 15521 8352 15555
rect 8300 15512 8352 15521
rect 8668 15512 8720 15564
rect 11796 15512 11848 15564
rect 14004 15512 14056 15564
rect 14740 15512 14792 15564
rect 15844 15555 15896 15564
rect 15844 15521 15853 15555
rect 15853 15521 15887 15555
rect 15887 15521 15896 15555
rect 15844 15512 15896 15521
rect 16856 15555 16908 15564
rect 16856 15521 16865 15555
rect 16865 15521 16899 15555
rect 16899 15521 16908 15555
rect 16856 15512 16908 15521
rect 18144 15512 18196 15564
rect 1216 15444 1268 15496
rect 2780 15444 2832 15496
rect 2964 15444 3016 15496
rect 5172 15444 5224 15496
rect 9404 15444 9456 15496
rect 9496 15444 9548 15496
rect 10508 15444 10560 15496
rect 11980 15444 12032 15496
rect 12992 15444 13044 15496
rect 13912 15444 13964 15496
rect 17224 15444 17276 15496
rect 6092 15376 6144 15428
rect 10784 15376 10836 15428
rect 12256 15376 12308 15428
rect 3056 15351 3108 15360
rect 3056 15317 3065 15351
rect 3065 15317 3099 15351
rect 3099 15317 3108 15351
rect 3056 15308 3108 15317
rect 3516 15351 3568 15360
rect 3516 15317 3525 15351
rect 3525 15317 3559 15351
rect 3559 15317 3568 15351
rect 3516 15308 3568 15317
rect 4528 15308 4580 15360
rect 12348 15308 12400 15360
rect 13636 15351 13688 15360
rect 13636 15317 13645 15351
rect 13645 15317 13679 15351
rect 13679 15317 13688 15351
rect 13636 15308 13688 15317
rect 17224 15308 17276 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2688 15104 2740 15156
rect 4528 15104 4580 15156
rect 8668 15104 8720 15156
rect 9036 15104 9088 15156
rect 9496 15104 9548 15156
rect 11796 15104 11848 15156
rect 12716 15104 12768 15156
rect 13360 15104 13412 15156
rect 14004 15104 14056 15156
rect 14740 15104 14792 15156
rect 17316 15104 17368 15156
rect 18144 15104 18196 15156
rect 2320 15036 2372 15088
rect 4252 15079 4304 15088
rect 4252 15045 4261 15079
rect 4261 15045 4295 15079
rect 4295 15045 4304 15079
rect 4252 15036 4304 15045
rect 5448 15036 5500 15088
rect 12348 15036 12400 15088
rect 15844 15036 15896 15088
rect 1584 15011 1636 15020
rect 1584 14977 1593 15011
rect 1593 14977 1627 15011
rect 1627 14977 1636 15011
rect 1584 14968 1636 14977
rect 3056 15011 3108 15020
rect 3056 14977 3065 15011
rect 3065 14977 3099 15011
rect 3099 14977 3108 15011
rect 3056 14968 3108 14977
rect 4712 14968 4764 15020
rect 5264 14968 5316 15020
rect 6736 14968 6788 15020
rect 2044 14832 2096 14884
rect 7104 14943 7156 14952
rect 7104 14909 7113 14943
rect 7113 14909 7147 14943
rect 7147 14909 7156 14943
rect 7104 14900 7156 14909
rect 7288 14943 7340 14952
rect 7288 14909 7297 14943
rect 7297 14909 7331 14943
rect 7331 14909 7340 14943
rect 7288 14900 7340 14909
rect 9956 14968 10008 15020
rect 8116 14943 8168 14952
rect 8116 14909 8125 14943
rect 8125 14909 8159 14943
rect 8159 14909 8168 14943
rect 8116 14900 8168 14909
rect 10692 14900 10744 14952
rect 13728 14968 13780 15020
rect 13912 14968 13964 15020
rect 11520 14900 11572 14952
rect 16028 14900 16080 14952
rect 16856 14900 16908 14952
rect 2688 14832 2740 14884
rect 3608 14832 3660 14884
rect 7472 14832 7524 14884
rect 10508 14875 10560 14884
rect 6736 14764 6788 14816
rect 7104 14807 7156 14816
rect 7104 14773 7113 14807
rect 7113 14773 7147 14807
rect 7147 14773 7156 14807
rect 7104 14764 7156 14773
rect 8300 14764 8352 14816
rect 9588 14807 9640 14816
rect 9588 14773 9597 14807
rect 9597 14773 9631 14807
rect 9631 14773 9640 14807
rect 9588 14764 9640 14773
rect 9680 14764 9732 14816
rect 10508 14841 10517 14875
rect 10517 14841 10551 14875
rect 10551 14841 10560 14875
rect 10508 14832 10560 14841
rect 11980 14832 12032 14884
rect 13636 14832 13688 14884
rect 14832 14832 14884 14884
rect 11520 14807 11572 14816
rect 11520 14773 11529 14807
rect 11529 14773 11563 14807
rect 11563 14773 11572 14807
rect 11520 14764 11572 14773
rect 12348 14764 12400 14816
rect 16212 14764 16264 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1676 14603 1728 14612
rect 1676 14569 1685 14603
rect 1685 14569 1719 14603
rect 1719 14569 1728 14603
rect 1676 14560 1728 14569
rect 2044 14603 2096 14612
rect 2044 14569 2053 14603
rect 2053 14569 2087 14603
rect 2087 14569 2096 14603
rect 2044 14560 2096 14569
rect 2780 14560 2832 14612
rect 4712 14560 4764 14612
rect 6368 14560 6420 14612
rect 6828 14560 6880 14612
rect 7012 14560 7064 14612
rect 2228 14535 2280 14544
rect 2228 14501 2237 14535
rect 2237 14501 2271 14535
rect 2271 14501 2280 14535
rect 2228 14492 2280 14501
rect 2504 14492 2556 14544
rect 3240 14492 3292 14544
rect 3700 14492 3752 14544
rect 5172 14492 5224 14544
rect 4252 14424 4304 14476
rect 5448 14467 5500 14476
rect 5448 14433 5457 14467
rect 5457 14433 5491 14467
rect 5491 14433 5500 14467
rect 5448 14424 5500 14433
rect 7932 14492 7984 14544
rect 9404 14603 9456 14612
rect 9404 14569 9413 14603
rect 9413 14569 9447 14603
rect 9447 14569 9456 14603
rect 9404 14560 9456 14569
rect 11612 14560 11664 14612
rect 12624 14603 12676 14612
rect 8760 14492 8812 14544
rect 6000 14424 6052 14476
rect 6184 14467 6236 14476
rect 6184 14433 6193 14467
rect 6193 14433 6227 14467
rect 6227 14433 6236 14467
rect 6184 14424 6236 14433
rect 6552 14467 6604 14476
rect 6552 14433 6561 14467
rect 6561 14433 6595 14467
rect 6595 14433 6604 14467
rect 6552 14424 6604 14433
rect 7288 14424 7340 14476
rect 10416 14492 10468 14544
rect 11336 14492 11388 14544
rect 12624 14569 12633 14603
rect 12633 14569 12667 14603
rect 12667 14569 12676 14603
rect 12624 14560 12676 14569
rect 12992 14603 13044 14612
rect 12992 14569 13001 14603
rect 13001 14569 13035 14603
rect 13035 14569 13044 14603
rect 12992 14560 13044 14569
rect 13176 14560 13228 14612
rect 13728 14560 13780 14612
rect 14556 14603 14608 14612
rect 14556 14569 14565 14603
rect 14565 14569 14599 14603
rect 14599 14569 14608 14603
rect 14556 14560 14608 14569
rect 16212 14603 16264 14612
rect 16212 14569 16221 14603
rect 16221 14569 16255 14603
rect 16255 14569 16264 14603
rect 16212 14560 16264 14569
rect 19524 14560 19576 14612
rect 20260 14560 20312 14612
rect 13636 14492 13688 14544
rect 13912 14535 13964 14544
rect 13912 14501 13921 14535
rect 13921 14501 13955 14535
rect 13955 14501 13964 14535
rect 13912 14492 13964 14501
rect 15476 14492 15528 14544
rect 15384 14424 15436 14476
rect 3792 14356 3844 14408
rect 6552 14288 6604 14340
rect 11796 14356 11848 14408
rect 18144 14356 18196 14408
rect 11980 14288 12032 14340
rect 14280 14263 14332 14272
rect 14280 14229 14289 14263
rect 14289 14229 14323 14263
rect 14323 14229 14332 14263
rect 14280 14220 14332 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 3148 14016 3200 14068
rect 1952 13880 2004 13932
rect 2228 13923 2280 13932
rect 2228 13889 2237 13923
rect 2237 13889 2271 13923
rect 2271 13889 2280 13923
rect 2228 13880 2280 13889
rect 3056 13855 3108 13864
rect 3056 13821 3065 13855
rect 3065 13821 3099 13855
rect 3099 13821 3108 13855
rect 3056 13812 3108 13821
rect 5448 14016 5500 14068
rect 6736 14016 6788 14068
rect 9956 14016 10008 14068
rect 10416 14059 10468 14068
rect 10416 14025 10425 14059
rect 10425 14025 10459 14059
rect 10459 14025 10468 14059
rect 10416 14016 10468 14025
rect 4988 13880 5040 13932
rect 9220 13948 9272 14000
rect 9588 13948 9640 14000
rect 10968 14016 11020 14068
rect 11888 14016 11940 14068
rect 13360 14059 13412 14068
rect 13360 14025 13369 14059
rect 13369 14025 13403 14059
rect 13403 14025 13412 14059
rect 13360 14016 13412 14025
rect 14832 14016 14884 14068
rect 15384 14016 15436 14068
rect 11520 13948 11572 14000
rect 13084 13948 13136 14000
rect 13452 13948 13504 14000
rect 5172 13855 5224 13864
rect 5172 13821 5181 13855
rect 5181 13821 5215 13855
rect 5215 13821 5224 13855
rect 5172 13812 5224 13821
rect 5540 13812 5592 13864
rect 6460 13812 6512 13864
rect 7012 13855 7064 13864
rect 7012 13821 7021 13855
rect 7021 13821 7055 13855
rect 7055 13821 7064 13855
rect 7012 13812 7064 13821
rect 7288 13855 7340 13864
rect 7288 13821 7297 13855
rect 7297 13821 7331 13855
rect 7331 13821 7340 13855
rect 7288 13812 7340 13821
rect 12624 13880 12676 13932
rect 9128 13855 9180 13864
rect 1676 13787 1728 13796
rect 1676 13753 1685 13787
rect 1685 13753 1719 13787
rect 1719 13753 1728 13787
rect 1676 13744 1728 13753
rect 2044 13744 2096 13796
rect 4252 13787 4304 13796
rect 4252 13753 4261 13787
rect 4261 13753 4295 13787
rect 4295 13753 4304 13787
rect 4252 13744 4304 13753
rect 6828 13744 6880 13796
rect 9128 13821 9137 13855
rect 9137 13821 9171 13855
rect 9171 13821 9180 13855
rect 9128 13812 9180 13821
rect 11888 13812 11940 13864
rect 14464 13880 14516 13932
rect 15476 13923 15528 13932
rect 15476 13889 15485 13923
rect 15485 13889 15519 13923
rect 15519 13889 15528 13923
rect 15476 13880 15528 13889
rect 15844 13948 15896 14000
rect 9312 13744 9364 13796
rect 2504 13719 2556 13728
rect 2504 13685 2513 13719
rect 2513 13685 2547 13719
rect 2547 13685 2556 13719
rect 2504 13676 2556 13685
rect 4528 13719 4580 13728
rect 4528 13685 4537 13719
rect 4537 13685 4571 13719
rect 4571 13685 4580 13719
rect 4528 13676 4580 13685
rect 6920 13719 6972 13728
rect 6920 13685 6929 13719
rect 6929 13685 6963 13719
rect 6963 13685 6972 13719
rect 6920 13676 6972 13685
rect 8760 13676 8812 13728
rect 8852 13676 8904 13728
rect 10968 13744 11020 13796
rect 11336 13744 11388 13796
rect 12532 13744 12584 13796
rect 13636 13787 13688 13796
rect 13636 13753 13645 13787
rect 13645 13753 13679 13787
rect 13679 13753 13688 13787
rect 13636 13744 13688 13753
rect 14280 13812 14332 13864
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1676 13515 1728 13524
rect 1676 13481 1685 13515
rect 1685 13481 1719 13515
rect 1719 13481 1728 13515
rect 1676 13472 1728 13481
rect 2504 13515 2556 13524
rect 2504 13481 2513 13515
rect 2513 13481 2547 13515
rect 2547 13481 2556 13515
rect 2504 13472 2556 13481
rect 3792 13515 3844 13524
rect 3792 13481 3801 13515
rect 3801 13481 3835 13515
rect 3835 13481 3844 13515
rect 3792 13472 3844 13481
rect 5264 13515 5316 13524
rect 5264 13481 5273 13515
rect 5273 13481 5307 13515
rect 5307 13481 5316 13515
rect 5264 13472 5316 13481
rect 5356 13472 5408 13524
rect 6092 13472 6144 13524
rect 6184 13472 6236 13524
rect 7288 13472 7340 13524
rect 7932 13515 7984 13524
rect 7932 13481 7941 13515
rect 7941 13481 7975 13515
rect 7975 13481 7984 13515
rect 7932 13472 7984 13481
rect 9128 13515 9180 13524
rect 9128 13481 9137 13515
rect 9137 13481 9171 13515
rect 9171 13481 9180 13515
rect 9128 13472 9180 13481
rect 11612 13515 11664 13524
rect 11612 13481 11621 13515
rect 11621 13481 11655 13515
rect 11655 13481 11664 13515
rect 11612 13472 11664 13481
rect 11980 13515 12032 13524
rect 11980 13481 11989 13515
rect 11989 13481 12023 13515
rect 12023 13481 12032 13515
rect 11980 13472 12032 13481
rect 12532 13515 12584 13524
rect 12532 13481 12541 13515
rect 12541 13481 12575 13515
rect 12575 13481 12584 13515
rect 12532 13472 12584 13481
rect 13268 13472 13320 13524
rect 15384 13515 15436 13524
rect 15384 13481 15393 13515
rect 15393 13481 15427 13515
rect 15427 13481 15436 13515
rect 15384 13472 15436 13481
rect 16948 13515 17000 13524
rect 16948 13481 16957 13515
rect 16957 13481 16991 13515
rect 16991 13481 17000 13515
rect 16948 13472 17000 13481
rect 5080 13404 5132 13456
rect 2964 13336 3016 13388
rect 3516 13336 3568 13388
rect 3976 13336 4028 13388
rect 5448 13379 5500 13388
rect 5448 13345 5457 13379
rect 5457 13345 5491 13379
rect 5491 13345 5500 13379
rect 5448 13336 5500 13345
rect 2136 13268 2188 13320
rect 3056 13268 3108 13320
rect 5356 13268 5408 13320
rect 5540 13268 5592 13320
rect 6828 13336 6880 13388
rect 7012 13336 7064 13388
rect 8024 13336 8076 13388
rect 8300 13404 8352 13456
rect 8392 13379 8444 13388
rect 8392 13345 8401 13379
rect 8401 13345 8435 13379
rect 8435 13345 8444 13379
rect 8392 13336 8444 13345
rect 11336 13404 11388 13456
rect 12348 13404 12400 13456
rect 13176 13404 13228 13456
rect 9864 13379 9916 13388
rect 9864 13345 9873 13379
rect 9873 13345 9907 13379
rect 9907 13345 9916 13379
rect 9864 13336 9916 13345
rect 10140 13336 10192 13388
rect 10692 13336 10744 13388
rect 11704 13336 11756 13388
rect 13084 13379 13136 13388
rect 13084 13345 13093 13379
rect 13093 13345 13127 13379
rect 13127 13345 13136 13379
rect 13084 13336 13136 13345
rect 13636 13336 13688 13388
rect 14096 13336 14148 13388
rect 15752 13379 15804 13388
rect 11980 13268 12032 13320
rect 12164 13311 12216 13320
rect 12164 13277 12173 13311
rect 12173 13277 12207 13311
rect 12207 13277 12216 13311
rect 12164 13268 12216 13277
rect 15752 13345 15761 13379
rect 15761 13345 15795 13379
rect 15795 13345 15804 13379
rect 15752 13336 15804 13345
rect 16856 13379 16908 13388
rect 16856 13345 16865 13379
rect 16865 13345 16899 13379
rect 16899 13345 16908 13379
rect 16856 13336 16908 13345
rect 17316 13379 17368 13388
rect 17316 13345 17325 13379
rect 17325 13345 17359 13379
rect 17359 13345 17368 13379
rect 17316 13336 17368 13345
rect 15844 13268 15896 13320
rect 2044 13200 2096 13252
rect 8852 13200 8904 13252
rect 9956 13200 10008 13252
rect 1952 13175 2004 13184
rect 1952 13141 1961 13175
rect 1961 13141 1995 13175
rect 1995 13141 2004 13175
rect 1952 13132 2004 13141
rect 2412 13132 2464 13184
rect 5080 13175 5132 13184
rect 5080 13141 5089 13175
rect 5089 13141 5123 13175
rect 5123 13141 5132 13175
rect 5080 13132 5132 13141
rect 13820 13175 13872 13184
rect 13820 13141 13829 13175
rect 13829 13141 13863 13175
rect 13863 13141 13872 13175
rect 13820 13132 13872 13141
rect 15292 13132 15344 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2964 12971 3016 12980
rect 2964 12937 2973 12971
rect 2973 12937 3007 12971
rect 3007 12937 3016 12971
rect 2964 12928 3016 12937
rect 3608 12971 3660 12980
rect 3608 12937 3617 12971
rect 3617 12937 3651 12971
rect 3651 12937 3660 12971
rect 3608 12928 3660 12937
rect 3976 12928 4028 12980
rect 5356 12971 5408 12980
rect 5356 12937 5365 12971
rect 5365 12937 5399 12971
rect 5399 12937 5408 12971
rect 5356 12928 5408 12937
rect 5448 12928 5500 12980
rect 8024 12971 8076 12980
rect 8024 12937 8033 12971
rect 8033 12937 8067 12971
rect 8067 12937 8076 12971
rect 8024 12928 8076 12937
rect 9588 12928 9640 12980
rect 10140 12971 10192 12980
rect 10140 12937 10149 12971
rect 10149 12937 10183 12971
rect 10183 12937 10192 12971
rect 10140 12928 10192 12937
rect 12532 12928 12584 12980
rect 15752 12928 15804 12980
rect 16856 12971 16908 12980
rect 16856 12937 16865 12971
rect 16865 12937 16899 12971
rect 16899 12937 16908 12971
rect 16856 12928 16908 12937
rect 2044 12835 2096 12844
rect 2044 12801 2053 12835
rect 2053 12801 2087 12835
rect 2087 12801 2096 12835
rect 2044 12792 2096 12801
rect 2504 12835 2556 12844
rect 2504 12801 2513 12835
rect 2513 12801 2547 12835
rect 2547 12801 2556 12835
rect 2504 12792 2556 12801
rect 3792 12792 3844 12844
rect 4528 12792 4580 12844
rect 9864 12860 9916 12912
rect 11704 12860 11756 12912
rect 14740 12860 14792 12912
rect 15292 12860 15344 12912
rect 3608 12724 3660 12776
rect 1676 12656 1728 12708
rect 6552 12724 6604 12776
rect 8484 12767 8536 12776
rect 5356 12656 5408 12708
rect 7012 12656 7064 12708
rect 8484 12733 8493 12767
rect 8493 12733 8527 12767
rect 8527 12733 8536 12767
rect 8484 12724 8536 12733
rect 9956 12792 10008 12844
rect 11244 12792 11296 12844
rect 12164 12792 12216 12844
rect 13820 12792 13872 12844
rect 17316 12860 17368 12912
rect 5448 12631 5500 12640
rect 5448 12597 5457 12631
rect 5457 12597 5491 12631
rect 5491 12597 5500 12631
rect 5448 12588 5500 12597
rect 7840 12588 7892 12640
rect 8852 12724 8904 12776
rect 11336 12767 11388 12776
rect 11336 12733 11345 12767
rect 11345 12733 11379 12767
rect 11379 12733 11388 12767
rect 11336 12724 11388 12733
rect 13360 12656 13412 12708
rect 13820 12699 13872 12708
rect 13820 12665 13829 12699
rect 13829 12665 13863 12699
rect 13863 12665 13872 12699
rect 13820 12656 13872 12665
rect 14188 12656 14240 12708
rect 16028 12699 16080 12708
rect 11060 12588 11112 12640
rect 14096 12631 14148 12640
rect 14096 12597 14105 12631
rect 14105 12597 14139 12631
rect 14139 12597 14148 12631
rect 14096 12588 14148 12597
rect 15200 12631 15252 12640
rect 15200 12597 15209 12631
rect 15209 12597 15243 12631
rect 15243 12597 15252 12631
rect 15200 12588 15252 12597
rect 16028 12665 16037 12699
rect 16037 12665 16071 12699
rect 16071 12665 16080 12699
rect 16028 12656 16080 12665
rect 15752 12588 15804 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1492 12384 1544 12436
rect 1952 12427 2004 12436
rect 1952 12393 1961 12427
rect 1961 12393 1995 12427
rect 1995 12393 2004 12427
rect 3792 12427 3844 12436
rect 1952 12384 2004 12393
rect 2044 12316 2096 12368
rect 2596 12359 2648 12368
rect 2596 12325 2605 12359
rect 2605 12325 2639 12359
rect 2639 12325 2648 12359
rect 2596 12316 2648 12325
rect 3792 12393 3801 12427
rect 3801 12393 3835 12427
rect 3835 12393 3844 12427
rect 3792 12384 3844 12393
rect 4620 12427 4672 12436
rect 4620 12393 4629 12427
rect 4629 12393 4663 12427
rect 4663 12393 4672 12427
rect 4620 12384 4672 12393
rect 5080 12427 5132 12436
rect 5080 12393 5089 12427
rect 5089 12393 5123 12427
rect 5123 12393 5132 12427
rect 5080 12384 5132 12393
rect 7012 12427 7064 12436
rect 7012 12393 7021 12427
rect 7021 12393 7055 12427
rect 7055 12393 7064 12427
rect 7012 12384 7064 12393
rect 7840 12384 7892 12436
rect 5356 12316 5408 12368
rect 8484 12384 8536 12436
rect 12808 12384 12860 12436
rect 13360 12427 13412 12436
rect 13360 12393 13369 12427
rect 13369 12393 13403 12427
rect 13403 12393 13412 12427
rect 13360 12384 13412 12393
rect 14832 12384 14884 12436
rect 16948 12384 17000 12436
rect 17132 12427 17184 12436
rect 17132 12393 17141 12427
rect 17141 12393 17175 12427
rect 17175 12393 17184 12427
rect 17132 12384 17184 12393
rect 10784 12359 10836 12368
rect 10784 12325 10793 12359
rect 10793 12325 10827 12359
rect 10827 12325 10836 12359
rect 10784 12316 10836 12325
rect 11428 12316 11480 12368
rect 11796 12316 11848 12368
rect 11888 12316 11940 12368
rect 13084 12359 13136 12368
rect 4436 12248 4488 12300
rect 5264 12248 5316 12300
rect 7932 12248 7984 12300
rect 8760 12291 8812 12300
rect 8760 12257 8769 12291
rect 8769 12257 8803 12291
rect 8803 12257 8812 12291
rect 8760 12248 8812 12257
rect 11980 12248 12032 12300
rect 13084 12325 13093 12359
rect 13093 12325 13127 12359
rect 13127 12325 13136 12359
rect 13084 12316 13136 12325
rect 13544 12316 13596 12368
rect 14188 12316 14240 12368
rect 14648 12316 14700 12368
rect 15384 12248 15436 12300
rect 15476 12248 15528 12300
rect 15936 12248 15988 12300
rect 17316 12291 17368 12300
rect 17316 12257 17325 12291
rect 17325 12257 17359 12291
rect 17359 12257 17368 12291
rect 17316 12248 17368 12257
rect 17592 12291 17644 12300
rect 17592 12257 17601 12291
rect 17601 12257 17635 12291
rect 17635 12257 17644 12291
rect 17592 12248 17644 12257
rect 2504 12223 2556 12232
rect 2504 12189 2513 12223
rect 2513 12189 2547 12223
rect 2547 12189 2556 12223
rect 2504 12180 2556 12189
rect 3148 12223 3200 12232
rect 3148 12189 3157 12223
rect 3157 12189 3191 12223
rect 3191 12189 3200 12223
rect 3148 12180 3200 12189
rect 10048 12180 10100 12232
rect 14188 12180 14240 12232
rect 15200 12180 15252 12232
rect 15844 12180 15896 12232
rect 16856 12112 16908 12164
rect 4712 12044 4764 12096
rect 8392 12044 8444 12096
rect 11060 12044 11112 12096
rect 15476 12044 15528 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 5356 11840 5408 11892
rect 7932 11840 7984 11892
rect 10784 11840 10836 11892
rect 11888 11840 11940 11892
rect 13544 11840 13596 11892
rect 14648 11883 14700 11892
rect 14648 11849 14657 11883
rect 14657 11849 14691 11883
rect 14691 11849 14700 11883
rect 14648 11840 14700 11849
rect 15752 11883 15804 11892
rect 15752 11849 15761 11883
rect 15761 11849 15795 11883
rect 15795 11849 15804 11883
rect 15752 11840 15804 11849
rect 15936 11840 15988 11892
rect 16580 11840 16632 11892
rect 17316 11840 17368 11892
rect 4436 11772 4488 11824
rect 8024 11772 8076 11824
rect 11980 11772 12032 11824
rect 15384 11772 15436 11824
rect 1952 11704 2004 11756
rect 2688 11704 2740 11756
rect 3148 11704 3200 11756
rect 5448 11704 5500 11756
rect 5540 11747 5592 11756
rect 5540 11713 5549 11747
rect 5549 11713 5583 11747
rect 5583 11713 5592 11747
rect 5540 11704 5592 11713
rect 8300 11704 8352 11756
rect 10048 11704 10100 11756
rect 10140 11704 10192 11756
rect 17132 11704 17184 11756
rect 6736 11636 6788 11688
rect 14832 11679 14884 11688
rect 14832 11645 14841 11679
rect 14841 11645 14875 11679
rect 14875 11645 14884 11679
rect 14832 11636 14884 11645
rect 17040 11679 17092 11688
rect 17040 11645 17049 11679
rect 17049 11645 17083 11679
rect 17083 11645 17092 11679
rect 17040 11636 17092 11645
rect 1676 11611 1728 11620
rect 1676 11577 1685 11611
rect 1685 11577 1719 11611
rect 1719 11577 1728 11611
rect 1676 11568 1728 11577
rect 3148 11611 3200 11620
rect 3148 11577 3157 11611
rect 3157 11577 3191 11611
rect 3191 11577 3200 11611
rect 3148 11568 3200 11577
rect 3240 11611 3292 11620
rect 3240 11577 3249 11611
rect 3249 11577 3283 11611
rect 3283 11577 3292 11611
rect 3240 11568 3292 11577
rect 5080 11568 5132 11620
rect 5632 11568 5684 11620
rect 2596 11543 2648 11552
rect 2596 11509 2605 11543
rect 2605 11509 2639 11543
rect 2639 11509 2648 11543
rect 2596 11500 2648 11509
rect 7840 11543 7892 11552
rect 7840 11509 7849 11543
rect 7849 11509 7883 11543
rect 7883 11509 7892 11543
rect 7840 11500 7892 11509
rect 8852 11611 8904 11620
rect 8852 11577 8861 11611
rect 8861 11577 8895 11611
rect 8895 11577 8904 11611
rect 8852 11568 8904 11577
rect 9220 11568 9272 11620
rect 10784 11568 10836 11620
rect 11888 11568 11940 11620
rect 12532 11568 12584 11620
rect 12716 11611 12768 11620
rect 12716 11577 12725 11611
rect 12725 11577 12759 11611
rect 12759 11577 12768 11611
rect 12716 11568 12768 11577
rect 13084 11568 13136 11620
rect 13360 11611 13412 11620
rect 13360 11577 13369 11611
rect 13369 11577 13403 11611
rect 13403 11577 13412 11611
rect 13360 11568 13412 11577
rect 14648 11568 14700 11620
rect 9128 11500 9180 11552
rect 14280 11500 14332 11552
rect 16764 11500 16816 11552
rect 17592 11500 17644 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1676 11339 1728 11348
rect 1676 11305 1685 11339
rect 1685 11305 1719 11339
rect 1719 11305 1728 11339
rect 1676 11296 1728 11305
rect 3148 11296 3200 11348
rect 5080 11296 5132 11348
rect 5632 11296 5684 11348
rect 6736 11339 6788 11348
rect 6736 11305 6745 11339
rect 6745 11305 6779 11339
rect 6779 11305 6788 11339
rect 6736 11296 6788 11305
rect 7840 11296 7892 11348
rect 8208 11296 8260 11348
rect 8852 11339 8904 11348
rect 8852 11305 8861 11339
rect 8861 11305 8895 11339
rect 8895 11305 8904 11339
rect 8852 11296 8904 11305
rect 10140 11296 10192 11348
rect 10784 11339 10836 11348
rect 10784 11305 10793 11339
rect 10793 11305 10827 11339
rect 10827 11305 10836 11339
rect 10784 11296 10836 11305
rect 12716 11296 12768 11348
rect 2228 11271 2280 11280
rect 2228 11237 2237 11271
rect 2237 11237 2271 11271
rect 2271 11237 2280 11271
rect 2228 11228 2280 11237
rect 2596 11228 2648 11280
rect 5356 11228 5408 11280
rect 6184 11228 6236 11280
rect 12808 11271 12860 11280
rect 12808 11237 12817 11271
rect 12817 11237 12851 11271
rect 12851 11237 12860 11271
rect 12808 11228 12860 11237
rect 13544 11296 13596 11348
rect 14464 11296 14516 11348
rect 14832 11228 14884 11280
rect 15476 11271 15528 11280
rect 15476 11237 15485 11271
rect 15485 11237 15519 11271
rect 15519 11237 15528 11271
rect 15476 11228 15528 11237
rect 16028 11271 16080 11280
rect 16028 11237 16037 11271
rect 16037 11237 16071 11271
rect 16071 11237 16080 11271
rect 16028 11228 16080 11237
rect 3240 11160 3292 11212
rect 4712 11203 4764 11212
rect 4712 11169 4721 11203
rect 4721 11169 4755 11203
rect 4755 11169 4764 11203
rect 4712 11160 4764 11169
rect 5264 11160 5316 11212
rect 6920 11160 6972 11212
rect 7104 11160 7156 11212
rect 14372 11160 14424 11212
rect 2136 11135 2188 11144
rect 2136 11101 2145 11135
rect 2145 11101 2179 11135
rect 2179 11101 2188 11135
rect 2136 11092 2188 11101
rect 2504 11092 2556 11144
rect 11244 11092 11296 11144
rect 12716 11135 12768 11144
rect 12716 11101 12725 11135
rect 12725 11101 12759 11135
rect 12759 11101 12768 11135
rect 12716 11092 12768 11101
rect 13360 11135 13412 11144
rect 13360 11101 13369 11135
rect 13369 11101 13403 11135
rect 13403 11101 13412 11135
rect 13360 11092 13412 11101
rect 14740 11092 14792 11144
rect 13820 11024 13872 11076
rect 15568 11092 15620 11144
rect 15752 11024 15804 11076
rect 3056 10999 3108 11008
rect 3056 10965 3065 10999
rect 3065 10965 3099 10999
rect 3099 10965 3108 10999
rect 3056 10956 3108 10965
rect 5356 10956 5408 11008
rect 9128 10999 9180 11008
rect 9128 10965 9137 10999
rect 9137 10965 9171 10999
rect 9171 10965 9180 10999
rect 9128 10956 9180 10965
rect 11336 10999 11388 11008
rect 11336 10965 11345 10999
rect 11345 10965 11379 10999
rect 11379 10965 11388 10999
rect 11336 10956 11388 10965
rect 11612 10999 11664 11008
rect 11612 10965 11621 10999
rect 11621 10965 11655 10999
rect 11655 10965 11664 10999
rect 11612 10956 11664 10965
rect 13544 10956 13596 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 4712 10795 4764 10804
rect 4712 10761 4721 10795
rect 4721 10761 4755 10795
rect 4755 10761 4764 10795
rect 4712 10752 4764 10761
rect 6184 10795 6236 10804
rect 6184 10761 6193 10795
rect 6193 10761 6227 10795
rect 6227 10761 6236 10795
rect 6184 10752 6236 10761
rect 6920 10752 6972 10804
rect 7104 10795 7156 10804
rect 7104 10761 7113 10795
rect 7113 10761 7147 10795
rect 7147 10761 7156 10795
rect 7104 10752 7156 10761
rect 10784 10752 10836 10804
rect 11336 10752 11388 10804
rect 14372 10752 14424 10804
rect 15476 10752 15528 10804
rect 15752 10795 15804 10804
rect 15752 10761 15761 10795
rect 15761 10761 15795 10795
rect 15795 10761 15804 10795
rect 15752 10752 15804 10761
rect 3148 10727 3200 10736
rect 3148 10693 3157 10727
rect 3157 10693 3191 10727
rect 3191 10693 3200 10727
rect 3148 10684 3200 10693
rect 7840 10684 7892 10736
rect 8300 10727 8352 10736
rect 8300 10693 8309 10727
rect 8309 10693 8343 10727
rect 8343 10693 8352 10727
rect 8300 10684 8352 10693
rect 11428 10727 11480 10736
rect 11428 10693 11437 10727
rect 11437 10693 11471 10727
rect 11471 10693 11480 10727
rect 11428 10684 11480 10693
rect 12716 10684 12768 10736
rect 2596 10659 2648 10668
rect 2596 10625 2605 10659
rect 2605 10625 2639 10659
rect 2639 10625 2648 10659
rect 2596 10616 2648 10625
rect 3056 10616 3108 10668
rect 9404 10616 9456 10668
rect 11612 10616 11664 10668
rect 13544 10616 13596 10668
rect 15568 10616 15620 10668
rect 16856 10591 16908 10600
rect 2136 10480 2188 10532
rect 2228 10412 2280 10464
rect 2872 10480 2924 10532
rect 5264 10523 5316 10532
rect 3976 10412 4028 10464
rect 5264 10489 5273 10523
rect 5273 10489 5307 10523
rect 5307 10489 5316 10523
rect 5264 10480 5316 10489
rect 5356 10523 5408 10532
rect 5356 10489 5365 10523
rect 5365 10489 5399 10523
rect 5399 10489 5408 10523
rect 5356 10480 5408 10489
rect 6000 10480 6052 10532
rect 7748 10523 7800 10532
rect 7748 10489 7757 10523
rect 7757 10489 7791 10523
rect 7791 10489 7800 10523
rect 7748 10480 7800 10489
rect 7840 10523 7892 10532
rect 7840 10489 7849 10523
rect 7849 10489 7883 10523
rect 7883 10489 7892 10523
rect 7840 10480 7892 10489
rect 9588 10480 9640 10532
rect 11336 10480 11388 10532
rect 13084 10480 13136 10532
rect 13820 10480 13872 10532
rect 14464 10523 14516 10532
rect 14464 10489 14473 10523
rect 14473 10489 14507 10523
rect 14507 10489 14516 10523
rect 14464 10480 14516 10489
rect 14740 10480 14792 10532
rect 15752 10480 15804 10532
rect 16856 10557 16865 10591
rect 16865 10557 16899 10591
rect 16899 10557 16908 10591
rect 16856 10548 16908 10557
rect 11244 10412 11296 10464
rect 14188 10412 14240 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2136 10208 2188 10260
rect 9128 10208 9180 10260
rect 9588 10208 9640 10260
rect 11244 10208 11296 10260
rect 12716 10208 12768 10260
rect 12808 10208 12860 10260
rect 13544 10251 13596 10260
rect 13544 10217 13553 10251
rect 13553 10217 13587 10251
rect 13587 10217 13596 10251
rect 13544 10208 13596 10217
rect 13636 10208 13688 10260
rect 14832 10208 14884 10260
rect 2872 10183 2924 10192
rect 2872 10149 2881 10183
rect 2881 10149 2915 10183
rect 2915 10149 2924 10183
rect 2872 10140 2924 10149
rect 6000 10183 6052 10192
rect 6000 10149 6009 10183
rect 6009 10149 6043 10183
rect 6043 10149 6052 10183
rect 6000 10140 6052 10149
rect 6276 10140 6328 10192
rect 6736 10140 6788 10192
rect 7840 10140 7892 10192
rect 8208 10183 8260 10192
rect 8208 10149 8217 10183
rect 8217 10149 8251 10183
rect 8251 10149 8260 10183
rect 8208 10140 8260 10149
rect 8944 10140 8996 10192
rect 9404 10140 9456 10192
rect 9864 10183 9916 10192
rect 9864 10149 9873 10183
rect 9873 10149 9907 10183
rect 9907 10149 9916 10183
rect 9864 10140 9916 10149
rect 14280 10140 14332 10192
rect 1676 10072 1728 10124
rect 2136 10072 2188 10124
rect 11520 10115 11572 10124
rect 11520 10081 11529 10115
rect 11529 10081 11563 10115
rect 11563 10081 11572 10115
rect 11520 10072 11572 10081
rect 5540 10004 5592 10056
rect 7564 10004 7616 10056
rect 9772 10047 9824 10056
rect 9772 10013 9781 10047
rect 9781 10013 9815 10047
rect 9815 10013 9824 10047
rect 9772 10004 9824 10013
rect 10048 10047 10100 10056
rect 10048 10013 10057 10047
rect 10057 10013 10091 10047
rect 10091 10013 10100 10047
rect 10048 10004 10100 10013
rect 11704 10004 11756 10056
rect 13084 10072 13136 10124
rect 13544 10072 13596 10124
rect 14096 10115 14148 10124
rect 14096 10081 14105 10115
rect 14105 10081 14139 10115
rect 14139 10081 14148 10115
rect 14096 10072 14148 10081
rect 15568 10072 15620 10124
rect 16856 10072 16908 10124
rect 17224 10072 17276 10124
rect 4068 9936 4120 9988
rect 5264 9936 5316 9988
rect 17316 9936 17368 9988
rect 4344 9868 4396 9920
rect 4896 9868 4948 9920
rect 10140 9868 10192 9920
rect 13728 9868 13780 9920
rect 17500 9911 17552 9920
rect 17500 9877 17509 9911
rect 17509 9877 17543 9911
rect 17543 9877 17552 9911
rect 17500 9868 17552 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2136 9707 2188 9716
rect 2136 9673 2145 9707
rect 2145 9673 2179 9707
rect 2179 9673 2188 9707
rect 2136 9664 2188 9673
rect 2596 9664 2648 9716
rect 3424 9664 3476 9716
rect 6276 9707 6328 9716
rect 6276 9673 6285 9707
rect 6285 9673 6319 9707
rect 6319 9673 6328 9707
rect 6276 9664 6328 9673
rect 8208 9664 8260 9716
rect 10692 9707 10744 9716
rect 10692 9673 10701 9707
rect 10701 9673 10735 9707
rect 10735 9673 10744 9707
rect 10692 9664 10744 9673
rect 11060 9664 11112 9716
rect 13544 9664 13596 9716
rect 17224 9664 17276 9716
rect 5540 9596 5592 9648
rect 6000 9596 6052 9648
rect 6368 9596 6420 9648
rect 3976 9460 4028 9512
rect 8024 9596 8076 9648
rect 8944 9639 8996 9648
rect 8944 9605 8953 9639
rect 8953 9605 8987 9639
rect 8987 9605 8996 9639
rect 8944 9596 8996 9605
rect 11520 9596 11572 9648
rect 12624 9596 12676 9648
rect 10692 9460 10744 9512
rect 5908 9435 5960 9444
rect 5908 9401 5917 9435
rect 5917 9401 5951 9435
rect 5951 9401 5960 9435
rect 5908 9392 5960 9401
rect 8208 9392 8260 9444
rect 8392 9435 8444 9444
rect 8392 9401 8401 9435
rect 8401 9401 8435 9435
rect 8435 9401 8444 9435
rect 8392 9392 8444 9401
rect 3148 9324 3200 9376
rect 4896 9367 4948 9376
rect 4896 9333 4905 9367
rect 4905 9333 4939 9367
rect 4939 9333 4948 9367
rect 4896 9324 4948 9333
rect 8760 9392 8812 9444
rect 9864 9392 9916 9444
rect 13728 9460 13780 9512
rect 15752 9460 15804 9512
rect 17040 9460 17092 9512
rect 11520 9435 11572 9444
rect 11520 9401 11529 9435
rect 11529 9401 11563 9435
rect 11563 9401 11572 9435
rect 11520 9392 11572 9401
rect 12532 9435 12584 9444
rect 12532 9401 12541 9435
rect 12541 9401 12575 9435
rect 12575 9401 12584 9435
rect 12532 9392 12584 9401
rect 13176 9435 13228 9444
rect 10140 9324 10192 9376
rect 12440 9324 12492 9376
rect 13176 9401 13185 9435
rect 13185 9401 13219 9435
rect 13219 9401 13228 9435
rect 13176 9392 13228 9401
rect 14924 9392 14976 9444
rect 14280 9367 14332 9376
rect 14280 9333 14289 9367
rect 14289 9333 14323 9367
rect 14323 9333 14332 9367
rect 14280 9324 14332 9333
rect 15384 9324 15436 9376
rect 15568 9367 15620 9376
rect 15568 9333 15577 9367
rect 15577 9333 15611 9367
rect 15611 9333 15620 9367
rect 15568 9324 15620 9333
rect 16856 9324 16908 9376
rect 17040 9324 17092 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2044 9120 2096 9172
rect 2412 9120 2464 9172
rect 4068 9120 4120 9172
rect 7564 9163 7616 9172
rect 7564 9129 7573 9163
rect 7573 9129 7607 9163
rect 7607 9129 7616 9163
rect 7564 9120 7616 9129
rect 8116 9163 8168 9172
rect 8116 9129 8125 9163
rect 8125 9129 8159 9163
rect 8159 9129 8168 9163
rect 8116 9120 8168 9129
rect 8208 9120 8260 9172
rect 9772 9120 9824 9172
rect 11704 9120 11756 9172
rect 12532 9120 12584 9172
rect 13728 9163 13780 9172
rect 1400 9052 1452 9104
rect 2596 8984 2648 9036
rect 5908 9052 5960 9104
rect 6552 9052 6604 9104
rect 2872 8984 2924 9036
rect 5172 8984 5224 9036
rect 5540 8916 5592 8968
rect 6368 8959 6420 8968
rect 6368 8925 6377 8959
rect 6377 8925 6411 8959
rect 6411 8925 6420 8959
rect 6368 8916 6420 8925
rect 6460 8916 6512 8968
rect 9496 8984 9548 9036
rect 11060 9052 11112 9104
rect 11888 9095 11940 9104
rect 11888 9061 11891 9095
rect 11891 9061 11925 9095
rect 11925 9061 11940 9095
rect 11888 9052 11940 9061
rect 12256 9052 12308 9104
rect 10140 8984 10192 9036
rect 11520 9027 11572 9036
rect 11520 8993 11529 9027
rect 11529 8993 11563 9027
rect 11563 8993 11572 9027
rect 11520 8984 11572 8993
rect 10692 8959 10744 8968
rect 10692 8925 10701 8959
rect 10701 8925 10735 8959
rect 10735 8925 10744 8959
rect 10692 8916 10744 8925
rect 13728 9129 13737 9163
rect 13737 9129 13771 9163
rect 13771 9129 13780 9163
rect 13728 9120 13780 9129
rect 15384 9052 15436 9104
rect 15752 9052 15804 9104
rect 13544 9027 13596 9036
rect 13544 8993 13553 9027
rect 13553 8993 13587 9027
rect 13587 8993 13596 9027
rect 13544 8984 13596 8993
rect 14096 8984 14148 9036
rect 14556 8984 14608 9036
rect 16856 9027 16908 9036
rect 16856 8993 16865 9027
rect 16865 8993 16899 9027
rect 16899 8993 16908 9027
rect 16856 8984 16908 8993
rect 14924 8916 14976 8968
rect 17040 8916 17092 8968
rect 848 8848 900 8900
rect 4436 8848 4488 8900
rect 6000 8848 6052 8900
rect 11152 8848 11204 8900
rect 12532 8848 12584 8900
rect 15936 8891 15988 8900
rect 8392 8780 8444 8832
rect 12440 8823 12492 8832
rect 12440 8789 12449 8823
rect 12449 8789 12483 8823
rect 12483 8789 12492 8823
rect 12440 8780 12492 8789
rect 14556 8823 14608 8832
rect 14556 8789 14565 8823
rect 14565 8789 14599 8823
rect 14599 8789 14608 8823
rect 14556 8780 14608 8789
rect 15936 8857 15945 8891
rect 15945 8857 15979 8891
rect 15979 8857 15988 8891
rect 15936 8848 15988 8857
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1584 8576 1636 8628
rect 2320 8576 2372 8628
rect 2872 8619 2924 8628
rect 2872 8585 2881 8619
rect 2881 8585 2915 8619
rect 2915 8585 2924 8619
rect 2872 8576 2924 8585
rect 3332 8619 3384 8628
rect 3332 8585 3341 8619
rect 3341 8585 3375 8619
rect 3375 8585 3384 8619
rect 3332 8576 3384 8585
rect 5172 8576 5224 8628
rect 6552 8619 6604 8628
rect 6552 8585 6561 8619
rect 6561 8585 6595 8619
rect 6595 8585 6604 8619
rect 6552 8576 6604 8585
rect 7748 8576 7800 8628
rect 7932 8576 7984 8628
rect 11060 8619 11112 8628
rect 11060 8585 11069 8619
rect 11069 8585 11103 8619
rect 11103 8585 11112 8619
rect 11060 8576 11112 8585
rect 15660 8576 15712 8628
rect 7564 8508 7616 8560
rect 13544 8508 13596 8560
rect 2688 8440 2740 8492
rect 8116 8440 8168 8492
rect 20 8372 72 8424
rect 2228 8372 2280 8424
rect 3332 8372 3384 8424
rect 6184 8415 6236 8424
rect 6184 8381 6193 8415
rect 6193 8381 6227 8415
rect 6227 8381 6236 8415
rect 6184 8372 6236 8381
rect 6828 8372 6880 8424
rect 10600 8440 10652 8492
rect 12256 8440 12308 8492
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 13176 8483 13228 8492
rect 13176 8449 13185 8483
rect 13185 8449 13219 8483
rect 13219 8449 13228 8483
rect 13176 8440 13228 8449
rect 13636 8440 13688 8492
rect 14556 8440 14608 8492
rect 14372 8415 14424 8424
rect 1676 8304 1728 8356
rect 5172 8304 5224 8356
rect 7932 8304 7984 8356
rect 9496 8304 9548 8356
rect 14372 8381 14381 8415
rect 14381 8381 14415 8415
rect 14415 8381 14424 8415
rect 14372 8372 14424 8381
rect 12348 8304 12400 8356
rect 5540 8279 5592 8288
rect 5540 8245 5549 8279
rect 5549 8245 5583 8279
rect 5583 8245 5592 8279
rect 5540 8236 5592 8245
rect 9128 8279 9180 8288
rect 9128 8245 9137 8279
rect 9137 8245 9171 8279
rect 9171 8245 9180 8279
rect 9128 8236 9180 8245
rect 10048 8279 10100 8288
rect 10048 8245 10057 8279
rect 10057 8245 10091 8279
rect 10091 8245 10100 8279
rect 10048 8236 10100 8245
rect 14280 8279 14332 8288
rect 14280 8245 14289 8279
rect 14289 8245 14323 8279
rect 14323 8245 14332 8279
rect 14280 8236 14332 8245
rect 15476 8236 15528 8288
rect 15752 8236 15804 8288
rect 15844 8236 15896 8288
rect 16856 8279 16908 8288
rect 16856 8245 16865 8279
rect 16865 8245 16899 8279
rect 16899 8245 16908 8279
rect 16856 8236 16908 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 6460 8032 6512 8084
rect 8392 8032 8444 8084
rect 9496 8075 9548 8084
rect 9496 8041 9505 8075
rect 9505 8041 9539 8075
rect 9539 8041 9548 8075
rect 9496 8032 9548 8041
rect 11520 8032 11572 8084
rect 12348 8075 12400 8084
rect 12348 8041 12357 8075
rect 12357 8041 12391 8075
rect 12391 8041 12400 8075
rect 12348 8032 12400 8041
rect 12624 8075 12676 8084
rect 12624 8041 12633 8075
rect 12633 8041 12667 8075
rect 12667 8041 12676 8075
rect 12624 8032 12676 8041
rect 14372 8032 14424 8084
rect 7932 7964 7984 8016
rect 6000 7896 6052 7948
rect 7472 7896 7524 7948
rect 7564 7896 7616 7948
rect 10048 7964 10100 8016
rect 12256 7964 12308 8016
rect 15476 8007 15528 8016
rect 15476 7973 15485 8007
rect 15485 7973 15519 8007
rect 15519 7973 15528 8007
rect 15476 7964 15528 7973
rect 15844 7964 15896 8016
rect 9956 7939 10008 7948
rect 9956 7905 9965 7939
rect 9965 7905 9999 7939
rect 9999 7905 10008 7939
rect 9956 7896 10008 7905
rect 10324 7939 10376 7948
rect 10324 7905 10333 7939
rect 10333 7905 10367 7939
rect 10367 7905 10376 7939
rect 10324 7896 10376 7905
rect 10692 7896 10744 7948
rect 11428 7939 11480 7948
rect 11428 7905 11437 7939
rect 11437 7905 11471 7939
rect 11471 7905 11480 7939
rect 11428 7896 11480 7905
rect 13268 7939 13320 7948
rect 13268 7905 13277 7939
rect 13277 7905 13311 7939
rect 13311 7905 13320 7939
rect 13268 7896 13320 7905
rect 8116 7828 8168 7880
rect 11336 7828 11388 7880
rect 14188 7896 14240 7948
rect 17132 7896 17184 7948
rect 10324 7760 10376 7812
rect 13820 7871 13872 7880
rect 13820 7837 13829 7871
rect 13829 7837 13863 7871
rect 13863 7837 13872 7871
rect 15384 7871 15436 7880
rect 13820 7828 13872 7837
rect 15384 7837 15393 7871
rect 15393 7837 15427 7871
rect 15427 7837 15436 7871
rect 15384 7828 15436 7837
rect 15936 7803 15988 7812
rect 15936 7769 15945 7803
rect 15945 7769 15979 7803
rect 15979 7769 15988 7803
rect 15936 7760 15988 7769
rect 7288 7735 7340 7744
rect 7288 7701 7297 7735
rect 7297 7701 7331 7735
rect 7331 7701 7340 7735
rect 7288 7692 7340 7701
rect 7748 7735 7800 7744
rect 7748 7701 7757 7735
rect 7757 7701 7791 7735
rect 7791 7701 7800 7735
rect 7748 7692 7800 7701
rect 14556 7735 14608 7744
rect 14556 7701 14565 7735
rect 14565 7701 14599 7735
rect 14599 7701 14608 7735
rect 14556 7692 14608 7701
rect 16488 7692 16540 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 6000 7488 6052 7540
rect 7288 7488 7340 7540
rect 10324 7488 10376 7540
rect 13268 7488 13320 7540
rect 14188 7488 14240 7540
rect 17132 7531 17184 7540
rect 17132 7497 17141 7531
rect 17141 7497 17175 7531
rect 17175 7497 17184 7531
rect 17132 7488 17184 7497
rect 9956 7420 10008 7472
rect 17040 7420 17092 7472
rect 9496 7352 9548 7404
rect 6184 7284 6236 7336
rect 7748 7216 7800 7268
rect 8760 7259 8812 7268
rect 8760 7225 8769 7259
rect 8769 7225 8803 7259
rect 8803 7225 8812 7259
rect 8760 7216 8812 7225
rect 11244 7284 11296 7336
rect 11888 7284 11940 7336
rect 12624 7327 12676 7336
rect 12624 7293 12633 7327
rect 12633 7293 12667 7327
rect 12667 7293 12676 7327
rect 12624 7284 12676 7293
rect 14188 7284 14240 7336
rect 16488 7352 16540 7404
rect 14556 7284 14608 7336
rect 15200 7259 15252 7268
rect 15200 7225 15209 7259
rect 15209 7225 15243 7259
rect 15243 7225 15252 7259
rect 15200 7216 15252 7225
rect 16120 7216 16172 7268
rect 16212 7259 16264 7268
rect 16212 7225 16221 7259
rect 16221 7225 16255 7259
rect 16255 7225 16264 7259
rect 16212 7216 16264 7225
rect 17776 7216 17828 7268
rect 7472 7191 7524 7200
rect 7472 7157 7481 7191
rect 7481 7157 7515 7191
rect 7515 7157 7524 7191
rect 7472 7148 7524 7157
rect 9680 7191 9732 7200
rect 9680 7157 9689 7191
rect 9689 7157 9723 7191
rect 9723 7157 9732 7191
rect 9680 7148 9732 7157
rect 12072 7148 12124 7200
rect 12256 7191 12308 7200
rect 12256 7157 12265 7191
rect 12265 7157 12299 7191
rect 12299 7157 12308 7191
rect 12256 7148 12308 7157
rect 12532 7191 12584 7200
rect 12532 7157 12541 7191
rect 12541 7157 12575 7191
rect 12575 7157 12584 7191
rect 12532 7148 12584 7157
rect 15476 7191 15528 7200
rect 15476 7157 15485 7191
rect 15485 7157 15519 7191
rect 15519 7157 15528 7191
rect 15476 7148 15528 7157
rect 15936 7191 15988 7200
rect 15936 7157 15945 7191
rect 15945 7157 15979 7191
rect 15979 7157 15988 7191
rect 15936 7148 15988 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 7564 6987 7616 6996
rect 7564 6953 7573 6987
rect 7573 6953 7607 6987
rect 7607 6953 7616 6987
rect 7564 6944 7616 6953
rect 7932 6987 7984 6996
rect 7932 6953 7941 6987
rect 7941 6953 7975 6987
rect 7975 6953 7984 6987
rect 7932 6944 7984 6953
rect 9496 6944 9548 6996
rect 11428 6987 11480 6996
rect 8116 6876 8168 6928
rect 8760 6919 8812 6928
rect 8760 6885 8769 6919
rect 8769 6885 8803 6919
rect 8803 6885 8812 6919
rect 8760 6876 8812 6885
rect 11428 6953 11437 6987
rect 11437 6953 11471 6987
rect 11471 6953 11480 6987
rect 11428 6944 11480 6953
rect 12256 6944 12308 6996
rect 14280 6944 14332 6996
rect 15384 6944 15436 6996
rect 15660 6987 15712 6996
rect 15660 6953 15669 6987
rect 15669 6953 15703 6987
rect 15703 6953 15712 6987
rect 15660 6944 15712 6953
rect 15936 6944 15988 6996
rect 16212 6987 16264 6996
rect 16212 6953 16221 6987
rect 16221 6953 16255 6987
rect 16255 6953 16264 6987
rect 16212 6944 16264 6953
rect 15844 6876 15896 6928
rect 7472 6808 7524 6860
rect 9680 6851 9732 6860
rect 9680 6817 9689 6851
rect 9689 6817 9723 6851
rect 9723 6817 9732 6851
rect 9680 6808 9732 6817
rect 11244 6808 11296 6860
rect 12532 6808 12584 6860
rect 15200 6808 15252 6860
rect 17040 6851 17092 6860
rect 17040 6817 17049 6851
rect 17049 6817 17083 6851
rect 17083 6817 17092 6851
rect 17040 6808 17092 6817
rect 17500 6851 17552 6860
rect 17500 6817 17509 6851
rect 17509 6817 17543 6851
rect 17543 6817 17552 6851
rect 17500 6808 17552 6817
rect 6644 6740 6696 6792
rect 15936 6740 15988 6792
rect 16120 6740 16172 6792
rect 6368 6672 6420 6724
rect 13268 6672 13320 6724
rect 18420 6672 18472 6724
rect 10600 6647 10652 6656
rect 10600 6613 10609 6647
rect 10609 6613 10643 6647
rect 10643 6613 10652 6647
rect 10600 6604 10652 6613
rect 12900 6647 12952 6656
rect 12900 6613 12909 6647
rect 12909 6613 12943 6647
rect 12943 6613 12952 6647
rect 12900 6604 12952 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 6644 6443 6696 6452
rect 6644 6409 6653 6443
rect 6653 6409 6687 6443
rect 6687 6409 6696 6443
rect 6644 6400 6696 6409
rect 9496 6443 9548 6452
rect 9496 6409 9505 6443
rect 9505 6409 9539 6443
rect 9539 6409 9548 6443
rect 9496 6400 9548 6409
rect 9772 6400 9824 6452
rect 10600 6443 10652 6452
rect 10600 6409 10609 6443
rect 10609 6409 10643 6443
rect 10643 6409 10652 6443
rect 10600 6400 10652 6409
rect 11244 6443 11296 6452
rect 11244 6409 11253 6443
rect 11253 6409 11287 6443
rect 11287 6409 11296 6443
rect 11244 6400 11296 6409
rect 12256 6400 12308 6452
rect 15936 6443 15988 6452
rect 15936 6409 15945 6443
rect 15945 6409 15979 6443
rect 15979 6409 15988 6443
rect 15936 6400 15988 6409
rect 17040 6400 17092 6452
rect 8116 6332 8168 6384
rect 9128 6332 9180 6384
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 10140 6307 10192 6316
rect 10140 6273 10149 6307
rect 10149 6273 10183 6307
rect 10183 6273 10192 6307
rect 10140 6264 10192 6273
rect 13176 6307 13228 6316
rect 13176 6273 13185 6307
rect 13185 6273 13219 6307
rect 13219 6273 13228 6307
rect 13176 6264 13228 6273
rect 14464 6264 14516 6316
rect 15844 6264 15896 6316
rect 16488 6307 16540 6316
rect 16488 6273 16497 6307
rect 16497 6273 16531 6307
rect 16531 6273 16540 6307
rect 16488 6264 16540 6273
rect 8208 6171 8260 6180
rect 8208 6137 8217 6171
rect 8217 6137 8251 6171
rect 8251 6137 8260 6171
rect 8208 6128 8260 6137
rect 9772 6171 9824 6180
rect 9772 6137 9781 6171
rect 9781 6137 9815 6171
rect 9815 6137 9824 6171
rect 9772 6128 9824 6137
rect 12532 6171 12584 6180
rect 12532 6137 12541 6171
rect 12541 6137 12575 6171
rect 12575 6137 12584 6171
rect 12532 6128 12584 6137
rect 12624 6171 12676 6180
rect 12624 6137 12633 6171
rect 12633 6137 12667 6171
rect 12667 6137 12676 6171
rect 12624 6128 12676 6137
rect 14280 6171 14332 6180
rect 14280 6137 14289 6171
rect 14289 6137 14323 6171
rect 14323 6137 14332 6171
rect 15568 6196 15620 6248
rect 14280 6128 14332 6137
rect 7472 6103 7524 6112
rect 7472 6069 7481 6103
rect 7481 6069 7515 6103
rect 7515 6069 7524 6103
rect 7472 6060 7524 6069
rect 15384 6060 15436 6112
rect 15568 6103 15620 6112
rect 15568 6069 15577 6103
rect 15577 6069 15611 6103
rect 15611 6069 15620 6103
rect 15568 6060 15620 6069
rect 17500 6103 17552 6112
rect 17500 6069 17509 6103
rect 17509 6069 17543 6103
rect 17543 6069 17552 6103
rect 17500 6060 17552 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 12532 5856 12584 5908
rect 14464 5899 14516 5908
rect 14464 5865 14473 5899
rect 14473 5865 14507 5899
rect 14507 5865 14516 5899
rect 14464 5856 14516 5865
rect 15292 5856 15344 5908
rect 16948 5899 17000 5908
rect 16948 5865 16957 5899
rect 16957 5865 16991 5899
rect 16991 5865 17000 5899
rect 16948 5856 17000 5865
rect 18512 5899 18564 5908
rect 18512 5865 18521 5899
rect 18521 5865 18555 5899
rect 18555 5865 18564 5899
rect 18512 5856 18564 5865
rect 7932 5788 7984 5840
rect 9864 5831 9916 5840
rect 9864 5797 9873 5831
rect 9873 5797 9907 5831
rect 9907 5797 9916 5831
rect 9864 5788 9916 5797
rect 12256 5788 12308 5840
rect 12900 5788 12952 5840
rect 13728 5788 13780 5840
rect 14188 5788 14240 5840
rect 6368 5763 6420 5772
rect 6368 5729 6377 5763
rect 6377 5729 6411 5763
rect 6411 5729 6420 5763
rect 6368 5720 6420 5729
rect 6460 5720 6512 5772
rect 9128 5763 9180 5772
rect 9128 5729 9137 5763
rect 9137 5729 9171 5763
rect 9171 5729 9180 5763
rect 9128 5720 9180 5729
rect 11336 5720 11388 5772
rect 14648 5720 14700 5772
rect 16396 5720 16448 5772
rect 16764 5720 16816 5772
rect 17040 5720 17092 5772
rect 17500 5788 17552 5840
rect 18420 5763 18472 5772
rect 18420 5729 18429 5763
rect 18429 5729 18463 5763
rect 18463 5729 18472 5763
rect 18420 5720 18472 5729
rect 18880 5763 18932 5772
rect 18880 5729 18889 5763
rect 18889 5729 18923 5763
rect 18923 5729 18932 5763
rect 18880 5720 18932 5729
rect 8024 5652 8076 5704
rect 9220 5652 9272 5704
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 10968 5652 11020 5704
rect 13268 5695 13320 5704
rect 13268 5661 13277 5695
rect 13277 5661 13311 5695
rect 13311 5661 13320 5695
rect 13268 5652 13320 5661
rect 13452 5652 13504 5704
rect 13084 5584 13136 5636
rect 14280 5584 14332 5636
rect 7564 5516 7616 5568
rect 8208 5516 8260 5568
rect 11428 5516 11480 5568
rect 12624 5516 12676 5568
rect 12992 5559 13044 5568
rect 12992 5525 13001 5559
rect 13001 5525 13035 5559
rect 13035 5525 13044 5559
rect 12992 5516 13044 5525
rect 15384 5516 15436 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 6368 5355 6420 5364
rect 6368 5321 6377 5355
rect 6377 5321 6411 5355
rect 6411 5321 6420 5355
rect 6368 5312 6420 5321
rect 6460 5312 6512 5364
rect 7932 5312 7984 5364
rect 7656 5244 7708 5296
rect 7840 5176 7892 5228
rect 9864 5312 9916 5364
rect 11336 5312 11388 5364
rect 13728 5355 13780 5364
rect 13728 5321 13737 5355
rect 13737 5321 13771 5355
rect 13771 5321 13780 5355
rect 13728 5312 13780 5321
rect 16396 5355 16448 5364
rect 16396 5321 16405 5355
rect 16405 5321 16439 5355
rect 16439 5321 16448 5355
rect 16396 5312 16448 5321
rect 17408 5355 17460 5364
rect 17408 5321 17417 5355
rect 17417 5321 17451 5355
rect 17451 5321 17460 5355
rect 17408 5312 17460 5321
rect 17776 5355 17828 5364
rect 17776 5321 17785 5355
rect 17785 5321 17819 5355
rect 17819 5321 17828 5355
rect 17776 5312 17828 5321
rect 18420 5312 18472 5364
rect 18880 5355 18932 5364
rect 18880 5321 18889 5355
rect 18889 5321 18923 5355
rect 18923 5321 18932 5355
rect 18880 5312 18932 5321
rect 10876 5244 10928 5296
rect 16580 5244 16632 5296
rect 9128 5219 9180 5228
rect 9128 5185 9137 5219
rect 9137 5185 9171 5219
rect 9171 5185 9180 5219
rect 9128 5176 9180 5185
rect 11244 5176 11296 5228
rect 13084 5219 13136 5228
rect 13084 5185 13093 5219
rect 13093 5185 13127 5219
rect 13127 5185 13136 5219
rect 13084 5176 13136 5185
rect 18512 5176 18564 5228
rect 9036 5040 9088 5092
rect 9220 5108 9272 5160
rect 9772 5040 9824 5092
rect 17408 5108 17460 5160
rect 17776 5108 17828 5160
rect 12164 5040 12216 5092
rect 10048 5015 10100 5024
rect 10048 4981 10057 5015
rect 10057 4981 10091 5015
rect 10091 4981 10100 5015
rect 10048 4972 10100 4981
rect 10140 4972 10192 5024
rect 12256 4972 12308 5024
rect 12716 4972 12768 5024
rect 12992 5040 13044 5092
rect 16764 5083 16816 5092
rect 16764 5049 16773 5083
rect 16773 5049 16807 5083
rect 16807 5049 16816 5083
rect 16764 5040 16816 5049
rect 14648 5015 14700 5024
rect 14648 4981 14657 5015
rect 14657 4981 14691 5015
rect 14691 4981 14700 5015
rect 14648 4972 14700 4981
rect 14740 4972 14792 5024
rect 15568 5015 15620 5024
rect 15568 4981 15577 5015
rect 15577 4981 15611 5015
rect 15611 4981 15620 5015
rect 15568 4972 15620 4981
rect 16120 5015 16172 5024
rect 16120 4981 16129 5015
rect 16129 4981 16163 5015
rect 16163 4981 16172 5015
rect 16120 4972 16172 4981
rect 16856 4972 16908 5024
rect 18420 4972 18472 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 7656 4811 7708 4820
rect 7656 4777 7665 4811
rect 7665 4777 7699 4811
rect 7699 4777 7708 4811
rect 7656 4768 7708 4777
rect 8024 4811 8076 4820
rect 8024 4777 8033 4811
rect 8033 4777 8067 4811
rect 8067 4777 8076 4811
rect 8024 4768 8076 4777
rect 9864 4768 9916 4820
rect 12256 4768 12308 4820
rect 12992 4768 13044 4820
rect 13268 4768 13320 4820
rect 15568 4768 15620 4820
rect 16028 4768 16080 4820
rect 17040 4768 17092 4820
rect 6828 4632 6880 4684
rect 9772 4700 9824 4752
rect 16120 4700 16172 4752
rect 17500 4700 17552 4752
rect 17776 4743 17828 4752
rect 17776 4709 17785 4743
rect 17785 4709 17819 4743
rect 17819 4709 17828 4743
rect 17776 4700 17828 4709
rect 8760 4632 8812 4684
rect 9036 4632 9088 4684
rect 9680 4675 9732 4684
rect 9680 4641 9689 4675
rect 9689 4641 9723 4675
rect 9723 4641 9732 4675
rect 9680 4632 9732 4641
rect 10968 4632 11020 4684
rect 14004 4632 14056 4684
rect 14648 4632 14700 4684
rect 16948 4632 17000 4684
rect 8300 4564 8352 4616
rect 9956 4564 10008 4616
rect 13636 4564 13688 4616
rect 17132 4607 17184 4616
rect 17132 4573 17141 4607
rect 17141 4573 17175 4607
rect 17175 4573 17184 4607
rect 17132 4564 17184 4573
rect 11888 4496 11940 4548
rect 6644 4428 6696 4480
rect 8852 4428 8904 4480
rect 9312 4428 9364 4480
rect 10876 4471 10928 4480
rect 10876 4437 10885 4471
rect 10885 4437 10919 4471
rect 10919 4437 10928 4471
rect 10876 4428 10928 4437
rect 12716 4428 12768 4480
rect 16028 4428 16080 4480
rect 16212 4471 16264 4480
rect 16212 4437 16221 4471
rect 16221 4437 16255 4471
rect 16255 4437 16264 4471
rect 16212 4428 16264 4437
rect 17868 4428 17920 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 8760 4267 8812 4276
rect 6644 4199 6696 4208
rect 6644 4165 6653 4199
rect 6653 4165 6687 4199
rect 6687 4165 6696 4199
rect 6644 4156 6696 4165
rect 8300 4156 8352 4208
rect 8760 4233 8769 4267
rect 8769 4233 8803 4267
rect 8803 4233 8812 4267
rect 8760 4224 8812 4233
rect 10048 4224 10100 4276
rect 13820 4224 13872 4276
rect 14004 4267 14056 4276
rect 14004 4233 14013 4267
rect 14013 4233 14047 4267
rect 14047 4233 14056 4267
rect 14004 4224 14056 4233
rect 14648 4267 14700 4276
rect 14648 4233 14657 4267
rect 14657 4233 14691 4267
rect 14691 4233 14700 4267
rect 14648 4224 14700 4233
rect 8944 4156 8996 4208
rect 10140 4156 10192 4208
rect 7564 4088 7616 4140
rect 8852 4088 8904 4140
rect 9036 4088 9088 4140
rect 9312 4131 9364 4140
rect 9312 4097 9321 4131
rect 9321 4097 9355 4131
rect 9355 4097 9364 4131
rect 9312 4088 9364 4097
rect 10876 4088 10928 4140
rect 10968 4131 11020 4140
rect 10968 4097 10977 4131
rect 10977 4097 11011 4131
rect 11011 4097 11020 4131
rect 10968 4088 11020 4097
rect 16856 4224 16908 4276
rect 16672 4156 16724 4208
rect 17500 4199 17552 4208
rect 17500 4165 17509 4199
rect 17509 4165 17543 4199
rect 17543 4165 17552 4199
rect 17500 4156 17552 4165
rect 13452 4020 13504 4072
rect 16580 4020 16632 4072
rect 19340 4088 19392 4140
rect 17684 4020 17736 4072
rect 7564 3995 7616 4004
rect 6828 3884 6880 3936
rect 7564 3961 7573 3995
rect 7573 3961 7607 3995
rect 7607 3961 7616 3995
rect 7564 3952 7616 3961
rect 7656 3952 7708 4004
rect 9036 3995 9088 4004
rect 9036 3961 9045 3995
rect 9045 3961 9079 3995
rect 9079 3961 9088 3995
rect 9036 3952 9088 3961
rect 8760 3884 8812 3936
rect 8852 3884 8904 3936
rect 10048 3952 10100 4004
rect 12256 3995 12308 4004
rect 12256 3961 12265 3995
rect 12265 3961 12299 3995
rect 12299 3961 12308 3995
rect 12256 3952 12308 3961
rect 14740 3952 14792 4004
rect 12440 3884 12492 3936
rect 15384 3952 15436 4004
rect 15844 3995 15896 4004
rect 15844 3961 15853 3995
rect 15853 3961 15887 3995
rect 15887 3961 15896 3995
rect 15844 3952 15896 3961
rect 16304 3952 16356 4004
rect 16120 3927 16172 3936
rect 16120 3893 16129 3927
rect 16129 3893 16163 3927
rect 16163 3893 16172 3927
rect 16120 3884 16172 3893
rect 16580 3884 16632 3936
rect 17224 3884 17276 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 3884 3680 3936 3732
rect 6000 3680 6052 3732
rect 7564 3723 7616 3732
rect 7564 3689 7573 3723
rect 7573 3689 7607 3723
rect 7607 3689 7616 3723
rect 7564 3680 7616 3689
rect 9036 3723 9088 3732
rect 9036 3689 9045 3723
rect 9045 3689 9079 3723
rect 9079 3689 9088 3723
rect 9036 3680 9088 3689
rect 9680 3680 9732 3732
rect 8116 3612 8168 3664
rect 8760 3612 8812 3664
rect 5448 3544 5500 3596
rect 6276 3544 6328 3596
rect 6644 3544 6696 3596
rect 5724 3408 5776 3460
rect 8852 3476 8904 3528
rect 9312 3476 9364 3528
rect 10324 3612 10376 3664
rect 12440 3680 12492 3732
rect 13452 3680 13504 3732
rect 11244 3655 11296 3664
rect 11244 3621 11253 3655
rect 11253 3621 11287 3655
rect 11287 3621 11296 3655
rect 11244 3612 11296 3621
rect 11888 3612 11940 3664
rect 12532 3612 12584 3664
rect 14096 3680 14148 3732
rect 13820 3655 13872 3664
rect 13820 3621 13829 3655
rect 13829 3621 13863 3655
rect 13863 3621 13872 3655
rect 15476 3655 15528 3664
rect 13820 3612 13872 3621
rect 15476 3621 15485 3655
rect 15485 3621 15519 3655
rect 15519 3621 15528 3655
rect 15476 3612 15528 3621
rect 16488 3680 16540 3732
rect 17224 3680 17276 3732
rect 16212 3612 16264 3664
rect 17408 3612 17460 3664
rect 17776 3612 17828 3664
rect 18604 3655 18656 3664
rect 18604 3621 18613 3655
rect 18613 3621 18647 3655
rect 18647 3621 18656 3655
rect 18604 3612 18656 3621
rect 16672 3544 16724 3596
rect 11244 3476 11296 3528
rect 14004 3519 14056 3528
rect 11980 3408 12032 3460
rect 14004 3485 14013 3519
rect 14013 3485 14047 3519
rect 14047 3485 14056 3519
rect 14004 3476 14056 3485
rect 15844 3519 15896 3528
rect 12716 3451 12768 3460
rect 12716 3417 12725 3451
rect 12725 3417 12759 3451
rect 12759 3417 12768 3451
rect 12716 3408 12768 3417
rect 15844 3485 15853 3519
rect 15853 3485 15887 3519
rect 15887 3485 15896 3519
rect 15844 3476 15896 3485
rect 16764 3476 16816 3528
rect 18512 3519 18564 3528
rect 18512 3485 18521 3519
rect 18521 3485 18555 3519
rect 18555 3485 18564 3519
rect 18512 3476 18564 3485
rect 17132 3408 17184 3460
rect 6920 3340 6972 3392
rect 8576 3340 8628 3392
rect 14556 3340 14608 3392
rect 16396 3383 16448 3392
rect 16396 3349 16405 3383
rect 16405 3349 16439 3383
rect 16439 3349 16448 3383
rect 16396 3340 16448 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 4252 3179 4304 3188
rect 4252 3145 4261 3179
rect 4261 3145 4295 3179
rect 4295 3145 4304 3179
rect 4252 3136 4304 3145
rect 8116 3136 8168 3188
rect 10324 3179 10376 3188
rect 10324 3145 10333 3179
rect 10333 3145 10367 3179
rect 10367 3145 10376 3179
rect 10324 3136 10376 3145
rect 11888 3179 11940 3188
rect 11888 3145 11897 3179
rect 11897 3145 11931 3179
rect 11931 3145 11940 3179
rect 11888 3136 11940 3145
rect 12348 3136 12400 3188
rect 12532 3136 12584 3188
rect 13820 3136 13872 3188
rect 15476 3136 15528 3188
rect 15660 3136 15712 3188
rect 17408 3179 17460 3188
rect 17408 3145 17417 3179
rect 17417 3145 17451 3179
rect 17451 3145 17460 3179
rect 17408 3136 17460 3145
rect 18512 3136 18564 3188
rect 7932 3068 7984 3120
rect 8392 3068 8444 3120
rect 6276 3043 6328 3052
rect 6276 3009 6285 3043
rect 6285 3009 6319 3043
rect 6319 3009 6328 3043
rect 6276 3000 6328 3009
rect 7012 3043 7064 3052
rect 7012 3009 7021 3043
rect 7021 3009 7055 3043
rect 7055 3009 7064 3043
rect 7012 3000 7064 3009
rect 7656 3043 7708 3052
rect 7656 3009 7665 3043
rect 7665 3009 7699 3043
rect 7699 3009 7708 3043
rect 7656 3000 7708 3009
rect 9220 3000 9272 3052
rect 4068 2932 4120 2984
rect 4252 2932 4304 2984
rect 5172 2864 5224 2916
rect 6000 2932 6052 2984
rect 8392 2932 8444 2984
rect 8576 2907 8628 2916
rect 5264 2839 5316 2848
rect 5264 2805 5273 2839
rect 5273 2805 5307 2839
rect 5307 2805 5316 2839
rect 5264 2796 5316 2805
rect 5448 2796 5500 2848
rect 6000 2796 6052 2848
rect 6644 2839 6696 2848
rect 6644 2805 6653 2839
rect 6653 2805 6687 2839
rect 6687 2805 6696 2839
rect 6644 2796 6696 2805
rect 8576 2873 8585 2907
rect 8585 2873 8619 2907
rect 8619 2873 8628 2907
rect 8576 2864 8628 2873
rect 12072 3068 12124 3120
rect 15752 3068 15804 3120
rect 12716 3000 12768 3052
rect 8116 2796 8168 2848
rect 8760 2796 8812 2848
rect 10784 2796 10836 2848
rect 11336 2864 11388 2916
rect 12072 2864 12124 2916
rect 12624 2907 12676 2916
rect 12624 2873 12633 2907
rect 12633 2873 12667 2907
rect 12667 2873 12676 2907
rect 12624 2864 12676 2873
rect 14556 2864 14608 2916
rect 15384 2864 15436 2916
rect 16120 2864 16172 2916
rect 16396 3068 16448 3120
rect 22100 3068 22152 3120
rect 16488 3043 16540 3052
rect 16488 3009 16497 3043
rect 16497 3009 16531 3043
rect 16531 3009 16540 3043
rect 16488 3000 16540 3009
rect 16764 3043 16816 3052
rect 16764 3009 16773 3043
rect 16773 3009 16807 3043
rect 16807 3009 16816 3043
rect 16764 3000 16816 3009
rect 17960 2932 18012 2984
rect 19524 2975 19576 2984
rect 19524 2941 19533 2975
rect 19533 2941 19567 2975
rect 19567 2941 19576 2975
rect 19524 2932 19576 2941
rect 20444 2975 20496 2984
rect 20444 2941 20453 2975
rect 20453 2941 20487 2975
rect 20487 2941 20496 2975
rect 20444 2932 20496 2941
rect 18604 2864 18656 2916
rect 16212 2796 16264 2848
rect 18144 2796 18196 2848
rect 25504 2796 25556 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 5540 2592 5592 2644
rect 7104 2592 7156 2644
rect 7196 2592 7248 2644
rect 5448 2456 5500 2508
rect 9036 2592 9088 2644
rect 10784 2635 10836 2644
rect 10784 2601 10793 2635
rect 10793 2601 10827 2635
rect 10827 2601 10836 2635
rect 10784 2592 10836 2601
rect 11980 2635 12032 2644
rect 11980 2601 11989 2635
rect 11989 2601 12023 2635
rect 12023 2601 12032 2635
rect 11980 2592 12032 2601
rect 12348 2635 12400 2644
rect 12348 2601 12357 2635
rect 12357 2601 12391 2635
rect 12391 2601 12400 2635
rect 12348 2592 12400 2601
rect 14096 2635 14148 2644
rect 14096 2601 14105 2635
rect 14105 2601 14139 2635
rect 14139 2601 14148 2635
rect 14096 2592 14148 2601
rect 7748 2524 7800 2576
rect 8024 2567 8076 2576
rect 8024 2533 8033 2567
rect 8033 2533 8067 2567
rect 8067 2533 8076 2567
rect 8024 2524 8076 2533
rect 8300 2567 8352 2576
rect 8300 2533 8309 2567
rect 8309 2533 8343 2567
rect 8343 2533 8352 2567
rect 8300 2524 8352 2533
rect 8668 2524 8720 2576
rect 8852 2567 8904 2576
rect 8852 2533 8861 2567
rect 8861 2533 8895 2567
rect 8895 2533 8904 2567
rect 8852 2524 8904 2533
rect 9496 2567 9548 2576
rect 9496 2533 9505 2567
rect 9505 2533 9539 2567
rect 9539 2533 9548 2567
rect 9496 2524 9548 2533
rect 12256 2524 12308 2576
rect 12716 2567 12768 2576
rect 12716 2533 12725 2567
rect 12725 2533 12759 2567
rect 12759 2533 12768 2567
rect 12716 2524 12768 2533
rect 12808 2567 12860 2576
rect 12808 2533 12817 2567
rect 12817 2533 12851 2567
rect 12851 2533 12860 2567
rect 12808 2524 12860 2533
rect 15660 2567 15712 2576
rect 15660 2533 15669 2567
rect 15669 2533 15703 2567
rect 15703 2533 15712 2567
rect 15660 2524 15712 2533
rect 16580 2567 16632 2576
rect 16580 2533 16589 2567
rect 16589 2533 16623 2567
rect 16623 2533 16632 2567
rect 16580 2524 16632 2533
rect 16764 2524 16816 2576
rect 7196 2320 7248 2372
rect 7932 2388 7984 2440
rect 9588 2456 9640 2508
rect 14280 2456 14332 2508
rect 11244 2388 11296 2440
rect 8116 2320 8168 2372
rect 11520 2320 11572 2372
rect 14004 2388 14056 2440
rect 20536 2592 20588 2644
rect 23480 2592 23532 2644
rect 18512 2524 18564 2576
rect 17868 2456 17920 2508
rect 19340 2456 19392 2508
rect 22376 2499 22428 2508
rect 22376 2465 22385 2499
rect 22385 2465 22419 2499
rect 22419 2465 22428 2499
rect 22376 2456 22428 2465
rect 24216 2456 24268 2508
rect 16120 2363 16172 2372
rect 16120 2329 16129 2363
rect 16129 2329 16163 2363
rect 16163 2329 16172 2363
rect 16120 2320 16172 2329
rect 17132 2320 17184 2372
rect 19156 2320 19208 2372
rect 21180 2320 21232 2372
rect 24124 2320 24176 2372
rect 27528 2320 27580 2372
rect 5172 2252 5224 2304
rect 5448 2252 5500 2304
rect 6092 2252 6144 2304
rect 9588 2252 9640 2304
rect 12716 2252 12768 2304
rect 14740 2252 14792 2304
rect 19524 2252 19576 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 5448 2048 5500 2100
rect 11060 2048 11112 2100
rect 6000 1980 6052 2032
rect 13084 1980 13136 2032
rect 5264 1912 5316 1964
rect 10140 1912 10192 1964
rect 2688 824 2740 876
rect 4804 824 4856 876
<< metal2 >>
rect 32 27526 336 27554
rect 32 8430 60 27526
rect 308 27418 336 27526
rect 386 27520 442 28000
rect 1122 27520 1178 28000
rect 1950 27520 2006 28000
rect 2056 27526 2360 27554
rect 400 27418 428 27520
rect 308 27390 428 27418
rect 1136 22642 1164 27520
rect 1964 27418 1992 27520
rect 2056 27418 2084 27526
rect 1964 27390 2084 27418
rect 1490 25392 1546 25401
rect 1490 25327 1546 25336
rect 1216 25152 1268 25158
rect 1216 25094 1268 25100
rect 1124 22636 1176 22642
rect 1124 22578 1176 22584
rect 112 22432 164 22438
rect 112 22374 164 22380
rect 124 21729 152 22374
rect 110 21720 166 21729
rect 110 21655 166 21664
rect 110 20360 166 20369
rect 110 20295 166 20304
rect 124 19281 152 20295
rect 110 19272 166 19281
rect 110 19207 166 19216
rect 112 16992 164 16998
rect 112 16934 164 16940
rect 124 16153 152 16934
rect 110 16144 166 16153
rect 110 16079 166 16088
rect 1228 15502 1256 25094
rect 1504 24410 1532 25327
rect 1584 24608 1636 24614
rect 1584 24550 1636 24556
rect 1492 24404 1544 24410
rect 1492 24346 1544 24352
rect 1596 24313 1624 24550
rect 1582 24304 1638 24313
rect 1582 24239 1638 24248
rect 1676 24268 1728 24274
rect 1676 24210 1728 24216
rect 1688 24070 1716 24210
rect 1676 24064 1728 24070
rect 1676 24006 1728 24012
rect 1688 23866 1716 24006
rect 1676 23860 1728 23866
rect 1676 23802 1728 23808
rect 1492 23112 1544 23118
rect 1492 23054 1544 23060
rect 1400 22568 1452 22574
rect 1400 22510 1452 22516
rect 1412 20602 1440 22510
rect 1400 20596 1452 20602
rect 1400 20538 1452 20544
rect 1504 18970 1532 23054
rect 1582 22536 1638 22545
rect 1582 22471 1638 22480
rect 1596 22234 1624 22471
rect 1584 22228 1636 22234
rect 1584 22170 1636 22176
rect 2332 22098 2360 27526
rect 2778 27520 2834 28000
rect 3514 27520 3570 28000
rect 4342 27520 4398 28000
rect 5170 27520 5226 28000
rect 5906 27520 5962 28000
rect 6734 27520 6790 28000
rect 7300 27526 7512 27554
rect 2502 26752 2558 26761
rect 2502 26687 2558 26696
rect 2412 24608 2464 24614
rect 2412 24550 2464 24556
rect 2424 23866 2452 24550
rect 2516 23866 2544 26687
rect 2792 25362 2820 27520
rect 2780 25356 2832 25362
rect 2780 25298 2832 25304
rect 2792 24954 2820 25298
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 2780 24948 2832 24954
rect 2780 24890 2832 24896
rect 2884 24682 2912 25094
rect 2872 24676 2924 24682
rect 2872 24618 2924 24624
rect 2964 24268 3016 24274
rect 2964 24210 3016 24216
rect 2412 23860 2464 23866
rect 2412 23802 2464 23808
rect 2504 23860 2556 23866
rect 2504 23802 2556 23808
rect 2976 23798 3004 24210
rect 2964 23792 3016 23798
rect 2964 23734 3016 23740
rect 2504 23180 2556 23186
rect 2504 23122 2556 23128
rect 2516 22778 2544 23122
rect 2504 22772 2556 22778
rect 2504 22714 2556 22720
rect 3424 22568 3476 22574
rect 3424 22510 3476 22516
rect 3436 22438 3464 22510
rect 3424 22432 3476 22438
rect 3424 22374 3476 22380
rect 2044 22092 2096 22098
rect 2044 22034 2096 22040
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 2056 21894 2084 22034
rect 2504 22024 2556 22030
rect 2504 21966 2556 21972
rect 2044 21888 2096 21894
rect 2044 21830 2096 21836
rect 1584 21412 1636 21418
rect 1584 21354 1636 21360
rect 1596 20806 1624 21354
rect 2056 21049 2084 21830
rect 2516 21690 2544 21966
rect 3240 21888 3292 21894
rect 3240 21830 3292 21836
rect 2504 21684 2556 21690
rect 2504 21626 2556 21632
rect 3252 21418 3280 21830
rect 2964 21412 3016 21418
rect 2964 21354 3016 21360
rect 3240 21412 3292 21418
rect 3240 21354 3292 21360
rect 3332 21412 3384 21418
rect 3332 21354 3384 21360
rect 2976 21078 3004 21354
rect 2412 21072 2464 21078
rect 2042 21040 2098 21049
rect 2412 21014 2464 21020
rect 2964 21072 3016 21078
rect 2964 21014 3016 21020
rect 2042 20975 2098 20984
rect 1584 20800 1636 20806
rect 1584 20742 1636 20748
rect 1676 20800 1728 20806
rect 1676 20742 1728 20748
rect 1596 19990 1624 20742
rect 1688 20398 1716 20742
rect 2424 20534 2452 21014
rect 2976 20913 3004 21014
rect 2962 20904 3018 20913
rect 2962 20839 3018 20848
rect 2780 20800 2832 20806
rect 2780 20742 2832 20748
rect 2228 20528 2280 20534
rect 2228 20470 2280 20476
rect 2412 20528 2464 20534
rect 2412 20470 2464 20476
rect 1676 20392 1728 20398
rect 1676 20334 1728 20340
rect 1584 19984 1636 19990
rect 1584 19926 1636 19932
rect 2240 19922 2268 20470
rect 2596 20392 2648 20398
rect 2648 20352 2728 20380
rect 2596 20334 2648 20340
rect 2228 19916 2280 19922
rect 2228 19858 2280 19864
rect 2240 19514 2268 19858
rect 2700 19718 2728 20352
rect 2688 19712 2740 19718
rect 2688 19654 2740 19660
rect 2228 19508 2280 19514
rect 2228 19450 2280 19456
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 1676 19168 1728 19174
rect 1676 19110 1728 19116
rect 1492 18964 1544 18970
rect 1492 18906 1544 18912
rect 1504 18290 1532 18906
rect 1492 18284 1544 18290
rect 1492 18226 1544 18232
rect 1688 18154 1716 19110
rect 2240 18902 2268 19246
rect 2700 19145 2728 19654
rect 2686 19136 2742 19145
rect 2686 19071 2742 19080
rect 2792 18902 2820 20742
rect 2872 20324 2924 20330
rect 2872 20266 2924 20272
rect 2884 19514 2912 20266
rect 3252 19825 3280 21354
rect 3344 19990 3372 21354
rect 3436 20058 3464 22374
rect 3528 22001 3556 27520
rect 3792 25152 3844 25158
rect 3792 25094 3844 25100
rect 3514 21992 3570 22001
rect 3514 21927 3570 21936
rect 3516 21344 3568 21350
rect 3516 21286 3568 21292
rect 3528 20330 3556 21286
rect 3804 21146 3832 25094
rect 4356 24614 4384 27520
rect 4528 25492 4580 25498
rect 4528 25434 4580 25440
rect 4540 24954 4568 25434
rect 4712 25152 4764 25158
rect 4712 25094 4764 25100
rect 4528 24948 4580 24954
rect 4528 24890 4580 24896
rect 4724 24818 4752 25094
rect 4712 24812 4764 24818
rect 4712 24754 4764 24760
rect 4988 24812 5040 24818
rect 4988 24754 5040 24760
rect 4528 24744 4580 24750
rect 4528 24686 4580 24692
rect 4344 24608 4396 24614
rect 4344 24550 4396 24556
rect 4540 24138 4568 24686
rect 4804 24676 4856 24682
rect 4804 24618 4856 24624
rect 4712 24336 4764 24342
rect 4712 24278 4764 24284
rect 4528 24132 4580 24138
rect 4528 24074 4580 24080
rect 4540 23798 4568 24074
rect 4724 23866 4752 24278
rect 4712 23860 4764 23866
rect 4712 23802 4764 23808
rect 4436 23792 4488 23798
rect 4436 23734 4488 23740
rect 4528 23792 4580 23798
rect 4528 23734 4580 23740
rect 4448 23526 4476 23734
rect 3976 23520 4028 23526
rect 3976 23462 4028 23468
rect 4436 23520 4488 23526
rect 4436 23462 4488 23468
rect 3988 23254 4016 23462
rect 3976 23248 4028 23254
rect 3976 23190 4028 23196
rect 4528 23248 4580 23254
rect 4528 23190 4580 23196
rect 4540 22982 4568 23190
rect 4712 23112 4764 23118
rect 4712 23054 4764 23060
rect 4528 22976 4580 22982
rect 4528 22918 4580 22924
rect 4540 22710 4568 22918
rect 4724 22778 4752 23054
rect 4712 22772 4764 22778
rect 4712 22714 4764 22720
rect 4528 22704 4580 22710
rect 4528 22646 4580 22652
rect 4252 22568 4304 22574
rect 4252 22510 4304 22516
rect 4264 22438 4292 22510
rect 4344 22500 4396 22506
rect 4344 22442 4396 22448
rect 4436 22500 4488 22506
rect 4436 22442 4488 22448
rect 4252 22432 4304 22438
rect 4252 22374 4304 22380
rect 4252 21412 4304 21418
rect 4252 21354 4304 21360
rect 3792 21140 3844 21146
rect 3792 21082 3844 21088
rect 3804 20942 3832 21082
rect 4160 21072 4212 21078
rect 4160 21014 4212 21020
rect 3792 20936 3844 20942
rect 3792 20878 3844 20884
rect 3516 20324 3568 20330
rect 3516 20266 3568 20272
rect 3424 20052 3476 20058
rect 3424 19994 3476 20000
rect 3332 19984 3384 19990
rect 3332 19926 3384 19932
rect 4172 19922 4200 21014
rect 4264 20942 4292 21354
rect 4356 21146 4384 22442
rect 4448 22166 4476 22442
rect 4436 22160 4488 22166
rect 4436 22102 4488 22108
rect 4448 21690 4476 22102
rect 4436 21684 4488 21690
rect 4436 21626 4488 21632
rect 4448 21350 4476 21626
rect 4540 21486 4568 22646
rect 4712 22568 4764 22574
rect 4712 22510 4764 22516
rect 4620 22024 4672 22030
rect 4620 21966 4672 21972
rect 4528 21480 4580 21486
rect 4528 21422 4580 21428
rect 4632 21418 4660 21966
rect 4724 21894 4752 22510
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4816 21690 4844 24618
rect 5000 24206 5028 24754
rect 4988 24200 5040 24206
rect 4988 24142 5040 24148
rect 5000 23798 5028 24142
rect 4988 23792 5040 23798
rect 4988 23734 5040 23740
rect 5000 23118 5028 23734
rect 5184 23474 5212 27520
rect 5920 25498 5948 27520
rect 5908 25492 5960 25498
rect 5908 25434 5960 25440
rect 6748 25362 6776 27520
rect 6000 25356 6052 25362
rect 6000 25298 6052 25304
rect 6736 25356 6788 25362
rect 6736 25298 6788 25304
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6012 24954 6040 25298
rect 7012 25220 7064 25226
rect 7012 25162 7064 25168
rect 6920 25152 6972 25158
rect 6920 25094 6972 25100
rect 6000 24948 6052 24954
rect 6000 24890 6052 24896
rect 5356 24608 5408 24614
rect 5356 24550 5408 24556
rect 5092 23446 5212 23474
rect 4988 23112 5040 23118
rect 4988 23054 5040 23060
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 4620 21412 4672 21418
rect 4620 21354 4672 21360
rect 4436 21344 4488 21350
rect 4436 21286 4488 21292
rect 4344 21140 4396 21146
rect 4344 21082 4396 21088
rect 4252 20936 4304 20942
rect 4252 20878 4304 20884
rect 4356 20398 4384 21082
rect 4344 20392 4396 20398
rect 4344 20334 4396 20340
rect 4896 20392 4948 20398
rect 4896 20334 4948 20340
rect 4160 19916 4212 19922
rect 4160 19858 4212 19864
rect 3238 19816 3294 19825
rect 3238 19751 3294 19760
rect 2964 19712 3016 19718
rect 2964 19654 3016 19660
rect 3608 19712 3660 19718
rect 3608 19654 3660 19660
rect 2872 19508 2924 19514
rect 2872 19450 2924 19456
rect 2884 19242 2912 19450
rect 2976 19310 3004 19654
rect 3148 19372 3200 19378
rect 3148 19314 3200 19320
rect 2964 19304 3016 19310
rect 2964 19246 3016 19252
rect 2872 19236 2924 19242
rect 2872 19178 2924 19184
rect 2228 18896 2280 18902
rect 2228 18838 2280 18844
rect 2780 18896 2832 18902
rect 2780 18838 2832 18844
rect 2240 18426 2268 18838
rect 2228 18420 2280 18426
rect 2228 18362 2280 18368
rect 1676 18148 1728 18154
rect 1676 18090 1728 18096
rect 1688 17882 1716 18090
rect 2240 17882 2268 18362
rect 2792 18290 2820 18838
rect 2884 18426 2912 19178
rect 3160 18970 3188 19314
rect 3148 18964 3200 18970
rect 3148 18906 3200 18912
rect 3620 18766 3648 19654
rect 4172 19514 4200 19858
rect 4160 19508 4212 19514
rect 4160 19450 4212 19456
rect 4356 18902 4384 20334
rect 4528 20256 4580 20262
rect 4528 20198 4580 20204
rect 4540 19378 4568 20198
rect 4528 19372 4580 19378
rect 4528 19314 4580 19320
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4632 18970 4660 19110
rect 4620 18964 4672 18970
rect 4620 18906 4672 18912
rect 4344 18896 4396 18902
rect 4344 18838 4396 18844
rect 4908 18766 4936 20334
rect 4986 19272 5042 19281
rect 4986 19207 5042 19216
rect 5000 19174 5028 19207
rect 4988 19168 5040 19174
rect 4988 19110 5040 19116
rect 3608 18760 3660 18766
rect 3608 18702 3660 18708
rect 4896 18760 4948 18766
rect 4896 18702 4948 18708
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 2780 18284 2832 18290
rect 2780 18226 2832 18232
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 2228 17876 2280 17882
rect 2228 17818 2280 17824
rect 2884 17814 2912 18362
rect 2872 17808 2924 17814
rect 2872 17750 2924 17756
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2136 17536 2188 17542
rect 2136 17478 2188 17484
rect 2148 17134 2176 17478
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 2136 17128 2188 17134
rect 2136 17070 2188 17076
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 1492 16516 1544 16522
rect 1492 16458 1544 16464
rect 1504 15978 1532 16458
rect 1676 16448 1728 16454
rect 1676 16390 1728 16396
rect 1688 15978 1716 16390
rect 1492 15972 1544 15978
rect 1492 15914 1544 15920
rect 1676 15972 1728 15978
rect 1676 15914 1728 15920
rect 1216 15496 1268 15502
rect 1216 15438 1268 15444
rect 1398 12744 1454 12753
rect 1398 12679 1454 12688
rect 1412 9110 1440 12679
rect 1504 12442 1532 15914
rect 1688 15638 1716 15914
rect 2056 15706 2084 16594
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 1676 15632 1728 15638
rect 1676 15574 1728 15580
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1492 12436 1544 12442
rect 1492 12378 1544 12384
rect 1400 9104 1452 9110
rect 1400 9046 1452 9052
rect 848 8900 900 8906
rect 848 8842 900 8848
rect 20 8424 72 8430
rect 20 8366 72 8372
rect 478 82 534 480
rect 860 82 888 8842
rect 1596 8634 1624 14962
rect 1688 14618 1716 15574
rect 2056 14890 2084 15642
rect 2044 14884 2096 14890
rect 2044 14826 2096 14832
rect 2056 14618 2084 14826
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 2044 14612 2096 14618
rect 2044 14554 2096 14560
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 1676 13796 1728 13802
rect 1676 13738 1728 13744
rect 1688 13530 1716 13738
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1964 13190 1992 13874
rect 2056 13802 2084 14554
rect 2148 13814 2176 17070
rect 2228 15972 2280 15978
rect 2228 15914 2280 15920
rect 2240 14550 2268 15914
rect 2320 15632 2372 15638
rect 2320 15574 2372 15580
rect 2332 15094 2360 15574
rect 2700 15162 2728 17274
rect 2792 16794 2820 17614
rect 2884 17338 2912 17750
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 2976 17066 3004 18566
rect 3332 18216 3384 18222
rect 3332 18158 3384 18164
rect 3344 17882 3372 18158
rect 3332 17876 3384 17882
rect 3332 17818 3384 17824
rect 3332 17536 3384 17542
rect 3332 17478 3384 17484
rect 2964 17060 3016 17066
rect 2964 17002 3016 17008
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2884 16182 2912 16594
rect 2872 16176 2924 16182
rect 2872 16118 2924 16124
rect 2976 15502 3004 17002
rect 3146 16960 3202 16969
rect 3146 16895 3202 16904
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2688 15156 2740 15162
rect 2688 15098 2740 15104
rect 2320 15088 2372 15094
rect 2320 15030 2372 15036
rect 2700 14890 2728 15098
rect 2688 14884 2740 14890
rect 2688 14826 2740 14832
rect 2792 14618 2820 15438
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 3068 15026 3096 15302
rect 3056 15020 3108 15026
rect 3056 14962 3108 14968
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 2228 14544 2280 14550
rect 2228 14486 2280 14492
rect 2504 14544 2556 14550
rect 2504 14486 2556 14492
rect 2240 13938 2268 14486
rect 2228 13932 2280 13938
rect 2228 13874 2280 13880
rect 2044 13796 2096 13802
rect 2148 13786 2360 13814
rect 2044 13738 2096 13744
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2044 13252 2096 13258
rect 2044 13194 2096 13200
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 2056 12850 2084 13194
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 1676 12708 1728 12714
rect 1676 12650 1728 12656
rect 1688 11626 1716 12650
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 1964 11762 1992 12378
rect 2056 12374 2084 12786
rect 2044 12368 2096 12374
rect 2044 12310 2096 12316
rect 2148 12220 2176 13262
rect 2056 12192 2176 12220
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 1676 11620 1728 11626
rect 1676 11562 1728 11568
rect 1688 11354 1716 11562
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1688 10130 1716 11290
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 2056 9178 2084 12192
rect 2228 11280 2280 11286
rect 2228 11222 2280 11228
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2148 10538 2176 11086
rect 2136 10532 2188 10538
rect 2136 10474 2188 10480
rect 2148 10266 2176 10474
rect 2240 10470 2268 11222
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2148 9722 2176 10066
rect 2136 9716 2188 9722
rect 2136 9658 2188 9664
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 2332 8634 2360 13786
rect 2516 13734 2544 14486
rect 3160 14074 3188 16895
rect 3344 15484 3372 17478
rect 3620 17066 3648 18702
rect 3884 18624 3936 18630
rect 3884 18566 3936 18572
rect 3608 17060 3660 17066
rect 3608 17002 3660 17008
rect 3516 16992 3568 16998
rect 3516 16934 3568 16940
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3436 16114 3464 16390
rect 3528 16114 3556 16934
rect 3620 16590 3648 17002
rect 3896 16726 3924 18566
rect 4908 18426 4936 18702
rect 4896 18420 4948 18426
rect 4896 18362 4948 18368
rect 4250 18320 4306 18329
rect 4250 18255 4306 18264
rect 4988 18284 5040 18290
rect 4264 17882 4292 18255
rect 4988 18226 5040 18232
rect 4344 18080 4396 18086
rect 4344 18022 4396 18028
rect 4252 17876 4304 17882
rect 4252 17818 4304 17824
rect 4356 16726 4384 18022
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4894 17640 4950 17649
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4540 16794 4568 16934
rect 4528 16788 4580 16794
rect 4528 16730 4580 16736
rect 3884 16720 3936 16726
rect 3884 16662 3936 16668
rect 4344 16720 4396 16726
rect 4344 16662 4396 16668
rect 3608 16584 3660 16590
rect 3608 16526 3660 16532
rect 4356 16250 4384 16662
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 3884 16176 3936 16182
rect 3884 16118 3936 16124
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 3436 15638 3464 16050
rect 3516 15972 3568 15978
rect 3516 15914 3568 15920
rect 3700 15972 3752 15978
rect 3700 15914 3752 15920
rect 3424 15632 3476 15638
rect 3424 15574 3476 15580
rect 3344 15456 3464 15484
rect 3240 14544 3292 14550
rect 3240 14486 3292 14492
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 2516 13530 2544 13670
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2964 13388 3016 13394
rect 2964 13330 3016 13336
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 2424 9178 2452 13126
rect 2976 12986 3004 13330
rect 3068 13326 3096 13806
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2516 12238 2544 12786
rect 2596 12368 2648 12374
rect 2596 12310 2648 12316
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2516 11150 2544 12174
rect 2608 11558 2636 12310
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 3160 11762 3188 12174
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 3148 11756 3200 11762
rect 3252 11744 3280 14486
rect 3252 11716 3372 11744
rect 3148 11698 3200 11704
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2608 11286 2636 11494
rect 2596 11280 2648 11286
rect 2596 11222 2648 11228
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2608 9722 2636 10610
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2596 9036 2648 9042
rect 2700 9024 2728 11698
rect 3148 11620 3200 11626
rect 3148 11562 3200 11568
rect 3240 11620 3292 11626
rect 3240 11562 3292 11568
rect 3160 11354 3188 11562
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 3056 11008 3108 11014
rect 3056 10950 3108 10956
rect 3068 10674 3096 10950
rect 3160 10742 3188 11290
rect 3252 11218 3280 11562
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 3148 10736 3200 10742
rect 3148 10678 3200 10684
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 2872 10532 2924 10538
rect 2872 10474 2924 10480
rect 2884 10198 2912 10474
rect 2872 10192 2924 10198
rect 2872 10134 2924 10140
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 2648 8996 2728 9024
rect 2596 8978 2648 8984
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2700 8498 2728 8996
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2884 8634 2912 8978
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2228 8424 2280 8430
rect 2280 8401 2360 8412
rect 2280 8392 2374 8401
rect 2280 8384 2318 8392
rect 2228 8366 2280 8372
rect 1676 8356 1728 8362
rect 2318 8327 2374 8336
rect 1676 8298 1728 8304
rect 478 54 888 82
rect 1398 82 1454 480
rect 1688 82 1716 8298
rect 2688 876 2740 882
rect 2688 818 2740 824
rect 1398 54 1716 82
rect 2410 82 2466 480
rect 2700 82 2728 818
rect 2410 54 2728 82
rect 3160 82 3188 9318
rect 3344 8634 3372 11716
rect 3436 9722 3464 15456
rect 3528 15366 3556 15914
rect 3516 15360 3568 15366
rect 3516 15302 3568 15308
rect 3528 13394 3556 15302
rect 3608 14884 3660 14890
rect 3608 14826 3660 14832
rect 3516 13388 3568 13394
rect 3516 13330 3568 13336
rect 3620 12986 3648 14826
rect 3712 14550 3740 15914
rect 3700 14544 3752 14550
rect 3700 14486 3752 14492
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3804 13530 3832 14350
rect 3792 13524 3844 13530
rect 3792 13466 3844 13472
rect 3608 12980 3660 12986
rect 3608 12922 3660 12928
rect 3620 12782 3648 12922
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3608 12776 3660 12782
rect 3608 12718 3660 12724
rect 3804 12442 3832 12786
rect 3792 12436 3844 12442
rect 3792 12378 3844 12384
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3344 8430 3372 8570
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3896 3738 3924 16118
rect 4356 16046 4384 16186
rect 4344 16040 4396 16046
rect 4344 15982 4396 15988
rect 4356 15706 4384 15982
rect 4632 15706 4660 17206
rect 4724 17134 4752 17614
rect 4894 17575 4950 17584
rect 4908 17542 4936 17575
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 4908 17134 4936 17478
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4724 16522 4752 17070
rect 4908 16794 4936 17070
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 4712 16516 4764 16522
rect 4712 16458 4764 16464
rect 4804 15972 4856 15978
rect 4804 15914 4856 15920
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 4252 15632 4304 15638
rect 4252 15574 4304 15580
rect 4264 15094 4292 15574
rect 4528 15360 4580 15366
rect 4528 15302 4580 15308
rect 4540 15162 4568 15302
rect 4528 15156 4580 15162
rect 4528 15098 4580 15104
rect 4252 15088 4304 15094
rect 4304 15036 4384 15042
rect 4252 15030 4384 15036
rect 4264 15014 4384 15030
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 3974 14240 4030 14249
rect 3974 14175 4030 14184
rect 3988 13394 4016 14175
rect 4264 13802 4292 14418
rect 4252 13796 4304 13802
rect 4252 13738 4304 13744
rect 4264 13705 4292 13738
rect 4250 13696 4306 13705
rect 4250 13631 4306 13640
rect 3976 13388 4028 13394
rect 3976 13330 4028 13336
rect 3988 12986 4016 13330
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3988 9518 4016 10406
rect 4068 9988 4120 9994
rect 4068 9930 4120 9936
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 4080 9178 4108 9930
rect 4356 9926 4384 15014
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4540 12850 4568 13670
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4632 12442 4660 15642
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4724 14618 4752 14962
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4448 11830 4476 12242
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4436 11824 4488 11830
rect 4436 11766 4488 11772
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4448 8906 4476 11766
rect 4724 11218 4752 12038
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4724 10810 4752 11154
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4436 8900 4488 8906
rect 4436 8842 4488 8848
rect 4250 6352 4306 6361
rect 4250 6287 4306 6296
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 4264 3194 4292 6287
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4264 2990 4292 3130
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 4080 2689 4108 2926
rect 4066 2680 4122 2689
rect 4066 2615 4122 2624
rect 4816 882 4844 15914
rect 5000 13938 5028 18226
rect 5092 16182 5120 23446
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 5276 19718 5304 20198
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 5170 19136 5226 19145
rect 5170 19071 5226 19080
rect 5184 18970 5212 19071
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 5172 17808 5224 17814
rect 5172 17750 5224 17756
rect 5184 17116 5212 17750
rect 5276 17610 5304 19654
rect 5264 17604 5316 17610
rect 5264 17546 5316 17552
rect 5264 17128 5316 17134
rect 5184 17088 5264 17116
rect 5184 16454 5212 17088
rect 5264 17070 5316 17076
rect 5172 16448 5224 16454
rect 5172 16390 5224 16396
rect 5080 16176 5132 16182
rect 5080 16118 5132 16124
rect 5184 15502 5212 16390
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 5276 15706 5304 15846
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5172 15496 5224 15502
rect 5172 15438 5224 15444
rect 5276 15026 5304 15642
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5172 14544 5224 14550
rect 5172 14486 5224 14492
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 5184 13870 5212 14486
rect 5172 13864 5224 13870
rect 5092 13812 5172 13814
rect 5092 13806 5224 13812
rect 5092 13786 5212 13806
rect 5092 13462 5120 13786
rect 5368 13530 5396 24550
rect 6932 24342 6960 25094
rect 7024 24818 7052 25162
rect 7196 25152 7248 25158
rect 7196 25094 7248 25100
rect 7012 24812 7064 24818
rect 7012 24754 7064 24760
rect 6920 24336 6972 24342
rect 6920 24278 6972 24284
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 6932 23866 6960 24278
rect 5448 23860 5500 23866
rect 5448 23802 5500 23808
rect 6920 23860 6972 23866
rect 6920 23802 6972 23808
rect 5460 23322 5488 23802
rect 5448 23316 5500 23322
rect 5448 23258 5500 23264
rect 5460 22234 5488 23258
rect 6276 23180 6328 23186
rect 6276 23122 6328 23128
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 6288 22778 6316 23122
rect 6276 22772 6328 22778
rect 6276 22714 6328 22720
rect 6920 22568 6972 22574
rect 6920 22510 6972 22516
rect 6092 22432 6144 22438
rect 6092 22374 6144 22380
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5448 20392 5500 20398
rect 5448 20334 5500 20340
rect 5460 19961 5488 20334
rect 5446 19952 5502 19961
rect 5446 19887 5502 19896
rect 5998 19952 6054 19961
rect 5998 19887 6054 19896
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5552 19174 5580 19654
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 5460 15570 5488 18158
rect 5552 17814 5580 19110
rect 6012 18834 6040 19887
rect 6000 18828 6052 18834
rect 6000 18770 6052 18776
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6012 18426 6040 18770
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 5540 17808 5592 17814
rect 5540 17750 5592 17756
rect 5632 17740 5684 17746
rect 5632 17682 5684 17688
rect 5644 17649 5672 17682
rect 5630 17640 5686 17649
rect 5630 17575 5686 17584
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5552 17270 5580 17478
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5540 17264 5592 17270
rect 5540 17206 5592 17212
rect 5552 17134 5580 17206
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5552 15994 5580 16594
rect 6000 16448 6052 16454
rect 6000 16390 6052 16396
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6012 16250 6040 16390
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5722 16008 5778 16017
rect 5552 15966 5722 15994
rect 5722 15943 5778 15952
rect 5736 15910 5764 15943
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 5908 15904 5960 15910
rect 5908 15846 5960 15852
rect 5920 15570 5948 15846
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5908 15564 5960 15570
rect 5960 15524 6040 15552
rect 5908 15506 5960 15512
rect 5460 15094 5488 15506
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5448 15088 5500 15094
rect 5448 15030 5500 15036
rect 5460 14482 5488 15030
rect 6012 14482 6040 15524
rect 6104 15434 6132 22374
rect 6552 22092 6604 22098
rect 6552 22034 6604 22040
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 6288 20058 6316 21830
rect 6564 21350 6592 22034
rect 6932 21894 6960 22510
rect 7024 22234 7052 24754
rect 7208 24342 7236 25094
rect 7196 24336 7248 24342
rect 7196 24278 7248 24284
rect 7208 23866 7236 24278
rect 7196 23860 7248 23866
rect 7196 23802 7248 23808
rect 7300 23186 7328 27526
rect 7484 27418 7512 27526
rect 7562 27520 7618 28000
rect 8298 27554 8354 28000
rect 8298 27526 8524 27554
rect 8298 27520 8354 27526
rect 7576 27418 7604 27520
rect 7484 27390 7604 27418
rect 7380 25356 7432 25362
rect 7380 25298 7432 25304
rect 8208 25356 8260 25362
rect 8208 25298 8260 25304
rect 7392 24682 7420 25298
rect 8024 25152 8076 25158
rect 8024 25094 8076 25100
rect 8036 24886 8064 25094
rect 8024 24880 8076 24886
rect 8024 24822 8076 24828
rect 7564 24812 7616 24818
rect 7564 24754 7616 24760
rect 7380 24676 7432 24682
rect 7380 24618 7432 24624
rect 7288 23180 7340 23186
rect 7288 23122 7340 23128
rect 7392 22778 7420 24618
rect 7576 24342 7604 24754
rect 7932 24676 7984 24682
rect 7932 24618 7984 24624
rect 7564 24336 7616 24342
rect 7564 24278 7616 24284
rect 7576 23474 7604 24278
rect 7656 24200 7708 24206
rect 7656 24142 7708 24148
rect 7668 23730 7696 24142
rect 7656 23724 7708 23730
rect 7656 23666 7708 23672
rect 7944 23594 7972 24618
rect 8220 24614 8248 25298
rect 8208 24608 8260 24614
rect 8208 24550 8260 24556
rect 8220 24342 8248 24550
rect 8208 24336 8260 24342
rect 8208 24278 8260 24284
rect 7932 23588 7984 23594
rect 7932 23530 7984 23536
rect 7484 23446 7604 23474
rect 8024 23520 8076 23526
rect 8024 23462 8076 23468
rect 7484 23118 7512 23446
rect 8036 23118 8064 23462
rect 8116 23248 8168 23254
rect 8116 23190 8168 23196
rect 7472 23112 7524 23118
rect 7472 23054 7524 23060
rect 8024 23112 8076 23118
rect 8024 23054 8076 23060
rect 7380 22772 7432 22778
rect 7380 22714 7432 22720
rect 7484 22234 7512 23054
rect 7932 22976 7984 22982
rect 7932 22918 7984 22924
rect 7012 22228 7064 22234
rect 7012 22170 7064 22176
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7288 22024 7340 22030
rect 7288 21966 7340 21972
rect 6920 21888 6972 21894
rect 6920 21830 6972 21836
rect 6644 21412 6696 21418
rect 6644 21354 6696 21360
rect 6552 21344 6604 21350
rect 6552 21286 6604 21292
rect 6276 20052 6328 20058
rect 6276 19994 6328 20000
rect 6460 19916 6512 19922
rect 6460 19858 6512 19864
rect 6472 19378 6500 19858
rect 6460 19372 6512 19378
rect 6460 19314 6512 19320
rect 6368 18828 6420 18834
rect 6368 18770 6420 18776
rect 6274 18456 6330 18465
rect 6274 18391 6330 18400
rect 6288 18358 6316 18391
rect 6276 18352 6328 18358
rect 6276 18294 6328 18300
rect 6380 17066 6408 18770
rect 6472 18290 6500 19314
rect 6564 18986 6592 21286
rect 6656 19174 6684 21354
rect 6932 21146 6960 21830
rect 7300 21350 7328 21966
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 7472 21344 7524 21350
rect 7472 21286 7524 21292
rect 7748 21344 7800 21350
rect 7748 21286 7800 21292
rect 6920 21140 6972 21146
rect 6920 21082 6972 21088
rect 7012 21004 7064 21010
rect 7012 20946 7064 20952
rect 6828 20800 6880 20806
rect 6828 20742 6880 20748
rect 6736 20256 6788 20262
rect 6736 20198 6788 20204
rect 6748 19990 6776 20198
rect 6736 19984 6788 19990
rect 6736 19926 6788 19932
rect 6748 19310 6776 19926
rect 6840 19922 6868 20742
rect 7024 20398 7052 20946
rect 7012 20392 7064 20398
rect 7012 20334 7064 20340
rect 7024 20058 7052 20334
rect 7300 20262 7328 21286
rect 7484 21010 7512 21286
rect 7472 21004 7524 21010
rect 7472 20946 7524 20952
rect 7656 21004 7708 21010
rect 7656 20946 7708 20952
rect 7484 20398 7512 20946
rect 7472 20392 7524 20398
rect 7472 20334 7524 20340
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6840 19514 6868 19858
rect 7288 19848 7340 19854
rect 7288 19790 7340 19796
rect 6828 19508 6880 19514
rect 6828 19450 6880 19456
rect 6736 19304 6788 19310
rect 6736 19246 6788 19252
rect 7300 19242 7328 19790
rect 7484 19514 7512 20334
rect 7668 20330 7696 20946
rect 7760 20534 7788 21286
rect 7748 20528 7800 20534
rect 7748 20470 7800 20476
rect 7656 20324 7708 20330
rect 7656 20266 7708 20272
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7472 19508 7524 19514
rect 7472 19450 7524 19456
rect 7380 19304 7432 19310
rect 7484 19292 7512 19450
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7432 19264 7512 19292
rect 7380 19246 7432 19252
rect 7288 19236 7340 19242
rect 7288 19178 7340 19184
rect 6644 19168 6696 19174
rect 6644 19110 6696 19116
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 6564 18958 6684 18986
rect 6460 18284 6512 18290
rect 6460 18226 6512 18232
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 6564 17610 6592 17682
rect 6552 17604 6604 17610
rect 6552 17546 6604 17552
rect 6368 17060 6420 17066
rect 6368 17002 6420 17008
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 6196 16454 6224 16594
rect 6184 16448 6236 16454
rect 6184 16390 6236 16396
rect 6196 15978 6224 16390
rect 6184 15972 6236 15978
rect 6184 15914 6236 15920
rect 6380 15570 6408 17002
rect 6564 16182 6592 17546
rect 6552 16176 6604 16182
rect 6552 16118 6604 16124
rect 6564 15706 6592 16118
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 6196 15473 6224 15506
rect 6182 15464 6238 15473
rect 6092 15428 6144 15434
rect 6182 15399 6238 15408
rect 6092 15370 6144 15376
rect 6196 14482 6224 15399
rect 6380 14618 6408 15506
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 6564 14482 6592 15642
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 6184 14476 6236 14482
rect 6552 14476 6604 14482
rect 6184 14418 6236 14424
rect 6472 14436 6552 14464
rect 5460 14074 5488 14418
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5080 13456 5132 13462
rect 5080 13398 5132 13404
rect 5092 13190 5120 13398
rect 5170 13288 5226 13297
rect 5170 13223 5226 13232
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 5092 12442 5120 13126
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 5080 11620 5132 11626
rect 5080 11562 5132 11568
rect 5092 11354 5120 11562
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 4908 9382 4936 9862
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4804 876 4856 882
rect 4804 818 4856 824
rect 3422 82 3478 480
rect 3160 54 3478 82
rect 478 0 534 54
rect 1398 0 1454 54
rect 2410 0 2466 54
rect 3422 0 3478 54
rect 4434 82 4490 480
rect 4908 82 4936 9318
rect 5184 9042 5212 13223
rect 5276 12306 5304 13466
rect 5460 13394 5488 14010
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5368 12986 5396 13262
rect 5460 12986 5488 13330
rect 5552 13326 5580 13806
rect 6196 13530 6224 14418
rect 6472 13870 6500 14436
rect 6552 14418 6604 14424
rect 6552 14340 6604 14346
rect 6552 14282 6604 14288
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 5368 12374 5396 12650
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 5276 11218 5304 12242
rect 5368 11898 5396 12310
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5368 11286 5396 11834
rect 5460 11762 5488 12582
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5356 11280 5408 11286
rect 5356 11222 5408 11228
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5368 10538 5396 10950
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5276 9994 5304 10474
rect 5354 10160 5410 10169
rect 5354 10095 5410 10104
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5184 8634 5212 8978
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5184 8362 5212 8570
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5172 2916 5224 2922
rect 5172 2858 5224 2864
rect 5184 2689 5212 2858
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 5170 2680 5226 2689
rect 5170 2615 5226 2624
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 5184 1601 5212 2246
rect 5276 1970 5304 2790
rect 5264 1964 5316 1970
rect 5264 1906 5316 1912
rect 5170 1592 5226 1601
rect 5170 1527 5226 1536
rect 4434 54 4936 82
rect 5368 82 5396 10095
rect 5552 10062 5580 11698
rect 5632 11620 5684 11626
rect 5632 11562 5684 11568
rect 5644 11354 5672 11562
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 6012 10198 6040 10474
rect 6000 10192 6052 10198
rect 6000 10134 6052 10140
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5552 9654 5580 9998
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6012 9654 6040 10134
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 5908 9444 5960 9450
rect 5908 9386 5960 9392
rect 5920 9110 5948 9386
rect 5908 9104 5960 9110
rect 5908 9046 5960 9052
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5552 8294 5580 8910
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5460 2854 5488 3538
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5552 2650 5580 8230
rect 6012 7954 6040 8842
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6012 7546 6040 7890
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6104 6225 6132 13466
rect 6564 12782 6592 14282
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6184 11280 6236 11286
rect 6184 11222 6236 11228
rect 6196 10810 6224 11222
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 6288 9722 6316 10134
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6380 8974 6408 9590
rect 6552 9104 6604 9110
rect 6552 9046 6604 9052
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6182 8528 6238 8537
rect 6182 8463 6238 8472
rect 6196 8430 6224 8463
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6196 7342 6224 8366
rect 6472 8090 6500 8910
rect 6564 8634 6592 9046
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6656 8514 6684 18958
rect 7104 18964 7156 18970
rect 7104 18906 7156 18912
rect 7116 18222 7144 18906
rect 7208 18222 7236 19110
rect 7484 18902 7512 19264
rect 7472 18896 7524 18902
rect 7472 18838 7524 18844
rect 7576 18630 7604 19314
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 7196 18216 7248 18222
rect 7196 18158 7248 18164
rect 7208 17882 7236 18158
rect 7196 17876 7248 17882
rect 7196 17818 7248 17824
rect 7472 17808 7524 17814
rect 7472 17750 7524 17756
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6840 17134 6868 17478
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 6840 16658 6868 17070
rect 7300 16726 7328 17070
rect 7484 16998 7512 17750
rect 7668 17134 7696 19654
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 7760 18970 7788 19246
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 7852 18290 7880 19110
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7288 16720 7340 16726
rect 7288 16662 7340 16668
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 7196 16584 7248 16590
rect 7196 16526 7248 16532
rect 7104 15972 7156 15978
rect 7104 15914 7156 15920
rect 7116 15609 7144 15914
rect 7102 15600 7158 15609
rect 7102 15535 7158 15544
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6748 14822 6776 14962
rect 7116 14958 7144 15535
rect 7104 14952 7156 14958
rect 7024 14912 7104 14940
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6748 14074 6776 14758
rect 7024 14618 7052 14912
rect 7104 14894 7156 14900
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6840 13802 6868 14554
rect 7024 13870 7052 14554
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 6828 13796 6880 13802
rect 6828 13738 6880 13744
rect 6840 13394 6868 13738
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6748 11354 6776 11630
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6748 10198 6776 11290
rect 6932 11218 6960 13670
rect 7024 13394 7052 13806
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 7024 12442 7052 12650
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 7116 11218 7144 14758
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 6932 10810 6960 11154
rect 7116 10810 7144 11154
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 6826 10704 6882 10713
rect 6826 10639 6882 10648
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 6840 8514 6868 10639
rect 6564 8486 6684 8514
rect 6748 8486 6868 8514
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6368 6724 6420 6730
rect 6368 6666 6420 6672
rect 6090 6216 6146 6225
rect 6090 6151 6146 6160
rect 6380 5778 6408 6666
rect 6472 5778 6500 8026
rect 6368 5772 6420 5778
rect 6368 5714 6420 5720
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6380 5370 6408 5714
rect 6472 5370 6500 5714
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5814 3496 5870 3505
rect 5724 3460 5776 3466
rect 5776 3440 5814 3448
rect 5776 3431 5870 3440
rect 5776 3420 5856 3431
rect 5724 3402 5776 3408
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6012 2990 6040 3674
rect 6274 3632 6330 3641
rect 6274 3567 6276 3576
rect 6328 3567 6330 3576
rect 6564 3584 6592 8486
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6656 6458 6684 6734
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6656 4214 6684 4422
rect 6644 4208 6696 4214
rect 6644 4150 6696 4156
rect 6644 3596 6696 3602
rect 6564 3556 6644 3584
rect 6276 3538 6328 3544
rect 6644 3538 6696 3544
rect 6288 3058 6316 3538
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6000 2984 6052 2990
rect 6052 2944 6132 2972
rect 6000 2926 6052 2932
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5460 2310 5488 2450
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 5460 2106 5488 2246
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5448 2100 5500 2106
rect 5448 2042 5500 2048
rect 6012 2038 6040 2790
rect 6104 2310 6132 2944
rect 6656 2854 6684 3538
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 6000 2032 6052 2038
rect 6656 2009 6684 2790
rect 6000 1974 6052 1980
rect 6642 2000 6698 2009
rect 6642 1935 6698 1944
rect 5446 82 5502 480
rect 5368 54 5502 82
rect 4434 0 4490 54
rect 5446 0 5502 54
rect 6458 82 6514 480
rect 6748 82 6776 8486
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6840 4690 6868 8366
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6840 3942 6868 4626
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6840 1329 6868 3878
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6932 3040 6960 3334
rect 7012 3052 7064 3058
rect 6932 3012 7012 3040
rect 7012 2994 7064 3000
rect 7102 2816 7158 2825
rect 7102 2751 7158 2760
rect 7116 2650 7144 2751
rect 7208 2650 7236 16526
rect 7300 16454 7328 16662
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7300 15706 7328 16390
rect 7484 15978 7512 16934
rect 7668 16658 7696 17070
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7564 16176 7616 16182
rect 7668 16164 7696 16594
rect 7616 16136 7696 16164
rect 7564 16118 7616 16124
rect 7472 15972 7524 15978
rect 7472 15914 7524 15920
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 7300 14958 7328 15642
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 7300 14482 7328 14894
rect 7484 14890 7512 15914
rect 7472 14884 7524 14890
rect 7472 14826 7524 14832
rect 7944 14550 7972 22918
rect 8128 22778 8156 23190
rect 8116 22772 8168 22778
rect 8116 22714 8168 22720
rect 8024 22500 8076 22506
rect 8024 22442 8076 22448
rect 8036 22166 8064 22442
rect 8128 22234 8156 22714
rect 8116 22228 8168 22234
rect 8116 22170 8168 22176
rect 8024 22160 8076 22166
rect 8024 22102 8076 22108
rect 8036 21418 8064 22102
rect 8496 21554 8524 27526
rect 9126 27520 9182 28000
rect 9954 27554 10010 28000
rect 9692 27526 10010 27554
rect 9140 25362 9168 27520
rect 9128 25356 9180 25362
rect 9128 25298 9180 25304
rect 8576 24744 8628 24750
rect 8852 24744 8904 24750
rect 8576 24686 8628 24692
rect 8772 24704 8852 24732
rect 8588 23254 8616 24686
rect 8576 23248 8628 23254
rect 8576 23190 8628 23196
rect 8576 22976 8628 22982
rect 8576 22918 8628 22924
rect 8588 21690 8616 22918
rect 8576 21684 8628 21690
rect 8576 21626 8628 21632
rect 8484 21548 8536 21554
rect 8484 21490 8536 21496
rect 8024 21412 8076 21418
rect 8024 21354 8076 21360
rect 8484 20936 8536 20942
rect 8484 20878 8536 20884
rect 8208 20392 8260 20398
rect 8208 20334 8260 20340
rect 8220 19718 8248 20334
rect 8208 19712 8260 19718
rect 8208 19654 8260 19660
rect 8114 18864 8170 18873
rect 8114 18799 8170 18808
rect 8208 18828 8260 18834
rect 8024 18624 8076 18630
rect 8024 18566 8076 18572
rect 8036 17785 8064 18566
rect 8022 17776 8078 17785
rect 8022 17711 8078 17720
rect 8128 17728 8156 18799
rect 8208 18770 8260 18776
rect 8220 18426 8248 18770
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 8496 18358 8524 20878
rect 8576 19916 8628 19922
rect 8576 19858 8628 19864
rect 8588 19174 8616 19858
rect 8668 19712 8720 19718
rect 8668 19654 8720 19660
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8484 18352 8536 18358
rect 8484 18294 8536 18300
rect 8208 17740 8260 17746
rect 8128 17700 8208 17728
rect 8128 16658 8156 17700
rect 8208 17682 8260 17688
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 8206 17232 8262 17241
rect 8206 17167 8262 17176
rect 8220 17134 8248 17167
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 8312 17066 8340 17614
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 8312 16794 8340 17002
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8024 16516 8076 16522
rect 8024 16458 8076 16464
rect 8036 16114 8064 16458
rect 8024 16108 8076 16114
rect 8024 16050 8076 16056
rect 8036 15706 8064 16050
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 8128 14958 8156 16594
rect 8390 16552 8446 16561
rect 8390 16487 8446 16496
rect 8404 16454 8432 16487
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8680 15570 8708 19654
rect 8772 15638 8800 24704
rect 8852 24686 8904 24692
rect 9692 23866 9720 27526
rect 9954 27520 10010 27526
rect 10690 27520 10746 28000
rect 11518 27554 11574 28000
rect 11518 27526 11836 27554
rect 11518 27520 11574 27526
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10140 25288 10192 25294
rect 10140 25230 10192 25236
rect 10048 24200 10100 24206
rect 10048 24142 10100 24148
rect 10060 23866 10088 24142
rect 9680 23860 9732 23866
rect 9680 23802 9732 23808
rect 10048 23860 10100 23866
rect 10048 23802 10100 23808
rect 9692 23662 9720 23802
rect 9772 23792 9824 23798
rect 9772 23734 9824 23740
rect 9680 23656 9732 23662
rect 9680 23598 9732 23604
rect 9404 23520 9456 23526
rect 9784 23474 9812 23734
rect 10060 23526 10088 23802
rect 10152 23798 10180 25230
rect 10704 24886 10732 27520
rect 11704 25356 11756 25362
rect 11704 25298 11756 25304
rect 11716 24954 11744 25298
rect 11704 24948 11756 24954
rect 11704 24890 11756 24896
rect 10692 24880 10744 24886
rect 10692 24822 10744 24828
rect 11808 24750 11836 27526
rect 12346 27520 12402 28000
rect 13082 27520 13138 28000
rect 13910 27520 13966 28000
rect 14738 27520 14794 28000
rect 15566 27554 15622 28000
rect 16302 27554 16358 28000
rect 15488 27526 15622 27554
rect 11796 24744 11848 24750
rect 10690 24712 10746 24721
rect 11796 24686 11848 24692
rect 10690 24647 10746 24656
rect 11980 24676 12032 24682
rect 10704 24614 10732 24647
rect 11980 24618 12032 24624
rect 10692 24608 10744 24614
rect 10692 24550 10744 24556
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10600 24336 10652 24342
rect 10600 24278 10652 24284
rect 10232 24064 10284 24070
rect 10232 24006 10284 24012
rect 10140 23792 10192 23798
rect 10140 23734 10192 23740
rect 10244 23644 10272 24006
rect 10612 23712 10640 24278
rect 10692 24268 10744 24274
rect 10692 24210 10744 24216
rect 11704 24268 11756 24274
rect 11704 24210 11756 24216
rect 10704 23866 10732 24210
rect 11716 23866 11744 24210
rect 10692 23860 10744 23866
rect 11704 23860 11756 23866
rect 10744 23820 10824 23848
rect 10692 23802 10744 23808
rect 10692 23724 10744 23730
rect 10612 23684 10692 23712
rect 10692 23666 10744 23672
rect 10152 23616 10272 23644
rect 9404 23462 9456 23468
rect 9312 22568 9364 22574
rect 9312 22510 9364 22516
rect 8942 21992 8998 22001
rect 9324 21962 9352 22510
rect 8942 21927 8998 21936
rect 9312 21956 9364 21962
rect 8852 18420 8904 18426
rect 8852 18362 8904 18368
rect 8864 18154 8892 18362
rect 8852 18148 8904 18154
rect 8852 18090 8904 18096
rect 8864 17882 8892 18090
rect 8852 17876 8904 17882
rect 8852 17818 8904 17824
rect 8760 15632 8812 15638
rect 8760 15574 8812 15580
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8668 15564 8720 15570
rect 8668 15506 8720 15512
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 8312 14822 8340 15506
rect 8680 15162 8708 15506
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 7932 14544 7984 14550
rect 7932 14486 7984 14492
rect 7288 14476 7340 14482
rect 7288 14418 7340 14424
rect 7300 13870 7328 14418
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7300 13530 7328 13806
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7852 12442 7880 12582
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 7852 11558 7880 12378
rect 7944 12306 7972 13466
rect 8312 13462 8340 14758
rect 8760 14544 8812 14550
rect 8760 14486 8812 14492
rect 8772 13734 8800 14486
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8852 13728 8904 13734
rect 8852 13670 8904 13676
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 8024 13388 8076 13394
rect 8024 13330 8076 13336
rect 8392 13388 8444 13394
rect 8392 13330 8444 13336
rect 8036 12986 8064 13330
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 8022 12744 8078 12753
rect 8022 12679 8078 12688
rect 7932 12300 7984 12306
rect 7932 12242 7984 12248
rect 7944 11898 7972 12242
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 8036 11830 8064 12679
rect 8404 12102 8432 13330
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8496 12442 8524 12718
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8772 12306 8800 13670
rect 8864 13258 8892 13670
rect 8852 13252 8904 13258
rect 8852 13194 8904 13200
rect 8864 12782 8892 13194
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8024 11824 8076 11830
rect 8024 11766 8076 11772
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7852 11354 7880 11494
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 7852 10742 7880 11290
rect 7840 10736 7892 10742
rect 7892 10696 7972 10724
rect 7840 10678 7892 10684
rect 7748 10532 7800 10538
rect 7748 10474 7800 10480
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7576 9178 7604 9998
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7576 8566 7604 9114
rect 7760 8634 7788 10474
rect 7852 10198 7880 10474
rect 7840 10192 7892 10198
rect 7840 10134 7892 10140
rect 7944 8634 7972 10696
rect 8036 9654 8064 11766
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8220 10198 8248 11290
rect 8312 10742 8340 11698
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8220 9722 8248 10134
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 8772 9450 8800 12242
rect 8852 11620 8904 11626
rect 8852 11562 8904 11568
rect 8864 11354 8892 11562
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8956 10282 8984 21927
rect 9312 21898 9364 21904
rect 9128 21344 9180 21350
rect 9128 21286 9180 21292
rect 9140 21078 9168 21286
rect 9128 21072 9180 21078
rect 9128 21014 9180 21020
rect 9220 21072 9272 21078
rect 9220 21014 9272 21020
rect 9036 21004 9088 21010
rect 9036 20946 9088 20952
rect 9048 20806 9076 20946
rect 9036 20800 9088 20806
rect 9036 20742 9088 20748
rect 9048 20466 9076 20742
rect 9036 20460 9088 20466
rect 9036 20402 9088 20408
rect 9048 20058 9076 20402
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 9140 19990 9168 21014
rect 9128 19984 9180 19990
rect 9128 19926 9180 19932
rect 9140 19718 9168 19926
rect 9232 19854 9260 21014
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 9128 19712 9180 19718
rect 9128 19654 9180 19660
rect 9036 18692 9088 18698
rect 9036 18634 9088 18640
rect 9048 18154 9076 18634
rect 9128 18624 9180 18630
rect 9128 18566 9180 18572
rect 9140 18290 9168 18566
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 9036 18148 9088 18154
rect 9036 18090 9088 18096
rect 9232 17184 9260 19790
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9324 17746 9352 18702
rect 9312 17740 9364 17746
rect 9312 17682 9364 17688
rect 9140 17156 9260 17184
rect 9416 17184 9444 23462
rect 9692 23446 9812 23474
rect 10048 23520 10100 23526
rect 10048 23462 10100 23468
rect 9692 23322 9720 23446
rect 9680 23316 9732 23322
rect 9680 23258 9732 23264
rect 10152 22624 10180 23616
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10704 23118 10732 23666
rect 10796 23254 10824 23820
rect 11704 23802 11756 23808
rect 10784 23248 10836 23254
rect 10784 23190 10836 23196
rect 11520 23248 11572 23254
rect 11520 23190 11572 23196
rect 10416 23112 10468 23118
rect 10416 23054 10468 23060
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10428 22642 10456 23054
rect 10796 22778 10824 23190
rect 11532 22778 11560 23190
rect 10784 22772 10836 22778
rect 10784 22714 10836 22720
rect 11520 22772 11572 22778
rect 11520 22714 11572 22720
rect 10060 22596 10180 22624
rect 10416 22636 10468 22642
rect 9956 22228 10008 22234
rect 9956 22170 10008 22176
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9784 21486 9812 21830
rect 9968 21622 9996 22170
rect 9956 21616 10008 21622
rect 9956 21558 10008 21564
rect 9496 21480 9548 21486
rect 9496 21422 9548 21428
rect 9772 21480 9824 21486
rect 9772 21422 9824 21428
rect 9508 19990 9536 21422
rect 9784 21146 9812 21422
rect 9968 21350 9996 21558
rect 9956 21344 10008 21350
rect 9956 21286 10008 21292
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9864 20256 9916 20262
rect 9864 20198 9916 20204
rect 9496 19984 9548 19990
rect 9496 19926 9548 19932
rect 9876 19922 9904 20198
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 9784 19281 9812 19654
rect 9876 19514 9904 19858
rect 9956 19780 10008 19786
rect 9956 19722 10008 19728
rect 9864 19508 9916 19514
rect 9864 19450 9916 19456
rect 9968 19378 9996 19722
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 9770 19272 9826 19281
rect 9770 19207 9826 19216
rect 9864 19236 9916 19242
rect 9784 18834 9812 19207
rect 9864 19178 9916 19184
rect 9772 18828 9824 18834
rect 9772 18770 9824 18776
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9508 17882 9536 18702
rect 9784 17882 9812 18770
rect 9876 18698 9904 19178
rect 9968 18834 9996 19314
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9968 18630 9996 18770
rect 9956 18624 10008 18630
rect 9956 18566 10008 18572
rect 10060 18408 10088 22596
rect 10416 22578 10468 22584
rect 10140 22500 10192 22506
rect 10140 22442 10192 22448
rect 10152 22234 10180 22442
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10140 22228 10192 22234
rect 10140 22170 10192 22176
rect 10796 21690 10824 22714
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 11152 22024 11204 22030
rect 11152 21966 11204 21972
rect 10784 21684 10836 21690
rect 10784 21626 10836 21632
rect 11164 21350 11192 21966
rect 11256 21418 11284 22034
rect 11532 21962 11560 22714
rect 11520 21956 11572 21962
rect 11520 21898 11572 21904
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 11244 21412 11296 21418
rect 11244 21354 11296 21360
rect 11152 21344 11204 21350
rect 11152 21286 11204 21292
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10324 21004 10376 21010
rect 10508 21004 10560 21010
rect 10376 20964 10456 20992
rect 10324 20946 10376 20952
rect 10428 20602 10456 20964
rect 10508 20946 10560 20952
rect 10784 21004 10836 21010
rect 10784 20946 10836 20952
rect 10416 20596 10468 20602
rect 10416 20538 10468 20544
rect 10428 20398 10456 20538
rect 10520 20534 10548 20946
rect 10508 20528 10560 20534
rect 10508 20470 10560 20476
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10140 19916 10192 19922
rect 10140 19858 10192 19864
rect 10152 19174 10180 19858
rect 10692 19848 10744 19854
rect 10692 19790 10744 19796
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10152 18834 10180 19110
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10416 18896 10468 18902
rect 10416 18838 10468 18844
rect 10140 18828 10192 18834
rect 10140 18770 10192 18776
rect 10152 18426 10180 18770
rect 9968 18380 10088 18408
rect 10140 18420 10192 18426
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9416 17156 9536 17184
rect 9140 15910 9168 17156
rect 9220 17060 9272 17066
rect 9220 17002 9272 17008
rect 9404 17060 9456 17066
rect 9404 17002 9456 17008
rect 9232 16590 9260 17002
rect 9220 16584 9272 16590
rect 9220 16526 9272 16532
rect 9416 16114 9444 17002
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9128 15904 9180 15910
rect 9128 15846 9180 15852
rect 9508 15502 9536 17156
rect 9864 16720 9916 16726
rect 9864 16662 9916 16668
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9784 16250 9812 16526
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9876 16046 9904 16662
rect 9864 16040 9916 16046
rect 9864 15982 9916 15988
rect 9968 15706 9996 18380
rect 10140 18362 10192 18368
rect 10324 18352 10376 18358
rect 10324 18294 10376 18300
rect 10048 18284 10100 18290
rect 10048 18226 10100 18232
rect 10060 17066 10088 18226
rect 10336 18154 10364 18294
rect 10428 18154 10456 18838
rect 10324 18148 10376 18154
rect 10324 18090 10376 18096
rect 10416 18148 10468 18154
rect 10416 18090 10468 18096
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 10152 17338 10180 17682
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10048 17060 10100 17066
rect 10048 17002 10100 17008
rect 10060 16590 10088 17002
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9588 15632 9640 15638
rect 9588 15574 9640 15580
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9496 15496 9548 15502
rect 9496 15438 9548 15444
rect 9036 15156 9088 15162
rect 9036 15098 9088 15104
rect 9048 13025 9076 15098
rect 9416 14618 9444 15438
rect 9508 15162 9536 15438
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9600 14822 9628 15574
rect 9968 15026 9996 15642
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 10520 14890 10548 15438
rect 10704 14958 10732 19790
rect 10796 19514 10824 20946
rect 11164 20466 11192 21286
rect 11152 20460 11204 20466
rect 11152 20402 11204 20408
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10980 19718 11008 20334
rect 10968 19712 11020 19718
rect 10968 19654 11020 19660
rect 10784 19508 10836 19514
rect 10784 19450 10836 19456
rect 10796 19417 10824 19450
rect 10876 19440 10928 19446
rect 10782 19408 10838 19417
rect 10876 19382 10928 19388
rect 10782 19343 10838 19352
rect 10888 18970 10916 19382
rect 10980 19310 11008 19654
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 10796 17134 10824 17478
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10796 16522 10824 17070
rect 10784 16516 10836 16522
rect 10784 16458 10836 16464
rect 10784 15428 10836 15434
rect 10784 15370 10836 15376
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10508 14884 10560 14890
rect 10508 14826 10560 14832
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9600 14006 9628 14758
rect 9220 14000 9272 14006
rect 9220 13942 9272 13948
rect 9588 14000 9640 14006
rect 9588 13942 9640 13948
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9140 13530 9168 13806
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9034 13016 9090 13025
rect 9034 12951 9090 12960
rect 9232 11626 9260 13942
rect 9692 13814 9720 14758
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10416 14544 10468 14550
rect 10416 14486 10468 14492
rect 10428 14074 10456 14486
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 9312 13796 9364 13802
rect 9312 13738 9364 13744
rect 9600 13786 9720 13814
rect 9324 13705 9352 13738
rect 9310 13696 9366 13705
rect 9310 13631 9366 13640
rect 9600 12986 9628 13786
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9140 11014 9168 11494
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 8956 10254 9076 10282
rect 9140 10266 9168 10950
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 8944 10192 8996 10198
rect 8944 10134 8996 10140
rect 8956 9654 8984 10134
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 8208 9444 8260 9450
rect 8208 9386 8260 9392
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8220 9178 8248 9386
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7564 8560 7616 8566
rect 7564 8502 7616 8508
rect 7944 8362 7972 8570
rect 8128 8498 8156 9114
rect 8404 8838 8432 9386
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 7944 8022 7972 8298
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7300 7546 7328 7686
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7484 7206 7512 7890
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7484 6866 7512 7142
rect 7576 7002 7604 7890
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7760 7274 7788 7686
rect 7748 7268 7800 7274
rect 7748 7210 7800 7216
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7484 6118 7512 6802
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7484 5273 7512 6054
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7470 5264 7526 5273
rect 7470 5199 7526 5208
rect 7576 4146 7604 5510
rect 7656 5296 7708 5302
rect 7656 5238 7708 5244
rect 7668 4826 7696 5238
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7576 4010 7604 4082
rect 7564 4004 7616 4010
rect 7564 3946 7616 3952
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 7576 3738 7604 3946
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7668 3058 7696 3946
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7760 2582 7788 7210
rect 7944 7002 7972 7958
rect 8128 7886 8156 8434
rect 8404 8090 8432 8774
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8760 7268 8812 7274
rect 8760 7210 8812 7216
rect 7932 6996 7984 7002
rect 7932 6938 7984 6944
rect 7944 5846 7972 6938
rect 8772 6934 8800 7210
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 8128 6390 8156 6870
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 7944 5370 7972 5782
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7852 5137 7880 5170
rect 7838 5128 7894 5137
rect 7838 5063 7894 5072
rect 8036 4826 8064 5646
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 8128 3670 8156 6326
rect 8772 6322 8800 6870
rect 9048 6610 9076 10254
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9416 10198 9444 10610
rect 9600 10538 9628 12922
rect 9876 12918 9904 13330
rect 9968 13258 9996 14010
rect 10796 13814 10824 15370
rect 10980 14074 11008 19246
rect 11072 18630 11100 19246
rect 11256 18834 11284 21354
rect 11520 21344 11572 21350
rect 11520 21286 11572 21292
rect 11532 21010 11560 21286
rect 11520 21004 11572 21010
rect 11520 20946 11572 20952
rect 11612 20936 11664 20942
rect 11612 20878 11664 20884
rect 11336 20392 11388 20398
rect 11336 20334 11388 20340
rect 11348 19281 11376 20334
rect 11428 19712 11480 19718
rect 11428 19654 11480 19660
rect 11440 19446 11468 19654
rect 11428 19440 11480 19446
rect 11428 19382 11480 19388
rect 11334 19272 11390 19281
rect 11334 19207 11390 19216
rect 11348 18834 11376 19207
rect 11624 18834 11652 20878
rect 11716 20874 11744 21830
rect 11796 21480 11848 21486
rect 11796 21422 11848 21428
rect 11704 20868 11756 20874
rect 11704 20810 11756 20816
rect 11808 20058 11836 21422
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11796 19916 11848 19922
rect 11796 19858 11848 19864
rect 11808 19514 11836 19858
rect 11796 19508 11848 19514
rect 11796 19450 11848 19456
rect 11244 18828 11296 18834
rect 11244 18770 11296 18776
rect 11336 18828 11388 18834
rect 11612 18828 11664 18834
rect 11388 18788 11468 18816
rect 11336 18770 11388 18776
rect 11336 18692 11388 18698
rect 11336 18634 11388 18640
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 11072 18465 11100 18566
rect 11058 18456 11114 18465
rect 11348 18426 11376 18634
rect 11440 18426 11468 18788
rect 11612 18770 11664 18776
rect 11058 18391 11114 18400
rect 11336 18420 11388 18426
rect 11336 18362 11388 18368
rect 11428 18420 11480 18426
rect 11428 18362 11480 18368
rect 11624 18154 11652 18770
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11612 18148 11664 18154
rect 11612 18090 11664 18096
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 11532 17746 11560 18022
rect 11624 17882 11652 18090
rect 11612 17876 11664 17882
rect 11612 17818 11664 17824
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11060 17060 11112 17066
rect 11060 17002 11112 17008
rect 11072 16726 11100 17002
rect 11716 16998 11744 17682
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10796 13786 10916 13814
rect 10980 13802 11008 14010
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 10152 12986 10180 13330
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 9588 10532 9640 10538
rect 9588 10474 9640 10480
rect 9600 10266 9628 10474
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9404 10192 9456 10198
rect 9404 10134 9456 10140
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9784 9178 9812 9998
rect 9876 9450 9904 10134
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9508 8362 9536 8978
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 8956 6582 9076 6610
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 8220 5574 8248 6122
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8312 4214 8340 4558
rect 8772 4282 8800 4626
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 8864 4146 8892 4422
rect 8956 4214 8984 6582
rect 9140 6390 9168 8230
rect 9508 8090 9536 8298
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9508 7410 9536 8026
rect 9968 7954 9996 12786
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 10060 11762 10088 12174
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10060 10062 10088 11698
rect 10152 11354 10180 11698
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 10140 9920 10192 9926
rect 10140 9862 10192 9868
rect 10152 9382 10180 9862
rect 10704 9722 10732 13330
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10796 11898 10824 12310
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10784 11620 10836 11626
rect 10784 11562 10836 11568
rect 10796 11354 10824 11562
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10796 10810 10824 11290
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10704 9518 10732 9658
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10152 9042 10180 9318
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10704 9092 10732 9454
rect 10612 9064 10732 9092
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 10060 8022 10088 8230
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 9956 7948 10008 7954
rect 10152 7936 10180 8978
rect 10612 8498 10640 9064
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 7954 10732 8910
rect 10324 7948 10376 7954
rect 10152 7908 10324 7936
rect 9956 7890 10008 7896
rect 10324 7890 10376 7896
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 9968 7478 9996 7890
rect 10336 7818 10364 7890
rect 10324 7812 10376 7818
rect 10324 7754 10376 7760
rect 10336 7546 10364 7754
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9508 6458 9536 6938
rect 9692 6866 9720 7142
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9128 6384 9180 6390
rect 9128 6326 9180 6332
rect 9784 6186 9812 6394
rect 9772 6180 9824 6186
rect 9772 6122 9824 6128
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9140 5234 9168 5714
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9232 5166 9260 5646
rect 9876 5370 9904 5782
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9036 5092 9088 5098
rect 9036 5034 9088 5040
rect 9048 4690 9076 5034
rect 9036 4684 9088 4690
rect 9036 4626 9088 4632
rect 8944 4208 8996 4214
rect 8944 4150 8996 4156
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8864 3942 8892 4082
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8772 3670 8800 3878
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 8128 3194 8156 3606
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 7944 2446 7972 3062
rect 8128 2854 8156 3130
rect 8392 3120 8444 3126
rect 8392 3062 8444 3068
rect 8404 2990 8432 3062
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8588 2922 8616 3334
rect 8576 2916 8628 2922
rect 8576 2858 8628 2864
rect 8116 2848 8168 2854
rect 8588 2825 8616 2858
rect 8760 2848 8812 2854
rect 8116 2790 8168 2796
rect 8574 2816 8630 2825
rect 8574 2751 8630 2760
rect 8680 2808 8760 2836
rect 8680 2582 8708 2808
rect 8760 2790 8812 2796
rect 8864 2582 8892 3470
rect 8956 2961 8984 4150
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 9048 4010 9076 4082
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 9048 3738 9076 3946
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9232 3058 9260 5102
rect 9772 5092 9824 5098
rect 9772 5034 9824 5040
rect 9784 4758 9812 5034
rect 9876 4826 9904 5306
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9324 4146 9352 4422
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9324 3534 9352 4082
rect 9692 3738 9720 4626
rect 9968 4622 9996 7414
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10612 6458 10640 6598
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10152 5710 10180 6258
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10888 5302 10916 13786
rect 10968 13796 11020 13802
rect 10968 13738 11020 13744
rect 11072 12646 11100 16050
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 11072 12102 11100 12582
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 11072 9722 11100 12038
rect 11060 9716 11112 9722
rect 11060 9658 11112 9664
rect 11072 9110 11100 9658
rect 11060 9104 11112 9110
rect 11060 9046 11112 9052
rect 11072 8634 11100 9046
rect 11164 8906 11192 16934
rect 11716 16658 11744 16934
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11520 15972 11572 15978
rect 11520 15914 11572 15920
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11256 12850 11284 15642
rect 11532 14958 11560 15914
rect 11716 15910 11744 16594
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11520 14952 11572 14958
rect 11520 14894 11572 14900
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11336 14544 11388 14550
rect 11336 14486 11388 14492
rect 11348 13802 11376 14486
rect 11532 14006 11560 14758
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11520 14000 11572 14006
rect 11520 13942 11572 13948
rect 11336 13796 11388 13802
rect 11336 13738 11388 13744
rect 11336 13456 11388 13462
rect 11336 13398 11388 13404
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11348 12782 11376 13398
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11428 12368 11480 12374
rect 11428 12310 11480 12316
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11256 10470 11284 11086
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11348 10810 11376 10950
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11348 10538 11376 10746
rect 11440 10742 11468 12310
rect 11428 10736 11480 10742
rect 11428 10678 11480 10684
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11256 10266 11284 10406
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11532 10130 11560 13942
rect 11624 13530 11652 14554
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11716 13394 11744 15846
rect 11808 15570 11836 18702
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11900 16250 11928 17138
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 11900 16046 11928 16186
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11808 15162 11836 15506
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11624 10674 11652 10950
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11532 9654 11560 10066
rect 11716 10062 11744 12854
rect 11808 12374 11836 14350
rect 11900 14074 11928 15982
rect 11992 15502 12020 24618
rect 12256 24608 12308 24614
rect 12256 24550 12308 24556
rect 12268 23474 12296 24550
rect 12360 24274 12388 27520
rect 12348 24268 12400 24274
rect 12348 24210 12400 24216
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 12176 23446 12296 23474
rect 12072 23044 12124 23050
rect 12072 22986 12124 22992
rect 12084 22166 12112 22986
rect 12176 22234 12204 23446
rect 12256 23112 12308 23118
rect 12256 23054 12308 23060
rect 12268 22642 12296 23054
rect 12360 22778 12388 23598
rect 12716 23520 12768 23526
rect 12716 23462 12768 23468
rect 12992 23520 13044 23526
rect 12992 23462 13044 23468
rect 12624 23316 12676 23322
rect 12624 23258 12676 23264
rect 12348 22772 12400 22778
rect 12348 22714 12400 22720
rect 12256 22636 12308 22642
rect 12256 22578 12308 22584
rect 12636 22574 12664 23258
rect 12728 22692 12756 23462
rect 12900 23112 12952 23118
rect 12900 23054 12952 23060
rect 12808 22704 12860 22710
rect 12728 22664 12808 22692
rect 12624 22568 12676 22574
rect 12624 22510 12676 22516
rect 12164 22228 12216 22234
rect 12164 22170 12216 22176
rect 12072 22160 12124 22166
rect 12072 22102 12124 22108
rect 12636 22098 12664 22510
rect 12728 22098 12756 22664
rect 12808 22646 12860 22652
rect 12912 22574 12940 23054
rect 13004 22982 13032 23462
rect 12992 22976 13044 22982
rect 12992 22918 13044 22924
rect 12900 22568 12952 22574
rect 12900 22510 12952 22516
rect 12912 22098 12940 22510
rect 13096 22098 13124 27520
rect 13360 25356 13412 25362
rect 13360 25298 13412 25304
rect 13176 25152 13228 25158
rect 13176 25094 13228 25100
rect 12624 22092 12676 22098
rect 12624 22034 12676 22040
rect 12716 22092 12768 22098
rect 12716 22034 12768 22040
rect 12900 22092 12952 22098
rect 12900 22034 12952 22040
rect 13084 22092 13136 22098
rect 13084 22034 13136 22040
rect 12636 21622 12664 22034
rect 12624 21616 12676 21622
rect 12624 21558 12676 21564
rect 12728 21078 12756 22034
rect 12912 21146 12940 22034
rect 12900 21140 12952 21146
rect 12900 21082 12952 21088
rect 12716 21072 12768 21078
rect 12716 21014 12768 21020
rect 12072 21004 12124 21010
rect 12072 20946 12124 20952
rect 12084 20262 12112 20946
rect 12072 20256 12124 20262
rect 12072 20198 12124 20204
rect 12084 19990 12112 20198
rect 12440 20052 12492 20058
rect 12440 19994 12492 20000
rect 12072 19984 12124 19990
rect 12072 19926 12124 19932
rect 12084 19310 12112 19926
rect 12452 19310 12480 19994
rect 12532 19780 12584 19786
rect 12532 19722 12584 19728
rect 12544 19310 12572 19722
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12256 19236 12308 19242
rect 12256 19178 12308 19184
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 12268 15434 12296 19178
rect 12544 18698 12572 19246
rect 12532 18692 12584 18698
rect 12532 18634 12584 18640
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12636 17921 12664 18158
rect 12900 18148 12952 18154
rect 12900 18090 12952 18096
rect 12622 17912 12678 17921
rect 12622 17847 12678 17856
rect 12532 17128 12584 17134
rect 12636 17116 12664 17847
rect 12716 17808 12768 17814
rect 12716 17750 12768 17756
rect 12584 17088 12664 17116
rect 12532 17070 12584 17076
rect 12440 17060 12492 17066
rect 12440 17002 12492 17008
rect 12452 16658 12480 17002
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12256 15428 12308 15434
rect 12256 15370 12308 15376
rect 12360 15366 12388 16594
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12348 15360 12400 15366
rect 12348 15302 12400 15308
rect 12360 15094 12388 15302
rect 12348 15088 12400 15094
rect 12348 15030 12400 15036
rect 11980 14884 12032 14890
rect 11980 14826 12032 14832
rect 11992 14346 12020 14826
rect 12360 14822 12388 15030
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 11980 14340 12032 14346
rect 11980 14282 12032 14288
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11900 13870 11928 14010
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11900 12374 11928 13806
rect 11992 13530 12020 14282
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 12360 13462 12388 14758
rect 12636 14618 12664 16526
rect 12728 16250 12756 17750
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 12820 16658 12848 17614
rect 12912 17134 12940 18090
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 12900 17128 12952 17134
rect 12900 17070 12952 17076
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12716 15632 12768 15638
rect 12716 15574 12768 15580
rect 12728 15162 12756 15574
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 13004 14618 13032 15438
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12992 14612 13044 14618
rect 12992 14554 13044 14560
rect 12636 13938 12664 14554
rect 13096 14006 13124 17274
rect 13188 14618 13216 25094
rect 13372 24886 13400 25298
rect 13544 25152 13596 25158
rect 13544 25094 13596 25100
rect 13360 24880 13412 24886
rect 13360 24822 13412 24828
rect 13452 22636 13504 22642
rect 13452 22578 13504 22584
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13372 21622 13400 21966
rect 13360 21616 13412 21622
rect 13360 21558 13412 21564
rect 13464 20448 13492 22578
rect 13556 20942 13584 25094
rect 13728 24608 13780 24614
rect 13728 24550 13780 24556
rect 13740 24313 13768 24550
rect 13726 24304 13782 24313
rect 13636 24268 13688 24274
rect 13726 24239 13782 24248
rect 13636 24210 13688 24216
rect 13648 23866 13676 24210
rect 13636 23860 13688 23866
rect 13636 23802 13688 23808
rect 13924 23730 13952 27520
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 14464 24608 14516 24614
rect 14464 24550 14516 24556
rect 13912 23724 13964 23730
rect 13912 23666 13964 23672
rect 13820 22024 13872 22030
rect 13820 21966 13872 21972
rect 13728 21888 13780 21894
rect 13728 21830 13780 21836
rect 13740 21554 13768 21830
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 13832 21418 13860 21966
rect 13820 21412 13872 21418
rect 13820 21354 13872 21360
rect 13544 20936 13596 20942
rect 13544 20878 13596 20884
rect 13556 20602 13584 20878
rect 14004 20800 14056 20806
rect 14004 20742 14056 20748
rect 13544 20596 13596 20602
rect 13544 20538 13596 20544
rect 14016 20505 14044 20742
rect 13372 20420 13492 20448
rect 14002 20496 14058 20505
rect 14002 20431 14058 20440
rect 13268 19916 13320 19922
rect 13268 19858 13320 19864
rect 13280 19514 13308 19858
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13268 18828 13320 18834
rect 13268 18770 13320 18776
rect 13280 17746 13308 18770
rect 13372 17796 13400 20420
rect 13452 20324 13504 20330
rect 13452 20266 13504 20272
rect 13464 20058 13492 20266
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 14004 19916 14056 19922
rect 14004 19858 14056 19864
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 13740 19378 13768 19790
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 14016 19174 14044 19858
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13372 17768 13584 17796
rect 13268 17740 13320 17746
rect 13320 17700 13400 17728
rect 13268 17682 13320 17688
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13280 16046 13308 17478
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 13372 15706 13400 17700
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 13464 15706 13492 16594
rect 13556 15978 13584 17768
rect 13740 17746 13768 18770
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 13924 18290 13952 18702
rect 13912 18284 13964 18290
rect 13912 18226 13964 18232
rect 14004 18080 14056 18086
rect 14004 18022 14056 18028
rect 13636 17740 13688 17746
rect 13636 17682 13688 17688
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 13648 17338 13676 17682
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13740 16794 13768 17138
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13740 16250 13768 16730
rect 13832 16522 13860 17274
rect 14016 17202 14044 18022
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 13912 17128 13964 17134
rect 13912 17070 13964 17076
rect 13924 16522 13952 17070
rect 14004 17060 14056 17066
rect 14004 17002 14056 17008
rect 13820 16516 13872 16522
rect 13820 16458 13872 16464
rect 13912 16516 13964 16522
rect 13912 16458 13964 16464
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13924 16114 13952 16458
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 13372 15552 13400 15642
rect 14016 15570 14044 17002
rect 14004 15564 14056 15570
rect 13372 15524 13492 15552
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13176 14612 13228 14618
rect 13228 14572 13308 14600
rect 13176 14554 13228 14560
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 13096 13814 13124 13942
rect 12532 13796 12584 13802
rect 13096 13786 13216 13814
rect 12532 13738 12584 13744
rect 12544 13530 12572 13738
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12348 13456 12400 13462
rect 12348 13398 12400 13404
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 11796 12368 11848 12374
rect 11796 12310 11848 12316
rect 11888 12368 11940 12374
rect 11888 12310 11940 12316
rect 11900 11898 11928 12310
rect 11992 12306 12020 13262
rect 12176 12850 12204 13262
rect 12544 12986 12572 13466
rect 13188 13462 13216 13786
rect 13280 13530 13308 14572
rect 13372 14074 13400 15098
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13176 13456 13228 13462
rect 13176 13398 13228 13404
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11992 11830 12020 12242
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 12544 11626 12572 12922
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 11888 11620 11940 11626
rect 11888 11562 11940 11568
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 12716 11620 12768 11626
rect 12716 11562 12768 11568
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11520 9648 11572 9654
rect 11520 9590 11572 9596
rect 11520 9444 11572 9450
rect 11520 9386 11572 9392
rect 11532 9042 11560 9386
rect 11716 9178 11744 9998
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11900 9110 11928 11562
rect 12728 11354 12756 11562
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12820 11286 12848 12378
rect 13096 12374 13124 13330
rect 13266 13016 13322 13025
rect 13266 12951 13322 12960
rect 13084 12368 13136 12374
rect 13084 12310 13136 12316
rect 13096 11626 13124 12310
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12728 10742 12756 11086
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12728 10266 12756 10678
rect 12820 10266 12848 11222
rect 13096 10538 13124 11562
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 13096 10130 13124 10474
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 12624 9648 12676 9654
rect 12624 9590 12676 9596
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11152 8900 11204 8906
rect 11152 8842 11204 8848
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 11242 8392 11298 8401
rect 11242 8327 11298 8336
rect 11256 7342 11284 8327
rect 11532 8090 11560 8978
rect 12268 8498 12296 9046
rect 12452 8838 12480 9318
rect 12544 9178 12572 9386
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 12268 8022 12296 8434
rect 12348 8356 12400 8362
rect 12348 8298 12400 8304
rect 12360 8090 12388 8298
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12256 8016 12308 8022
rect 12256 7958 12308 7964
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 11256 6458 11284 6802
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11348 5778 11376 7822
rect 11440 7002 11468 7890
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10876 5296 10928 5302
rect 10876 5238 10928 5244
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 10060 4282 10088 4966
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 10060 4010 10088 4218
rect 10152 4214 10180 4966
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10980 4690 11008 5646
rect 11348 5370 11376 5714
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 10140 4208 10192 4214
rect 10140 4150 10192 4156
rect 10888 4146 10916 4422
rect 10980 4146 11008 4626
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 11256 3670 11284 5170
rect 11440 4154 11468 5510
rect 11900 4554 11928 7278
rect 12268 7206 12296 7958
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 11888 4548 11940 4554
rect 11888 4490 11940 4496
rect 11348 4126 11468 4154
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 11244 3664 11296 3670
rect 11244 3606 11296 3612
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 10336 3194 10364 3606
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 8942 2952 8998 2961
rect 8942 2887 8998 2896
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 9494 2680 9550 2689
rect 9036 2644 9088 2650
rect 10289 2672 10585 2692
rect 10796 2650 10824 2790
rect 9494 2615 9550 2624
rect 10784 2644 10836 2650
rect 9036 2586 9088 2592
rect 8024 2576 8076 2582
rect 8300 2576 8352 2582
rect 8076 2536 8300 2564
rect 8024 2518 8076 2524
rect 8300 2518 8352 2524
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 8852 2576 8904 2582
rect 8852 2518 8904 2524
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 7196 2372 7248 2378
rect 7196 2314 7248 2320
rect 8116 2372 8168 2378
rect 8116 2314 8168 2320
rect 6826 1320 6882 1329
rect 6826 1255 6882 1264
rect 6458 54 6776 82
rect 7208 82 7236 2314
rect 7470 82 7526 480
rect 7208 54 7526 82
rect 8128 82 8156 2314
rect 8390 82 8446 480
rect 8128 54 8446 82
rect 9048 82 9076 2586
rect 9508 2582 9536 2615
rect 10784 2586 10836 2592
rect 9496 2576 9548 2582
rect 9496 2518 9548 2524
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 9600 2310 9628 2450
rect 11256 2446 11284 3470
rect 11348 2922 11376 4126
rect 11888 3664 11940 3670
rect 11888 3606 11940 3612
rect 11900 3194 11928 3606
rect 11980 3460 12032 3466
rect 11980 3402 12032 3408
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11336 2916 11388 2922
rect 11336 2858 11388 2864
rect 11992 2650 12020 3402
rect 12084 3126 12112 7142
rect 12268 7002 12296 7142
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12268 6458 12296 6938
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12268 5846 12296 6394
rect 12256 5840 12308 5846
rect 12256 5782 12308 5788
rect 12164 5092 12216 5098
rect 12164 5034 12216 5040
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 12084 2922 12112 3062
rect 12072 2916 12124 2922
rect 12072 2858 12124 2864
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 11610 2408 11666 2417
rect 11520 2372 11572 2378
rect 11572 2352 11610 2360
rect 11572 2343 11666 2352
rect 11572 2332 11652 2343
rect 11520 2314 11572 2320
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 11060 2100 11112 2106
rect 11060 2042 11112 2048
rect 10140 1964 10192 1970
rect 10140 1906 10192 1912
rect 9402 82 9458 480
rect 9048 54 9458 82
rect 10152 82 10180 1906
rect 10414 82 10470 480
rect 10152 54 10470 82
rect 11072 82 11100 2042
rect 11426 82 11482 480
rect 11072 54 11482 82
rect 12176 82 12204 5034
rect 12256 5024 12308 5030
rect 12256 4966 12308 4972
rect 12268 4826 12296 4966
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 12268 4010 12296 4762
rect 12256 4004 12308 4010
rect 12256 3946 12308 3952
rect 12254 3496 12310 3505
rect 12254 3431 12310 3440
rect 12268 2582 12296 3431
rect 12360 3194 12388 8026
rect 12452 4154 12480 8774
rect 12544 8498 12572 8842
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12636 8090 12664 9590
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 13188 8498 13216 9386
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12636 7342 12664 8026
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12544 6866 12572 7142
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12544 5914 12572 6122
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 12636 5574 12664 6122
rect 12912 5846 12940 6598
rect 13188 6322 13216 8434
rect 13280 7954 13308 12951
rect 13372 12714 13400 14010
rect 13464 14006 13492 15524
rect 14004 15506 14056 15512
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13648 14890 13676 15302
rect 13924 15026 13952 15438
rect 14016 15162 14044 15506
rect 14004 15156 14056 15162
rect 14004 15098 14056 15104
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 13636 14884 13688 14890
rect 13556 14844 13636 14872
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 13360 12708 13412 12714
rect 13360 12650 13412 12656
rect 13372 12442 13400 12650
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 13556 12374 13584 14844
rect 13636 14826 13688 14832
rect 13740 14618 13768 14962
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13924 14550 13952 14962
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13912 14544 13964 14550
rect 13912 14486 13964 14492
rect 13648 13802 13676 14486
rect 13636 13796 13688 13802
rect 13636 13738 13688 13744
rect 13648 13394 13676 13738
rect 14108 13394 14136 24550
rect 14280 24404 14332 24410
rect 14280 24346 14332 24352
rect 14188 24200 14240 24206
rect 14188 24142 14240 24148
rect 14200 23662 14228 24142
rect 14292 23798 14320 24346
rect 14476 23866 14504 24550
rect 14752 24274 14780 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14740 24268 14792 24274
rect 14740 24210 14792 24216
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14464 23860 14516 23866
rect 14464 23802 14516 23808
rect 14280 23792 14332 23798
rect 14280 23734 14332 23740
rect 14476 23662 14504 23802
rect 14188 23656 14240 23662
rect 14188 23598 14240 23604
rect 14464 23656 14516 23662
rect 14464 23598 14516 23604
rect 14200 23322 14228 23598
rect 14188 23316 14240 23322
rect 14188 23258 14240 23264
rect 14200 22982 14228 23258
rect 14476 23186 14504 23598
rect 14556 23588 14608 23594
rect 14556 23530 14608 23536
rect 14464 23180 14516 23186
rect 14464 23122 14516 23128
rect 14188 22976 14240 22982
rect 14188 22918 14240 22924
rect 14200 22574 14228 22918
rect 14476 22778 14504 23122
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 14280 22704 14332 22710
rect 14280 22646 14332 22652
rect 14292 22574 14320 22646
rect 14476 22574 14504 22714
rect 14188 22568 14240 22574
rect 14188 22510 14240 22516
rect 14280 22568 14332 22574
rect 14280 22510 14332 22516
rect 14464 22568 14516 22574
rect 14464 22510 14516 22516
rect 14292 22234 14320 22510
rect 14280 22228 14332 22234
rect 14280 22170 14332 22176
rect 14464 22024 14516 22030
rect 14464 21966 14516 21972
rect 14476 21690 14504 21966
rect 14464 21684 14516 21690
rect 14464 21626 14516 21632
rect 14372 21412 14424 21418
rect 14372 21354 14424 21360
rect 14188 21072 14240 21078
rect 14188 21014 14240 21020
rect 14200 20788 14228 21014
rect 14384 20942 14412 21354
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 14372 20800 14424 20806
rect 14200 20760 14372 20788
rect 14372 20742 14424 20748
rect 14384 20262 14412 20742
rect 14372 20256 14424 20262
rect 14372 20198 14424 20204
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 14200 17882 14228 19110
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 14384 16726 14412 20198
rect 14464 19236 14516 19242
rect 14464 19178 14516 19184
rect 14476 18698 14504 19178
rect 14464 18692 14516 18698
rect 14464 18634 14516 18640
rect 14464 16992 14516 16998
rect 14464 16934 14516 16940
rect 14372 16720 14424 16726
rect 14372 16662 14424 16668
rect 14384 16454 14412 16662
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 14384 16250 14412 16390
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14370 16144 14426 16153
rect 14370 16079 14426 16088
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 14292 15706 14320 15982
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14292 13870 14320 14214
rect 14280 13864 14332 13870
rect 14280 13806 14332 13812
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13832 12850 13860 13126
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13820 12708 13872 12714
rect 13820 12650 13872 12656
rect 13544 12368 13596 12374
rect 13544 12310 13596 12316
rect 13556 11898 13584 12310
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13360 11620 13412 11626
rect 13360 11562 13412 11568
rect 13372 11150 13400 11562
rect 13556 11354 13584 11834
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13832 11082 13860 12650
rect 14108 12646 14136 13330
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13544 11008 13596 11014
rect 13544 10950 13596 10956
rect 13556 10674 13584 10950
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13556 10266 13584 10610
rect 13832 10538 13860 11018
rect 14108 10713 14136 12582
rect 14200 12374 14228 12650
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 14188 12232 14240 12238
rect 14240 12192 14320 12220
rect 14188 12174 14240 12180
rect 14292 11558 14320 12192
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14094 10704 14150 10713
rect 14094 10639 14150 10648
rect 13820 10532 13872 10538
rect 13820 10474 13872 10480
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13556 9722 13584 10066
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13556 8566 13584 8978
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13648 8498 13676 10202
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13740 9518 13768 9862
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13740 9178 13768 9454
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 14108 9042 14136 10066
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 14200 7954 14228 10406
rect 14292 10198 14320 11494
rect 14384 11218 14412 16079
rect 14476 13938 14504 16934
rect 14568 14618 14596 23530
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14740 22704 14792 22710
rect 14740 22646 14792 22652
rect 14648 22092 14700 22098
rect 14648 22034 14700 22040
rect 14660 21690 14688 22034
rect 14648 21684 14700 21690
rect 14648 21626 14700 21632
rect 14648 21344 14700 21350
rect 14648 21286 14700 21292
rect 14660 18902 14688 21286
rect 14648 18896 14700 18902
rect 14648 18838 14700 18844
rect 14660 18358 14688 18838
rect 14648 18352 14700 18358
rect 14648 18294 14700 18300
rect 14752 16590 14780 22646
rect 15304 22438 15332 23122
rect 15292 22432 15344 22438
rect 15292 22374 15344 22380
rect 15200 22160 15252 22166
rect 15200 22102 15252 22108
rect 15212 21876 15240 22102
rect 15304 22001 15332 22374
rect 15384 22024 15436 22030
rect 15290 21992 15346 22001
rect 15384 21966 15436 21972
rect 15290 21927 15346 21936
rect 15212 21848 15332 21876
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15304 21690 15332 21848
rect 15396 21690 15424 21966
rect 14832 21684 14884 21690
rect 14832 21626 14884 21632
rect 15292 21684 15344 21690
rect 15292 21626 15344 21632
rect 15384 21684 15436 21690
rect 15384 21626 15436 21632
rect 14844 20330 14872 21626
rect 15384 21412 15436 21418
rect 15384 21354 15436 21360
rect 15396 20806 15424 21354
rect 15384 20800 15436 20806
rect 15384 20742 15436 20748
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 14832 20324 14884 20330
rect 14832 20266 14884 20272
rect 14844 17270 14872 20266
rect 15304 20262 15332 20538
rect 15384 20392 15436 20398
rect 15384 20334 15436 20340
rect 15286 20256 15338 20262
rect 15286 20198 15338 20204
rect 15298 20139 15332 20198
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 19496 15332 20139
rect 15396 19718 15424 20334
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 15212 19468 15332 19496
rect 15212 19156 15240 19468
rect 15292 19168 15344 19174
rect 15212 19128 15292 19156
rect 15292 19110 15344 19116
rect 15304 18850 15332 19110
rect 15396 18970 15424 19654
rect 15488 19514 15516 27526
rect 15566 27520 15622 27526
rect 16132 27526 16358 27554
rect 16028 22432 16080 22438
rect 16028 22374 16080 22380
rect 15844 22024 15896 22030
rect 15844 21966 15896 21972
rect 15660 21412 15712 21418
rect 15660 21354 15712 21360
rect 15672 20466 15700 21354
rect 15856 20942 15884 21966
rect 15936 21072 15988 21078
rect 16040 21049 16068 22374
rect 15936 21014 15988 21020
rect 16026 21040 16082 21049
rect 15844 20936 15896 20942
rect 15844 20878 15896 20884
rect 15948 20602 15976 21014
rect 16026 20975 16082 20984
rect 15936 20596 15988 20602
rect 15936 20538 15988 20544
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15672 19854 15700 20402
rect 15936 20392 15988 20398
rect 15936 20334 15988 20340
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15568 19712 15620 19718
rect 15568 19654 15620 19660
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 15580 19310 15608 19654
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 15660 19236 15712 19242
rect 15660 19178 15712 19184
rect 15384 18964 15436 18970
rect 15384 18906 15436 18912
rect 15672 18850 15700 19178
rect 15304 18822 15700 18850
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15304 17796 15332 18822
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 15396 18086 15424 18702
rect 15568 18352 15620 18358
rect 15568 18294 15620 18300
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15476 17808 15528 17814
rect 15304 17768 15476 17796
rect 15476 17750 15528 17756
rect 15292 17604 15344 17610
rect 15292 17546 15344 17552
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15304 17270 15332 17546
rect 14832 17264 14884 17270
rect 14832 17206 14884 17212
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 14844 16250 14872 17206
rect 15488 16998 15516 17750
rect 15580 17066 15608 18294
rect 15856 17542 15884 19654
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 15948 17354 15976 20334
rect 16132 19922 16160 27526
rect 16302 27520 16358 27526
rect 16776 27526 17080 27554
rect 16396 22568 16448 22574
rect 16396 22510 16448 22516
rect 16408 20913 16436 22510
rect 16580 21548 16632 21554
rect 16580 21490 16632 21496
rect 16592 21146 16620 21490
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 16488 20936 16540 20942
rect 16394 20904 16450 20913
rect 16488 20878 16540 20884
rect 16394 20839 16450 20848
rect 16500 20602 16528 20878
rect 16488 20596 16540 20602
rect 16488 20538 16540 20544
rect 16580 20256 16632 20262
rect 16580 20198 16632 20204
rect 16592 20058 16620 20198
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16396 19984 16448 19990
rect 16396 19926 16448 19932
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 16040 19446 16068 19790
rect 16408 19514 16436 19926
rect 16396 19508 16448 19514
rect 16396 19450 16448 19456
rect 16028 19440 16080 19446
rect 16028 19382 16080 19388
rect 16040 18902 16068 19382
rect 16776 19174 16804 27526
rect 17052 27418 17080 27526
rect 17130 27520 17186 28000
rect 17958 27520 18014 28000
rect 18694 27520 18750 28000
rect 19522 27520 19578 28000
rect 20350 27554 20406 28000
rect 19996 27526 20406 27554
rect 17144 27418 17172 27520
rect 17052 27390 17172 27418
rect 17972 24614 18000 27520
rect 17960 24608 18012 24614
rect 17960 24550 18012 24556
rect 18708 24410 18736 27520
rect 18696 24404 18748 24410
rect 18696 24346 18748 24352
rect 18420 23656 18472 23662
rect 18420 23598 18472 23604
rect 16856 21888 16908 21894
rect 16856 21830 16908 21836
rect 16868 21418 16896 21830
rect 16856 21412 16908 21418
rect 16856 21354 16908 21360
rect 16868 20874 16896 21354
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 16856 20868 16908 20874
rect 16856 20810 16908 20816
rect 16868 19786 16896 20810
rect 16960 19961 16988 21286
rect 17500 21004 17552 21010
rect 17500 20946 17552 20952
rect 17512 20262 17540 20946
rect 17682 20496 17738 20505
rect 17682 20431 17738 20440
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 16946 19952 17002 19961
rect 16946 19887 17002 19896
rect 16856 19780 16908 19786
rect 16856 19722 16908 19728
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16028 18896 16080 18902
rect 16028 18838 16080 18844
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 16488 18624 16540 18630
rect 16488 18566 16540 18572
rect 16120 18216 16172 18222
rect 16120 18158 16172 18164
rect 15672 17326 15976 17354
rect 15568 17060 15620 17066
rect 15568 17002 15620 17008
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15580 16794 15608 17002
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 15396 15978 15424 16186
rect 15384 15972 15436 15978
rect 15384 15914 15436 15920
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 14740 15564 14792 15570
rect 14740 15506 14792 15512
rect 14752 15162 14780 15506
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14752 13025 14780 15098
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14844 14074 14872 14826
rect 15396 14482 15424 15642
rect 15476 14544 15528 14550
rect 15476 14486 15528 14492
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15396 14074 15424 14418
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15488 13938 15516 14486
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14738 13016 14794 13025
rect 14956 13008 15252 13028
rect 14738 12951 14794 12960
rect 15304 12918 15332 13126
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 15292 12912 15344 12918
rect 15292 12854 15344 12860
rect 14648 12368 14700 12374
rect 14648 12310 14700 12316
rect 14660 11898 14688 12310
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 14660 11626 14688 11834
rect 14648 11620 14700 11626
rect 14648 11562 14700 11568
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 14384 10810 14412 11154
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14476 10538 14504 11290
rect 14752 11150 14780 12854
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 14832 12436 14884 12442
rect 14832 12378 14884 12384
rect 14844 11694 14872 12378
rect 15212 12238 15240 12582
rect 15396 12306 15424 13466
rect 15488 12306 15516 13874
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15396 11830 15424 12242
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15384 11824 15436 11830
rect 15384 11766 15436 11772
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 15488 11286 15516 12038
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15580 11234 15608 15846
rect 15672 13297 15700 17326
rect 15844 16720 15896 16726
rect 15844 16662 15896 16668
rect 15856 16182 15884 16662
rect 16132 16658 16160 18158
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 16224 17814 16252 18022
rect 16212 17808 16264 17814
rect 16212 17750 16264 17756
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 15934 16552 15990 16561
rect 16028 16516 16080 16522
rect 15990 16496 16028 16504
rect 15934 16487 16028 16496
rect 15948 16476 16028 16487
rect 16028 16458 16080 16464
rect 16316 16250 16344 18566
rect 16500 18290 16528 18566
rect 16868 18290 16896 19722
rect 17224 18828 17276 18834
rect 17408 18828 17460 18834
rect 17276 18788 17356 18816
rect 17224 18770 17276 18776
rect 16488 18284 16540 18290
rect 16488 18226 16540 18232
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 16500 17270 16528 18226
rect 17328 18086 17356 18788
rect 17408 18770 17460 18776
rect 16672 18080 16724 18086
rect 16672 18022 16724 18028
rect 17316 18080 17368 18086
rect 17316 18022 17368 18028
rect 16684 17882 16712 18022
rect 16762 17912 16818 17921
rect 16672 17876 16724 17882
rect 16762 17847 16818 17856
rect 16672 17818 16724 17824
rect 16488 17264 16540 17270
rect 16488 17206 16540 17212
rect 16500 16726 16528 17206
rect 16488 16720 16540 16726
rect 16488 16662 16540 16668
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16304 16244 16356 16250
rect 16304 16186 16356 16192
rect 15844 16176 15896 16182
rect 15844 16118 15896 16124
rect 16592 15910 16620 16526
rect 16776 16046 16804 17847
rect 17040 17672 17092 17678
rect 17040 17614 17092 17620
rect 17052 17338 17080 17614
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16868 16794 16896 17138
rect 16856 16788 16908 16794
rect 16856 16730 16908 16736
rect 16764 16040 16816 16046
rect 16764 15982 16816 15988
rect 17222 16008 17278 16017
rect 17222 15943 17278 15952
rect 16580 15904 16632 15910
rect 16580 15846 16632 15852
rect 15844 15564 15896 15570
rect 15844 15506 15896 15512
rect 15856 15094 15884 15506
rect 15844 15088 15896 15094
rect 15844 15030 15896 15036
rect 15856 14006 15884 15030
rect 16028 14952 16080 14958
rect 16028 14894 16080 14900
rect 15844 14000 15896 14006
rect 15844 13942 15896 13948
rect 15856 13814 15884 13942
rect 15764 13786 15884 13814
rect 15764 13394 15792 13786
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15658 13288 15714 13297
rect 15658 13223 15714 13232
rect 15764 12986 15792 13330
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 15764 11898 15792 12582
rect 15856 12238 15884 13262
rect 16040 12714 16068 14894
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16224 14618 16252 14758
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16028 12708 16080 12714
rect 16028 12650 16080 12656
rect 15936 12300 15988 12306
rect 15936 12242 15988 12248
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15948 11898 15976 12242
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15936 11892 15988 11898
rect 15936 11834 15988 11840
rect 16040 11286 16068 12650
rect 16592 11898 16620 15846
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 16868 14958 16896 15506
rect 17236 15502 17264 15943
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16868 12986 16896 13330
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16960 12442 16988 13466
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 17132 12436 17184 12442
rect 17132 12378 17184 12384
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16028 11280 16080 11286
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 14752 10538 14780 11086
rect 14464 10532 14516 10538
rect 14464 10474 14516 10480
rect 14740 10532 14792 10538
rect 14740 10474 14792 10480
rect 14844 10266 14872 11222
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15488 10810 15516 11222
rect 15580 11206 15700 11234
rect 16028 11222 16080 11228
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15580 10674 15608 11086
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 14280 10192 14332 10198
rect 14280 10134 14332 10140
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14924 9444 14976 9450
rect 14924 9386 14976 9392
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14292 8294 14320 9318
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 14568 8838 14596 8978
rect 14936 8974 14964 9386
rect 15580 9382 15608 10066
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15396 9110 15424 9318
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14568 8498 14596 8774
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 13280 7546 13308 7890
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13280 6730 13308 7482
rect 13268 6724 13320 6730
rect 13268 6666 13320 6672
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 12900 5840 12952 5846
rect 12900 5782 12952 5788
rect 13188 5692 13216 6258
rect 13728 5840 13780 5846
rect 13728 5782 13780 5788
rect 13268 5704 13320 5710
rect 13188 5664 13268 5692
rect 13268 5646 13320 5652
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13084 5636 13136 5642
rect 13084 5578 13136 5584
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 13004 5098 13032 5510
rect 13096 5234 13124 5578
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 12992 5092 13044 5098
rect 12992 5034 13044 5040
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12728 4486 12756 4966
rect 13004 4826 13032 5034
rect 13280 4826 13308 5646
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12452 4126 12572 4154
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12452 3738 12480 3878
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12544 3670 12572 4126
rect 12532 3664 12584 3670
rect 12532 3606 12584 3612
rect 12544 3194 12572 3606
rect 12728 3466 12756 4422
rect 13464 4078 13492 5646
rect 13740 5370 13768 5782
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13636 4616 13688 4622
rect 13832 4604 13860 7822
rect 14200 7546 14228 7890
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14200 7342 14228 7482
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 14200 5846 14228 7278
rect 14292 7002 14320 8230
rect 14384 8090 14412 8366
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14568 7750 14596 8434
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15488 8022 15516 8230
rect 15476 8016 15528 8022
rect 15476 7958 15528 7964
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14568 7342 14596 7686
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 15200 7268 15252 7274
rect 15200 7210 15252 7216
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14292 6186 14320 6938
rect 15212 6866 15240 7210
rect 15396 7002 15424 7822
rect 15488 7206 15516 7958
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 15200 6860 15252 6866
rect 15252 6820 15332 6848
rect 15200 6802 15252 6808
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 14280 6180 14332 6186
rect 14280 6122 14332 6128
rect 14476 5914 14504 6258
rect 15304 5914 15332 6820
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 14188 5840 14240 5846
rect 14188 5782 14240 5788
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 14280 5636 14332 5642
rect 14280 5578 14332 5584
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 13688 4576 13860 4604
rect 13636 4558 13688 4564
rect 13832 4282 13860 4576
rect 14016 4282 14044 4626
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13464 3738 13492 4014
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 12716 3460 12768 3466
rect 12716 3402 12768 3408
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12360 2904 12388 3130
rect 12728 3058 12756 3402
rect 13832 3194 13860 3606
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 12716 3052 12768 3058
rect 12716 2994 12768 3000
rect 12624 2916 12676 2922
rect 12360 2876 12624 2904
rect 12360 2650 12388 2876
rect 12676 2876 12848 2904
rect 12624 2858 12676 2864
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 12820 2582 12848 2876
rect 12256 2576 12308 2582
rect 12256 2518 12308 2524
rect 12716 2576 12768 2582
rect 12716 2518 12768 2524
rect 12808 2576 12860 2582
rect 12808 2518 12860 2524
rect 12728 2310 12756 2518
rect 14016 2446 14044 3470
rect 14108 2650 14136 3674
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 14292 2514 14320 5578
rect 14660 5137 14688 5714
rect 15396 5574 15424 6054
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14646 5128 14702 5137
rect 14646 5063 14702 5072
rect 14660 5030 14688 5063
rect 14648 5024 14700 5030
rect 14648 4966 14700 4972
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14660 4282 14688 4626
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14752 4010 14780 4966
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15396 4010 15424 5510
rect 14740 4004 14792 4010
rect 14740 3946 14792 3952
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 15290 3632 15346 3641
rect 15290 3567 15346 3576
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14568 2922 14596 3334
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14556 2916 14608 2922
rect 14556 2858 14608 2864
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 12716 2304 12768 2310
rect 12716 2246 12768 2252
rect 13084 2032 13136 2038
rect 13084 1974 13136 1980
rect 12438 82 12494 480
rect 12176 54 12494 82
rect 13096 82 13124 1974
rect 14568 1601 14596 2858
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 14554 1592 14610 1601
rect 14554 1527 14610 1536
rect 13450 82 13506 480
rect 13096 54 13506 82
rect 6458 0 6514 54
rect 7470 0 7526 54
rect 8390 0 8446 54
rect 9402 0 9458 54
rect 10414 0 10470 54
rect 11426 0 11482 54
rect 12438 0 12494 54
rect 13450 0 13506 54
rect 14462 82 14518 480
rect 14752 82 14780 2246
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14462 54 14780 82
rect 15304 82 15332 3567
rect 15396 2922 15424 3946
rect 15488 3670 15516 7142
rect 15580 6361 15608 9318
rect 15672 8634 15700 11206
rect 15752 11076 15804 11082
rect 15752 11018 15804 11024
rect 15764 10810 15792 11018
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15752 10532 15804 10538
rect 15752 10474 15804 10480
rect 15764 10033 15792 10474
rect 15750 10024 15806 10033
rect 15750 9959 15806 9968
rect 15764 9518 15792 9959
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15752 9104 15804 9110
rect 15752 9046 15804 9052
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15764 8294 15792 9046
rect 15936 8900 15988 8906
rect 15936 8842 15988 8848
rect 15752 8288 15804 8294
rect 15752 8230 15804 8236
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15566 6352 15622 6361
rect 15566 6287 15622 6296
rect 15568 6248 15620 6254
rect 15672 6236 15700 6938
rect 15620 6208 15700 6236
rect 15568 6190 15620 6196
rect 15580 6118 15608 6190
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15580 5030 15608 6054
rect 15568 5024 15620 5030
rect 15568 4966 15620 4972
rect 15580 4826 15608 4966
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15476 3664 15528 3670
rect 15476 3606 15528 3612
rect 15488 3194 15516 3606
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15384 2916 15436 2922
rect 15384 2858 15436 2864
rect 15672 2582 15700 3130
rect 15764 3126 15792 8230
rect 15856 8022 15884 8230
rect 15844 8016 15896 8022
rect 15844 7958 15896 7964
rect 15856 7313 15884 7958
rect 15948 7818 15976 8842
rect 15936 7812 15988 7818
rect 15936 7754 15988 7760
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16500 7410 16528 7686
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 15842 7304 15898 7313
rect 15842 7239 15898 7248
rect 16120 7268 16172 7274
rect 16120 7210 16172 7216
rect 16212 7268 16264 7274
rect 16212 7210 16264 7216
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 15948 7002 15976 7142
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 15844 6928 15896 6934
rect 15844 6870 15896 6876
rect 15856 6322 15884 6870
rect 16132 6798 16160 7210
rect 16224 7002 16252 7210
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 15948 6458 15976 6734
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 16500 6322 16528 7346
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16776 5778 16804 11494
rect 16868 10606 16896 12106
rect 17144 11762 17172 12378
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 17040 11688 17092 11694
rect 17040 11630 17092 11636
rect 17052 11121 17080 11630
rect 17038 11112 17094 11121
rect 17038 11047 17094 11056
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16868 9382 16896 10066
rect 17052 9518 17080 11047
rect 17236 10130 17264 15302
rect 17328 15162 17356 18022
rect 17420 17882 17448 18770
rect 17408 17876 17460 17882
rect 17408 17818 17460 17824
rect 17408 17740 17460 17746
rect 17408 17682 17460 17688
rect 17420 16998 17448 17682
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 17328 12918 17356 13330
rect 17316 12912 17368 12918
rect 17316 12854 17368 12860
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17328 11898 17356 12242
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17236 9722 17264 10066
rect 17328 9994 17356 11834
rect 17316 9988 17368 9994
rect 17316 9930 17368 9936
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 16868 9042 16896 9318
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16868 8294 16896 8978
rect 17052 8974 17080 9318
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 16764 5772 16816 5778
rect 16764 5714 16816 5720
rect 16408 5370 16436 5714
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16580 5296 16632 5302
rect 16580 5238 16632 5244
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 16040 4604 16068 4762
rect 16132 4758 16160 4966
rect 16120 4752 16172 4758
rect 16120 4694 16172 4700
rect 16040 4576 16160 4604
rect 16028 4480 16080 4486
rect 16028 4422 16080 4428
rect 15844 4004 15896 4010
rect 15844 3946 15896 3952
rect 15856 3534 15884 3946
rect 15844 3528 15896 3534
rect 16040 3505 16068 4422
rect 16132 3942 16160 4576
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 16132 3516 16160 3878
rect 16224 3670 16252 4422
rect 16592 4078 16620 5238
rect 16776 5098 16804 5714
rect 16868 5681 16896 8230
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 17144 7546 17172 7890
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 17040 7472 17092 7478
rect 17040 7414 17092 7420
rect 17052 6866 17080 7414
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 17052 6458 17080 6802
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 16854 5672 16910 5681
rect 16854 5607 16910 5616
rect 16764 5092 16816 5098
rect 16764 5034 16816 5040
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16868 4282 16896 4966
rect 16960 4690 16988 5850
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 17052 4826 17080 5714
rect 17420 5370 17448 16934
rect 17512 10169 17540 20198
rect 17696 19360 17724 20431
rect 17776 19916 17828 19922
rect 17776 19858 17828 19864
rect 17788 19514 17816 19858
rect 17776 19508 17828 19514
rect 17776 19450 17828 19456
rect 18326 19408 18382 19417
rect 17776 19372 17828 19378
rect 17696 19332 17776 19360
rect 18326 19343 18382 19352
rect 17776 19314 17828 19320
rect 17788 19174 17816 19314
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 17592 12300 17644 12306
rect 17788 12288 17816 19110
rect 18156 18970 18184 19246
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 18340 18834 18368 19343
rect 18328 18828 18380 18834
rect 18328 18770 18380 18776
rect 18340 18426 18368 18770
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18326 17776 18382 17785
rect 18326 17711 18382 17720
rect 18340 17678 18368 17711
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18340 17338 18368 17614
rect 18328 17332 18380 17338
rect 18328 17274 18380 17280
rect 18236 15904 18288 15910
rect 18236 15846 18288 15852
rect 18144 15564 18196 15570
rect 18144 15506 18196 15512
rect 18156 15162 18184 15506
rect 18248 15473 18276 15846
rect 18432 15638 18460 23598
rect 18512 20392 18564 20398
rect 18512 20334 18564 20340
rect 18524 20262 18552 20334
rect 18512 20256 18564 20262
rect 18512 20198 18564 20204
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 18524 19854 18552 20198
rect 18512 19848 18564 19854
rect 18616 19825 18644 20198
rect 18788 19916 18840 19922
rect 18788 19858 18840 19864
rect 18512 19790 18564 19796
rect 18602 19816 18658 19825
rect 18524 17270 18552 19790
rect 18602 19751 18658 19760
rect 18800 19310 18828 19858
rect 18972 19712 19024 19718
rect 18972 19654 19024 19660
rect 18788 19304 18840 19310
rect 18786 19272 18788 19281
rect 18840 19272 18842 19281
rect 18786 19207 18842 19216
rect 18984 18873 19012 19654
rect 18970 18864 19026 18873
rect 18970 18799 19026 18808
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 18512 17264 18564 17270
rect 18616 17241 18644 18566
rect 18696 17536 18748 17542
rect 18696 17478 18748 17484
rect 18512 17206 18564 17212
rect 18602 17232 18658 17241
rect 18602 17167 18658 17176
rect 18604 16652 18656 16658
rect 18604 16594 18656 16600
rect 18616 16250 18644 16594
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 18420 15632 18472 15638
rect 18708 15609 18736 17478
rect 19536 16250 19564 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19524 16244 19576 16250
rect 19524 16186 19576 16192
rect 19996 16182 20024 27526
rect 20350 27520 20406 27526
rect 21086 27520 21142 28000
rect 21914 27554 21970 28000
rect 21652 27526 21970 27554
rect 20720 24268 20772 24274
rect 20720 24210 20772 24216
rect 20732 23730 20760 24210
rect 21100 23866 21128 27520
rect 21088 23860 21140 23866
rect 21088 23802 21140 23808
rect 21652 23798 21680 27526
rect 21914 27520 21970 27526
rect 22742 27520 22798 28000
rect 23478 27520 23534 28000
rect 23952 27526 24256 27554
rect 22756 23866 22784 27520
rect 23492 24410 23520 27520
rect 23480 24404 23532 24410
rect 23480 24346 23532 24352
rect 22744 23860 22796 23866
rect 22744 23802 22796 23808
rect 21640 23792 21692 23798
rect 21640 23734 21692 23740
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 20260 23656 20312 23662
rect 20260 23598 20312 23604
rect 19984 16176 20036 16182
rect 19984 16118 20036 16124
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 18420 15574 18472 15580
rect 18694 15600 18750 15609
rect 18694 15535 18750 15544
rect 18234 15464 18290 15473
rect 18234 15399 18290 15408
rect 18144 15156 18196 15162
rect 18144 15098 18196 15104
rect 18156 14414 18184 15098
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 20272 14618 20300 23598
rect 20732 16153 20760 23666
rect 21364 23656 21416 23662
rect 21364 23598 21416 23604
rect 23480 23656 23532 23662
rect 23480 23598 23532 23604
rect 21376 20466 21404 23598
rect 22284 22568 22336 22574
rect 22284 22510 22336 22516
rect 22296 22234 22324 22510
rect 22284 22228 22336 22234
rect 22284 22170 22336 22176
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 20718 16144 20774 16153
rect 20718 16079 20774 16088
rect 23492 16017 23520 23598
rect 23952 22778 23980 27526
rect 24228 27418 24256 27526
rect 24306 27520 24362 28000
rect 25134 27520 25190 28000
rect 25870 27520 25926 28000
rect 26698 27520 26754 28000
rect 27526 27520 27582 28000
rect 24320 27418 24348 27520
rect 24228 27390 24348 27418
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 25148 24721 25176 27520
rect 25134 24712 25190 24721
rect 25134 24647 25190 24656
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 23940 22772 23992 22778
rect 23940 22714 23992 22720
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 25884 21690 25912 27520
rect 26712 24313 26740 27520
rect 26698 24304 26754 24313
rect 26698 24239 26754 24248
rect 27540 23866 27568 27520
rect 27528 23860 27580 23866
rect 27528 23802 27580 23808
rect 25872 21684 25924 21690
rect 25872 21626 25924 21632
rect 23940 21480 23992 21486
rect 23940 21422 23992 21428
rect 23952 20398 23980 21422
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 23940 20392 23992 20398
rect 23940 20334 23992 20340
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 23478 16008 23534 16017
rect 23478 15943 23534 15952
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 20260 14612 20312 14618
rect 20260 14554 20312 14560
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 19536 12753 19564 14554
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 19522 12744 19578 12753
rect 19522 12679 19578 12688
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 17644 12260 17816 12288
rect 17592 12242 17644 12248
rect 17604 11558 17632 12242
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 17498 10160 17554 10169
rect 17498 10095 17554 10104
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 17512 6866 17540 9862
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17512 6118 17540 6802
rect 17500 6112 17552 6118
rect 17500 6054 17552 6060
rect 17512 5846 17540 6054
rect 17500 5840 17552 5846
rect 17500 5782 17552 5788
rect 17788 5370 17816 7210
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 18420 6724 18472 6730
rect 18420 6666 18472 6672
rect 17958 6216 18014 6225
rect 17958 6151 18014 6160
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 17420 5166 17448 5306
rect 17788 5166 17816 5306
rect 17408 5160 17460 5166
rect 17408 5102 17460 5108
rect 17776 5160 17828 5166
rect 17776 5102 17828 5108
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 16948 4684 17000 4690
rect 16948 4626 17000 4632
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16672 4208 16724 4214
rect 16672 4150 16724 4156
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16304 4004 16356 4010
rect 16304 3946 16356 3952
rect 16212 3664 16264 3670
rect 16212 3606 16264 3612
rect 15844 3470 15896 3476
rect 16026 3496 16082 3505
rect 16132 3488 16252 3516
rect 16026 3431 16082 3440
rect 15752 3120 15804 3126
rect 15752 3062 15804 3068
rect 16120 2916 16172 2922
rect 16120 2858 16172 2864
rect 15660 2576 15712 2582
rect 15660 2518 15712 2524
rect 16132 2378 16160 2858
rect 16224 2854 16252 3488
rect 16212 2848 16264 2854
rect 16212 2790 16264 2796
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 15382 82 15438 480
rect 15304 54 15438 82
rect 16316 82 16344 3946
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16408 3126 16436 3334
rect 16396 3120 16448 3126
rect 16396 3062 16448 3068
rect 16500 3058 16528 3674
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16592 2582 16620 3878
rect 16684 3602 16712 4150
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16776 3058 16804 3470
rect 17144 3466 17172 4558
rect 17420 4154 17448 5102
rect 17788 4758 17816 5102
rect 17500 4752 17552 4758
rect 17500 4694 17552 4700
rect 17776 4752 17828 4758
rect 17776 4694 17828 4700
rect 17512 4214 17540 4694
rect 17328 4126 17448 4154
rect 17500 4208 17552 4214
rect 17500 4150 17552 4156
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 17236 3738 17264 3878
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17132 3460 17184 3466
rect 17132 3402 17184 3408
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 16776 2582 16804 2994
rect 16580 2576 16632 2582
rect 16580 2518 16632 2524
rect 16764 2576 16816 2582
rect 16764 2518 16816 2524
rect 17144 2378 17172 3402
rect 17328 3097 17356 4126
rect 17684 4072 17736 4078
rect 17684 4014 17736 4020
rect 17408 3664 17460 3670
rect 17408 3606 17460 3612
rect 17420 3194 17448 3606
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17314 3088 17370 3097
rect 17314 3023 17370 3032
rect 17132 2372 17184 2378
rect 17132 2314 17184 2320
rect 16394 82 16450 480
rect 16316 54 16450 82
rect 14462 0 14518 54
rect 15382 0 15438 54
rect 16394 0 16450 54
rect 17406 82 17462 480
rect 17696 82 17724 4014
rect 17788 3670 17816 4694
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17776 3664 17828 3670
rect 17776 3606 17828 3612
rect 17880 2514 17908 4422
rect 17972 2990 18000 6151
rect 18432 5778 18460 6666
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18420 5772 18472 5778
rect 18420 5714 18472 5720
rect 18432 5370 18460 5714
rect 18420 5364 18472 5370
rect 18420 5306 18472 5312
rect 18524 5234 18552 5850
rect 18880 5772 18932 5778
rect 18880 5714 18932 5720
rect 18892 5370 18920 5714
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 18880 5364 18932 5370
rect 18880 5306 18932 5312
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 18420 5024 18472 5030
rect 18420 4966 18472 4972
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 17868 2508 17920 2514
rect 17868 2450 17920 2456
rect 17406 54 17724 82
rect 18156 82 18184 2790
rect 18432 2564 18460 4966
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 18604 3664 18656 3670
rect 18604 3606 18656 3612
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18524 3194 18552 3470
rect 18512 3188 18564 3194
rect 18512 3130 18564 3136
rect 18616 2922 18644 3606
rect 18604 2916 18656 2922
rect 18604 2858 18656 2864
rect 18512 2576 18564 2582
rect 18432 2536 18512 2564
rect 18512 2518 18564 2524
rect 19352 2514 19380 4082
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 24214 3496 24270 3505
rect 24214 3431 24270 3440
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 19524 2984 19576 2990
rect 19524 2926 19576 2932
rect 20444 2984 20496 2990
rect 20444 2926 20496 2932
rect 19340 2508 19392 2514
rect 19340 2450 19392 2456
rect 19156 2372 19208 2378
rect 19156 2314 19208 2320
rect 18418 82 18474 480
rect 18156 54 18474 82
rect 19168 82 19196 2314
rect 19536 2310 19564 2926
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19524 2304 19576 2310
rect 19524 2246 19576 2252
rect 20456 2009 20484 2926
rect 20536 2644 20588 2650
rect 20536 2586 20588 2592
rect 20442 2000 20498 2009
rect 20442 1935 20498 1944
rect 19430 82 19486 480
rect 19168 54 19486 82
rect 17406 0 17462 54
rect 18418 0 18474 54
rect 19430 0 19486 54
rect 20442 82 20498 480
rect 20548 82 20576 2586
rect 21180 2372 21232 2378
rect 21180 2314 21232 2320
rect 20442 54 20576 82
rect 21192 82 21220 2314
rect 21454 82 21510 480
rect 21192 54 21510 82
rect 22112 82 22140 3062
rect 22374 2952 22430 2961
rect 22374 2887 22430 2896
rect 22388 2514 22416 2887
rect 23480 2644 23532 2650
rect 23480 2586 23532 2592
rect 22376 2508 22428 2514
rect 22376 2450 22428 2456
rect 22374 82 22430 480
rect 22112 54 22430 82
rect 20442 0 20498 54
rect 21454 0 21510 54
rect 22374 0 22430 54
rect 23386 82 23442 480
rect 23492 82 23520 2586
rect 24228 2514 24256 3431
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 25504 2848 25556 2854
rect 25504 2790 25556 2796
rect 24216 2508 24268 2514
rect 24216 2450 24268 2456
rect 24124 2372 24176 2378
rect 24124 2314 24176 2320
rect 23386 54 23520 82
rect 24136 82 24164 2314
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24398 82 24454 480
rect 24136 54 24454 82
rect 23386 0 23442 54
rect 24398 0 24454 54
rect 25410 82 25466 480
rect 25516 82 25544 2790
rect 26146 2408 26202 2417
rect 26146 2343 26202 2352
rect 27528 2372 27580 2378
rect 25410 54 25544 82
rect 26160 82 26188 2343
rect 27528 2314 27580 2320
rect 26422 82 26478 480
rect 26160 54 26478 82
rect 25410 0 25466 54
rect 26422 0 26478 54
rect 27434 82 27490 480
rect 27540 82 27568 2314
rect 27434 54 27568 82
rect 27434 0 27490 54
<< via2 >>
rect 1490 25336 1546 25392
rect 110 21664 166 21720
rect 110 20304 166 20360
rect 110 19216 166 19272
rect 110 16088 166 16144
rect 1582 24248 1638 24304
rect 1582 22480 1638 22536
rect 2502 26696 2558 26752
rect 2042 20984 2098 21040
rect 2962 20848 3018 20904
rect 2686 19080 2742 19136
rect 3514 21936 3570 21992
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 3238 19760 3294 19816
rect 4986 19216 5042 19272
rect 1398 12688 1454 12744
rect 3146 16904 3202 16960
rect 4250 18264 4306 18320
rect 2318 8336 2374 8392
rect 4894 17584 4950 17640
rect 3974 14184 4030 14240
rect 4250 13640 4306 13696
rect 4250 6296 4306 6352
rect 4066 2624 4122 2680
rect 5170 19080 5226 19136
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5446 19896 5502 19952
rect 5998 19896 6054 19952
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5630 17584 5686 17640
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5722 15952 5778 16008
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 6274 18400 6330 18456
rect 6182 15408 6238 15464
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5170 13232 5226 13288
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5354 10104 5410 10160
rect 5170 2624 5226 2680
rect 5170 1536 5226 1592
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 6182 8472 6238 8528
rect 7102 15544 7158 15600
rect 6826 10648 6882 10704
rect 6090 6160 6146 6216
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5814 3440 5870 3496
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 6274 3596 6330 3632
rect 6274 3576 6276 3596
rect 6276 3576 6328 3596
rect 6328 3576 6330 3596
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6642 1944 6698 2000
rect 7102 2760 7158 2816
rect 8114 18808 8170 18864
rect 8022 17720 8078 17776
rect 8206 17176 8262 17232
rect 8390 16496 8446 16552
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10690 24656 10746 24712
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 8942 21936 8998 21992
rect 8022 12688 8078 12744
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 9770 19216 9826 19272
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10782 19352 10838 19408
rect 9034 12960 9090 13016
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 9310 13640 9366 13696
rect 7470 5208 7526 5264
rect 7838 5072 7894 5128
rect 11334 19216 11390 19272
rect 11058 18400 11114 18456
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 8574 2760 8630 2816
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 12622 17856 12678 17912
rect 13726 24248 13782 24304
rect 14002 20440 14058 20496
rect 13266 12960 13322 13016
rect 11242 8336 11298 8392
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 8942 2896 8998 2952
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 9494 2624 9550 2680
rect 6826 1264 6882 1320
rect 11610 2352 11666 2408
rect 12254 3440 12310 3496
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14370 16088 14426 16144
rect 14094 10648 14150 10704
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 15290 21936 15346 21992
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 16026 20984 16082 21040
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 16394 20848 16450 20904
rect 17682 20440 17738 20496
rect 16946 19896 17002 19952
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14738 12960 14794 13016
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 15934 16496 15990 16552
rect 16762 17856 16818 17912
rect 17222 15952 17278 16008
rect 15658 13232 15714 13288
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14646 5072 14702 5128
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15290 3576 15346 3632
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14554 1536 14610 1592
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15750 9968 15806 10024
rect 15566 6296 15622 6352
rect 15842 7248 15898 7304
rect 17038 11056 17094 11112
rect 16854 5616 16910 5672
rect 18326 19352 18382 19408
rect 18326 17720 18382 17776
rect 18602 19760 18658 19816
rect 18786 19252 18788 19272
rect 18788 19252 18840 19272
rect 18840 19252 18842 19272
rect 18786 19216 18842 19252
rect 18970 18808 19026 18864
rect 18602 17176 18658 17232
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 18694 15544 18750 15600
rect 18234 15408 18290 15464
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 20718 16088 20774 16144
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 25134 24656 25190 24712
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 26698 24248 26754 24304
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 23478 15952 23534 16008
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 19522 12688 19578 12744
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 17498 10104 17554 10160
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 17958 6160 18014 6216
rect 16026 3440 16082 3496
rect 17314 3032 17370 3088
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 24214 3440 24270 3496
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20442 1944 20498 2000
rect 22374 2896 22430 2952
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 26146 2352 26202 2408
<< metal3 >>
rect 0 27208 480 27328
rect 62 26754 122 27208
rect 2497 26754 2563 26757
rect 62 26752 2563 26754
rect 62 26696 2502 26752
rect 2558 26696 2563 26752
rect 62 26694 2563 26696
rect 2497 26691 2563 26694
rect 0 25848 480 25968
rect 62 25394 122 25848
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 1485 25394 1551 25397
rect 62 25392 1551 25394
rect 62 25336 1490 25392
rect 1546 25336 1551 25392
rect 62 25334 1551 25336
rect 1485 25331 1551 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 10685 24714 10751 24717
rect 25129 24714 25195 24717
rect 10685 24712 25195 24714
rect 10685 24656 10690 24712
rect 10746 24656 25134 24712
rect 25190 24656 25195 24712
rect 10685 24654 25195 24656
rect 10685 24651 10751 24654
rect 25129 24651 25195 24654
rect 0 24580 480 24608
rect 0 24516 60 24580
rect 124 24516 480 24580
rect 0 24488 480 24516
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 54 24244 60 24308
rect 124 24306 130 24308
rect 1577 24306 1643 24309
rect 124 24304 1643 24306
rect 124 24248 1582 24304
rect 1638 24248 1643 24304
rect 124 24246 1643 24248
rect 124 24244 130 24246
rect 1577 24243 1643 24246
rect 13721 24306 13787 24309
rect 26693 24306 26759 24309
rect 13721 24304 26759 24306
rect 13721 24248 13726 24304
rect 13782 24248 26698 24304
rect 26754 24248 26759 24304
rect 13721 24246 26759 24248
rect 13721 24243 13787 24246
rect 26693 24243 26759 24246
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 0 22992 480 23112
rect 62 22538 122 22992
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 1577 22538 1643 22541
rect 62 22536 1643 22538
rect 62 22480 1582 22536
rect 1638 22480 1643 22536
rect 62 22478 1643 22480
rect 1577 22475 1643 22478
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 3509 21994 3575 21997
rect 8937 21994 9003 21997
rect 15285 21994 15351 21997
rect 3509 21992 15351 21994
rect 3509 21936 3514 21992
rect 3570 21936 8942 21992
rect 8998 21936 15290 21992
rect 15346 21936 15351 21992
rect 3509 21934 15351 21936
rect 3509 21931 3575 21934
rect 8937 21931 9003 21934
rect 15285 21931 15351 21934
rect 5610 21792 5930 21793
rect 0 21720 480 21752
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 0 21664 110 21720
rect 166 21664 480 21720
rect 0 21632 480 21664
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 2037 21042 2103 21045
rect 16021 21042 16087 21045
rect 2037 21040 16087 21042
rect 2037 20984 2042 21040
rect 2098 20984 16026 21040
rect 16082 20984 16087 21040
rect 2037 20982 16087 20984
rect 2037 20979 2103 20982
rect 16021 20979 16087 20982
rect 2957 20906 3023 20909
rect 16389 20906 16455 20909
rect 2957 20904 16455 20906
rect 2957 20848 2962 20904
rect 3018 20848 16394 20904
rect 16450 20848 16455 20904
rect 2957 20846 16455 20848
rect 2957 20843 3023 20846
rect 16389 20843 16455 20846
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 13997 20498 14063 20501
rect 17677 20498 17743 20501
rect 13997 20496 17743 20498
rect 13997 20440 14002 20496
rect 14058 20440 17682 20496
rect 17738 20440 17743 20496
rect 13997 20438 17743 20440
rect 13997 20435 14063 20438
rect 17677 20435 17743 20438
rect 0 20360 480 20392
rect 0 20304 110 20360
rect 166 20304 480 20360
rect 0 20272 480 20304
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 5441 19954 5507 19957
rect 5993 19954 6059 19957
rect 16941 19954 17007 19957
rect 5441 19952 17007 19954
rect 5441 19896 5446 19952
rect 5502 19896 5998 19952
rect 6054 19896 16946 19952
rect 17002 19896 17007 19952
rect 5441 19894 17007 19896
rect 5441 19891 5507 19894
rect 5993 19891 6059 19894
rect 16941 19891 17007 19894
rect 3233 19818 3299 19821
rect 18597 19818 18663 19821
rect 3233 19816 18663 19818
rect 3233 19760 3238 19816
rect 3294 19760 18602 19816
rect 18658 19760 18663 19816
rect 3233 19758 18663 19760
rect 3233 19755 3299 19758
rect 18597 19755 18663 19758
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 10777 19410 10843 19413
rect 18321 19410 18387 19413
rect 10777 19408 18387 19410
rect 10777 19352 10782 19408
rect 10838 19352 18326 19408
rect 18382 19352 18387 19408
rect 10777 19350 18387 19352
rect 10777 19347 10843 19350
rect 18321 19347 18387 19350
rect 105 19274 171 19277
rect 4981 19274 5047 19277
rect 105 19272 5047 19274
rect 105 19216 110 19272
rect 166 19216 4986 19272
rect 5042 19216 5047 19272
rect 105 19214 5047 19216
rect 105 19211 171 19214
rect 4981 19211 5047 19214
rect 9765 19274 9831 19277
rect 11329 19274 11395 19277
rect 18781 19274 18847 19277
rect 9765 19272 18847 19274
rect 9765 19216 9770 19272
rect 9826 19216 11334 19272
rect 11390 19216 18786 19272
rect 18842 19216 18847 19272
rect 9765 19214 18847 19216
rect 9765 19211 9831 19214
rect 11329 19211 11395 19214
rect 18781 19211 18847 19214
rect 2681 19138 2747 19141
rect 5165 19138 5231 19141
rect 2681 19136 5231 19138
rect 2681 19080 2686 19136
rect 2742 19080 5170 19136
rect 5226 19080 5231 19136
rect 2681 19078 5231 19080
rect 2681 19075 2747 19078
rect 5165 19075 5231 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 0 18776 480 18896
rect 8109 18866 8175 18869
rect 18965 18866 19031 18869
rect 8109 18864 19031 18866
rect 8109 18808 8114 18864
rect 8170 18808 18970 18864
rect 19026 18808 19031 18864
rect 8109 18806 19031 18808
rect 8109 18803 8175 18806
rect 18965 18803 19031 18806
rect 62 18322 122 18776
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 6269 18458 6335 18461
rect 11053 18458 11119 18461
rect 6269 18456 11119 18458
rect 6269 18400 6274 18456
rect 6330 18400 11058 18456
rect 11114 18400 11119 18456
rect 6269 18398 11119 18400
rect 6269 18395 6335 18398
rect 11053 18395 11119 18398
rect 4245 18322 4311 18325
rect 62 18320 4311 18322
rect 62 18264 4250 18320
rect 4306 18264 4311 18320
rect 62 18262 4311 18264
rect 4245 18259 4311 18262
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 12617 17914 12683 17917
rect 16757 17914 16823 17917
rect 12617 17912 16823 17914
rect 12617 17856 12622 17912
rect 12678 17856 16762 17912
rect 16818 17856 16823 17912
rect 12617 17854 16823 17856
rect 12617 17851 12683 17854
rect 16757 17851 16823 17854
rect 8017 17778 8083 17781
rect 18321 17778 18387 17781
rect 8017 17776 18387 17778
rect 8017 17720 8022 17776
rect 8078 17720 18326 17776
rect 18382 17720 18387 17776
rect 8017 17718 18387 17720
rect 8017 17715 8083 17718
rect 18321 17715 18387 17718
rect 4889 17642 4955 17645
rect 5625 17642 5691 17645
rect 4889 17640 5691 17642
rect 4889 17584 4894 17640
rect 4950 17584 5630 17640
rect 5686 17584 5691 17640
rect 4889 17582 5691 17584
rect 4889 17579 4955 17582
rect 5625 17579 5691 17582
rect 0 17416 480 17536
rect 5610 17440 5930 17441
rect 62 16962 122 17416
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 8201 17234 8267 17237
rect 18597 17234 18663 17237
rect 8201 17232 18663 17234
rect 8201 17176 8206 17232
rect 8262 17176 18602 17232
rect 18658 17176 18663 17232
rect 8201 17174 18663 17176
rect 8201 17171 8267 17174
rect 18597 17171 18663 17174
rect 3141 16962 3207 16965
rect 62 16960 3207 16962
rect 62 16904 3146 16960
rect 3202 16904 3207 16960
rect 62 16902 3207 16904
rect 3141 16899 3207 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 8385 16554 8451 16557
rect 15929 16554 15995 16557
rect 8385 16552 15995 16554
rect 8385 16496 8390 16552
rect 8446 16496 15934 16552
rect 15990 16496 15995 16552
rect 8385 16494 15995 16496
rect 8385 16491 8451 16494
rect 15929 16491 15995 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 0 16144 480 16176
rect 14365 16146 14431 16149
rect 20713 16146 20779 16149
rect 0 16088 110 16144
rect 166 16088 480 16144
rect 0 16056 480 16088
rect 13770 16144 20779 16146
rect 13770 16088 14370 16144
rect 14426 16088 20718 16144
rect 20774 16088 20779 16144
rect 13770 16086 20779 16088
rect 5717 16010 5783 16013
rect 13770 16010 13830 16086
rect 14365 16083 14431 16086
rect 20713 16083 20779 16086
rect 5717 16008 13830 16010
rect 5717 15952 5722 16008
rect 5778 15952 13830 16008
rect 5717 15950 13830 15952
rect 17217 16010 17283 16013
rect 23473 16010 23539 16013
rect 17217 16008 23539 16010
rect 17217 15952 17222 16008
rect 17278 15952 23478 16008
rect 23534 15952 23539 16008
rect 17217 15950 23539 15952
rect 5717 15947 5783 15950
rect 17217 15947 17283 15950
rect 23473 15947 23539 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 7097 15602 7163 15605
rect 18689 15602 18755 15605
rect 7097 15600 18755 15602
rect 7097 15544 7102 15600
rect 7158 15544 18694 15600
rect 18750 15544 18755 15600
rect 7097 15542 18755 15544
rect 7097 15539 7163 15542
rect 18689 15539 18755 15542
rect 6177 15466 6243 15469
rect 18229 15466 18295 15469
rect 6177 15464 18295 15466
rect 6177 15408 6182 15464
rect 6238 15408 18234 15464
rect 18290 15408 18295 15464
rect 6177 15406 18295 15408
rect 6177 15403 6243 15406
rect 18229 15403 18295 15406
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 0 14696 480 14816
rect 10277 14720 10597 14721
rect 62 14242 122 14696
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 3969 14242 4035 14245
rect 62 14240 4035 14242
rect 62 14184 3974 14240
rect 4030 14184 4035 14240
rect 62 14182 4035 14184
rect 3969 14179 4035 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 4245 13698 4311 13701
rect 9305 13698 9371 13701
rect 4245 13696 9371 13698
rect 4245 13640 4250 13696
rect 4306 13640 9310 13696
rect 9366 13640 9371 13696
rect 4245 13638 9371 13640
rect 4245 13635 4311 13638
rect 9305 13635 9371 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 0 13200 480 13320
rect 5165 13290 5231 13293
rect 15653 13290 15719 13293
rect 5165 13288 15719 13290
rect 5165 13232 5170 13288
rect 5226 13232 15658 13288
rect 15714 13232 15719 13288
rect 5165 13230 15719 13232
rect 5165 13227 5231 13230
rect 15653 13227 15719 13230
rect 62 12746 122 13200
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 9029 13018 9095 13021
rect 13261 13018 13327 13021
rect 14733 13018 14799 13021
rect 9029 13016 14799 13018
rect 9029 12960 9034 13016
rect 9090 12960 13266 13016
rect 13322 12960 14738 13016
rect 14794 12960 14799 13016
rect 9029 12958 14799 12960
rect 9029 12955 9095 12958
rect 13261 12955 13327 12958
rect 14733 12955 14799 12958
rect 1393 12746 1459 12749
rect 62 12744 1459 12746
rect 62 12688 1398 12744
rect 1454 12688 1459 12744
rect 62 12686 1459 12688
rect 1393 12683 1459 12686
rect 8017 12746 8083 12749
rect 19517 12746 19583 12749
rect 8017 12744 19583 12746
rect 8017 12688 8022 12744
rect 8078 12688 19522 12744
rect 19578 12688 19583 12744
rect 8017 12686 19583 12688
rect 8017 12683 8083 12686
rect 19517 12683 19583 12686
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 5610 12000 5930 12001
rect 0 11840 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 62 11114 122 11840
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 17033 11114 17099 11117
rect 62 11112 17099 11114
rect 62 11056 17038 11112
rect 17094 11056 17099 11112
rect 62 11054 17099 11056
rect 17033 11051 17099 11054
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 6821 10706 6887 10709
rect 14089 10706 14155 10709
rect 6821 10704 14155 10706
rect 6821 10648 6826 10704
rect 6882 10648 14094 10704
rect 14150 10648 14155 10704
rect 6821 10646 14155 10648
rect 6821 10643 6887 10646
rect 14089 10643 14155 10646
rect 0 10480 480 10600
rect 62 10026 122 10480
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 5349 10162 5415 10165
rect 17493 10162 17559 10165
rect 5349 10160 17559 10162
rect 5349 10104 5354 10160
rect 5410 10104 17498 10160
rect 17554 10104 17559 10160
rect 5349 10102 17559 10104
rect 5349 10099 5415 10102
rect 17493 10099 17559 10102
rect 15745 10026 15811 10029
rect 62 10024 15811 10026
rect 62 9968 15750 10024
rect 15806 9968 15811 10024
rect 62 9966 15811 9968
rect 15745 9963 15811 9966
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 0 8984 480 9104
rect 62 8530 122 8984
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 6177 8530 6243 8533
rect 62 8528 6243 8530
rect 62 8472 6182 8528
rect 6238 8472 6243 8528
rect 62 8470 6243 8472
rect 6177 8467 6243 8470
rect 2313 8394 2379 8397
rect 11237 8394 11303 8397
rect 2313 8392 11303 8394
rect 2313 8336 2318 8392
rect 2374 8336 11242 8392
rect 11298 8336 11303 8392
rect 2313 8334 11303 8336
rect 2313 8331 2379 8334
rect 11237 8331 11303 8334
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 0 7624 480 7744
rect 5610 7648 5930 7649
rect 62 7306 122 7624
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 15837 7306 15903 7309
rect 62 7304 15903 7306
rect 62 7248 15842 7304
rect 15898 7248 15903 7304
rect 62 7246 15903 7248
rect 15837 7243 15903 7246
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 0 6264 480 6384
rect 4245 6354 4311 6357
rect 15561 6354 15627 6357
rect 4245 6352 15627 6354
rect 4245 6296 4250 6352
rect 4306 6296 15566 6352
rect 15622 6296 15627 6352
rect 4245 6294 15627 6296
rect 4245 6291 4311 6294
rect 15561 6291 15627 6294
rect 62 5674 122 6264
rect 6085 6218 6151 6221
rect 17953 6218 18019 6221
rect 6085 6216 18019 6218
rect 6085 6160 6090 6216
rect 6146 6160 17958 6216
rect 18014 6160 18019 6216
rect 6085 6158 18019 6160
rect 6085 6155 6151 6158
rect 17953 6155 18019 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 16849 5674 16915 5677
rect 62 5672 16915 5674
rect 62 5616 16854 5672
rect 16910 5616 16915 5672
rect 62 5614 16915 5616
rect 16849 5611 16915 5614
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 7465 5266 7531 5269
rect 62 5264 7531 5266
rect 62 5208 7470 5264
rect 7526 5208 7531 5264
rect 62 5206 7531 5208
rect 62 4888 122 5206
rect 7465 5203 7531 5206
rect 7833 5130 7899 5133
rect 14641 5130 14707 5133
rect 7833 5128 14707 5130
rect 7833 5072 7838 5128
rect 7894 5072 14646 5128
rect 14702 5072 14707 5128
rect 7833 5070 14707 5072
rect 7833 5067 7899 5070
rect 14641 5067 14707 5070
rect 10277 4928 10597 4929
rect 0 4768 480 4888
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 6269 3634 6335 3637
rect 15285 3634 15351 3637
rect 6269 3632 15351 3634
rect 6269 3576 6274 3632
rect 6330 3576 15290 3632
rect 15346 3576 15351 3632
rect 6269 3574 15351 3576
rect 6269 3571 6335 3574
rect 15285 3571 15351 3574
rect 0 3408 480 3528
rect 5809 3498 5875 3501
rect 12249 3498 12315 3501
rect 5809 3496 12315 3498
rect 5809 3440 5814 3496
rect 5870 3440 12254 3496
rect 12310 3440 12315 3496
rect 5809 3438 12315 3440
rect 5809 3435 5875 3438
rect 12249 3435 12315 3438
rect 16021 3498 16087 3501
rect 24209 3498 24275 3501
rect 16021 3496 24275 3498
rect 16021 3440 16026 3496
rect 16082 3440 24214 3496
rect 24270 3440 24275 3496
rect 16021 3438 24275 3440
rect 16021 3435 16087 3438
rect 24209 3435 24275 3438
rect 62 3090 122 3408
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 17309 3090 17375 3093
rect 62 3088 17375 3090
rect 62 3032 17314 3088
rect 17370 3032 17375 3088
rect 62 3030 17375 3032
rect 17309 3027 17375 3030
rect 8937 2954 9003 2957
rect 22369 2954 22435 2957
rect 8937 2952 22435 2954
rect 8937 2896 8942 2952
rect 8998 2896 22374 2952
rect 22430 2896 22435 2952
rect 8937 2894 22435 2896
rect 8937 2891 9003 2894
rect 22369 2891 22435 2894
rect 7097 2818 7163 2821
rect 8569 2818 8635 2821
rect 7097 2816 8635 2818
rect 7097 2760 7102 2816
rect 7158 2760 8574 2816
rect 8630 2760 8635 2816
rect 7097 2758 8635 2760
rect 7097 2755 7163 2758
rect 8569 2755 8635 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 4061 2682 4127 2685
rect 62 2680 4127 2682
rect 62 2624 4066 2680
rect 4122 2624 4127 2680
rect 62 2622 4127 2624
rect 62 2168 122 2622
rect 4061 2619 4127 2622
rect 5165 2682 5231 2685
rect 9489 2682 9555 2685
rect 5165 2680 9555 2682
rect 5165 2624 5170 2680
rect 5226 2624 9494 2680
rect 9550 2624 9555 2680
rect 5165 2622 9555 2624
rect 5165 2619 5231 2622
rect 9489 2619 9555 2622
rect 11605 2410 11671 2413
rect 26141 2410 26207 2413
rect 11605 2408 26207 2410
rect 11605 2352 11610 2408
rect 11666 2352 26146 2408
rect 26202 2352 26207 2408
rect 11605 2350 26207 2352
rect 11605 2347 11671 2350
rect 26141 2347 26207 2350
rect 5610 2208 5930 2209
rect 0 2048 480 2168
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 6637 2002 6703 2005
rect 20437 2002 20503 2005
rect 6637 2000 20503 2002
rect 6637 1944 6642 2000
rect 6698 1944 20442 2000
rect 20498 1944 20503 2000
rect 6637 1942 20503 1944
rect 6637 1939 6703 1942
rect 20437 1939 20503 1942
rect 5165 1594 5231 1597
rect 14549 1594 14615 1597
rect 5165 1592 14615 1594
rect 5165 1536 5170 1592
rect 5226 1536 14554 1592
rect 14610 1536 14615 1592
rect 5165 1534 14615 1536
rect 5165 1531 5231 1534
rect 14549 1531 14615 1534
rect 6821 1322 6887 1325
rect 62 1320 6887 1322
rect 62 1264 6826 1320
rect 6882 1264 6887 1320
rect 62 1262 6887 1264
rect 62 808 122 1262
rect 6821 1259 6887 1262
rect 0 688 480 808
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 60 24516 124 24580
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 60 24244 124 24308
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 59 24580 125 24581
rect 59 24516 60 24580
rect 124 24516 125 24580
rect 59 24515 125 24516
rect 62 24309 122 24515
rect 59 24308 125 24309
rect 59 24244 60 24308
rect 124 24244 125 24308
rect 59 24243 125 24244
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_15 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_0_23 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_19 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2944 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_35
timestamp 1586364061
transform 1 0 4324 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_31
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_32 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_4  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_42
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_43
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_46
timestamp 1586364061
transform 1 0 5336 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_47
timestamp 1586364061
transform 1 0 5428 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_68
timestamp 1586364061
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7084 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6900 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_76
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_72
timestamp 1586364061
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_89
timestamp 1586364061
transform 1 0 9292 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_97
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_93
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _232_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_101
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_102
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_142
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_138
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_142
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_1  FILLER_1_146
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14352 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_158
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_162
timestamp 1586364061
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_169
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_165
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_173
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_187
timestamp 1586364061
transform 1 0 18308 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 18400 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_191
timestamp 1586364061
transform 1 0 18676 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_192
timestamp 1586364061
transform 1 0 18768 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 18952 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _237_
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 20056 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_204
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_198
timestamp 1586364061
transform 1 0 19320 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_202
timestamp 1586364061
transform 1 0 19688 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_214
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 20976 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _235_
timestamp 1586364061
transform 1 0 21252 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_227
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_223
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 21804 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _234_
timestamp 1586364061
transform 1 0 22356 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_230
timestamp 1586364061
transform 1 0 22264 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_218
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_0_239
timestamp 1586364061
transform 1 0 23092 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_235
timestamp 1586364061
transform 1 0 22724 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 22908 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_249
timestamp 1586364061
transform 1 0 24012 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_242
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_249 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_0_247
timestamp 1586364061
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _233_
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _231_
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_259
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_263
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_253
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_265
timestamp 1586364061
transform 1 0 25484 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4968 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5980 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_40
timestamp 1586364061
transform 1 0 4784 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_45
timestamp 1586364061
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_49
timestamp 1586364061
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_52
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_2  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_71
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10304 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_97
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_8  FILLER_2_111
timestamp 1586364061
transform 1 0 11316 0 -1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_128
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_132
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_151
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_180
timestamp 1586364061
transform 1 0 17664 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_184
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_197
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_213
timestamp 1586364061
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_47
timestamp 1586364061
transform 1 0 5428 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6992 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_66
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8924 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 8740 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_81
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_94
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_4_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_111
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_115
timestamp 1586364061
transform 1 0 11684 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_134
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_138
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_142
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_148
timestamp 1586364061
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17480 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_161
timestamp 1586364061
transform 1 0 15916 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_165
timestamp 1586364061
transform 1 0 16284 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_172
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_176
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_180
timestamp 1586364061
transform 1 0 17664 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_187
timestamp 1586364061
transform 1 0 18308 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_191
timestamp 1586364061
transform 1 0 18676 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_198
timestamp 1586364061
transform 1 0 19320 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_202
timestamp 1586364061
transform 1 0 19688 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_214
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_226
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_3_238
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 7544 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_62
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_66
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _160_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7912 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_72
timestamp 1586364061
transform 1 0 7728 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_83
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_87
timestamp 1586364061
transform 1 0 9108 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_104
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_4_108
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_116
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13708 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13524 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_133
timestamp 1586364061
transform 1 0 13340 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_140
timestamp 1586364061
transform 1 0 13984 0 -1 4896
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_152
timestamp 1586364061
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_165
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_12  FILLER_4_182
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_194
timestamp 1586364061
transform 1 0 18952 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 6256 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 6992 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_55
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_58
timestamp 1586364061
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_66
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9108 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_79
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_83
timestamp 1586364061
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_102
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_109
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_113
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_117
timestamp 1586364061
transform 1 0 11868 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_121
timestamp 1586364061
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_139
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_145
timestamp 1586364061
transform 1 0 14444 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_149
timestamp 1586364061
transform 1 0 14812 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_164
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_168
timestamp 1586364061
transform 1 0 16560 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 18492 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_187
timestamp 1586364061
transform 1 0 18308 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_191
timestamp 1586364061
transform 1 0 18676 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_195
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_207
timestamp 1586364061
transform 1 0 20148 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_219
timestamp 1586364061
transform 1 0 21252 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_231
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_243
timestamp 1586364061
transform 1 0 23460 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_67
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_69
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_65
timestamp 1586364061
transform 1 0 7084 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _208_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6992 0 1 5984
box -38 -48 314 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_89
timestamp 1586364061
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_84
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_88
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_101
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_105
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_110
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _207_
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_120
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_123
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_127
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_140
timestamp 1586364061
transform 1 0 13984 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_136
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_150
timestamp 1586364061
transform 1 0 14904 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_146
timestamp 1586364061
transform 1 0 14536 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_155
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 14352 0 1 5984
box -38 -48 1050 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_4  FILLER_6_167
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15916 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_176
timestamp 1586364061
transform 1 0 17296 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_172
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 17480 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_180
timestamp 1586364061
transform 1 0 17664 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_180
timestamp 1586364061
transform 1 0 17664 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_197
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_6_209
timestamp 1586364061
transform 1 0 20332 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_213
timestamp 1586364061
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_67
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_71
timestamp 1586364061
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_104
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 11960 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_114
timestamp 1586364061
transform 1 0 11592 0 -1 7072
box -38 -48 406 592
use scs8hd_conb_1  _209_
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 590 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 17020 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_165
timestamp 1586364061
transform 1 0 16284 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_182
timestamp 1586364061
transform 1 0 17848 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_194
timestamp 1586364061
transform 1 0 18952 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6992 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_67
timestamp 1586364061
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_84
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_88
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_101
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_105
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _138_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_109
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_140
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 314 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 14444 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_154
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_158
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_1  _156_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_50
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_54
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_65
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_69
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 9844 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_104
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_123
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_127
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_140
timestamp 1586364061
transform 1 0 13984 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_144
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_147
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_151
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_167
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_174
timestamp 1586364061
transform 1 0 17112 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_186
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_198
timestamp 1586364061
transform 1 0 19320 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_210
timestamp 1586364061
transform 1 0 20424 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_6
timestamp 1586364061
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_10
timestamp 1586364061
transform 1 0 2024 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_17
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_21
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_25
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_37
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_41
timestamp 1586364061
transform 1 0 4876 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_44
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_69
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_73
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_88
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 9936 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 9752 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_92
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_105
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_109
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 406 592
use scs8hd_decap_4  FILLER_11_115
timestamp 1586364061
transform 1 0 11684 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_119
timestamp 1586364061
transform 1 0 12052 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_136
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_140
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_155
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_166
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_170
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_173
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_181
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2668 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_9
timestamp 1586364061
transform 1 0 1932 0 -1 9248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_20
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_28
timestamp 1586364061
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4968 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_12_40
timestamp 1586364061
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_45
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_62
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_71
timestamp 1586364061
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 9936 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11500 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_109
timestamp 1586364061
transform 1 0 11132 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_112
timestamp 1586364061
transform 1 0 11408 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_124
timestamp 1586364061
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_128
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_132
timestamp 1586364061
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_143
timestamp 1586364061
transform 1 0 14260 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_147
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_174
timestamp 1586364061
transform 1 0 17112 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_198
timestamp 1586364061
transform 1 0 19320 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_6  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 590 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_9
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 2024 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 314 592
use scs8hd_inv_8  _192_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_19
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_26
timestamp 1586364061
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_30
timestamp 1586364061
transform 1 0 3864 0 1 9248
box -38 -48 590 592
use scs8hd_decap_8  FILLER_14_20
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_28
timestamp 1586364061
transform 1 0 3680 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_40
timestamp 1586364061
transform 1 0 4784 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_43
timestamp 1586364061
transform 1 0 5060 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_36
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 4508 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4876 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_48
timestamp 1586364061
transform 1 0 5520 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_61
timestamp 1586364061
transform 1 0 6716 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_69
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_70
timestamp 1586364061
transform 1 0 7544 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7268 0 1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8280 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7728 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_87
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_73
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_90
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_94
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_91
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_102
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_124
timestamp 1586364061
transform 1 0 12512 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_119
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12328 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_132
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_128
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_138
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_157
timestamp 1586364061
transform 1 0 15548 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_4  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_155
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_14_168
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_166
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16100 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_178
timestamp 1586364061
transform 1 0 17480 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_174
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_170
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _148_
timestamp 1586364061
transform 1 0 17296 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_182
timestamp 1586364061
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_187
timestamp 1586364061
transform 1 0 18308 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_191
timestamp 1586364061
transform 1 0 18676 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_179
timestamp 1586364061
transform 1 0 17572 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_191
timestamp 1586364061
transform 1 0 18676 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_203
timestamp 1586364061
transform 1 0 19780 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_203
timestamp 1586364061
transform 1 0 19780 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_211
timestamp 1586364061
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_215
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_227
timestamp 1586364061
transform 1 0 21988 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_239
timestamp 1586364061
transform 1 0 23092 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_243
timestamp 1586364061
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_conb_1  _215_
timestamp 1586364061
transform 1 0 1472 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2024 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_12
timestamp 1586364061
transform 1 0 2208 0 1 10336
box -38 -48 314 592
use scs8hd_conb_1  _219_
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_24
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_28
timestamp 1586364061
transform 1 0 3680 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_32
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_40
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_67
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_80
timestamp 1586364061
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_84
timestamp 1586364061
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_97
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_103
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13708 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_139
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_152
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _137_
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16284 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 17296 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_163
timestamp 1586364061
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_167
timestamp 1586364061
transform 1 0 16468 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_174
timestamp 1586364061
transform 1 0 17112 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_178
timestamp 1586364061
transform 1 0 17480 0 1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_182
timestamp 1586364061
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_19
timestamp 1586364061
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_41
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_46
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_50
timestamp 1586364061
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_16_62
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_81
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_85
timestamp 1586364061
transform 1 0 8924 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_89
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 10396 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_112
timestamp 1586364061
transform 1 0 11408 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_116
timestamp 1586364061
transform 1 0 11776 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_122
timestamp 1586364061
transform 1 0 12328 0 -1 11424
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_134
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_149
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use scs8hd_conb_1  _220_
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_16_174
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_198
timestamp 1586364061
transform 1 0 19320 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_13
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_17
timestamp 1586364061
transform 1 0 2668 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3036 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_30
timestamp 1586364061
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_34
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_40
timestamp 1586364061
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 590 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_79
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_91
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_95
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_134
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_138
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_142
timestamp 1586364061
transform 1 0 14168 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_146
timestamp 1586364061
transform 1 0 14536 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_160
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_164
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_30
timestamp 1586364061
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_35
timestamp 1586364061
transform 1 0 4324 0 -1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 4968 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__D
timestamp 1586364061
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_40
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 6900 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_55
timestamp 1586364061
transform 1 0 6164 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_6  FILLER_18_65
timestamp 1586364061
transform 1 0 7084 0 -1 12512
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_101
timestamp 1586364061
transform 1 0 10396 0 -1 12512
box -38 -48 222 592
use scs8hd_or2_4  _136_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12144 0 -1 12512
box -38 -48 682 592
use scs8hd_decap_8  FILLER_18_112
timestamp 1586364061
transform 1 0 11408 0 -1 12512
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_127
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_131
timestamp 1586364061
transform 1 0 13156 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_135
timestamp 1586364061
transform 1 0 13524 0 -1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_151
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _099_
timestamp 1586364061
transform 1 0 17020 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_18_165
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_182
timestamp 1586364061
transform 1 0 17848 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_194
timestamp 1586364061
transform 1 0 18952 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_11
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 866 592
use scs8hd_inv_8  _189_
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_25
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_21
timestamp 1586364061
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_22
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_18
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_35
timestamp 1586364061
transform 1 0 4324 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__D
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_20_39
timestamp 1586364061
transform 1 0 4692 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_43
timestamp 1586364061
transform 1 0 5060 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 4968 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 4508 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_50
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 5244 0 1 12512
box -38 -48 222 592
use scs8hd_conb_1  _216_
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 314 592
use scs8hd_nor4_4  _169_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_20_61
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_58
timestamp 1586364061
transform 1 0 6440 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_54
timestamp 1586364061
transform 1 0 6072 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_69
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_65
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 6900 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_76
timestamp 1586364061
transform 1 0 8096 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_72
timestamp 1586364061
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_89
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_86
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_82
timestamp 1586364061
transform 1 0 8648 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8464 0 1 12512
box -38 -48 1050 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_95
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_91
timestamp 1586364061
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_20_107
timestamp 1586364061
transform 1 0 10948 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_19_99
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12144 0 -1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_113
timestamp 1586364061
transform 1 0 11500 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_116
timestamp 1586364061
transform 1 0 11776 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_131
timestamp 1586364061
transform 1 0 13156 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_127
timestamp 1586364061
transform 1 0 12788 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_142
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_135
timestamp 1586364061
transform 1 0 13524 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_139
timestamp 1586364061
transform 1 0 13892 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13892 0 -1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_20_150
timestamp 1586364061
transform 1 0 14904 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_150
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_143
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_167
timestamp 1586364061
transform 1 0 16468 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_167
timestamp 1586364061
transform 1 0 16468 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_163
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_177
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_173
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_192
timestamp 1586364061
transform 1 0 18768 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_204
timestamp 1586364061
transform 1 0 19872 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_212
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_263
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_13
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_17
timestamp 1586364061
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 3036 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_25
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_31
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_35
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 130 592
use scs8hd_nor4_4  _170_
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_nor4_4  _174_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__174__C
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_79
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_83
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use scs8hd_or2_4  _093_
timestamp 1586364061
transform 1 0 10856 0 1 13600
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_98
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_102
timestamp 1586364061
transform 1 0 10488 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 11684 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_113
timestamp 1586364061
transform 1 0 11500 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_117
timestamp 1586364061
transform 1 0 11868 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_134
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_138
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_153
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_157
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_170
timestamp 1586364061
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_174
timestamp 1586364061
transform 1 0 17112 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_182
timestamp 1586364061
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_1  _094_
timestamp 1586364061
transform 1 0 4140 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__168__D
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_20
timestamp 1586364061
transform 1 0 2944 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_24
timestamp 1586364061
transform 1 0 3312 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_28
timestamp 1586364061
transform 1 0 3680 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 130 592
use scs8hd_nor4_4  _168_
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 4600 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 4968 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_36
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_40
timestamp 1586364061
transform 1 0 4784 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__D
timestamp 1586364061
transform 1 0 6900 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_61
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_65
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_69
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_73
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_106
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 866 592
use scs8hd_fill_2  FILLER_22_123
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_127
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_140
timestamp 1586364061
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_144
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_148
timestamp 1586364061
transform 1 0 14720 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_152
timestamp 1586364061
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_165
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_177
timestamp 1586364061
transform 1 0 17388 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_189
timestamp 1586364061
transform 1 0 18492 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_201
timestamp 1586364061
transform 1 0 19596 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_213
timestamp 1586364061
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_13
timestamp 1586364061
transform 1 0 2300 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_17
timestamp 1586364061
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3036 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_32
timestamp 1586364061
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_36
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use scs8hd_nor4_4  _175_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__175__C
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_55
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_79
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_83
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_87
timestamp 1586364061
transform 1 0 9108 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_91
timestamp 1586364061
transform 1 0 9476 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_103
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_107
timestamp 1586364061
transform 1 0 10948 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _088_
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 314 592
use scs8hd_buf_1  _127_
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 12880 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_126
timestamp 1586364061
transform 1 0 12696 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_130
timestamp 1586364061
transform 1 0 13064 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_134
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15088 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_144
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_148
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_161
timestamp 1586364061
transform 1 0 15916 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_165
timestamp 1586364061
transform 1 0 16284 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_169
timestamp 1586364061
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_173
timestamp 1586364061
transform 1 0 17020 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_177
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18216 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_188
timestamp 1586364061
transform 1 0 18400 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_200
timestamp 1586364061
transform 1 0 19504 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_212
timestamp 1586364061
transform 1 0 20608 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_224
timestamp 1586364061
transform 1 0 21712 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_23_236
timestamp 1586364061
transform 1 0 22816 0 1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_13
timestamp 1586364061
transform 1 0 2300 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_17
timestamp 1586364061
transform 1 0 2668 0 -1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3036 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_35
timestamp 1586364061
transform 1 0 4324 0 -1 15776
box -38 -48 314 592
use scs8hd_nor4_4  _166_
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 4968 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_40
timestamp 1586364061
transform 1 0 4784 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__D
timestamp 1586364061
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_61
timestamp 1586364061
transform 1 0 6716 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_65
timestamp 1586364061
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_69
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_2  FILLER_24_73
timestamp 1586364061
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 774 592
use scs8hd_buf_1  _105_
timestamp 1586364061
transform 1 0 11500 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 11960 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_110
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_116
timestamp 1586364061
transform 1 0 11776 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_120
timestamp 1586364061
transform 1 0 12144 0 -1 15776
box -38 -48 406 592
use scs8hd_buf_1  _117_
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13892 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_133
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_137
timestamp 1586364061
transform 1 0 13708 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_144
timestamp 1586364061
transform 1 0 14352 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_152
timestamp 1586364061
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_24_174
timestamp 1586364061
transform 1 0 17112 0 -1 15776
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_189
timestamp 1586364061
transform 1 0 18492 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_201
timestamp 1586364061
transform 1 0 19596 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_213
timestamp 1586364061
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_12
timestamp 1586364061
transform 1 0 2208 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_16
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_29
timestamp 1586364061
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_33
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use scs8hd_inv_8  _198_
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5612 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_46
timestamp 1586364061
transform 1 0 5336 0 1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__C
timestamp 1586364061
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__D
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_66
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_82
timestamp 1586364061
transform 1 0 8648 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use scs8hd_or2_4  _126_
timestamp 1586364061
transform 1 0 10948 0 1 15776
box -38 -48 682 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_99
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_103
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 13156 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 12972 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 12604 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_127
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_140
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15180 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_144
timestamp 1586364061
transform 1 0 14352 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_149
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 222 592
use scs8hd_buf_1  _144_
timestamp 1586364061
transform 1 0 16744 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_162
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_166
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_173
timestamp 1586364061
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_177
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 590 592
use scs8hd_buf_1  _164_
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 18492 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_187
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_191
timestamp 1586364061
transform 1 0 18676 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_195
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_207
timestamp 1586364061
transform 1 0 20148 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_219
timestamp 1586364061
transform 1 0 21252 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_231
timestamp 1586364061
transform 1 0 22356 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_243
timestamp 1586364061
transform 1 0 23460 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _230_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_27_14
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_11
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_16
timestamp 1586364061
transform 1 0 2576 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_12
timestamp 1586364061
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2392 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2760 0 -1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_32
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_28
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__D
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__C
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use scs8hd_nor4_4  _178_
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 1602 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__179__C
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_46
timestamp 1586364061
transform 1 0 5336 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_52
timestamp 1586364061
transform 1 0 5888 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_nor4_4  _176_
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1602 592
use scs8hd_nor4_4  _177_
timestamp 1586364061
transform 1 0 6624 0 -1 16864
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__176__C
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__D
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 6072 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__B
timestamp 1586364061
transform 1 0 6440 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_79
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_77
timestamp 1586364061
transform 1 0 8188 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 8372 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_83
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_89
timestamp 1586364061
transform 1 0 9292 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_85
timestamp 1586364061
transform 1 0 8924 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_81
timestamp 1586364061
transform 1 0 8556 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_96
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_100
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_106
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__C
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 10488 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_or3_4  _155_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10672 0 1 16864
box -38 -48 866 592
use scs8hd_decap_3  FILLER_27_113
timestamp 1586364061
transform 1 0 11500 0 1 16864
box -38 -48 314 592
use scs8hd_decap_6  FILLER_26_110
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_116
timestamp 1586364061
transform 1 0 11776 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_or2_4  _116_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 682 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13892 0 1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 13340 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_126
timestamp 1586364061
transform 1 0 12696 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_130
timestamp 1586364061
transform 1 0 13064 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_27_130
timestamp 1586364061
transform 1 0 13064 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_150
timestamp 1586364061
transform 1 0 14904 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_149
timestamp 1586364061
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_154
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 15088 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_167
timestamp 1586364061
transform 1 0 16468 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_167
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_174
timestamp 1586364061
transform 1 0 17112 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17480 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _221_
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_187
timestamp 1586364061
transform 1 0 18308 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_180
timestamp 1586364061
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_buf_1  _173_
timestamp 1586364061
transform 1 0 17848 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_1  _146_
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_191
timestamp 1586364061
transform 1 0 18676 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 18492 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_195
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_185
timestamp 1586364061
transform 1 0 18124 0 -1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_197
timestamp 1586364061
transform 1 0 19228 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_26_209
timestamp 1586364061
transform 1 0 20332 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_213
timestamp 1586364061
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_207
timestamp 1586364061
transform 1 0 20148 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_219
timestamp 1586364061
transform 1 0 21252 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_231
timestamp 1586364061
transform 1 0 22356 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_243
timestamp 1586364061
transform 1 0 23460 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 1050 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 1932 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_11
timestamp 1586364061
transform 1 0 2116 0 -1 17952
box -38 -48 130 592
use scs8hd_buf_2  _228_
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__178__B
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use scs8hd_nor4_4  _179_
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__181__D
timestamp 1586364061
transform 1 0 4968 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__D
timestamp 1586364061
transform 1 0 4600 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_36
timestamp 1586364061
transform 1 0 4416 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_40
timestamp 1586364061
transform 1 0 4784 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_61
timestamp 1586364061
transform 1 0 6716 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_67
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_71
timestamp 1586364061
transform 1 0 7636 0 -1 17952
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7728 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 8924 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_83
timestamp 1586364061
transform 1 0 8740 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_87
timestamp 1586364061
transform 1 0 9108 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_8  _145_
timestamp 1586364061
transform 1 0 10120 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__C
timestamp 1586364061
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_97
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_107
timestamp 1586364061
transform 1 0 10948 0 -1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 12052 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 11316 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_113
timestamp 1586364061
transform 1 0 11500 0 -1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_128
timestamp 1586364061
transform 1 0 12880 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_133
timestamp 1586364061
transform 1 0 13340 0 -1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15732 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_4  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_158
timestamp 1586364061
transform 1 0 15640 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 16928 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_170
timestamp 1586364061
transform 1 0 16744 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_174
timestamp 1586364061
transform 1 0 17112 0 -1 17952
box -38 -48 406 592
use scs8hd_buf_1  _172_
timestamp 1586364061
transform 1 0 18492 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_181
timestamp 1586364061
transform 1 0 17756 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_12  FILLER_28_192
timestamp 1586364061
transform 1 0 18768 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_204
timestamp 1586364061
transform 1 0 19872 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_212
timestamp 1586364061
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_12
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_16
timestamp 1586364061
transform 1 0 2576 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3312 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2760 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_20
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_35
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 314 592
use scs8hd_inv_8  _171_
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__181__B
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__C
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_40
timestamp 1586364061
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_or3_4  _101_
timestamp 1586364061
transform 1 0 7084 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_78
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_91
timestamp 1586364061
transform 1 0 9476 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_96
timestamp 1586364061
transform 1 0 9936 0 1 17952
box -38 -48 314 592
use scs8hd_or2_4  _089_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 11684 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_108
timestamp 1586364061
transform 1 0 11040 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_113
timestamp 1586364061
transform 1 0 11500 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_117
timestamp 1586364061
transform 1 0 11868 0 1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 13892 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_130
timestamp 1586364061
transform 1 0 13064 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_134
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_150
timestamp 1586364061
transform 1 0 14904 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_156
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_160
timestamp 1586364061
transform 1 0 15824 0 1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 18400 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 406 592
use scs8hd_decap_4  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_29_190
timestamp 1586364061
transform 1 0 18584 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_202
timestamp 1586364061
transform 1 0 19688 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_214
timestamp 1586364061
transform 1 0 20792 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_226
timestamp 1586364061
transform 1 0 21896 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_29_238
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 590 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3036 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_19
timestamp 1586364061
transform 1 0 2852 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_35
timestamp 1586364061
transform 1 0 4324 0 -1 19040
box -38 -48 222 592
use scs8hd_nor4_4  _181_
timestamp 1586364061
transform 1 0 5060 0 -1 19040
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_39
timestamp 1586364061
transform 1 0 4692 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__C
timestamp 1586364061
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__B
timestamp 1586364061
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_60
timestamp 1586364061
transform 1 0 6624 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_64
timestamp 1586364061
transform 1 0 6992 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_67
timestamp 1586364061
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_71
timestamp 1586364061
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 8004 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_88
timestamp 1586364061
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use scs8hd_or3_4  _097_
timestamp 1586364061
transform 1 0 9752 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_103
timestamp 1586364061
transform 1 0 10580 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_107
timestamp 1586364061
transform 1 0 10948 0 -1 19040
box -38 -48 222 592
use scs8hd_or3_4  _104_
timestamp 1586364061
transform 1 0 11316 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 11132 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_120
timestamp 1586364061
transform 1 0 12144 0 -1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 13156 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_125
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_140
timestamp 1586364061
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_144
timestamp 1586364061
transform 1 0 14352 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_152
timestamp 1586364061
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 16836 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_163
timestamp 1586364061
transform 1 0 16100 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_168
timestamp 1586364061
transform 1 0 16560 0 -1 19040
box -38 -48 314 592
use scs8hd_buf_1  _165_
timestamp 1586364061
transform 1 0 18400 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 18032 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_180
timestamp 1586364061
transform 1 0 17664 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_186
timestamp 1586364061
transform 1 0 18216 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_191
timestamp 1586364061
transform 1 0 18676 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_203
timestamp 1586364061
transform 1 0 19780 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_211
timestamp 1586364061
transform 1 0 20516 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_inv_8  _197_
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_12
timestamp 1586364061
transform 1 0 2208 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_16
timestamp 1586364061
transform 1 0 2576 0 1 19040
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3036 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 4232 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_32
timestamp 1586364061
transform 1 0 4048 0 1 19040
box -38 -48 222 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__188__B
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__C
timestamp 1586364061
transform 1 0 5428 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_36
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_44
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_49
timestamp 1586364061
transform 1 0 5612 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_nor4_4  _187_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__187__D
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__D
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_inv_8  _084_
timestamp 1586364061
transform 1 0 9200 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_79
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_83
timestamp 1586364061
transform 1 0 8740 0 1 19040
box -38 -48 314 592
use scs8hd_or3_4  _147_
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__C
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_97
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_101
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use scs8hd_or3_4  _107_
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_buf_1  _108_
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_132
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_136
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15456 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 14444 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 14812 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_143
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_151
timestamp 1586364061
transform 1 0 14996 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_167
timestamp 1586364061
transform 1 0 16468 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_193
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_197
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_209
timestamp 1586364061
transform 1 0 20332 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_221
timestamp 1586364061
transform 1 0 21436 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_233
timestamp 1586364061
transform 1 0 22540 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_31_241
timestamp 1586364061
transform 1 0 23276 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_inv_8  _199_
timestamp 1586364061
transform 1 0 1564 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2576 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_14
timestamp 1586364061
transform 1 0 2392 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 2944 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_18
timestamp 1586364061
transform 1 0 2760 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_22
timestamp 1586364061
transform 1 0 3128 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_26
timestamp 1586364061
transform 1 0 3496 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__187__C
timestamp 1586364061
transform 1 0 5980 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__D
timestamp 1586364061
transform 1 0 5060 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 5612 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_41
timestamp 1586364061
transform 1 0 4876 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_45
timestamp 1586364061
transform 1 0 5244 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_51
timestamp 1586364061
transform 1 0 5796 0 -1 20128
box -38 -48 222 592
use scs8hd_nor4_4  _188_
timestamp 1586364061
transform 1 0 6164 0 -1 20128
box -38 -48 1602 592
use scs8hd_buf_1  _102_
timestamp 1586364061
transform 1 0 8556 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__185__C
timestamp 1586364061
transform 1 0 7912 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__B
timestamp 1586364061
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 8280 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_72
timestamp 1586364061
transform 1 0 7728 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_76
timestamp 1586364061
transform 1 0 8096 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_88
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use scs8hd_or3_4  _087_
timestamp 1586364061
transform 1 0 9936 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__147__C
timestamp 1586364061
transform 1 0 10948 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__D
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_8  _085_
timestamp 1586364061
transform 1 0 11500 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__107__C
timestamp 1586364061
transform 1 0 12512 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 11316 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_109
timestamp 1586364061
transform 1 0 11132 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_122
timestamp 1586364061
transform 1 0 12328 0 -1 20128
box -38 -48 222 592
use scs8hd_or3_4  _110_
timestamp 1586364061
transform 1 0 13064 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_126
timestamp 1586364061
transform 1 0 12696 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_139
timestamp 1586364061
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14904 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_143
timestamp 1586364061
transform 1 0 14260 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_149
timestamp 1586364061
transform 1 0 14812 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_158
timestamp 1586364061
transform 1 0 15640 0 -1 20128
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_173
timestamp 1586364061
transform 1 0 17020 0 -1 20128
box -38 -48 774 592
use scs8hd_buf_1  _111_
timestamp 1586364061
transform 1 0 17756 0 -1 20128
box -38 -48 314 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 18768 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_184
timestamp 1586364061
transform 1 0 18032 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_32_195
timestamp 1586364061
transform 1 0 19044 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_32_207
timestamp 1586364061
transform 1 0 20148 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_213
timestamp 1586364061
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_34_7
timestamp 1586364061
transform 1 0 1748 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_6
timestamp 1586364061
transform 1 0 1656 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_10
timestamp 1586364061
transform 1 0 2024 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2024 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2208 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 -1 21216
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2392 0 1 20128
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_34_25
timestamp 1586364061
transform 1 0 3404 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_21
timestamp 1586364061
transform 1 0 3036 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_25
timestamp 1586364061
transform 1 0 3404 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_32
timestamp 1586364061
transform 1 0 4048 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_29
timestamp 1586364061
transform 1 0 3772 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__C
timestamp 1586364061
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__B
timestamp 1586364061
transform 1 0 4232 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 866 592
use scs8hd_nor4_4  _182_
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 1602 592
use scs8hd_conb_1  _217_
timestamp 1586364061
transform 1 0 5612 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 5060 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_41
timestamp 1586364061
transform 1 0 4876 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_45
timestamp 1586364061
transform 1 0 5244 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_52
timestamp 1586364061
transform 1 0 5888 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 6072 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__B
timestamp 1586364061
transform 1 0 6440 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__C
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__D
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__185__D
timestamp 1586364061
transform 1 0 7176 0 1 20128
box -38 -48 222 592
use scs8hd_nor4_4  _186_
timestamp 1586364061
transform 1 0 6624 0 -1 21216
box -38 -48 1602 592
use scs8hd_nor4_4  _185_
timestamp 1586364061
transform 1 0 7360 0 1 20128
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__184__C
timestamp 1586364061
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_85
timestamp 1586364061
transform 1 0 8924 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_89
timestamp 1586364061
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_77
timestamp 1586364061
transform 1 0 8188 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_85
timestamp 1586364061
transform 1 0 8924 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_88
timestamp 1586364061
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use scs8hd_nor4_4  _183_
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1602 592
use scs8hd_nor4_4  _184_
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__183__D
timestamp 1586364061
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__B
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_114
timestamp 1586364061
transform 1 0 11592 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_110
timestamp 1586364061
transform 1 0 11224 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 11408 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__C
timestamp 1586364061
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_120
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_inv_8  _100_
timestamp 1586364061
transform 1 0 11960 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_131
timestamp 1586364061
transform 1 0 13156 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_127
timestamp 1586364061
transform 1 0 12788 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_129
timestamp 1586364061
transform 1 0 12972 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13156 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 13340 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_135
timestamp 1586364061
transform 1 0 13524 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_142
timestamp 1586364061
transform 1 0 14168 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_8  FILLER_34_145
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_146
timestamp 1586364061
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_158
timestamp 1586364061
transform 1 0 15640 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 -1 21216
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 14904 0 1 20128
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_34_168
timestamp 1586364061
transform 1 0 16560 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_165
timestamp 1586364061
transform 1 0 16284 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_161
timestamp 1586364061
transform 1 0 15916 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_176
timestamp 1586364061
transform 1 0 17296 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_172
timestamp 1586364061
transform 1 0 16928 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17480 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17296 0 -1 21216
box -38 -48 314 592
use scs8hd_buf_1  _163_
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 18492 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_180
timestamp 1586364061
transform 1 0 17664 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_187
timestamp 1586364061
transform 1 0 18308 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_191
timestamp 1586364061
transform 1 0 18676 0 1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_179
timestamp 1586364061
transform 1 0 17572 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_191
timestamp 1586364061
transform 1 0 18676 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_198
timestamp 1586364061
transform 1 0 19320 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_202
timestamp 1586364061
transform 1 0 19688 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_214
timestamp 1586364061
transform 1 0 20792 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_203
timestamp 1586364061
transform 1 0 19780 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_34_211
timestamp 1586364061
transform 1 0 20516 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_226
timestamp 1586364061
transform 1 0 21896 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_33_238
timestamp 1586364061
transform 1 0 23000 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 866 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2392 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_12
timestamp 1586364061
transform 1 0 2208 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_16
timestamp 1586364061
transform 1 0 2576 0 1 21216
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3128 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 4140 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_31
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_35
timestamp 1586364061
transform 1 0 4324 0 1 21216
box -38 -48 222 592
use scs8hd_inv_8  _206_
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4508 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5704 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_48
timestamp 1586364061
transform 1 0 5520 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_52
timestamp 1586364061
transform 1 0 5888 0 1 21216
box -38 -48 590 592
use scs8hd_buf_1  _092_
timestamp 1586364061
transform 1 0 7544 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__B
timestamp 1586364061
transform 1 0 7360 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_58
timestamp 1586364061
transform 1 0 6440 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_66
timestamp 1586364061
transform 1 0 7176 0 1 21216
box -38 -48 222 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 8556 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_73
timestamp 1586364061
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_77
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_84
timestamp 1586364061
transform 1 0 8832 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_88
timestamp 1586364061
transform 1 0 9200 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9568 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_103
timestamp 1586364061
transform 1 0 10580 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_107
timestamp 1586364061
transform 1 0 10948 0 1 21216
box -38 -48 222 592
use scs8hd_buf_1  _086_
timestamp 1586364061
transform 1 0 11316 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_114
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13064 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_128
timestamp 1586364061
transform 1 0 12880 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_132
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15180 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_145
timestamp 1586364061
transform 1 0 14444 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_149
timestamp 1586364061
transform 1 0 14812 0 1 21216
box -38 -48 222 592
use scs8hd_buf_1  _135_
timestamp 1586364061
transform 1 0 16744 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_162
timestamp 1586364061
transform 1 0 16008 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_166
timestamp 1586364061
transform 1 0 16376 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_173
timestamp 1586364061
transform 1 0 17020 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_177
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_181
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _242_
timestamp 1586364061
transform 1 0 23920 0 1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 24472 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_252
timestamp 1586364061
transform 1 0 24288 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_256
timestamp 1586364061
transform 1 0 24656 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_268
timestamp 1586364061
transform 1 0 25760 0 1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_35_276
timestamp 1586364061
transform 1 0 26496 0 1 21216
box -38 -48 130 592
use scs8hd_conb_1  _211_
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 314 592
use scs8hd_buf_2  _225_
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__225__A
timestamp 1586364061
transform 1 0 1932 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_7
timestamp 1586364061
transform 1 0 1748 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_11
timestamp 1586364061
transform 1 0 2116 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4324 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_18
timestamp 1586364061
transform 1 0 2760 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_6  FILLER_36_24
timestamp 1586364061
transform 1 0 3312 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_30
timestamp 1586364061
transform 1 0 3864 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4508 0 -1 22304
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_36_48
timestamp 1586364061
transform 1 0 5520 0 -1 22304
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 22304
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6532 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_62
timestamp 1586364061
transform 1 0 6808 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_66
timestamp 1586364061
transform 1 0 7176 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_81
timestamp 1586364061
transform 1 0 8556 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_36_89
timestamp 1586364061
transform 1 0 9292 0 -1 22304
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_104
timestamp 1586364061
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use scs8hd_buf_1  _098_
timestamp 1586364061
transform 1 0 11500 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_108
timestamp 1586364061
transform 1 0 11040 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_112
timestamp 1586364061
transform 1 0 11408 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_116
timestamp 1586364061
transform 1 0 11776 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_120
timestamp 1586364061
transform 1 0 12144 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_124
timestamp 1586364061
transform 1 0 12512 0 -1 22304
box -38 -48 130 592
use scs8hd_or3_4  _134_
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_134
timestamp 1586364061
transform 1 0 13432 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_138
timestamp 1586364061
transform 1 0 13800 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_149
timestamp 1586364061
transform 1 0 14812 0 -1 22304
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17296 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_163
timestamp 1586364061
transform 1 0 16100 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_175
timestamp 1586364061
transform 1 0 17204 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_179
timestamp 1586364061
transform 1 0 17572 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_191
timestamp 1586364061
transform 1 0 18676 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_203
timestamp 1586364061
transform 1 0 19780 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  FILLER_36_211
timestamp 1586364061
transform 1 0 20516 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_buf_1  _180_
timestamp 1586364061
transform 1 0 2668 0 1 22304
box -38 -48 314 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 2392 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_11
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_37_16
timestamp 1586364061
transform 1 0 2576 0 1 22304
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3680 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 3128 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3496 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_20
timestamp 1586364061
transform 1 0 2944 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_24
timestamp 1586364061
transform 1 0 3312 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_31
timestamp 1586364061
transform 1 0 3956 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_35
timestamp 1586364061
transform 1 0 4324 0 1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4508 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_50
timestamp 1586364061
transform 1 0 5704 0 1 22304
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_54
timestamp 1586364061
transform 1 0 6072 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 8648 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 8464 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_73
timestamp 1586364061
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_77
timestamp 1586364061
transform 1 0 8188 0 1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_91
timestamp 1586364061
transform 1 0 9476 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_95
timestamp 1586364061
transform 1 0 9844 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_108
timestamp 1586364061
transform 1 0 11040 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_114
timestamp 1586364061
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_118
timestamp 1586364061
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 222 592
use scs8hd_or3_4  _114_
timestamp 1586364061
transform 1 0 12604 0 1 22304
box -38 -48 866 592
use scs8hd_or3_4  _125_
timestamp 1586364061
transform 1 0 14168 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 13984 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 13616 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_134
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_138
timestamp 1586364061
transform 1 0 13800 0 1 22304
box -38 -48 222 592
use scs8hd_buf_1  _115_
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_151
timestamp 1586364061
transform 1 0 14996 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_156
timestamp 1586364061
transform 1 0 15456 0 1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 16192 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_162
timestamp 1586364061
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_166
timestamp 1586364061
transform 1 0 16376 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_173
timestamp 1586364061
transform 1 0 17020 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_177
timestamp 1586364061
transform 1 0 17388 0 1 22304
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_buf_2  _244_
timestamp 1586364061
transform 1 0 22264 0 1 22304
box -38 -48 406 592
use scs8hd_decap_8  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_228
timestamp 1586364061
transform 1 0 22080 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__244__A
timestamp 1586364061
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_234
timestamp 1586364061
transform 1 0 22632 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_238
timestamp 1586364061
transform 1 0 23000 0 1 22304
box -38 -48 590 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_inv_8  _205_
timestamp 1586364061
transform 1 0 2392 0 -1 23392
box -38 -48 866 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_6
timestamp 1586364061
transform 1 0 1656 0 -1 23392
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_23
timestamp 1586364061
transform 1 0 3220 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_4  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4416 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_47
timestamp 1586364061
transform 1 0 5428 0 -1 23392
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 -1 23392
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6532 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_62
timestamp 1586364061
transform 1 0 6808 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_8  FILLER_38_79
timestamp 1586364061
transform 1 0 8372 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_38_87
timestamp 1586364061
transform 1 0 9108 0 -1 23392
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_97
timestamp 1586364061
transform 1 0 10028 0 -1 23392
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_38_109
timestamp 1586364061
transform 1 0 11132 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 13432 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__C
timestamp 1586364061
transform 1 0 12880 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_126
timestamp 1586364061
transform 1 0 12696 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_130
timestamp 1586364061
transform 1 0 13064 0 -1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__C
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_143
timestamp 1586364061
transform 1 0 14260 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_147
timestamp 1586364061
transform 1 0 14628 0 -1 23392
box -38 -48 590 592
use scs8hd_decap_12  FILLER_38_157
timestamp 1586364061
transform 1 0 15548 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_169
timestamp 1586364061
transform 1 0 16652 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_181
timestamp 1586364061
transform 1 0 17756 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_193
timestamp 1586364061
transform 1 0 18860 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_205
timestamp 1586364061
transform 1 0 19964 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_38_213
timestamp 1586364061
transform 1 0 20700 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_7
timestamp 1586364061
transform 1 0 1748 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_39_7
timestamp 1586364061
transform 1 0 1748 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__223__A
timestamp 1586364061
transform 1 0 1564 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_buf_2  _223_
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_17
timestamp 1586364061
transform 1 0 2668 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__222__A
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 314 592
use scs8hd_buf_2  _222_
timestamp 1586364061
transform 1 0 2300 0 1 23392
box -38 -48 406 592
use scs8hd_decap_6  FILLER_39_21
timestamp 1586364061
transform 1 0 3036 0 1 23392
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_30
timestamp 1586364061
transform 1 0 3864 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_29
timestamp 1586364061
transform 1 0 3772 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3956 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_18
timestamp 1586364061
transform 1 0 2760 0 -1 24480
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 1 23392
box -38 -48 866 592
use scs8hd_conb_1  _214_
timestamp 1586364061
transform 1 0 5704 0 1 23392
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 -1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_42
timestamp 1586364061
transform 1 0 4968 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_46
timestamp 1586364061
transform 1 0 5336 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_40_36
timestamp 1586364061
transform 1 0 4416 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_46
timestamp 1586364061
transform 1 0 5336 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_58
timestamp 1586364061
transform 1 0 6440 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_71
timestamp 1586364061
transform 1 0 7636 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_66
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 -1 24480
box -38 -48 866 592
use scs8hd_conb_1  _213_
timestamp 1586364061
transform 1 0 8372 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9108 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_79
timestamp 1586364061
transform 1 0 8372 0 1 23392
box -38 -48 774 592
use scs8hd_decap_4  FILLER_40_75
timestamp 1586364061
transform 1 0 8004 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_8  FILLER_40_82
timestamp 1586364061
transform 1 0 8648 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_90
timestamp 1586364061
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_94
timestamp 1586364061
transform 1 0 9752 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_90
timestamp 1586364061
transform 1 0 9384 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9568 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_106
timestamp 1586364061
transform 1 0 10856 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_107
timestamp 1586364061
transform 1 0 10948 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 866 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 10028 0 -1 24480
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11592 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 11132 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_111
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_39_116
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_40_139
timestamp 1586364061
transform 1 0 13892 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_138
timestamp 1586364061
transform 1 0 13800 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_134
timestamp 1586364061
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 13616 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 14168 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 13984 0 1 23392
box -38 -48 222 592
use scs8hd_inv_8  _124_
timestamp 1586364061
transform 1 0 12604 0 1 23392
box -38 -48 866 592
use scs8hd_or3_4  _091_
timestamp 1586364061
transform 1 0 14168 0 1 23392
box -38 -48 866 592
use scs8hd_inv_8  _090_
timestamp 1586364061
transform 1 0 13064 0 -1 24480
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 14536 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_151
timestamp 1586364061
transform 1 0 14996 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_144
timestamp 1586364061
transform 1 0 14352 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_148
timestamp 1586364061
transform 1 0 14720 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_152
timestamp 1586364061
transform 1 0 15088 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16192 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_162
timestamp 1586364061
transform 1 0 16008 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_166
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_39_178
timestamp 1586364061
transform 1 0 17480 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _248_
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_182
timestamp 1586364061
transform 1 0 17848 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _247_
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__247__A
timestamp 1586364061
transform 1 0 20792 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__248__A
timestamp 1586364061
transform 1 0 19688 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_200
timestamp 1586364061
transform 1 0 19504 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_204
timestamp 1586364061
transform 1 0 19872 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_212
timestamp 1586364061
transform 1 0 20608 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_221
timestamp 1586364061
transform 1 0 21436 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_6  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 590 592
use scs8hd_decap_4  FILLER_39_216
timestamp 1586364061
transform 1 0 20976 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _246_
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _245_
timestamp 1586364061
transform 1 0 21528 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_228
timestamp 1586364061
transform 1 0 22080 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_224
timestamp 1586364061
transform 1 0 21712 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__245__A
timestamp 1586364061
transform 1 0 22264 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__246__A
timestamp 1586364061
transform 1 0 21896 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_226
timestamp 1586364061
transform 1 0 21896 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_232
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_238
timestamp 1586364061
transform 1 0 23000 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _240_
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_250
timestamp 1586364061
transform 1 0 24104 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_262
timestamp 1586364061
transform 1 0 25208 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_275
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_274
timestamp 1586364061
transform 1 0 26312 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_2  _224_
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 406 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__224__A
timestamp 1586364061
transform 1 0 2300 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_7
timestamp 1586364061
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_11
timestamp 1586364061
transform 1 0 2116 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3220 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3680 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_19
timestamp 1586364061
transform 1 0 2852 0 1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_41_22
timestamp 1586364061
transform 1 0 3128 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_26
timestamp 1586364061
transform 1 0 3496 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_30
timestamp 1586364061
transform 1 0 3864 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_34
timestamp 1586364061
transform 1 0 4232 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_47
timestamp 1586364061
transform 1 0 5428 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_53
timestamp 1586364061
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_57
timestamp 1586364061
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 314 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 8648 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 8464 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8096 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_78
timestamp 1586364061
transform 1 0 8280 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 10212 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 10764 0 1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_41_91
timestamp 1586364061
transform 1 0 9476 0 1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_41_103
timestamp 1586364061
transform 1 0 10580 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_107
timestamp 1586364061
transform 1 0 10948 0 1 24480
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_114
timestamp 1586364061
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_118
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 14076 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_126
timestamp 1586364061
transform 1 0 12696 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_130
timestamp 1586364061
transform 1 0 13064 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_134
timestamp 1586364061
transform 1 0 13432 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_139
timestamp 1586364061
transform 1 0 13892 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_143
timestamp 1586364061
transform 1 0 14260 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_155
timestamp 1586364061
transform 1 0 15364 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_167
timestamp 1586364061
transform 1 0 16468 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_41_179
timestamp 1586364061
transform 1 0 17572 0 1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_6
timestamp 1586364061
transform 1 0 1656 0 -1 25568
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_18
timestamp 1586364061
transform 1 0 2760 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_23
timestamp 1586364061
transform 1 0 3220 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_4  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5796 0 -1 25568
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4508 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4968 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_36
timestamp 1586364061
transform 1 0 4416 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_40
timestamp 1586364061
transform 1 0 4784 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_1  FILLER_42_50
timestamp 1586364061
transform 1 0 5704 0 -1 25568
box -38 -48 130 592
use scs8hd_inv_8  _204_
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_54
timestamp 1586364061
transform 1 0 6072 0 -1 25568
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_72
timestamp 1586364061
transform 1 0 7728 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_76
timestamp 1586364061
transform 1 0 8096 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_8  FILLER_42_85
timestamp 1586364061
transform 1 0 8924 0 -1 25568
box -38 -48 774 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 10028 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_100
timestamp 1586364061
transform 1 0 10304 0 -1 25568
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_42_112
timestamp 1586364061
transform 1 0 11408 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_116
timestamp 1586364061
transform 1 0 11776 0 -1 25568
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13156 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_6  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_134
timestamp 1586364061
transform 1 0 13432 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_146
timestamp 1586364061
transform 1 0 14536 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_42_154
timestamp 1586364061
transform 1 0 15272 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 15566 27520 15622 28000 6 address[0]
port 0 nsew default input
rlabel metal2 s 16302 27520 16358 28000 6 address[1]
port 1 nsew default input
rlabel metal2 s 17130 27520 17186 28000 6 address[2]
port 2 nsew default input
rlabel metal2 s 17958 27520 18014 28000 6 address[3]
port 3 nsew default input
rlabel metal2 s 18694 27520 18750 28000 6 address[4]
port 4 nsew default input
rlabel metal2 s 19522 27520 19578 28000 6 address[5]
port 5 nsew default input
rlabel metal2 s 20350 27520 20406 28000 6 address[6]
port 6 nsew default input
rlabel metal2 s 9402 0 9458 480 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal2 s 15382 0 15438 480 6 bottom_right_grid_pin_11_
port 8 nsew default input
rlabel metal2 s 16394 0 16450 480 6 bottom_right_grid_pin_13_
port 9 nsew default input
rlabel metal2 s 17406 0 17462 480 6 bottom_right_grid_pin_15_
port 10 nsew default input
rlabel metal2 s 10414 0 10470 480 6 bottom_right_grid_pin_1_
port 11 nsew default input
rlabel metal2 s 11426 0 11482 480 6 bottom_right_grid_pin_3_
port 12 nsew default input
rlabel metal2 s 12438 0 12494 480 6 bottom_right_grid_pin_5_
port 13 nsew default input
rlabel metal2 s 13450 0 13506 480 6 bottom_right_grid_pin_7_
port 14 nsew default input
rlabel metal2 s 14462 0 14518 480 6 bottom_right_grid_pin_9_
port 15 nsew default input
rlabel metal3 s 0 688 480 808 6 chanx_left_in[0]
port 16 nsew default input
rlabel metal3 s 0 2048 480 2168 6 chanx_left_in[1]
port 17 nsew default input
rlabel metal3 s 0 3408 480 3528 6 chanx_left_in[2]
port 18 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[3]
port 19 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chanx_left_in[4]
port 20 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[5]
port 21 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[6]
port 22 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[7]
port 23 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[8]
port 24 nsew default input
rlabel metal3 s 0 16056 480 16176 6 chanx_left_out[0]
port 25 nsew default tristate
rlabel metal3 s 0 17416 480 17536 6 chanx_left_out[1]
port 26 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chanx_left_out[2]
port 27 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chanx_left_out[3]
port 28 nsew default tristate
rlabel metal3 s 0 21632 480 21752 6 chanx_left_out[4]
port 29 nsew default tristate
rlabel metal3 s 0 22992 480 23112 6 chanx_left_out[5]
port 30 nsew default tristate
rlabel metal3 s 0 24488 480 24608 6 chanx_left_out[6]
port 31 nsew default tristate
rlabel metal3 s 0 25848 480 25968 6 chanx_left_out[7]
port 32 nsew default tristate
rlabel metal3 s 0 27208 480 27328 6 chanx_left_out[8]
port 33 nsew default tristate
rlabel metal2 s 478 0 534 480 6 chany_bottom_in[0]
port 34 nsew default input
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_in[1]
port 35 nsew default input
rlabel metal2 s 2410 0 2466 480 6 chany_bottom_in[2]
port 36 nsew default input
rlabel metal2 s 3422 0 3478 480 6 chany_bottom_in[3]
port 37 nsew default input
rlabel metal2 s 4434 0 4490 480 6 chany_bottom_in[4]
port 38 nsew default input
rlabel metal2 s 5446 0 5502 480 6 chany_bottom_in[5]
port 39 nsew default input
rlabel metal2 s 6458 0 6514 480 6 chany_bottom_in[6]
port 40 nsew default input
rlabel metal2 s 7470 0 7526 480 6 chany_bottom_in[7]
port 41 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_in[8]
port 42 nsew default input
rlabel metal2 s 19430 0 19486 480 6 chany_bottom_out[0]
port 43 nsew default tristate
rlabel metal2 s 20442 0 20498 480 6 chany_bottom_out[1]
port 44 nsew default tristate
rlabel metal2 s 21454 0 21510 480 6 chany_bottom_out[2]
port 45 nsew default tristate
rlabel metal2 s 22374 0 22430 480 6 chany_bottom_out[3]
port 46 nsew default tristate
rlabel metal2 s 23386 0 23442 480 6 chany_bottom_out[4]
port 47 nsew default tristate
rlabel metal2 s 24398 0 24454 480 6 chany_bottom_out[5]
port 48 nsew default tristate
rlabel metal2 s 25410 0 25466 480 6 chany_bottom_out[6]
port 49 nsew default tristate
rlabel metal2 s 26422 0 26478 480 6 chany_bottom_out[7]
port 50 nsew default tristate
rlabel metal2 s 27434 0 27490 480 6 chany_bottom_out[8]
port 51 nsew default tristate
rlabel metal2 s 386 27520 442 28000 6 chany_top_in[0]
port 52 nsew default input
rlabel metal2 s 1122 27520 1178 28000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 1950 27520 2006 28000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 2778 27520 2834 28000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 3514 27520 3570 28000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 4342 27520 4398 28000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 5170 27520 5226 28000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 5906 27520 5962 28000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 6734 27520 6790 28000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 21086 27520 21142 28000 6 chany_top_out[0]
port 61 nsew default tristate
rlabel metal2 s 21914 27520 21970 28000 6 chany_top_out[1]
port 62 nsew default tristate
rlabel metal2 s 22742 27520 22798 28000 6 chany_top_out[2]
port 63 nsew default tristate
rlabel metal2 s 23478 27520 23534 28000 6 chany_top_out[3]
port 64 nsew default tristate
rlabel metal2 s 24306 27520 24362 28000 6 chany_top_out[4]
port 65 nsew default tristate
rlabel metal2 s 25134 27520 25190 28000 6 chany_top_out[5]
port 66 nsew default tristate
rlabel metal2 s 25870 27520 25926 28000 6 chany_top_out[6]
port 67 nsew default tristate
rlabel metal2 s 26698 27520 26754 28000 6 chany_top_out[7]
port 68 nsew default tristate
rlabel metal2 s 27526 27520 27582 28000 6 chany_top_out[8]
port 69 nsew default tristate
rlabel metal2 s 18418 0 18474 480 6 data_in
port 70 nsew default input
rlabel metal2 s 14738 27520 14794 28000 6 enable
port 71 nsew default input
rlabel metal3 s 0 14696 480 14816 6 left_bottom_grid_pin_12_
port 72 nsew default input
rlabel metal3 s 0 13200 480 13320 6 left_top_grid_pin_10_
port 73 nsew default input
rlabel metal2 s 7562 27520 7618 28000 6 top_left_grid_pin_13_
port 74 nsew default input
rlabel metal2 s 12346 27520 12402 28000 6 top_right_grid_pin_11_
port 75 nsew default input
rlabel metal2 s 13082 27520 13138 28000 6 top_right_grid_pin_13_
port 76 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 top_right_grid_pin_15_
port 77 nsew default input
rlabel metal2 s 8298 27520 8354 28000 6 top_right_grid_pin_1_
port 78 nsew default input
rlabel metal2 s 9126 27520 9182 28000 6 top_right_grid_pin_3_
port 79 nsew default input
rlabel metal2 s 9954 27520 10010 28000 6 top_right_grid_pin_5_
port 80 nsew default input
rlabel metal2 s 10690 27520 10746 28000 6 top_right_grid_pin_7_
port 81 nsew default input
rlabel metal2 s 11518 27520 11574 28000 6 top_right_grid_pin_9_
port 82 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 83 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 84 nsew default input
<< end >>
