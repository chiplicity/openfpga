magic
tech EFS8A
magscale 1 2
timestamp 1604430918
<< locali >>
rect 6377 13719 6411 14025
rect 6469 12699 6503 12937
rect 20729 12631 20763 12733
rect 16037 10455 16071 10761
rect 3249 10047 3283 10149
rect 6469 7327 6503 7497
<< viali >>
rect 12357 21097 12391 21131
rect 17417 21097 17451 21131
rect 26709 21097 26743 21131
rect 12173 20961 12207 20995
rect 17233 20961 17267 20995
rect 18613 20961 18647 20995
rect 18705 20961 18739 20995
rect 26525 20961 26559 20995
rect 18797 20893 18831 20927
rect 5089 20757 5123 20791
rect 12633 20757 12667 20791
rect 18245 20757 18279 20791
rect 1593 20553 1627 20587
rect 2605 20553 2639 20587
rect 7021 20553 7055 20587
rect 9321 20553 9355 20587
rect 14657 20553 14691 20587
rect 16865 20553 16899 20587
rect 20361 20553 20395 20587
rect 24409 20553 24443 20587
rect 26893 20553 26927 20587
rect 11529 20485 11563 20519
rect 12449 20485 12483 20519
rect 25421 20485 25455 20519
rect 5457 20417 5491 20451
rect 5549 20417 5583 20451
rect 12265 20417 12299 20451
rect 13001 20417 13035 20451
rect 18705 20417 18739 20451
rect 1409 20349 1443 20383
rect 2421 20349 2455 20383
rect 2881 20349 2915 20383
rect 4905 20349 4939 20383
rect 6837 20349 6871 20383
rect 9137 20349 9171 20383
rect 12817 20349 12851 20383
rect 14473 20349 14507 20383
rect 14933 20349 14967 20383
rect 16681 20349 16715 20383
rect 17785 20349 17819 20383
rect 20177 20349 20211 20383
rect 24225 20349 24259 20383
rect 25237 20349 25271 20383
rect 5365 20281 5399 20315
rect 11805 20281 11839 20315
rect 18613 20281 18647 20315
rect 1961 20213 1995 20247
rect 4445 20213 4479 20247
rect 4997 20213 5031 20247
rect 7389 20213 7423 20247
rect 9689 20213 9723 20247
rect 12909 20213 12943 20247
rect 16589 20213 16623 20247
rect 17509 20213 17543 20247
rect 18153 20213 18187 20247
rect 18521 20213 18555 20247
rect 19165 20213 19199 20247
rect 19625 20213 19659 20247
rect 20729 20213 20763 20247
rect 24777 20213 24811 20247
rect 25789 20213 25823 20247
rect 26433 20213 26467 20247
rect 4445 20009 4479 20043
rect 5273 20009 5307 20043
rect 5641 20009 5675 20043
rect 12357 20009 12391 20043
rect 16681 20009 16715 20043
rect 17233 20009 17267 20043
rect 17601 20009 17635 20043
rect 18797 20009 18831 20043
rect 18245 19941 18279 19975
rect 4261 19873 4295 19907
rect 11805 19873 11839 19907
rect 12265 19873 12299 19907
rect 19165 19873 19199 19907
rect 26893 19873 26927 19907
rect 5733 19805 5767 19839
rect 5825 19805 5859 19839
rect 11437 19805 11471 19839
rect 12449 19805 12483 19839
rect 17693 19805 17727 19839
rect 17785 19805 17819 19839
rect 19257 19805 19291 19839
rect 19349 19805 19383 19839
rect 26985 19805 27019 19839
rect 27169 19805 27203 19839
rect 11897 19737 11931 19771
rect 3525 19669 3559 19703
rect 5089 19669 5123 19703
rect 6285 19669 6319 19703
rect 10885 19669 10919 19703
rect 13001 19669 13035 19703
rect 15117 19669 15151 19703
rect 18613 19669 18647 19703
rect 19809 19669 19843 19703
rect 25421 19669 25455 19703
rect 26525 19669 26559 19703
rect 4997 19465 5031 19499
rect 6009 19465 6043 19499
rect 10793 19465 10827 19499
rect 13921 19465 13955 19499
rect 16589 19465 16623 19499
rect 18981 19465 19015 19499
rect 3341 19329 3375 19363
rect 3985 19329 4019 19363
rect 5549 19329 5583 19363
rect 6377 19329 6411 19363
rect 11345 19329 11379 19363
rect 15577 19329 15611 19363
rect 2973 19261 3007 19295
rect 3801 19261 3835 19295
rect 5457 19261 5491 19295
rect 8861 19261 8895 19295
rect 9321 19261 9355 19295
rect 9873 19261 9907 19295
rect 11253 19261 11287 19295
rect 12548 19261 12582 19295
rect 14841 19261 14875 19295
rect 18429 19261 18463 19295
rect 19533 19261 19567 19295
rect 25329 19261 25363 19295
rect 25585 19261 25619 19295
rect 27997 19261 28031 19295
rect 10333 19193 10367 19227
rect 11161 19193 11195 19227
rect 12786 19193 12820 19227
rect 15393 19193 15427 19227
rect 16957 19193 16991 19227
rect 17877 19193 17911 19227
rect 19800 19193 19834 19227
rect 3433 19125 3467 19159
rect 3893 19125 3927 19159
rect 4445 19125 4479 19159
rect 4813 19125 4847 19159
rect 5365 19125 5399 19159
rect 6837 19125 6871 19159
rect 9045 19125 9079 19159
rect 10609 19125 10643 19159
rect 11897 19125 11931 19159
rect 15025 19125 15059 19159
rect 15485 19125 15519 19159
rect 17325 19125 17359 19159
rect 18521 19125 18555 19159
rect 19441 19125 19475 19159
rect 20913 19125 20947 19159
rect 25145 19125 25179 19159
rect 26709 19125 26743 19159
rect 27261 19125 27295 19159
rect 27629 19125 27663 19159
rect 2421 18921 2455 18955
rect 3893 18921 3927 18955
rect 6101 18921 6135 18955
rect 7205 18921 7239 18955
rect 7665 18921 7699 18955
rect 9781 18921 9815 18955
rect 10149 18921 10183 18955
rect 12725 18921 12759 18955
rect 13277 18921 13311 18955
rect 14197 18921 14231 18955
rect 18429 18921 18463 18955
rect 18797 18921 18831 18955
rect 18981 18921 19015 18955
rect 20913 18921 20947 18955
rect 22661 18921 22695 18955
rect 24869 18921 24903 18955
rect 26341 18921 26375 18955
rect 26985 18921 27019 18955
rect 4629 18853 4663 18887
rect 4966 18853 5000 18887
rect 11590 18853 11624 18887
rect 20361 18853 20395 18887
rect 2237 18785 2271 18819
rect 2697 18785 2731 18819
rect 7573 18785 7607 18819
rect 9505 18785 9539 18819
rect 10241 18785 10275 18819
rect 11345 18785 11379 18819
rect 16764 18785 16798 18819
rect 19349 18785 19383 18819
rect 21281 18785 21315 18819
rect 22477 18785 22511 18819
rect 25237 18785 25271 18819
rect 25329 18785 25363 18819
rect 25973 18785 26007 18819
rect 26893 18785 26927 18819
rect 4721 18717 4755 18751
rect 7757 18717 7791 18751
rect 10333 18717 10367 18751
rect 16497 18717 16531 18751
rect 19441 18717 19475 18751
rect 19533 18717 19567 18751
rect 21373 18717 21407 18751
rect 21465 18717 21499 18751
rect 25421 18717 25455 18751
rect 27077 18717 27111 18751
rect 24777 18649 24811 18683
rect 26525 18649 26559 18683
rect 1869 18581 1903 18615
rect 3433 18581 3467 18615
rect 6929 18581 6963 18615
rect 8585 18581 8619 18615
rect 8953 18581 8987 18615
rect 10793 18581 10827 18615
rect 15025 18581 15059 18615
rect 17877 18581 17911 18615
rect 19993 18581 20027 18615
rect 22017 18581 22051 18615
rect 27537 18581 27571 18615
rect 3341 18377 3375 18411
rect 4905 18377 4939 18411
rect 7849 18377 7883 18411
rect 10793 18377 10827 18411
rect 12449 18377 12483 18411
rect 18061 18377 18095 18411
rect 19625 18377 19659 18411
rect 24041 18377 24075 18411
rect 26985 18377 27019 18411
rect 6837 18309 6871 18343
rect 9873 18309 9907 18343
rect 10609 18309 10643 18343
rect 16957 18309 16991 18343
rect 17877 18309 17911 18343
rect 25881 18309 25915 18343
rect 26525 18309 26559 18343
rect 27997 18309 28031 18343
rect 3893 18241 3927 18275
rect 5549 18241 5583 18275
rect 5917 18241 5951 18275
rect 7389 18241 7423 18275
rect 9045 18241 9079 18275
rect 10241 18241 10275 18275
rect 11437 18241 11471 18275
rect 11897 18241 11931 18275
rect 13093 18241 13127 18275
rect 13461 18241 13495 18275
rect 17509 18241 17543 18275
rect 18521 18241 18555 18275
rect 18613 18241 18647 18275
rect 20085 18241 20119 18275
rect 20177 18241 20211 18275
rect 22109 18241 22143 18275
rect 27537 18241 27571 18275
rect 1409 18173 1443 18207
rect 3709 18173 3743 18207
rect 11161 18173 11195 18207
rect 12817 18173 12851 18207
rect 14197 18173 14231 18207
rect 18429 18173 18463 18207
rect 19993 18173 20027 18207
rect 21465 18173 21499 18207
rect 21925 18173 21959 18207
rect 24501 18173 24535 18207
rect 2053 18105 2087 18139
rect 5273 18105 5307 18139
rect 7297 18105 7331 18139
rect 8953 18105 8987 18139
rect 12173 18105 12207 18139
rect 14442 18105 14476 18139
rect 19073 18105 19107 18139
rect 22937 18105 22971 18139
rect 24746 18105 24780 18139
rect 1593 18037 1627 18071
rect 2421 18037 2455 18071
rect 2789 18037 2823 18071
rect 3249 18037 3283 18071
rect 3801 18037 3835 18071
rect 4353 18037 4387 18071
rect 4813 18037 4847 18071
rect 5365 18037 5399 18071
rect 6561 18037 6595 18071
rect 7205 18037 7239 18071
rect 8309 18037 8343 18071
rect 8493 18037 8527 18071
rect 8861 18037 8895 18071
rect 11253 18037 11287 18071
rect 12909 18037 12943 18071
rect 14105 18037 14139 18071
rect 15577 18037 15611 18071
rect 16497 18037 16531 18071
rect 19441 18037 19475 18071
rect 20913 18037 20947 18071
rect 21557 18037 21591 18071
rect 22017 18037 22051 18071
rect 22661 18037 22695 18071
rect 24317 18037 24351 18071
rect 27353 18037 27387 18071
rect 27445 18037 27479 18071
rect 1777 17833 1811 17867
rect 3433 17833 3467 17867
rect 4353 17833 4387 17867
rect 4721 17833 4755 17867
rect 6377 17833 6411 17867
rect 7665 17833 7699 17867
rect 8033 17833 8067 17867
rect 9413 17833 9447 17867
rect 11621 17833 11655 17867
rect 12173 17833 12207 17867
rect 13645 17833 13679 17867
rect 17233 17833 17267 17867
rect 19717 17833 19751 17867
rect 20269 17833 20303 17867
rect 20913 17833 20947 17867
rect 24961 17833 24995 17867
rect 26157 17833 26191 17867
rect 26525 17833 26559 17867
rect 5242 17765 5276 17799
rect 6929 17765 6963 17799
rect 8401 17765 8435 17799
rect 14105 17765 14139 17799
rect 18245 17765 18279 17799
rect 18604 17765 18638 17799
rect 20729 17765 20763 17799
rect 22722 17765 22756 17799
rect 26985 17765 27019 17799
rect 2145 17697 2179 17731
rect 4997 17697 5031 17731
rect 7389 17697 7423 17731
rect 9689 17697 9723 17731
rect 9945 17697 9979 17731
rect 14013 17697 14047 17731
rect 16109 17697 16143 17731
rect 21281 17697 21315 17731
rect 25421 17697 25455 17731
rect 26893 17697 26927 17731
rect 2237 17629 2271 17663
rect 2329 17629 2363 17663
rect 8493 17629 8527 17663
rect 8677 17629 8711 17663
rect 12725 17629 12759 17663
rect 14197 17629 14231 17663
rect 15853 17629 15887 17663
rect 18337 17629 18371 17663
rect 21373 17629 21407 17663
rect 21465 17629 21499 17663
rect 22477 17629 22511 17663
rect 27169 17629 27203 17663
rect 1685 17561 1719 17595
rect 11989 17561 12023 17595
rect 2789 17493 2823 17527
rect 11069 17493 11103 17527
rect 13001 17493 13035 17527
rect 21925 17493 21959 17527
rect 23857 17493 23891 17527
rect 24593 17493 24627 17527
rect 25329 17493 25363 17527
rect 27629 17493 27663 17527
rect 3157 17289 3191 17323
rect 5641 17289 5675 17323
rect 6193 17289 6227 17323
rect 6653 17289 6687 17323
rect 7849 17289 7883 17323
rect 9689 17289 9723 17323
rect 10609 17289 10643 17323
rect 10793 17289 10827 17323
rect 11805 17289 11839 17323
rect 12449 17289 12483 17323
rect 13737 17289 13771 17323
rect 16405 17289 16439 17323
rect 16957 17289 16991 17323
rect 18337 17289 18371 17323
rect 19809 17289 19843 17323
rect 20637 17289 20671 17323
rect 25697 17289 25731 17323
rect 28089 17289 28123 17323
rect 10241 17221 10275 17255
rect 25053 17221 25087 17255
rect 11345 17153 11379 17187
rect 13001 17153 13035 17187
rect 14013 17153 14047 17187
rect 18981 17153 19015 17187
rect 25973 17153 26007 17187
rect 1685 17085 1719 17119
rect 1777 17085 1811 17119
rect 2044 17085 2078 17119
rect 4261 17085 4295 17119
rect 4517 17085 4551 17119
rect 8309 17085 8343 17119
rect 11161 17085 11195 17119
rect 12817 17085 12851 17119
rect 15025 17085 15059 17119
rect 17785 17085 17819 17119
rect 18797 17085 18831 17119
rect 21097 17085 21131 17119
rect 23029 17085 23063 17119
rect 23397 17085 23431 17119
rect 23673 17085 23707 17119
rect 26157 17085 26191 17119
rect 4169 17017 4203 17051
rect 7113 17017 7147 17051
rect 8576 17017 8610 17051
rect 11253 17017 11287 17051
rect 15292 17017 15326 17051
rect 20269 17017 20303 17051
rect 21364 17017 21398 17051
rect 23940 17017 23974 17051
rect 26402 17017 26436 17051
rect 3709 16949 3743 16983
rect 7389 16949 7423 16983
rect 8217 16949 8251 16983
rect 12265 16949 12299 16983
rect 12909 16949 12943 16983
rect 14473 16949 14507 16983
rect 14933 16949 14967 16983
rect 17509 16949 17543 16983
rect 18705 16949 18739 16983
rect 19441 16949 19475 16983
rect 20913 16949 20947 16983
rect 22477 16949 22511 16983
rect 27537 16949 27571 16983
rect 1685 16745 1719 16779
rect 4997 16745 5031 16779
rect 7941 16745 7975 16779
rect 9689 16745 9723 16779
rect 11253 16745 11287 16779
rect 12817 16745 12851 16779
rect 13737 16745 13771 16779
rect 15301 16745 15335 16779
rect 17325 16745 17359 16779
rect 18429 16745 18463 16779
rect 20729 16745 20763 16779
rect 23029 16745 23063 16779
rect 24685 16745 24719 16779
rect 24869 16745 24903 16779
rect 25329 16745 25363 16779
rect 26525 16745 26559 16779
rect 3341 16677 3375 16711
rect 5632 16677 5666 16711
rect 8401 16677 8435 16711
rect 9137 16677 9171 16711
rect 10149 16677 10183 16711
rect 15761 16677 15795 16711
rect 20361 16677 20395 16711
rect 25237 16677 25271 16711
rect 2053 16609 2087 16643
rect 5365 16609 5399 16643
rect 7573 16609 7607 16643
rect 8493 16609 8527 16643
rect 9505 16609 9539 16643
rect 10057 16609 10091 16643
rect 11693 16609 11727 16643
rect 15025 16609 15059 16643
rect 15669 16609 15703 16643
rect 16681 16609 16715 16643
rect 17233 16609 17267 16643
rect 18797 16609 18831 16643
rect 21364 16609 21398 16643
rect 23581 16609 23615 16643
rect 26893 16609 26927 16643
rect 26985 16609 27019 16643
rect 2145 16541 2179 16575
rect 2329 16541 2363 16575
rect 4077 16541 4111 16575
rect 8585 16541 8619 16575
rect 10241 16541 10275 16575
rect 11437 16541 11471 16575
rect 14289 16541 14323 16575
rect 15853 16541 15887 16575
rect 17417 16541 17451 16575
rect 18889 16541 18923 16575
rect 19073 16541 19107 16575
rect 21097 16541 21131 16575
rect 25421 16541 25455 16575
rect 27077 16541 27111 16575
rect 8033 16473 8067 16507
rect 16865 16473 16899 16507
rect 24133 16473 24167 16507
rect 2697 16405 2731 16439
rect 3709 16405 3743 16439
rect 4537 16405 4571 16439
rect 6745 16405 6779 16439
rect 10885 16405 10919 16439
rect 16405 16405 16439 16439
rect 18153 16405 18187 16439
rect 22477 16405 22511 16439
rect 23489 16405 23523 16439
rect 26249 16405 26283 16439
rect 2881 16201 2915 16235
rect 4721 16201 4755 16235
rect 5365 16201 5399 16235
rect 5733 16201 5767 16235
rect 8125 16201 8159 16235
rect 9597 16201 9631 16235
rect 10793 16201 10827 16235
rect 11805 16201 11839 16235
rect 12449 16201 12483 16235
rect 13461 16201 13495 16235
rect 15577 16201 15611 16235
rect 17233 16201 17267 16235
rect 21373 16201 21407 16235
rect 24593 16201 24627 16235
rect 25605 16201 25639 16235
rect 28089 16201 28123 16235
rect 16221 16133 16255 16167
rect 20821 16133 20855 16167
rect 24501 16133 24535 16167
rect 25973 16133 26007 16167
rect 2421 16065 2455 16099
rect 7389 16065 7423 16099
rect 11345 16065 11379 16099
rect 12265 16065 12299 16099
rect 13093 16065 13127 16099
rect 22017 16065 22051 16099
rect 25145 16065 25179 16099
rect 3157 15997 3191 16031
rect 3341 15997 3375 16031
rect 3597 15997 3631 16031
rect 8217 15997 8251 16031
rect 14197 15997 14231 16031
rect 14464 15997 14498 16031
rect 18061 15997 18095 16031
rect 18317 15997 18351 16031
rect 21833 15997 21867 16031
rect 22753 15997 22787 16031
rect 24961 15997 24995 16031
rect 26157 15997 26191 16031
rect 26424 15997 26458 16031
rect 1685 15929 1719 15963
rect 2145 15929 2179 15963
rect 8462 15929 8496 15963
rect 10701 15929 10735 15963
rect 12817 15929 12851 15963
rect 14105 15929 14139 15963
rect 16865 15929 16899 15963
rect 21741 15929 21775 15963
rect 23121 15929 23155 15963
rect 24133 15929 24167 15963
rect 25053 15929 25087 15963
rect 1777 15861 1811 15895
rect 2237 15861 2271 15895
rect 6101 15861 6135 15895
rect 7757 15861 7791 15895
rect 10241 15861 10275 15895
rect 11161 15861 11195 15895
rect 11253 15861 11287 15895
rect 12909 15861 12943 15895
rect 16589 15861 16623 15895
rect 17785 15861 17819 15895
rect 19441 15861 19475 15895
rect 19993 15861 20027 15895
rect 21097 15861 21131 15895
rect 22385 15861 22419 15895
rect 27537 15861 27571 15895
rect 4077 15657 4111 15691
rect 4537 15657 4571 15691
rect 8217 15657 8251 15691
rect 8585 15657 8619 15691
rect 9689 15657 9723 15691
rect 13185 15657 13219 15691
rect 14473 15657 14507 15691
rect 17233 15657 17267 15691
rect 17785 15657 17819 15691
rect 21097 15657 21131 15691
rect 22109 15657 22143 15691
rect 23213 15657 23247 15691
rect 24777 15657 24811 15691
rect 25881 15657 25915 15691
rect 27537 15657 27571 15691
rect 7941 15589 7975 15623
rect 9137 15589 9171 15623
rect 9505 15589 9539 15623
rect 12050 15589 12084 15623
rect 15568 15589 15602 15623
rect 1501 15521 1535 15555
rect 1768 15521 1802 15555
rect 4445 15521 4479 15555
rect 5273 15521 5307 15555
rect 6000 15521 6034 15555
rect 10057 15521 10091 15555
rect 18501 15521 18535 15555
rect 21465 15521 21499 15555
rect 23581 15521 23615 15555
rect 24685 15521 24719 15555
rect 25145 15521 25179 15555
rect 26893 15521 26927 15555
rect 4629 15453 4663 15487
rect 5733 15453 5767 15487
rect 10149 15453 10183 15487
rect 10333 15453 10367 15487
rect 11529 15453 11563 15487
rect 11805 15453 11839 15487
rect 15301 15453 15335 15487
rect 18245 15453 18279 15487
rect 21557 15453 21591 15487
rect 21741 15453 21775 15487
rect 23673 15453 23707 15487
rect 23857 15453 23891 15487
rect 25237 15453 25271 15487
rect 25421 15453 25455 15487
rect 26157 15453 26191 15487
rect 26985 15453 27019 15487
rect 27169 15453 27203 15487
rect 2881 15385 2915 15419
rect 3525 15317 3559 15351
rect 3893 15317 3927 15351
rect 5641 15317 5675 15351
rect 7113 15317 7147 15351
rect 10793 15317 10827 15351
rect 13829 15317 13863 15351
rect 16681 15317 16715 15351
rect 18061 15317 18095 15351
rect 19625 15317 19659 15351
rect 20269 15317 20303 15351
rect 20729 15317 20763 15351
rect 24317 15317 24351 15351
rect 26525 15317 26559 15351
rect 1961 15113 1995 15147
rect 6193 15113 6227 15147
rect 7849 15113 7883 15147
rect 8953 15113 8987 15147
rect 11529 15113 11563 15147
rect 12173 15113 12207 15147
rect 16037 15113 16071 15147
rect 20085 15113 20119 15147
rect 21649 15113 21683 15147
rect 3525 15045 3559 15079
rect 7665 15045 7699 15079
rect 9229 15045 9263 15079
rect 12909 15045 12943 15079
rect 13921 15045 13955 15079
rect 15853 15045 15887 15079
rect 2605 14977 2639 15011
rect 4077 14977 4111 15011
rect 4537 14977 4571 15011
rect 5825 14977 5859 15011
rect 7297 14977 7331 15011
rect 8401 14977 8435 15011
rect 9413 14977 9447 15011
rect 11897 14977 11931 15011
rect 13553 14977 13587 15011
rect 14289 14977 14323 15011
rect 14933 14977 14967 15011
rect 15117 14977 15151 15011
rect 16589 14977 16623 15011
rect 19165 14977 19199 15011
rect 19625 14977 19659 15011
rect 20729 14977 20763 15011
rect 22201 14977 22235 15011
rect 23213 14977 23247 15011
rect 27353 14977 27387 15011
rect 1869 14909 1903 14943
rect 2329 14909 2363 14943
rect 5089 14909 5123 14943
rect 8217 14909 8251 14943
rect 13277 14909 13311 14943
rect 14841 14909 14875 14943
rect 15577 14909 15611 14943
rect 21189 14909 21223 14943
rect 22017 14909 22051 14943
rect 24317 14909 24351 14943
rect 27261 14909 27295 14943
rect 2421 14841 2455 14875
rect 5549 14841 5583 14875
rect 9658 14841 9692 14875
rect 13369 14841 13403 14875
rect 16405 14841 16439 14875
rect 18429 14841 18463 14875
rect 18889 14841 18923 14875
rect 24562 14841 24596 14875
rect 28181 14841 28215 14875
rect 2973 14773 3007 14807
rect 3433 14773 3467 14807
rect 3893 14773 3927 14807
rect 3985 14773 4019 14807
rect 5181 14773 5215 14807
rect 5641 14773 5675 14807
rect 6561 14773 6595 14807
rect 6837 14773 6871 14807
rect 8309 14773 8343 14807
rect 10793 14773 10827 14807
rect 12817 14773 12851 14807
rect 14473 14773 14507 14807
rect 16497 14773 16531 14807
rect 17049 14773 17083 14807
rect 17417 14773 17451 14807
rect 17877 14773 17911 14807
rect 18521 14773 18555 14807
rect 18981 14773 19015 14807
rect 19901 14773 19935 14807
rect 20453 14773 20487 14807
rect 20545 14773 20579 14807
rect 21465 14773 21499 14807
rect 22109 14773 22143 14807
rect 22937 14773 22971 14807
rect 24225 14773 24259 14807
rect 25697 14773 25731 14807
rect 26617 14773 26651 14807
rect 26801 14773 26835 14807
rect 27169 14773 27203 14807
rect 27813 14773 27847 14807
rect 1961 14569 1995 14603
rect 2973 14569 3007 14603
rect 3617 14569 3651 14603
rect 4629 14569 4663 14603
rect 5273 14569 5307 14603
rect 8401 14569 8435 14603
rect 8493 14569 8527 14603
rect 12449 14569 12483 14603
rect 13093 14569 13127 14603
rect 13645 14569 13679 14603
rect 14105 14569 14139 14603
rect 15301 14569 15335 14603
rect 17141 14569 17175 14603
rect 18245 14569 18279 14603
rect 19625 14569 19659 14603
rect 20361 14569 20395 14603
rect 20729 14569 20763 14603
rect 22845 14569 22879 14603
rect 23489 14569 23523 14603
rect 23765 14569 23799 14603
rect 25973 14569 26007 14603
rect 27537 14569 27571 14603
rect 5702 14501 5736 14535
rect 16405 14501 16439 14535
rect 18981 14501 19015 14535
rect 26341 14501 26375 14535
rect 2329 14433 2363 14467
rect 4077 14433 4111 14467
rect 5457 14433 5491 14467
rect 9965 14433 9999 14467
rect 11336 14433 11370 14467
rect 14013 14433 14047 14467
rect 15669 14433 15703 14467
rect 15761 14433 15795 14467
rect 17509 14433 17543 14467
rect 19717 14433 19751 14467
rect 21732 14433 21766 14467
rect 24205 14433 24239 14467
rect 26893 14433 26927 14467
rect 2421 14365 2455 14399
rect 2605 14365 2639 14399
rect 8677 14365 8711 14399
rect 11069 14365 11103 14399
rect 14197 14365 14231 14399
rect 15853 14365 15887 14399
rect 17601 14365 17635 14399
rect 17785 14365 17819 14399
rect 19901 14365 19935 14399
rect 21465 14365 21499 14399
rect 23949 14365 23983 14399
rect 26985 14365 27019 14399
rect 27077 14365 27111 14399
rect 1685 14297 1719 14331
rect 7389 14297 7423 14331
rect 8033 14297 8067 14331
rect 13461 14297 13495 14331
rect 15025 14297 15059 14331
rect 4261 14229 4295 14263
rect 6837 14229 6871 14263
rect 7849 14229 7883 14263
rect 9137 14229 9171 14263
rect 9505 14229 9539 14263
rect 10333 14229 10367 14263
rect 10885 14229 10919 14263
rect 16681 14229 16715 14263
rect 18521 14229 18555 14263
rect 19257 14229 19291 14263
rect 21097 14229 21131 14263
rect 25329 14229 25363 14263
rect 26525 14229 26559 14263
rect 2053 14025 2087 14059
rect 2421 14025 2455 14059
rect 4629 14025 4663 14059
rect 6193 14025 6227 14059
rect 6377 14025 6411 14059
rect 6561 14025 6595 14059
rect 8309 14025 8343 14059
rect 9229 14025 9263 14059
rect 10793 14025 10827 14059
rect 14749 14025 14783 14059
rect 16497 14025 16531 14059
rect 20085 14025 20119 14059
rect 23489 14025 23523 14059
rect 24225 14025 24259 14059
rect 25329 14025 25363 14059
rect 27721 14025 27755 14059
rect 1593 13957 1627 13991
rect 5181 13957 5215 13991
rect 2605 13889 2639 13923
rect 5825 13889 5859 13923
rect 1409 13821 1443 13855
rect 5549 13821 5583 13855
rect 2872 13753 2906 13787
rect 6837 13957 6871 13991
rect 10609 13957 10643 13991
rect 13829 13957 13863 13991
rect 14933 13957 14967 13991
rect 19441 13957 19475 13991
rect 28089 13957 28123 13991
rect 7481 13889 7515 13923
rect 7849 13889 7883 13923
rect 9045 13889 9079 13923
rect 9873 13889 9907 13923
rect 11345 13889 11379 13923
rect 14473 13889 14507 13923
rect 15577 13889 15611 13923
rect 20637 13889 20671 13923
rect 24777 13889 24811 13923
rect 7297 13821 7331 13855
rect 8585 13821 8619 13855
rect 11253 13821 11287 13855
rect 11897 13821 11931 13855
rect 12265 13821 12299 13855
rect 12449 13821 12483 13855
rect 15393 13821 15427 13855
rect 16037 13821 16071 13855
rect 16773 13821 16807 13855
rect 17509 13821 17543 13855
rect 18061 13821 18095 13855
rect 21097 13821 21131 13855
rect 21353 13821 21387 13855
rect 23121 13821 23155 13855
rect 24685 13821 24719 13855
rect 25789 13821 25823 13855
rect 26045 13821 26079 13855
rect 9597 13753 9631 13787
rect 9689 13753 9723 13787
rect 12716 13753 12750 13787
rect 18306 13753 18340 13787
rect 25605 13753 25639 13787
rect 3985 13685 4019 13719
rect 5089 13685 5123 13719
rect 5641 13685 5675 13719
rect 6377 13685 6411 13719
rect 7205 13685 7239 13719
rect 10241 13685 10275 13719
rect 11161 13685 11195 13719
rect 15301 13685 15335 13719
rect 16957 13685 16991 13719
rect 17785 13685 17819 13719
rect 20913 13685 20947 13719
rect 22477 13685 22511 13719
rect 23949 13685 23983 13719
rect 24593 13685 24627 13719
rect 27169 13685 27203 13719
rect 4077 13481 4111 13515
rect 4537 13481 4571 13515
rect 6285 13481 6319 13515
rect 9689 13481 9723 13515
rect 10057 13481 10091 13515
rect 11253 13481 11287 13515
rect 11529 13481 11563 13515
rect 11897 13481 11931 13515
rect 13553 13481 13587 13515
rect 14105 13481 14139 13515
rect 19165 13481 19199 13515
rect 20269 13481 20303 13515
rect 21189 13481 21223 13515
rect 22753 13481 22787 13515
rect 23121 13481 23155 13515
rect 24133 13481 24167 13515
rect 24777 13481 24811 13515
rect 25881 13481 25915 13515
rect 27629 13481 27663 13515
rect 3893 13413 3927 13447
rect 7380 13413 7414 13447
rect 14933 13413 14967 13447
rect 19625 13413 19659 13447
rect 22661 13413 22695 13447
rect 1501 13345 1535 13379
rect 1768 13345 1802 13379
rect 4445 13345 4479 13379
rect 5641 13345 5675 13379
rect 7113 13345 7147 13379
rect 9045 13345 9079 13379
rect 9505 13345 9539 13379
rect 10149 13345 10183 13379
rect 14013 13345 14047 13379
rect 15485 13345 15519 13379
rect 16764 13345 16798 13379
rect 21557 13345 21591 13379
rect 23765 13345 23799 13379
rect 24685 13345 24719 13379
rect 26893 13345 26927 13379
rect 4721 13277 4755 13311
rect 5273 13277 5307 13311
rect 10333 13277 10367 13311
rect 11989 13277 12023 13311
rect 12081 13277 12115 13311
rect 14197 13277 14231 13311
rect 16497 13277 16531 13311
rect 19717 13277 19751 13311
rect 19809 13277 19843 13311
rect 21649 13277 21683 13311
rect 21833 13277 21867 13311
rect 23213 13277 23247 13311
rect 23305 13277 23339 13311
rect 24961 13277 24995 13311
rect 26985 13277 27019 13311
rect 27169 13277 27203 13311
rect 2881 13209 2915 13243
rect 3525 13209 3559 13243
rect 12909 13209 12943 13243
rect 19257 13209 19291 13243
rect 20729 13209 20763 13243
rect 26249 13209 26283 13243
rect 5825 13141 5859 13175
rect 6929 13141 6963 13175
rect 8493 13141 8527 13175
rect 10885 13141 10919 13175
rect 12633 13141 12667 13175
rect 13645 13141 13679 13175
rect 15945 13141 15979 13175
rect 16313 13141 16347 13175
rect 17877 13141 17911 13175
rect 18429 13141 18463 13175
rect 22201 13141 22235 13175
rect 24317 13141 24351 13175
rect 25329 13141 25363 13175
rect 26525 13141 26559 13175
rect 4537 12937 4571 12971
rect 4813 12937 4847 12971
rect 6469 12937 6503 12971
rect 6561 12937 6595 12971
rect 8585 12937 8619 12971
rect 11253 12937 11287 12971
rect 13737 12937 13771 12971
rect 14841 12937 14875 12971
rect 17509 12937 17543 12971
rect 19993 12937 20027 12971
rect 22385 12937 22419 12971
rect 23029 12937 23063 12971
rect 24869 12937 24903 12971
rect 25697 12937 25731 12971
rect 28089 12937 28123 12971
rect 6285 12869 6319 12903
rect 1685 12801 1719 12835
rect 4169 12801 4203 12835
rect 5733 12801 5767 12835
rect 5549 12733 5583 12767
rect 10149 12869 10183 12903
rect 11805 12869 11839 12903
rect 12173 12869 12207 12903
rect 14749 12869 14783 12903
rect 16405 12869 16439 12903
rect 19441 12869 19475 12903
rect 25973 12869 26007 12903
rect 7665 12801 7699 12835
rect 8769 12801 8803 12835
rect 11345 12801 11379 12835
rect 13001 12801 13035 12835
rect 15301 12801 15335 12835
rect 15485 12801 15519 12835
rect 15945 12801 15979 12835
rect 17049 12801 17083 12835
rect 23489 12801 23523 12835
rect 24225 12801 24259 12835
rect 24409 12801 24443 12835
rect 7573 12733 7607 12767
rect 8125 12733 8159 12767
rect 9025 12733 9059 12767
rect 12909 12733 12943 12767
rect 14013 12733 14047 12767
rect 15209 12733 15243 12767
rect 16773 12733 16807 12767
rect 17877 12733 17911 12767
rect 18061 12733 18095 12767
rect 18328 12733 18362 12767
rect 20729 12733 20763 12767
rect 21005 12733 21039 12767
rect 24133 12733 24167 12767
rect 26157 12733 26191 12767
rect 26424 12733 26458 12767
rect 1952 12665 1986 12699
rect 5641 12665 5675 12699
rect 6469 12665 6503 12699
rect 7481 12665 7515 12699
rect 16865 12665 16899 12699
rect 20453 12665 20487 12699
rect 21250 12665 21284 12699
rect 25145 12665 25179 12699
rect 3065 12597 3099 12631
rect 3617 12597 3651 12631
rect 5181 12597 5215 12631
rect 7113 12597 7147 12631
rect 10793 12597 10827 12631
rect 12449 12597 12483 12631
rect 12817 12597 12851 12631
rect 16313 12597 16347 12631
rect 20729 12597 20763 12631
rect 20821 12597 20855 12631
rect 23765 12597 23799 12631
rect 27537 12597 27571 12631
rect 1961 12393 1995 12427
rect 2237 12393 2271 12427
rect 7021 12393 7055 12427
rect 7113 12393 7147 12427
rect 8861 12393 8895 12427
rect 9965 12393 9999 12427
rect 11989 12393 12023 12427
rect 12633 12393 12667 12427
rect 14013 12393 14047 12427
rect 14933 12393 14967 12427
rect 15577 12393 15611 12427
rect 16037 12393 16071 12427
rect 16681 12393 16715 12427
rect 17049 12393 17083 12427
rect 18521 12393 18555 12427
rect 19349 12393 19383 12427
rect 19717 12393 19751 12427
rect 21281 12393 21315 12427
rect 21833 12393 21867 12427
rect 22845 12393 22879 12427
rect 26985 12393 27019 12427
rect 9137 12325 9171 12359
rect 10876 12325 10910 12359
rect 13737 12325 13771 12359
rect 21925 12325 21959 12359
rect 26157 12325 26191 12359
rect 2789 12257 2823 12291
rect 2881 12257 2915 12291
rect 3433 12257 3467 12291
rect 4077 12257 4111 12291
rect 5825 12257 5859 12291
rect 7481 12257 7515 12291
rect 7573 12257 7607 12291
rect 15945 12257 15979 12291
rect 17141 12257 17175 12291
rect 17408 12257 17442 12291
rect 23121 12257 23155 12291
rect 23653 12257 23687 12291
rect 25329 12257 25363 12291
rect 26893 12257 26927 12291
rect 1409 12189 1443 12223
rect 3065 12189 3099 12223
rect 5917 12189 5951 12223
rect 6101 12189 6135 12223
rect 7665 12189 7699 12223
rect 10609 12189 10643 12223
rect 16221 12189 16255 12223
rect 22017 12189 22051 12223
rect 23397 12189 23431 12223
rect 27169 12189 27203 12223
rect 5273 12121 5307 12155
rect 6653 12121 6687 12155
rect 20729 12121 20763 12155
rect 21465 12121 21499 12155
rect 2421 12053 2455 12087
rect 3893 12053 3927 12087
rect 4261 12053 4295 12087
rect 4629 12053 4663 12087
rect 5457 12053 5491 12087
rect 8125 12053 8159 12087
rect 10241 12053 10275 12087
rect 20085 12053 20119 12087
rect 24777 12053 24811 12087
rect 25789 12053 25823 12087
rect 26525 12053 26559 12087
rect 1685 11849 1719 11883
rect 4169 11849 4203 11883
rect 5089 11849 5123 11883
rect 6285 11849 6319 11883
rect 6653 11849 6687 11883
rect 7849 11849 7883 11883
rect 8401 11849 8435 11883
rect 9413 11849 9447 11883
rect 10057 11849 10091 11883
rect 11161 11849 11195 11883
rect 15301 11849 15335 11883
rect 15945 11849 15979 11883
rect 16405 11849 16439 11883
rect 17417 11849 17451 11883
rect 17785 11849 17819 11883
rect 21373 11849 21407 11883
rect 21925 11849 21959 11883
rect 23121 11849 23155 11883
rect 24041 11849 24075 11883
rect 26617 11849 26651 11883
rect 26985 11849 27019 11883
rect 28089 11849 28123 11883
rect 9965 11781 9999 11815
rect 11437 11781 11471 11815
rect 22385 11781 22419 11815
rect 25605 11781 25639 11815
rect 4721 11713 4755 11747
rect 5733 11713 5767 11747
rect 7389 11713 7423 11747
rect 8309 11713 8343 11747
rect 8953 11713 8987 11747
rect 10609 11713 10643 11747
rect 17049 11713 17083 11747
rect 18337 11713 18371 11747
rect 19073 11713 19107 11747
rect 24501 11713 24535 11747
rect 24593 11713 24627 11747
rect 25513 11713 25547 11747
rect 26157 11713 26191 11747
rect 2053 11645 2087 11679
rect 2145 11645 2179 11679
rect 7205 11645 7239 11679
rect 7297 11645 7331 11679
rect 10425 11645 10459 11679
rect 19993 11645 20027 11679
rect 22477 11645 22511 11679
rect 25973 11645 26007 11679
rect 27169 11645 27203 11679
rect 27721 11645 27755 11679
rect 2390 11577 2424 11611
rect 5641 11577 5675 11611
rect 8769 11577 8803 11611
rect 11805 11577 11839 11611
rect 15669 11577 15703 11611
rect 18797 11577 18831 11611
rect 19441 11577 19475 11611
rect 20238 11577 20272 11611
rect 23397 11577 23431 11611
rect 25145 11577 25179 11611
rect 26065 11577 26099 11611
rect 3525 11509 3559 11543
rect 5181 11509 5215 11543
rect 5549 11509 5583 11543
rect 6837 11509 6871 11543
rect 8861 11509 8895 11543
rect 10517 11509 10551 11543
rect 16773 11509 16807 11543
rect 16865 11509 16899 11543
rect 18429 11509 18463 11543
rect 18889 11509 18923 11543
rect 19809 11509 19843 11543
rect 22661 11509 22695 11543
rect 23857 11509 23891 11543
rect 24409 11509 24443 11543
rect 27353 11509 27387 11543
rect 2421 11305 2455 11339
rect 3525 11305 3559 11339
rect 6837 11305 6871 11339
rect 7481 11305 7515 11339
rect 8401 11305 8435 11339
rect 9321 11305 9355 11339
rect 10241 11305 10275 11339
rect 11253 11305 11287 11339
rect 11805 11305 11839 11339
rect 12265 11305 12299 11339
rect 16037 11305 16071 11339
rect 16129 11305 16163 11339
rect 17141 11305 17175 11339
rect 17693 11305 17727 11339
rect 18797 11305 18831 11339
rect 19257 11305 19291 11339
rect 21281 11305 21315 11339
rect 23489 11305 23523 11339
rect 23581 11305 23615 11339
rect 24041 11305 24075 11339
rect 24685 11305 24719 11339
rect 24961 11305 24995 11339
rect 26341 11305 26375 11339
rect 26525 11305 26559 11339
rect 1685 11237 1719 11271
rect 2789 11237 2823 11271
rect 7757 11237 7791 11271
rect 12173 11237 12207 11271
rect 16497 11237 16531 11271
rect 19165 11237 19199 11271
rect 21373 11237 21407 11271
rect 26985 11237 27019 11271
rect 4077 11169 4111 11203
rect 5724 11169 5758 11203
rect 8309 11169 8343 11203
rect 8953 11169 8987 11203
rect 10609 11169 10643 11203
rect 16589 11169 16623 11203
rect 18061 11169 18095 11203
rect 19625 11169 19659 11203
rect 19717 11169 19751 11203
rect 23949 11169 23983 11203
rect 25329 11169 25363 11203
rect 26893 11169 26927 11203
rect 2881 11101 2915 11135
rect 2973 11101 3007 11135
rect 5457 11101 5491 11135
rect 8493 11101 8527 11135
rect 10701 11101 10735 11135
rect 10885 11101 10919 11135
rect 12357 11101 12391 11135
rect 16773 11101 16807 11135
rect 17601 11101 17635 11135
rect 18153 11101 18187 11135
rect 18245 11101 18279 11135
rect 19809 11101 19843 11135
rect 21557 11101 21591 11135
rect 22477 11101 22511 11135
rect 24225 11101 24259 11135
rect 27077 11101 27111 11135
rect 3893 11033 3927 11067
rect 4261 11033 4295 11067
rect 7941 11033 7975 11067
rect 10149 11033 10183 11067
rect 20361 11033 20395 11067
rect 20913 11033 20947 11067
rect 22017 11033 22051 11067
rect 25513 11033 25547 11067
rect 2237 10965 2271 10999
rect 4721 10965 4755 10999
rect 4997 10965 5031 10999
rect 15669 10965 15703 10999
rect 2697 10761 2731 10795
rect 3709 10761 3743 10795
rect 4169 10761 4203 10795
rect 6837 10761 6871 10795
rect 10241 10761 10275 10795
rect 11253 10761 11287 10795
rect 11805 10761 11839 10795
rect 12265 10761 12299 10795
rect 12633 10761 12667 10795
rect 15393 10761 15427 10795
rect 15761 10761 15795 10795
rect 16037 10761 16071 10795
rect 16221 10761 16255 10795
rect 18061 10761 18095 10795
rect 19349 10761 19383 10795
rect 21833 10761 21867 10795
rect 22109 10761 22143 10795
rect 22477 10761 22511 10795
rect 23397 10761 23431 10795
rect 25053 10761 25087 10795
rect 25605 10761 25639 10795
rect 26249 10761 26283 10795
rect 26433 10761 26467 10795
rect 2237 10693 2271 10727
rect 9413 10693 9447 10727
rect 3341 10625 3375 10659
rect 7389 10625 7423 10659
rect 7849 10625 7883 10659
rect 10057 10625 10091 10659
rect 10885 10625 10919 10659
rect 1409 10557 1443 10591
rect 2605 10557 2639 10591
rect 3065 10557 3099 10591
rect 4261 10557 4295 10591
rect 4528 10557 4562 10591
rect 6653 10557 6687 10591
rect 7297 10557 7331 10591
rect 8401 10557 8435 10591
rect 9045 10557 9079 10591
rect 10609 10557 10643 10591
rect 7205 10489 7239 10523
rect 9781 10489 9815 10523
rect 16405 10693 16439 10727
rect 17877 10693 17911 10727
rect 27445 10693 27479 10727
rect 16957 10625 16991 10659
rect 18613 10625 18647 10659
rect 23121 10625 23155 10659
rect 26893 10625 26927 10659
rect 27077 10625 27111 10659
rect 28181 10625 28215 10659
rect 17417 10557 17451 10591
rect 18429 10557 18463 10591
rect 19809 10557 19843 10591
rect 20076 10557 20110 10591
rect 23673 10557 23707 10591
rect 23940 10557 23974 10591
rect 26801 10557 26835 10591
rect 27813 10557 27847 10591
rect 16773 10489 16807 10523
rect 18521 10489 18555 10523
rect 1593 10421 1627 10455
rect 3157 10421 3191 10455
rect 5641 10421 5675 10455
rect 6193 10421 6227 10455
rect 8309 10421 8343 10455
rect 8585 10421 8619 10455
rect 10701 10421 10735 10455
rect 16037 10421 16071 10455
rect 16865 10421 16899 10455
rect 19717 10421 19751 10455
rect 21189 10421 21223 10455
rect 1961 10217 1995 10251
rect 2329 10217 2363 10251
rect 3525 10217 3559 10251
rect 4445 10217 4479 10251
rect 5089 10217 5123 10251
rect 5457 10217 5491 10251
rect 5641 10217 5675 10251
rect 6009 10217 6043 10251
rect 6929 10217 6963 10251
rect 8953 10217 8987 10251
rect 9321 10217 9355 10251
rect 10609 10217 10643 10251
rect 16037 10217 16071 10251
rect 16497 10217 16531 10251
rect 17141 10217 17175 10251
rect 18429 10217 18463 10251
rect 19257 10217 19291 10251
rect 20269 10217 20303 10251
rect 20913 10217 20947 10251
rect 21281 10217 21315 10251
rect 24041 10217 24075 10251
rect 24409 10217 24443 10251
rect 26249 10217 26283 10251
rect 26525 10217 26559 10251
rect 26985 10217 27019 10251
rect 1409 10149 1443 10183
rect 3249 10149 3283 10183
rect 6101 10149 6135 10183
rect 18153 10149 18187 10183
rect 19717 10149 19751 10183
rect 21373 10149 21407 10183
rect 23121 10149 23155 10183
rect 2789 10081 2823 10115
rect 7573 10081 7607 10115
rect 8585 10081 8619 10115
rect 17049 10081 17083 10115
rect 19165 10081 19199 10115
rect 19625 10081 19659 10115
rect 23765 10081 23799 10115
rect 24225 10081 24259 10115
rect 25329 10081 25363 10115
rect 26893 10081 26927 10115
rect 2881 10013 2915 10047
rect 2973 10013 3007 10047
rect 3249 10013 3283 10047
rect 4537 10013 4571 10047
rect 4721 10013 4755 10047
rect 6193 10013 6227 10047
rect 7665 10013 7699 10047
rect 7849 10013 7883 10047
rect 10333 10013 10367 10047
rect 17325 10013 17359 10047
rect 17785 10013 17819 10047
rect 19901 10013 19935 10047
rect 21557 10013 21591 10047
rect 23213 10013 23247 10047
rect 27169 10013 27203 10047
rect 2421 9945 2455 9979
rect 4077 9945 4111 9979
rect 7205 9945 7239 9979
rect 8217 9945 8251 9979
rect 3893 9877 3927 9911
rect 16681 9877 16715 9911
rect 25513 9877 25547 9911
rect 4537 9673 4571 9707
rect 6285 9673 6319 9707
rect 21281 9673 21315 9707
rect 21741 9673 21775 9707
rect 24133 9673 24167 9707
rect 25237 9673 25271 9707
rect 27353 9673 27387 9707
rect 2697 9605 2731 9639
rect 5181 9605 5215 9639
rect 8861 9605 8895 9639
rect 16313 9605 16347 9639
rect 18889 9605 18923 9639
rect 25513 9605 25547 9639
rect 26341 9605 26375 9639
rect 2053 9537 2087 9571
rect 2237 9537 2271 9571
rect 5549 9537 5583 9571
rect 15945 9537 15979 9571
rect 16865 9537 16899 9571
rect 17049 9537 17083 9571
rect 3065 9469 3099 9503
rect 3157 9469 3191 9503
rect 5641 9469 5675 9503
rect 6929 9469 6963 9503
rect 18521 9469 18555 9503
rect 19349 9469 19383 9503
rect 19605 9469 19639 9503
rect 24225 9469 24259 9503
rect 24777 9469 24811 9503
rect 25329 9469 25363 9503
rect 25881 9469 25915 9503
rect 26433 9469 26467 9503
rect 27537 9469 27571 9503
rect 28089 9469 28123 9503
rect 1961 9401 1995 9435
rect 3424 9401 3458 9435
rect 7174 9401 7208 9435
rect 15577 9401 15611 9435
rect 16773 9401 16807 9435
rect 26985 9401 27019 9435
rect 1593 9333 1627 9367
rect 5825 9333 5859 9367
rect 6561 9333 6595 9367
rect 8309 9333 8343 9367
rect 16405 9333 16439 9367
rect 17417 9333 17451 9367
rect 17785 9333 17819 9367
rect 19257 9333 19291 9367
rect 20729 9333 20763 9367
rect 22109 9333 22143 9367
rect 24409 9333 24443 9367
rect 26617 9333 26651 9367
rect 27721 9333 27755 9367
rect 1685 9129 1719 9163
rect 3249 9129 3283 9163
rect 4353 9129 4387 9163
rect 6101 9129 6135 9163
rect 7573 9129 7607 9163
rect 7665 9129 7699 9163
rect 15485 9129 15519 9163
rect 19073 9129 19107 9163
rect 21373 9129 21407 9163
rect 27169 9129 27203 9163
rect 2329 9061 2363 9095
rect 2421 9061 2455 9095
rect 21281 9061 21315 9095
rect 3893 8993 3927 9027
rect 4988 8993 5022 9027
rect 16405 8993 16439 9027
rect 16764 8993 16798 9027
rect 19625 8993 19659 9027
rect 25329 8993 25363 9027
rect 26525 8993 26559 9027
rect 2605 8925 2639 8959
rect 4721 8925 4755 8959
rect 7021 8925 7055 8959
rect 7849 8925 7883 8959
rect 16497 8925 16531 8959
rect 19717 8925 19751 8959
rect 19901 8925 19935 8959
rect 21557 8925 21591 8959
rect 7205 8857 7239 8891
rect 20913 8857 20947 8891
rect 1961 8789 1995 8823
rect 8401 8789 8435 8823
rect 17877 8789 17911 8823
rect 18797 8789 18831 8823
rect 19257 8789 19291 8823
rect 20269 8789 20303 8823
rect 25513 8789 25547 8823
rect 26709 8789 26743 8823
rect 1593 8585 1627 8619
rect 3801 8585 3835 8619
rect 6009 8585 6043 8619
rect 6837 8585 6871 8619
rect 7849 8585 7883 8619
rect 16313 8585 16347 8619
rect 20729 8585 20763 8619
rect 22201 8585 22235 8619
rect 25237 8585 25271 8619
rect 25881 8585 25915 8619
rect 27353 8585 27387 8619
rect 27721 8585 27755 8619
rect 2789 8517 2823 8551
rect 5549 8517 5583 8551
rect 8401 8517 8435 8551
rect 9413 8517 9447 8551
rect 15945 8517 15979 8551
rect 21189 8517 21223 8551
rect 26617 8517 26651 8551
rect 2237 8449 2271 8483
rect 2421 8449 2455 8483
rect 3709 8449 3743 8483
rect 4261 8449 4295 8483
rect 4445 8449 4479 8483
rect 7297 8449 7331 8483
rect 7481 8449 7515 8483
rect 8953 8449 8987 8483
rect 15577 8449 15611 8483
rect 16865 8449 16899 8483
rect 17049 8449 17083 8483
rect 17785 8449 17819 8483
rect 18613 8449 18647 8483
rect 19349 8449 19383 8483
rect 20085 8449 20119 8483
rect 20269 8449 20303 8483
rect 21741 8449 21775 8483
rect 3157 8381 3191 8415
rect 5365 8381 5399 8415
rect 6653 8381 6687 8415
rect 7205 8381 7239 8415
rect 8309 8381 8343 8415
rect 8861 8381 8895 8415
rect 16773 8381 16807 8415
rect 19993 8381 20027 8415
rect 21557 8381 21591 8415
rect 21649 8381 21683 8415
rect 25329 8381 25363 8415
rect 26433 8381 26467 8415
rect 26985 8381 27019 8415
rect 27537 8381 27571 8415
rect 28089 8381 28123 8415
rect 2145 8313 2179 8347
rect 4169 8313 4203 8347
rect 4905 8313 4939 8347
rect 17509 8313 17543 8347
rect 18521 8313 18555 8347
rect 21097 8313 21131 8347
rect 1777 8245 1811 8279
rect 5273 8245 5307 8279
rect 8769 8245 8803 8279
rect 16405 8245 16439 8279
rect 18061 8245 18095 8279
rect 18429 8245 18463 8279
rect 19625 8245 19659 8279
rect 25513 8245 25547 8279
rect 1685 8041 1719 8075
rect 1961 8041 1995 8075
rect 3801 8041 3835 8075
rect 4077 8041 4111 8075
rect 4445 8041 4479 8075
rect 6377 8041 6411 8075
rect 6837 8041 6871 8075
rect 7389 8041 7423 8075
rect 16221 8041 16255 8075
rect 16589 8041 16623 8075
rect 18797 8041 18831 8075
rect 19717 8041 19751 8075
rect 21281 8041 21315 8075
rect 21557 8041 21591 8075
rect 21925 8041 21959 8075
rect 3341 7973 3375 8007
rect 4537 7973 4571 8007
rect 19625 7973 19659 8007
rect 20269 7973 20303 8007
rect 2329 7905 2363 7939
rect 6745 7905 6779 7939
rect 16773 7905 16807 7939
rect 17040 7905 17074 7939
rect 26525 7905 26559 7939
rect 2421 7837 2455 7871
rect 2513 7837 2547 7871
rect 3065 7837 3099 7871
rect 4721 7837 4755 7871
rect 6285 7837 6319 7871
rect 7021 7837 7055 7871
rect 19073 7837 19107 7871
rect 19901 7837 19935 7871
rect 19257 7769 19291 7803
rect 7757 7701 7791 7735
rect 8401 7701 8435 7735
rect 18153 7701 18187 7735
rect 26709 7701 26743 7735
rect 2421 7497 2455 7531
rect 3525 7497 3559 7531
rect 3801 7497 3835 7531
rect 4261 7497 4295 7531
rect 4537 7497 4571 7531
rect 5365 7497 5399 7531
rect 6469 7497 6503 7531
rect 6561 7497 6595 7531
rect 6929 7497 6963 7531
rect 7941 7497 7975 7531
rect 15945 7497 15979 7531
rect 17417 7497 17451 7531
rect 17877 7497 17911 7531
rect 19257 7497 19291 7531
rect 19349 7497 19383 7531
rect 20361 7497 20395 7531
rect 26985 7497 27019 7531
rect 4905 7429 4939 7463
rect 5917 7429 5951 7463
rect 6285 7361 6319 7395
rect 18521 7429 18555 7463
rect 26341 7429 26375 7463
rect 7573 7361 7607 7395
rect 16313 7361 16347 7395
rect 17049 7361 17083 7395
rect 19901 7361 19935 7395
rect 1409 7293 1443 7327
rect 2513 7293 2547 7327
rect 3065 7293 3099 7327
rect 3617 7293 3651 7327
rect 4721 7293 4755 7327
rect 6469 7293 6503 7327
rect 7389 7293 7423 7327
rect 16773 7293 16807 7327
rect 16865 7293 16899 7327
rect 19809 7293 19843 7327
rect 26433 7293 26467 7327
rect 27537 7293 27571 7327
rect 28089 7293 28123 7327
rect 2053 7225 2087 7259
rect 18889 7225 18923 7259
rect 19717 7225 19751 7259
rect 1593 7157 1627 7191
rect 2697 7157 2731 7191
rect 7297 7157 7331 7191
rect 16405 7157 16439 7191
rect 26617 7157 26651 7191
rect 27721 7157 27755 7191
rect 4353 6953 4387 6987
rect 6377 6953 6411 6987
rect 16773 6953 16807 6987
rect 19441 6953 19475 6987
rect 19717 6953 19751 6987
rect 1409 6817 1443 6851
rect 2329 6817 2363 6851
rect 2513 6817 2547 6851
rect 3065 6817 3099 6851
rect 3525 6817 3559 6851
rect 15393 6817 15427 6851
rect 16497 6817 16531 6851
rect 26525 6817 26559 6851
rect 1961 6749 1995 6783
rect 2697 6681 2731 6715
rect 1593 6613 1627 6647
rect 6929 6613 6963 6647
rect 15577 6613 15611 6647
rect 26709 6613 26743 6647
rect 1593 6409 1627 6443
rect 3065 6409 3099 6443
rect 15485 6409 15519 6443
rect 26525 6409 26559 6443
rect 2053 6341 2087 6375
rect 2421 6273 2455 6307
rect 1409 6205 1443 6239
rect 2513 6205 2547 6239
rect 2697 6069 2731 6103
rect 2053 5865 2087 5899
rect 2605 5865 2639 5899
rect 1409 5729 1443 5763
rect 1593 5525 1627 5559
rect 1593 5321 1627 5355
rect 26433 5117 26467 5151
rect 26985 5117 27019 5151
rect 26617 4981 26651 5015
rect 2053 3145 2087 3179
rect 1409 2941 1443 2975
rect 26433 2941 26467 2975
rect 26985 2941 27019 2975
rect 1593 2805 1627 2839
rect 26617 2805 26651 2839
rect 6377 2601 6411 2635
rect 8585 2601 8619 2635
rect 6745 2465 6779 2499
rect 7472 2465 7506 2499
rect 7205 2397 7239 2431
<< metal1 >>
rect 3510 22788 3516 22840
rect 3568 22828 3574 22840
rect 10594 22828 10600 22840
rect 3568 22800 10600 22828
rect 3568 22788 3574 22800
rect 10594 22788 10600 22800
rect 10652 22788 10658 22840
rect 3418 22516 3424 22568
rect 3476 22556 3482 22568
rect 7466 22556 7472 22568
rect 3476 22528 7472 22556
rect 3476 22516 3482 22528
rect 7466 22516 7472 22528
rect 7524 22516 7530 22568
rect 1104 21786 28888 21808
rect 1104 21734 5982 21786
rect 6034 21734 6046 21786
rect 6098 21734 6110 21786
rect 6162 21734 6174 21786
rect 6226 21734 15982 21786
rect 16034 21734 16046 21786
rect 16098 21734 16110 21786
rect 16162 21734 16174 21786
rect 16226 21734 25982 21786
rect 26034 21734 26046 21786
rect 26098 21734 26110 21786
rect 26162 21734 26174 21786
rect 26226 21734 28888 21786
rect 1104 21712 28888 21734
rect 3786 21632 3792 21684
rect 3844 21672 3850 21684
rect 4798 21672 4804 21684
rect 3844 21644 4804 21672
rect 3844 21632 3850 21644
rect 4798 21632 4804 21644
rect 4856 21632 4862 21684
rect 1104 21242 28888 21264
rect 1104 21190 10982 21242
rect 11034 21190 11046 21242
rect 11098 21190 11110 21242
rect 11162 21190 11174 21242
rect 11226 21190 20982 21242
rect 21034 21190 21046 21242
rect 21098 21190 21110 21242
rect 21162 21190 21174 21242
rect 21226 21190 28888 21242
rect 1104 21168 28888 21190
rect 12345 21131 12403 21137
rect 12345 21097 12357 21131
rect 12391 21128 12403 21131
rect 13998 21128 14004 21140
rect 12391 21100 14004 21128
rect 12391 21097 12403 21100
rect 12345 21091 12403 21097
rect 13998 21088 14004 21100
rect 14056 21088 14062 21140
rect 17405 21131 17463 21137
rect 17405 21097 17417 21131
rect 17451 21128 17463 21131
rect 19610 21128 19616 21140
rect 17451 21100 19616 21128
rect 17451 21097 17463 21100
rect 17405 21091 17463 21097
rect 19610 21088 19616 21100
rect 19668 21088 19674 21140
rect 26697 21131 26755 21137
rect 26697 21097 26709 21131
rect 26743 21128 26755 21131
rect 28994 21128 29000 21140
rect 26743 21100 29000 21128
rect 26743 21097 26755 21100
rect 26697 21091 26755 21097
rect 28994 21088 29000 21100
rect 29052 21088 29058 21140
rect 12158 20992 12164 21004
rect 12119 20964 12164 20992
rect 12158 20952 12164 20964
rect 12216 20952 12222 21004
rect 17126 20952 17132 21004
rect 17184 20992 17190 21004
rect 17221 20995 17279 21001
rect 17221 20992 17233 20995
rect 17184 20964 17233 20992
rect 17184 20952 17190 20964
rect 17221 20961 17233 20964
rect 17267 20961 17279 20995
rect 17221 20955 17279 20961
rect 17954 20952 17960 21004
rect 18012 20992 18018 21004
rect 18601 20995 18659 21001
rect 18601 20992 18613 20995
rect 18012 20964 18613 20992
rect 18012 20952 18018 20964
rect 18601 20961 18613 20964
rect 18647 20961 18659 20995
rect 18601 20955 18659 20961
rect 18693 20995 18751 21001
rect 18693 20961 18705 20995
rect 18739 20992 18751 20995
rect 19610 20992 19616 21004
rect 18739 20964 19616 20992
rect 18739 20961 18751 20964
rect 18693 20955 18751 20961
rect 19610 20952 19616 20964
rect 19668 20952 19674 21004
rect 24026 20952 24032 21004
rect 24084 20992 24090 21004
rect 26513 20995 26571 21001
rect 26513 20992 26525 20995
rect 24084 20964 26525 20992
rect 24084 20952 24090 20964
rect 26513 20961 26525 20964
rect 26559 20992 26571 20995
rect 26878 20992 26884 21004
rect 26559 20964 26884 20992
rect 26559 20961 26571 20964
rect 26513 20955 26571 20961
rect 26878 20952 26884 20964
rect 26936 20952 26942 21004
rect 18785 20927 18843 20933
rect 18785 20893 18797 20927
rect 18831 20893 18843 20927
rect 18785 20887 18843 20893
rect 4062 20816 4068 20868
rect 4120 20856 4126 20868
rect 5626 20856 5632 20868
rect 4120 20828 5632 20856
rect 4120 20816 4126 20828
rect 5626 20816 5632 20828
rect 5684 20816 5690 20868
rect 18690 20816 18696 20868
rect 18748 20856 18754 20868
rect 18800 20856 18828 20887
rect 18748 20828 18828 20856
rect 18748 20816 18754 20828
rect 21726 20816 21732 20868
rect 21784 20856 21790 20868
rect 25682 20856 25688 20868
rect 21784 20828 25688 20856
rect 21784 20816 21790 20828
rect 25682 20816 25688 20828
rect 25740 20816 25746 20868
rect 5074 20788 5080 20800
rect 5035 20760 5080 20788
rect 5074 20748 5080 20760
rect 5132 20748 5138 20800
rect 9766 20748 9772 20800
rect 9824 20788 9830 20800
rect 12621 20791 12679 20797
rect 12621 20788 12633 20791
rect 9824 20760 12633 20788
rect 9824 20748 9830 20760
rect 12621 20757 12633 20760
rect 12667 20788 12679 20791
rect 12802 20788 12808 20800
rect 12667 20760 12808 20788
rect 12667 20757 12679 20760
rect 12621 20751 12679 20757
rect 12802 20748 12808 20760
rect 12860 20748 12866 20800
rect 18230 20788 18236 20800
rect 18191 20760 18236 20788
rect 18230 20748 18236 20760
rect 18288 20748 18294 20800
rect 21266 20748 21272 20800
rect 21324 20788 21330 20800
rect 25774 20788 25780 20800
rect 21324 20760 25780 20788
rect 21324 20748 21330 20760
rect 25774 20748 25780 20760
rect 25832 20748 25838 20800
rect 1104 20698 28888 20720
rect 1104 20646 5982 20698
rect 6034 20646 6046 20698
rect 6098 20646 6110 20698
rect 6162 20646 6174 20698
rect 6226 20646 15982 20698
rect 16034 20646 16046 20698
rect 16098 20646 16110 20698
rect 16162 20646 16174 20698
rect 16226 20646 25982 20698
rect 26034 20646 26046 20698
rect 26098 20646 26110 20698
rect 26162 20646 26174 20698
rect 26226 20646 28888 20698
rect 1104 20624 28888 20646
rect 934 20544 940 20596
rect 992 20584 998 20596
rect 1581 20587 1639 20593
rect 1581 20584 1593 20587
rect 992 20556 1593 20584
rect 992 20544 998 20556
rect 1581 20553 1593 20556
rect 1627 20553 1639 20587
rect 1581 20547 1639 20553
rect 2593 20587 2651 20593
rect 2593 20553 2605 20587
rect 2639 20584 2651 20587
rect 2682 20584 2688 20596
rect 2639 20556 2688 20584
rect 2639 20553 2651 20556
rect 2593 20547 2651 20553
rect 2682 20544 2688 20556
rect 2740 20544 2746 20596
rect 7009 20587 7067 20593
rect 7009 20553 7021 20587
rect 7055 20584 7067 20587
rect 8202 20584 8208 20596
rect 7055 20556 8208 20584
rect 7055 20553 7067 20556
rect 7009 20547 7067 20553
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 9309 20587 9367 20593
rect 9309 20553 9321 20587
rect 9355 20584 9367 20587
rect 10226 20584 10232 20596
rect 9355 20556 10232 20584
rect 9355 20553 9367 20556
rect 9309 20547 9367 20553
rect 10226 20544 10232 20556
rect 10284 20544 10290 20596
rect 14645 20587 14703 20593
rect 14645 20553 14657 20587
rect 14691 20584 14703 20587
rect 15838 20584 15844 20596
rect 14691 20556 15844 20584
rect 14691 20553 14703 20556
rect 14645 20547 14703 20553
rect 15838 20544 15844 20556
rect 15896 20544 15902 20596
rect 16853 20587 16911 20593
rect 16853 20553 16865 20587
rect 16899 20584 16911 20587
rect 17770 20584 17776 20596
rect 16899 20556 17776 20584
rect 16899 20553 16911 20556
rect 16853 20547 16911 20553
rect 17770 20544 17776 20556
rect 17828 20544 17834 20596
rect 20346 20584 20352 20596
rect 20307 20556 20352 20584
rect 20346 20544 20352 20556
rect 20404 20544 20410 20596
rect 24397 20587 24455 20593
rect 24397 20553 24409 20587
rect 24443 20584 24455 20587
rect 25222 20584 25228 20596
rect 24443 20556 25228 20584
rect 24443 20553 24455 20556
rect 24397 20547 24455 20553
rect 25222 20544 25228 20556
rect 25280 20544 25286 20596
rect 26878 20584 26884 20596
rect 26839 20556 26884 20584
rect 26878 20544 26884 20556
rect 26936 20544 26942 20596
rect 11517 20519 11575 20525
rect 11517 20485 11529 20519
rect 11563 20516 11575 20519
rect 12158 20516 12164 20528
rect 11563 20488 12164 20516
rect 11563 20485 11575 20488
rect 11517 20479 11575 20485
rect 12158 20476 12164 20488
rect 12216 20516 12222 20528
rect 12437 20519 12495 20525
rect 12437 20516 12449 20519
rect 12216 20488 12449 20516
rect 12216 20476 12222 20488
rect 12437 20485 12449 20488
rect 12483 20485 12495 20519
rect 25406 20516 25412 20528
rect 25367 20488 25412 20516
rect 12437 20479 12495 20485
rect 25406 20476 25412 20488
rect 25464 20476 25470 20528
rect 5074 20408 5080 20460
rect 5132 20448 5138 20460
rect 5445 20451 5503 20457
rect 5445 20448 5457 20451
rect 5132 20420 5457 20448
rect 5132 20408 5138 20420
rect 5445 20417 5457 20420
rect 5491 20417 5503 20451
rect 5445 20411 5503 20417
rect 5537 20451 5595 20457
rect 5537 20417 5549 20451
rect 5583 20417 5595 20451
rect 5537 20411 5595 20417
rect 12253 20451 12311 20457
rect 12253 20417 12265 20451
rect 12299 20448 12311 20451
rect 12989 20451 13047 20457
rect 12989 20448 13001 20451
rect 12299 20420 13001 20448
rect 12299 20417 12311 20420
rect 12253 20411 12311 20417
rect 12989 20417 13001 20420
rect 13035 20448 13047 20451
rect 13630 20448 13636 20460
rect 13035 20420 13636 20448
rect 13035 20417 13047 20420
rect 12989 20411 13047 20417
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 1443 20352 1992 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 1964 20253 1992 20352
rect 2038 20340 2044 20392
rect 2096 20380 2102 20392
rect 2409 20383 2467 20389
rect 2409 20380 2421 20383
rect 2096 20352 2421 20380
rect 2096 20340 2102 20352
rect 2409 20349 2421 20352
rect 2455 20380 2467 20383
rect 2869 20383 2927 20389
rect 2869 20380 2881 20383
rect 2455 20352 2881 20380
rect 2455 20349 2467 20352
rect 2409 20343 2467 20349
rect 2869 20349 2881 20352
rect 2915 20349 2927 20383
rect 4890 20380 4896 20392
rect 4803 20352 4896 20380
rect 2869 20343 2927 20349
rect 4890 20340 4896 20352
rect 4948 20380 4954 20392
rect 5552 20380 5580 20411
rect 13630 20408 13636 20420
rect 13688 20408 13694 20460
rect 18690 20448 18696 20460
rect 18651 20420 18696 20448
rect 18690 20408 18696 20420
rect 18748 20408 18754 20460
rect 4948 20352 5580 20380
rect 6825 20383 6883 20389
rect 4948 20340 4954 20352
rect 6825 20349 6837 20383
rect 6871 20380 6883 20383
rect 9125 20383 9183 20389
rect 6871 20352 7420 20380
rect 6871 20349 6883 20352
rect 6825 20343 6883 20349
rect 5353 20315 5411 20321
rect 5353 20312 5365 20315
rect 4448 20284 5365 20312
rect 1949 20247 2007 20253
rect 1949 20213 1961 20247
rect 1995 20244 2007 20247
rect 2314 20244 2320 20256
rect 1995 20216 2320 20244
rect 1995 20213 2007 20216
rect 1949 20207 2007 20213
rect 2314 20204 2320 20216
rect 2372 20204 2378 20256
rect 4154 20204 4160 20256
rect 4212 20244 4218 20256
rect 4448 20253 4476 20284
rect 5353 20281 5365 20284
rect 5399 20281 5411 20315
rect 5353 20275 5411 20281
rect 7392 20256 7420 20352
rect 9125 20349 9137 20383
rect 9171 20380 9183 20383
rect 12618 20380 12624 20392
rect 9171 20352 9720 20380
rect 9171 20349 9183 20352
rect 9125 20343 9183 20349
rect 9692 20256 9720 20352
rect 11808 20352 12624 20380
rect 10778 20272 10784 20324
rect 10836 20312 10842 20324
rect 11808 20321 11836 20352
rect 12618 20340 12624 20352
rect 12676 20340 12682 20392
rect 12802 20380 12808 20392
rect 12763 20352 12808 20380
rect 12802 20340 12808 20352
rect 12860 20340 12866 20392
rect 13814 20340 13820 20392
rect 13872 20380 13878 20392
rect 14461 20383 14519 20389
rect 14461 20380 14473 20383
rect 13872 20352 14473 20380
rect 13872 20340 13878 20352
rect 14461 20349 14473 20352
rect 14507 20380 14519 20383
rect 14921 20383 14979 20389
rect 14921 20380 14933 20383
rect 14507 20352 14933 20380
rect 14507 20349 14519 20352
rect 14461 20343 14519 20349
rect 14921 20349 14933 20352
rect 14967 20349 14979 20383
rect 16666 20380 16672 20392
rect 16627 20352 16672 20380
rect 14921 20343 14979 20349
rect 16666 20340 16672 20352
rect 16724 20340 16730 20392
rect 17770 20380 17776 20392
rect 17731 20352 17776 20380
rect 17770 20340 17776 20352
rect 17828 20340 17834 20392
rect 20165 20383 20223 20389
rect 20165 20349 20177 20383
rect 20211 20380 20223 20383
rect 24213 20383 24271 20389
rect 20211 20352 20760 20380
rect 20211 20349 20223 20352
rect 20165 20343 20223 20349
rect 11793 20315 11851 20321
rect 11793 20312 11805 20315
rect 10836 20284 11805 20312
rect 10836 20272 10842 20284
rect 11793 20281 11805 20284
rect 11839 20281 11851 20315
rect 11793 20275 11851 20281
rect 18322 20272 18328 20324
rect 18380 20312 18386 20324
rect 18601 20315 18659 20321
rect 18601 20312 18613 20315
rect 18380 20284 18613 20312
rect 18380 20272 18386 20284
rect 18601 20281 18613 20284
rect 18647 20281 18659 20315
rect 18601 20275 18659 20281
rect 4433 20247 4491 20253
rect 4433 20244 4445 20247
rect 4212 20216 4445 20244
rect 4212 20204 4218 20216
rect 4433 20213 4445 20216
rect 4479 20213 4491 20247
rect 4982 20244 4988 20256
rect 4943 20216 4988 20244
rect 4433 20207 4491 20213
rect 4982 20204 4988 20216
rect 5040 20204 5046 20256
rect 7374 20244 7380 20256
rect 7335 20216 7380 20244
rect 7374 20204 7380 20216
rect 7432 20204 7438 20256
rect 9674 20244 9680 20256
rect 9635 20216 9680 20244
rect 9674 20204 9680 20216
rect 9732 20204 9738 20256
rect 12618 20204 12624 20256
rect 12676 20244 12682 20256
rect 12897 20247 12955 20253
rect 12897 20244 12909 20247
rect 12676 20216 12909 20244
rect 12676 20204 12682 20216
rect 12897 20213 12909 20216
rect 12943 20213 12955 20247
rect 12897 20207 12955 20213
rect 16577 20247 16635 20253
rect 16577 20213 16589 20247
rect 16623 20244 16635 20247
rect 17126 20244 17132 20256
rect 16623 20216 17132 20244
rect 16623 20213 16635 20216
rect 16577 20207 16635 20213
rect 17126 20204 17132 20216
rect 17184 20204 17190 20256
rect 17494 20244 17500 20256
rect 17455 20216 17500 20244
rect 17494 20204 17500 20216
rect 17552 20204 17558 20256
rect 18138 20244 18144 20256
rect 18099 20216 18144 20244
rect 18138 20204 18144 20216
rect 18196 20204 18202 20256
rect 18414 20204 18420 20256
rect 18472 20244 18478 20256
rect 18509 20247 18567 20253
rect 18509 20244 18521 20247
rect 18472 20216 18521 20244
rect 18472 20204 18478 20216
rect 18509 20213 18521 20216
rect 18555 20244 18567 20247
rect 19153 20247 19211 20253
rect 19153 20244 19165 20247
rect 18555 20216 19165 20244
rect 18555 20213 18567 20216
rect 18509 20207 18567 20213
rect 19153 20213 19165 20216
rect 19199 20213 19211 20247
rect 19610 20244 19616 20256
rect 19523 20216 19616 20244
rect 19153 20207 19211 20213
rect 19610 20204 19616 20216
rect 19668 20244 19674 20256
rect 20530 20244 20536 20256
rect 19668 20216 20536 20244
rect 19668 20204 19674 20216
rect 20530 20204 20536 20216
rect 20588 20204 20594 20256
rect 20732 20253 20760 20352
rect 24213 20349 24225 20383
rect 24259 20380 24271 20383
rect 25225 20383 25283 20389
rect 24259 20352 24808 20380
rect 24259 20349 24271 20352
rect 24213 20343 24271 20349
rect 24780 20256 24808 20352
rect 25225 20349 25237 20383
rect 25271 20380 25283 20383
rect 25271 20352 25820 20380
rect 25271 20349 25283 20352
rect 25225 20343 25283 20349
rect 25792 20256 25820 20352
rect 20717 20247 20775 20253
rect 20717 20213 20729 20247
rect 20763 20244 20775 20247
rect 21818 20244 21824 20256
rect 20763 20216 21824 20244
rect 20763 20213 20775 20216
rect 20717 20207 20775 20213
rect 21818 20204 21824 20216
rect 21876 20204 21882 20256
rect 24762 20244 24768 20256
rect 24723 20216 24768 20244
rect 24762 20204 24768 20216
rect 24820 20204 24826 20256
rect 25774 20244 25780 20256
rect 25735 20216 25780 20244
rect 25774 20204 25780 20216
rect 25832 20204 25838 20256
rect 26421 20247 26479 20253
rect 26421 20213 26433 20247
rect 26467 20244 26479 20247
rect 26694 20244 26700 20256
rect 26467 20216 26700 20244
rect 26467 20213 26479 20216
rect 26421 20207 26479 20213
rect 26694 20204 26700 20216
rect 26752 20204 26758 20256
rect 1104 20154 28888 20176
rect 1104 20102 10982 20154
rect 11034 20102 11046 20154
rect 11098 20102 11110 20154
rect 11162 20102 11174 20154
rect 11226 20102 20982 20154
rect 21034 20102 21046 20154
rect 21098 20102 21110 20154
rect 21162 20102 21174 20154
rect 21226 20102 28888 20154
rect 1104 20080 28888 20102
rect 4430 20040 4436 20052
rect 4391 20012 4436 20040
rect 4430 20000 4436 20012
rect 4488 20000 4494 20052
rect 5074 20000 5080 20052
rect 5132 20040 5138 20052
rect 5261 20043 5319 20049
rect 5261 20040 5273 20043
rect 5132 20012 5273 20040
rect 5132 20000 5138 20012
rect 5261 20009 5273 20012
rect 5307 20009 5319 20043
rect 5626 20040 5632 20052
rect 5587 20012 5632 20040
rect 5261 20003 5319 20009
rect 5626 20000 5632 20012
rect 5684 20000 5690 20052
rect 11790 20000 11796 20052
rect 11848 20040 11854 20052
rect 12345 20043 12403 20049
rect 12345 20040 12357 20043
rect 11848 20012 12357 20040
rect 11848 20000 11854 20012
rect 12345 20009 12357 20012
rect 12391 20009 12403 20043
rect 16666 20040 16672 20052
rect 16627 20012 16672 20040
rect 12345 20003 12403 20009
rect 16666 20000 16672 20012
rect 16724 20040 16730 20052
rect 17221 20043 17279 20049
rect 17221 20040 17233 20043
rect 16724 20012 17233 20040
rect 16724 20000 16730 20012
rect 17221 20009 17233 20012
rect 17267 20009 17279 20043
rect 17586 20040 17592 20052
rect 17499 20012 17592 20040
rect 17221 20003 17279 20009
rect 17586 20000 17592 20012
rect 17644 20040 17650 20052
rect 18785 20043 18843 20049
rect 18785 20040 18797 20043
rect 17644 20012 18797 20040
rect 17644 20000 17650 20012
rect 18785 20009 18797 20012
rect 18831 20009 18843 20043
rect 18785 20003 18843 20009
rect 17494 19932 17500 19984
rect 17552 19972 17558 19984
rect 18233 19975 18291 19981
rect 18233 19972 18245 19975
rect 17552 19944 18245 19972
rect 17552 19932 17558 19944
rect 18233 19941 18245 19944
rect 18279 19972 18291 19975
rect 18690 19972 18696 19984
rect 18279 19944 18696 19972
rect 18279 19941 18291 19944
rect 18233 19935 18291 19941
rect 18690 19932 18696 19944
rect 18748 19932 18754 19984
rect 4062 19864 4068 19916
rect 4120 19904 4126 19916
rect 4249 19907 4307 19913
rect 4249 19904 4261 19907
rect 4120 19876 4261 19904
rect 4120 19864 4126 19876
rect 4249 19873 4261 19876
rect 4295 19873 4307 19907
rect 4249 19867 4307 19873
rect 11793 19907 11851 19913
rect 11793 19873 11805 19907
rect 11839 19904 11851 19907
rect 12158 19904 12164 19916
rect 11839 19876 12164 19904
rect 11839 19873 11851 19876
rect 11793 19867 11851 19873
rect 12158 19864 12164 19876
rect 12216 19904 12222 19916
rect 12253 19907 12311 19913
rect 12253 19904 12265 19907
rect 12216 19876 12265 19904
rect 12216 19864 12222 19876
rect 12253 19873 12265 19876
rect 12299 19873 12311 19907
rect 12253 19867 12311 19873
rect 19153 19907 19211 19913
rect 19153 19873 19165 19907
rect 19199 19904 19211 19907
rect 19610 19904 19616 19916
rect 19199 19876 19616 19904
rect 19199 19873 19211 19876
rect 19153 19867 19211 19873
rect 19610 19864 19616 19876
rect 19668 19864 19674 19916
rect 26881 19907 26939 19913
rect 26881 19873 26893 19907
rect 26927 19904 26939 19907
rect 27246 19904 27252 19916
rect 26927 19876 27252 19904
rect 26927 19873 26939 19876
rect 26881 19867 26939 19873
rect 27246 19864 27252 19876
rect 27304 19864 27310 19916
rect 5718 19836 5724 19848
rect 5679 19808 5724 19836
rect 5718 19796 5724 19808
rect 5776 19796 5782 19848
rect 5813 19839 5871 19845
rect 5813 19805 5825 19839
rect 5859 19805 5871 19839
rect 11422 19836 11428 19848
rect 11335 19808 11428 19836
rect 5813 19799 5871 19805
rect 5828 19768 5856 19799
rect 11422 19796 11428 19808
rect 11480 19836 11486 19848
rect 12437 19839 12495 19845
rect 12437 19836 12449 19839
rect 11480 19808 12449 19836
rect 11480 19796 11486 19808
rect 12437 19805 12449 19808
rect 12483 19805 12495 19839
rect 17678 19836 17684 19848
rect 17639 19808 17684 19836
rect 12437 19799 12495 19805
rect 17678 19796 17684 19808
rect 17736 19796 17742 19848
rect 17770 19796 17776 19848
rect 17828 19836 17834 19848
rect 19242 19836 19248 19848
rect 17828 19808 17873 19836
rect 19203 19808 19248 19836
rect 17828 19796 17834 19808
rect 19242 19796 19248 19808
rect 19300 19796 19306 19848
rect 19337 19839 19395 19845
rect 19337 19805 19349 19839
rect 19383 19805 19395 19839
rect 26970 19836 26976 19848
rect 26931 19808 26976 19836
rect 19337 19799 19395 19805
rect 5368 19740 5856 19768
rect 5368 19712 5396 19740
rect 10962 19728 10968 19780
rect 11020 19768 11026 19780
rect 11885 19771 11943 19777
rect 11885 19768 11897 19771
rect 11020 19740 11897 19768
rect 11020 19728 11026 19740
rect 11885 19737 11897 19740
rect 11931 19737 11943 19771
rect 11885 19731 11943 19737
rect 19150 19728 19156 19780
rect 19208 19768 19214 19780
rect 19352 19768 19380 19799
rect 26970 19796 26976 19808
rect 27028 19796 27034 19848
rect 27157 19839 27215 19845
rect 27157 19805 27169 19839
rect 27203 19836 27215 19839
rect 27430 19836 27436 19848
rect 27203 19808 27436 19836
rect 27203 19805 27215 19808
rect 27157 19799 27215 19805
rect 27430 19796 27436 19808
rect 27488 19796 27494 19848
rect 19208 19740 19380 19768
rect 19208 19728 19214 19740
rect 3513 19703 3571 19709
rect 3513 19669 3525 19703
rect 3559 19700 3571 19703
rect 3878 19700 3884 19712
rect 3559 19672 3884 19700
rect 3559 19669 3571 19672
rect 3513 19663 3571 19669
rect 3878 19660 3884 19672
rect 3936 19660 3942 19712
rect 5077 19703 5135 19709
rect 5077 19669 5089 19703
rect 5123 19700 5135 19703
rect 5350 19700 5356 19712
rect 5123 19672 5356 19700
rect 5123 19669 5135 19672
rect 5077 19663 5135 19669
rect 5350 19660 5356 19672
rect 5408 19660 5414 19712
rect 5534 19660 5540 19712
rect 5592 19700 5598 19712
rect 6273 19703 6331 19709
rect 6273 19700 6285 19703
rect 5592 19672 6285 19700
rect 5592 19660 5598 19672
rect 6273 19669 6285 19672
rect 6319 19669 6331 19703
rect 10870 19700 10876 19712
rect 10831 19672 10876 19700
rect 6273 19663 6331 19669
rect 10870 19660 10876 19672
rect 10928 19660 10934 19712
rect 12986 19700 12992 19712
rect 12947 19672 12992 19700
rect 12986 19660 12992 19672
rect 13044 19660 13050 19712
rect 15102 19700 15108 19712
rect 15015 19672 15108 19700
rect 15102 19660 15108 19672
rect 15160 19700 15166 19712
rect 15562 19700 15568 19712
rect 15160 19672 15568 19700
rect 15160 19660 15166 19672
rect 15562 19660 15568 19672
rect 15620 19660 15626 19712
rect 18322 19660 18328 19712
rect 18380 19700 18386 19712
rect 18601 19703 18659 19709
rect 18601 19700 18613 19703
rect 18380 19672 18613 19700
rect 18380 19660 18386 19672
rect 18601 19669 18613 19672
rect 18647 19669 18659 19703
rect 18601 19663 18659 19669
rect 19610 19660 19616 19712
rect 19668 19700 19674 19712
rect 19797 19703 19855 19709
rect 19797 19700 19809 19703
rect 19668 19672 19809 19700
rect 19668 19660 19674 19672
rect 19797 19669 19809 19672
rect 19843 19669 19855 19703
rect 25406 19700 25412 19712
rect 25367 19672 25412 19700
rect 19797 19663 19855 19669
rect 25406 19660 25412 19672
rect 25464 19660 25470 19712
rect 26510 19700 26516 19712
rect 26471 19672 26516 19700
rect 26510 19660 26516 19672
rect 26568 19660 26574 19712
rect 1104 19610 28888 19632
rect 1104 19558 5982 19610
rect 6034 19558 6046 19610
rect 6098 19558 6110 19610
rect 6162 19558 6174 19610
rect 6226 19558 15982 19610
rect 16034 19558 16046 19610
rect 16098 19558 16110 19610
rect 16162 19558 16174 19610
rect 16226 19558 25982 19610
rect 26034 19558 26046 19610
rect 26098 19558 26110 19610
rect 26162 19558 26174 19610
rect 26226 19558 28888 19610
rect 1104 19536 28888 19558
rect 4985 19499 5043 19505
rect 4985 19465 4997 19499
rect 5031 19496 5043 19499
rect 5074 19496 5080 19508
rect 5031 19468 5080 19496
rect 5031 19465 5043 19468
rect 4985 19459 5043 19465
rect 5074 19456 5080 19468
rect 5132 19456 5138 19508
rect 5626 19456 5632 19508
rect 5684 19496 5690 19508
rect 5997 19499 6055 19505
rect 5997 19496 6009 19499
rect 5684 19468 6009 19496
rect 5684 19456 5690 19468
rect 5997 19465 6009 19468
rect 6043 19496 6055 19499
rect 6730 19496 6736 19508
rect 6043 19468 6736 19496
rect 6043 19465 6055 19468
rect 5997 19459 6055 19465
rect 6730 19456 6736 19468
rect 6788 19456 6794 19508
rect 10778 19496 10784 19508
rect 10739 19468 10784 19496
rect 10778 19456 10784 19468
rect 10836 19456 10842 19508
rect 13630 19456 13636 19508
rect 13688 19496 13694 19508
rect 13906 19496 13912 19508
rect 13688 19468 13912 19496
rect 13688 19456 13694 19468
rect 13906 19456 13912 19468
rect 13964 19456 13970 19508
rect 16577 19499 16635 19505
rect 16577 19465 16589 19499
rect 16623 19496 16635 19499
rect 17586 19496 17592 19508
rect 16623 19468 17592 19496
rect 16623 19465 16635 19468
rect 16577 19459 16635 19465
rect 17586 19456 17592 19468
rect 17644 19456 17650 19508
rect 18690 19456 18696 19508
rect 18748 19496 18754 19508
rect 18969 19499 19027 19505
rect 18969 19496 18981 19499
rect 18748 19468 18981 19496
rect 18748 19456 18754 19468
rect 18969 19465 18981 19468
rect 19015 19465 19027 19499
rect 18969 19459 19027 19465
rect 3329 19363 3387 19369
rect 3329 19329 3341 19363
rect 3375 19360 3387 19363
rect 3694 19360 3700 19372
rect 3375 19332 3700 19360
rect 3375 19329 3387 19332
rect 3329 19323 3387 19329
rect 3694 19320 3700 19332
rect 3752 19360 3758 19372
rect 3973 19363 4031 19369
rect 3973 19360 3985 19363
rect 3752 19332 3985 19360
rect 3752 19320 3758 19332
rect 3973 19329 3985 19332
rect 4019 19329 4031 19363
rect 4982 19360 4988 19372
rect 3973 19323 4031 19329
rect 4080 19332 4988 19360
rect 2961 19295 3019 19301
rect 2961 19261 2973 19295
rect 3007 19292 3019 19295
rect 3789 19295 3847 19301
rect 3789 19292 3801 19295
rect 3007 19264 3801 19292
rect 3007 19261 3019 19264
rect 2961 19255 3019 19261
rect 3789 19261 3801 19264
rect 3835 19292 3847 19295
rect 4080 19292 4108 19332
rect 4982 19320 4988 19332
rect 5040 19320 5046 19372
rect 5350 19320 5356 19372
rect 5408 19360 5414 19372
rect 5537 19363 5595 19369
rect 5537 19360 5549 19363
rect 5408 19332 5549 19360
rect 5408 19320 5414 19332
rect 5537 19329 5549 19332
rect 5583 19360 5595 19363
rect 6365 19363 6423 19369
rect 6365 19360 6377 19363
rect 5583 19332 6377 19360
rect 5583 19329 5595 19332
rect 5537 19323 5595 19329
rect 6365 19329 6377 19332
rect 6411 19329 6423 19363
rect 6365 19323 6423 19329
rect 10870 19320 10876 19372
rect 10928 19360 10934 19372
rect 11330 19360 11336 19372
rect 10928 19332 11100 19360
rect 11291 19332 11336 19360
rect 10928 19320 10934 19332
rect 5442 19292 5448 19304
rect 3835 19264 4108 19292
rect 5403 19264 5448 19292
rect 3835 19261 3847 19264
rect 3789 19255 3847 19261
rect 5442 19252 5448 19264
rect 5500 19252 5506 19304
rect 8294 19252 8300 19304
rect 8352 19292 8358 19304
rect 8849 19295 8907 19301
rect 8849 19292 8861 19295
rect 8352 19264 8861 19292
rect 8352 19252 8358 19264
rect 8849 19261 8861 19264
rect 8895 19292 8907 19295
rect 9309 19295 9367 19301
rect 9309 19292 9321 19295
rect 8895 19264 9321 19292
rect 8895 19261 8907 19264
rect 8849 19255 8907 19261
rect 9309 19261 9321 19264
rect 9355 19261 9367 19295
rect 9309 19255 9367 19261
rect 9861 19295 9919 19301
rect 9861 19261 9873 19295
rect 9907 19292 9919 19295
rect 10134 19292 10140 19304
rect 9907 19264 10140 19292
rect 9907 19261 9919 19264
rect 9861 19255 9919 19261
rect 10134 19252 10140 19264
rect 10192 19292 10198 19304
rect 10962 19292 10968 19304
rect 10192 19264 10968 19292
rect 10192 19252 10198 19264
rect 10962 19252 10968 19264
rect 11020 19252 11026 19304
rect 11072 19292 11100 19332
rect 11330 19320 11336 19332
rect 11388 19320 11394 19372
rect 15562 19360 15568 19372
rect 15523 19332 15568 19360
rect 15562 19320 15568 19332
rect 15620 19320 15626 19372
rect 11241 19295 11299 19301
rect 11241 19292 11253 19295
rect 11072 19264 11253 19292
rect 11241 19261 11253 19264
rect 11287 19292 11299 19295
rect 11882 19292 11888 19304
rect 11287 19264 11888 19292
rect 11287 19261 11299 19264
rect 11241 19255 11299 19261
rect 11882 19252 11888 19264
rect 11940 19252 11946 19304
rect 12526 19252 12532 19304
rect 12584 19301 12590 19304
rect 12584 19292 12594 19301
rect 14826 19292 14832 19304
rect 12584 19264 12629 19292
rect 14739 19264 14832 19292
rect 12584 19255 12594 19264
rect 12584 19252 12590 19255
rect 14826 19252 14832 19264
rect 14884 19292 14890 19304
rect 18417 19295 18475 19301
rect 14884 19264 15516 19292
rect 14884 19252 14890 19264
rect 4062 19224 4068 19236
rect 3436 19196 4068 19224
rect 3436 19165 3464 19196
rect 4062 19184 4068 19196
rect 4120 19184 4126 19236
rect 5718 19224 5724 19236
rect 4448 19196 5724 19224
rect 4448 19168 4476 19196
rect 5718 19184 5724 19196
rect 5776 19184 5782 19236
rect 10321 19227 10379 19233
rect 10321 19193 10333 19227
rect 10367 19224 10379 19227
rect 11149 19227 11207 19233
rect 11149 19224 11161 19227
rect 10367 19196 11161 19224
rect 10367 19193 10379 19196
rect 10321 19187 10379 19193
rect 11149 19193 11161 19196
rect 11195 19224 11207 19227
rect 12250 19224 12256 19236
rect 11195 19196 12256 19224
rect 11195 19193 11207 19196
rect 11149 19187 11207 19193
rect 12250 19184 12256 19196
rect 12308 19184 12314 19236
rect 12710 19184 12716 19236
rect 12768 19233 12774 19236
rect 12768 19227 12832 19233
rect 12768 19193 12786 19227
rect 12820 19193 12832 19227
rect 12768 19187 12832 19193
rect 12768 19184 12774 19187
rect 14918 19184 14924 19236
rect 14976 19224 14982 19236
rect 15381 19227 15439 19233
rect 15381 19224 15393 19227
rect 14976 19196 15393 19224
rect 14976 19184 14982 19196
rect 15381 19193 15393 19196
rect 15427 19193 15439 19227
rect 15381 19187 15439 19193
rect 3421 19159 3479 19165
rect 3421 19125 3433 19159
rect 3467 19125 3479 19159
rect 3878 19156 3884 19168
rect 3839 19128 3884 19156
rect 3421 19119 3479 19125
rect 3878 19116 3884 19128
rect 3936 19116 3942 19168
rect 4430 19156 4436 19168
rect 4391 19128 4436 19156
rect 4430 19116 4436 19128
rect 4488 19116 4494 19168
rect 4614 19116 4620 19168
rect 4672 19156 4678 19168
rect 4801 19159 4859 19165
rect 4801 19156 4813 19159
rect 4672 19128 4813 19156
rect 4672 19116 4678 19128
rect 4801 19125 4813 19128
rect 4847 19156 4859 19159
rect 5353 19159 5411 19165
rect 5353 19156 5365 19159
rect 4847 19128 5365 19156
rect 4847 19125 4859 19128
rect 4801 19119 4859 19125
rect 5353 19125 5365 19128
rect 5399 19125 5411 19159
rect 6822 19156 6828 19168
rect 6783 19128 6828 19156
rect 5353 19119 5411 19125
rect 6822 19116 6828 19128
rect 6880 19116 6886 19168
rect 9030 19156 9036 19168
rect 8991 19128 9036 19156
rect 9030 19116 9036 19128
rect 9088 19116 9094 19168
rect 10410 19116 10416 19168
rect 10468 19156 10474 19168
rect 10597 19159 10655 19165
rect 10597 19156 10609 19159
rect 10468 19128 10609 19156
rect 10468 19116 10474 19128
rect 10597 19125 10609 19128
rect 10643 19156 10655 19159
rect 11330 19156 11336 19168
rect 10643 19128 11336 19156
rect 10643 19125 10655 19128
rect 10597 19119 10655 19125
rect 11330 19116 11336 19128
rect 11388 19116 11394 19168
rect 11790 19116 11796 19168
rect 11848 19156 11854 19168
rect 11885 19159 11943 19165
rect 11885 19156 11897 19159
rect 11848 19128 11897 19156
rect 11848 19116 11854 19128
rect 11885 19125 11897 19128
rect 11931 19125 11943 19159
rect 11885 19119 11943 19125
rect 12526 19116 12532 19168
rect 12584 19156 12590 19168
rect 12986 19156 12992 19168
rect 12584 19128 12992 19156
rect 12584 19116 12590 19128
rect 12986 19116 12992 19128
rect 13044 19116 13050 19168
rect 15010 19156 15016 19168
rect 14971 19128 15016 19156
rect 15010 19116 15016 19128
rect 15068 19116 15074 19168
rect 15488 19165 15516 19264
rect 18417 19261 18429 19295
rect 18463 19292 18475 19295
rect 18598 19292 18604 19304
rect 18463 19264 18604 19292
rect 18463 19261 18475 19264
rect 18417 19255 18475 19261
rect 18598 19252 18604 19264
rect 18656 19292 18662 19304
rect 19150 19292 19156 19304
rect 18656 19264 19156 19292
rect 18656 19252 18662 19264
rect 19150 19252 19156 19264
rect 19208 19252 19214 19304
rect 19521 19295 19579 19301
rect 19521 19261 19533 19295
rect 19567 19261 19579 19295
rect 25317 19295 25375 19301
rect 25317 19292 25329 19295
rect 19521 19255 19579 19261
rect 25148 19264 25329 19292
rect 16945 19227 17003 19233
rect 16945 19193 16957 19227
rect 16991 19224 17003 19227
rect 17678 19224 17684 19236
rect 16991 19196 17684 19224
rect 16991 19193 17003 19196
rect 16945 19187 17003 19193
rect 17678 19184 17684 19196
rect 17736 19184 17742 19236
rect 17865 19227 17923 19233
rect 17865 19193 17877 19227
rect 17911 19224 17923 19227
rect 19242 19224 19248 19236
rect 17911 19196 19248 19224
rect 17911 19193 17923 19196
rect 17865 19187 17923 19193
rect 19242 19184 19248 19196
rect 19300 19184 19306 19236
rect 15473 19159 15531 19165
rect 15473 19125 15485 19159
rect 15519 19156 15531 19159
rect 16390 19156 16396 19168
rect 15519 19128 16396 19156
rect 15519 19125 15531 19128
rect 15473 19119 15531 19125
rect 16390 19116 16396 19128
rect 16448 19116 16454 19168
rect 17313 19159 17371 19165
rect 17313 19125 17325 19159
rect 17359 19156 17371 19159
rect 17770 19156 17776 19168
rect 17359 19128 17776 19156
rect 17359 19125 17371 19128
rect 17313 19119 17371 19125
rect 17770 19116 17776 19128
rect 17828 19116 17834 19168
rect 18509 19159 18567 19165
rect 18509 19125 18521 19159
rect 18555 19156 18567 19159
rect 18874 19156 18880 19168
rect 18555 19128 18880 19156
rect 18555 19125 18567 19128
rect 18509 19119 18567 19125
rect 18874 19116 18880 19128
rect 18932 19116 18938 19168
rect 19429 19159 19487 19165
rect 19429 19125 19441 19159
rect 19475 19156 19487 19159
rect 19536 19156 19564 19255
rect 19794 19233 19800 19236
rect 19788 19224 19800 19233
rect 19755 19196 19800 19224
rect 19788 19187 19800 19196
rect 19794 19184 19800 19187
rect 19852 19184 19858 19236
rect 19886 19156 19892 19168
rect 19475 19128 19892 19156
rect 19475 19125 19487 19128
rect 19429 19119 19487 19125
rect 19886 19116 19892 19128
rect 19944 19116 19950 19168
rect 20714 19116 20720 19168
rect 20772 19156 20778 19168
rect 20901 19159 20959 19165
rect 20901 19156 20913 19159
rect 20772 19128 20913 19156
rect 20772 19116 20778 19128
rect 20901 19125 20913 19128
rect 20947 19125 20959 19159
rect 20901 19119 20959 19125
rect 24302 19116 24308 19168
rect 24360 19156 24366 19168
rect 25148 19165 25176 19264
rect 25317 19261 25329 19264
rect 25363 19261 25375 19295
rect 25317 19255 25375 19261
rect 25406 19252 25412 19304
rect 25464 19292 25470 19304
rect 25573 19295 25631 19301
rect 25573 19292 25585 19295
rect 25464 19264 25585 19292
rect 25464 19252 25470 19264
rect 25573 19261 25585 19264
rect 25619 19292 25631 19295
rect 25866 19292 25872 19304
rect 25619 19264 25872 19292
rect 25619 19261 25631 19264
rect 25573 19255 25631 19261
rect 25866 19252 25872 19264
rect 25924 19252 25930 19304
rect 27430 19252 27436 19304
rect 27488 19292 27494 19304
rect 27985 19295 28043 19301
rect 27985 19292 27997 19295
rect 27488 19264 27997 19292
rect 27488 19252 27494 19264
rect 27985 19261 27997 19264
rect 28031 19261 28043 19295
rect 27985 19255 28043 19261
rect 25133 19159 25191 19165
rect 25133 19156 25145 19159
rect 24360 19128 25145 19156
rect 24360 19116 24366 19128
rect 25133 19125 25145 19128
rect 25179 19125 25191 19159
rect 25133 19119 25191 19125
rect 25406 19116 25412 19168
rect 25464 19156 25470 19168
rect 26697 19159 26755 19165
rect 26697 19156 26709 19159
rect 25464 19128 26709 19156
rect 25464 19116 25470 19128
rect 26697 19125 26709 19128
rect 26743 19125 26755 19159
rect 27246 19156 27252 19168
rect 27207 19128 27252 19156
rect 26697 19119 26755 19125
rect 27246 19116 27252 19128
rect 27304 19116 27310 19168
rect 27614 19156 27620 19168
rect 27575 19128 27620 19156
rect 27614 19116 27620 19128
rect 27672 19116 27678 19168
rect 1104 19066 28888 19088
rect 1104 19014 10982 19066
rect 11034 19014 11046 19066
rect 11098 19014 11110 19066
rect 11162 19014 11174 19066
rect 11226 19014 20982 19066
rect 21034 19014 21046 19066
rect 21098 19014 21110 19066
rect 21162 19014 21174 19066
rect 21226 19014 28888 19066
rect 1104 18992 28888 19014
rect 2406 18952 2412 18964
rect 2367 18924 2412 18952
rect 2406 18912 2412 18924
rect 2464 18912 2470 18964
rect 3881 18955 3939 18961
rect 3881 18921 3893 18955
rect 3927 18952 3939 18955
rect 4062 18952 4068 18964
rect 3927 18924 4068 18952
rect 3927 18921 3939 18924
rect 3881 18915 3939 18921
rect 4062 18912 4068 18924
rect 4120 18912 4126 18964
rect 5626 18912 5632 18964
rect 5684 18952 5690 18964
rect 6086 18952 6092 18964
rect 5684 18924 6092 18952
rect 5684 18912 5690 18924
rect 6086 18912 6092 18924
rect 6144 18912 6150 18964
rect 7190 18952 7196 18964
rect 7151 18924 7196 18952
rect 7190 18912 7196 18924
rect 7248 18912 7254 18964
rect 7650 18952 7656 18964
rect 7611 18924 7656 18952
rect 7650 18912 7656 18924
rect 7708 18912 7714 18964
rect 9766 18952 9772 18964
rect 9727 18924 9772 18952
rect 9766 18912 9772 18924
rect 9824 18912 9830 18964
rect 10134 18952 10140 18964
rect 10095 18924 10140 18952
rect 10134 18912 10140 18924
rect 10192 18912 10198 18964
rect 11330 18912 11336 18964
rect 11388 18952 11394 18964
rect 12710 18952 12716 18964
rect 11388 18924 12716 18952
rect 11388 18912 11394 18924
rect 12710 18912 12716 18924
rect 12768 18952 12774 18964
rect 13265 18955 13323 18961
rect 13265 18952 13277 18955
rect 12768 18924 13277 18952
rect 12768 18912 12774 18924
rect 13265 18921 13277 18924
rect 13311 18921 13323 18955
rect 13265 18915 13323 18921
rect 13906 18912 13912 18964
rect 13964 18952 13970 18964
rect 14185 18955 14243 18961
rect 14185 18952 14197 18955
rect 13964 18924 14197 18952
rect 13964 18912 13970 18924
rect 14185 18921 14197 18924
rect 14231 18921 14243 18955
rect 14185 18915 14243 18921
rect 18230 18912 18236 18964
rect 18288 18952 18294 18964
rect 18417 18955 18475 18961
rect 18417 18952 18429 18955
rect 18288 18924 18429 18952
rect 18288 18912 18294 18924
rect 18417 18921 18429 18924
rect 18463 18921 18475 18955
rect 18417 18915 18475 18921
rect 18690 18912 18696 18964
rect 18748 18952 18754 18964
rect 18785 18955 18843 18961
rect 18785 18952 18797 18955
rect 18748 18924 18797 18952
rect 18748 18912 18754 18924
rect 18785 18921 18797 18924
rect 18831 18921 18843 18955
rect 18785 18915 18843 18921
rect 18969 18955 19027 18961
rect 18969 18921 18981 18955
rect 19015 18952 19027 18955
rect 19242 18952 19248 18964
rect 19015 18924 19248 18952
rect 19015 18921 19027 18924
rect 18969 18915 19027 18921
rect 4617 18887 4675 18893
rect 4617 18853 4629 18887
rect 4663 18884 4675 18887
rect 4890 18884 4896 18896
rect 4663 18856 4896 18884
rect 4663 18853 4675 18856
rect 4617 18847 4675 18853
rect 4890 18844 4896 18856
rect 4948 18893 4954 18896
rect 4948 18887 5012 18893
rect 4948 18853 4966 18887
rect 5000 18884 5012 18887
rect 5534 18884 5540 18896
rect 5000 18856 5540 18884
rect 5000 18853 5012 18856
rect 4948 18847 5012 18853
rect 4948 18844 4954 18847
rect 5534 18844 5540 18856
rect 5592 18844 5598 18896
rect 11422 18844 11428 18896
rect 11480 18884 11486 18896
rect 11578 18887 11636 18893
rect 11578 18884 11590 18887
rect 11480 18856 11590 18884
rect 11480 18844 11486 18856
rect 11578 18853 11590 18856
rect 11624 18853 11636 18887
rect 18800 18884 18828 18915
rect 19242 18912 19248 18924
rect 19300 18912 19306 18964
rect 20530 18912 20536 18964
rect 20588 18952 20594 18964
rect 20901 18955 20959 18961
rect 20901 18952 20913 18955
rect 20588 18924 20913 18952
rect 20588 18912 20594 18924
rect 20901 18921 20913 18924
rect 20947 18921 20959 18955
rect 20901 18915 20959 18921
rect 22649 18955 22707 18961
rect 22649 18921 22661 18955
rect 22695 18952 22707 18955
rect 23382 18952 23388 18964
rect 22695 18924 23388 18952
rect 22695 18921 22707 18924
rect 22649 18915 22707 18921
rect 23382 18912 23388 18924
rect 23440 18912 23446 18964
rect 24854 18952 24860 18964
rect 24815 18924 24860 18952
rect 24854 18912 24860 18924
rect 24912 18912 24918 18964
rect 26329 18955 26387 18961
rect 26329 18921 26341 18955
rect 26375 18952 26387 18955
rect 26510 18952 26516 18964
rect 26375 18924 26516 18952
rect 26375 18921 26387 18924
rect 26329 18915 26387 18921
rect 26510 18912 26516 18924
rect 26568 18952 26574 18964
rect 26973 18955 27031 18961
rect 26973 18952 26985 18955
rect 26568 18924 26985 18952
rect 26568 18912 26574 18924
rect 26973 18921 26985 18924
rect 27019 18921 27031 18955
rect 26973 18915 27031 18921
rect 19794 18884 19800 18896
rect 18800 18856 19800 18884
rect 11578 18847 11636 18853
rect 2222 18816 2228 18828
rect 2183 18788 2228 18816
rect 2222 18776 2228 18788
rect 2280 18816 2286 18828
rect 2685 18819 2743 18825
rect 2685 18816 2697 18819
rect 2280 18788 2697 18816
rect 2280 18776 2286 18788
rect 2685 18785 2697 18788
rect 2731 18785 2743 18819
rect 7558 18816 7564 18828
rect 7519 18788 7564 18816
rect 2685 18779 2743 18785
rect 7558 18776 7564 18788
rect 7616 18776 7622 18828
rect 9493 18819 9551 18825
rect 9493 18785 9505 18819
rect 9539 18816 9551 18819
rect 10226 18816 10232 18828
rect 9539 18788 10232 18816
rect 9539 18785 9551 18788
rect 9493 18779 9551 18785
rect 10226 18776 10232 18788
rect 10284 18776 10290 18828
rect 11333 18819 11391 18825
rect 11333 18785 11345 18819
rect 11379 18816 11391 18819
rect 12526 18816 12532 18828
rect 11379 18788 12532 18816
rect 11379 18785 11391 18788
rect 11333 18779 11391 18785
rect 12526 18776 12532 18788
rect 12584 18776 12590 18828
rect 16758 18825 16764 18828
rect 16752 18816 16764 18825
rect 16719 18788 16764 18816
rect 16752 18779 16764 18788
rect 16758 18776 16764 18779
rect 16816 18776 16822 18828
rect 19058 18776 19064 18828
rect 19116 18816 19122 18828
rect 19337 18819 19395 18825
rect 19337 18816 19349 18819
rect 19116 18788 19349 18816
rect 19116 18776 19122 18788
rect 19337 18785 19349 18788
rect 19383 18785 19395 18819
rect 19337 18779 19395 18785
rect 4706 18748 4712 18760
rect 4667 18720 4712 18748
rect 4706 18708 4712 18720
rect 4764 18708 4770 18760
rect 6914 18708 6920 18760
rect 6972 18748 6978 18760
rect 7745 18751 7803 18757
rect 7745 18748 7757 18751
rect 6972 18720 7757 18748
rect 6972 18708 6978 18720
rect 7745 18717 7757 18720
rect 7791 18748 7803 18751
rect 7834 18748 7840 18760
rect 7791 18720 7840 18748
rect 7791 18717 7803 18720
rect 7745 18711 7803 18717
rect 7834 18708 7840 18720
rect 7892 18708 7898 18760
rect 10318 18748 10324 18760
rect 10279 18720 10324 18748
rect 10318 18708 10324 18720
rect 10376 18708 10382 18760
rect 16482 18748 16488 18760
rect 16443 18720 16488 18748
rect 16482 18708 16488 18720
rect 16540 18708 16546 18760
rect 19426 18748 19432 18760
rect 19387 18720 19432 18748
rect 19426 18708 19432 18720
rect 19484 18708 19490 18760
rect 19536 18757 19564 18856
rect 19794 18844 19800 18856
rect 19852 18884 19858 18896
rect 20162 18884 20168 18896
rect 19852 18856 20168 18884
rect 19852 18844 19858 18856
rect 20162 18844 20168 18856
rect 20220 18884 20226 18896
rect 20349 18887 20407 18893
rect 20349 18884 20361 18887
rect 20220 18856 20361 18884
rect 20220 18844 20226 18856
rect 20349 18853 20361 18856
rect 20395 18853 20407 18887
rect 20349 18847 20407 18853
rect 21269 18819 21327 18825
rect 21269 18785 21281 18819
rect 21315 18816 21327 18819
rect 22462 18816 22468 18828
rect 21315 18788 22324 18816
rect 22423 18788 22468 18816
rect 21315 18785 21327 18788
rect 21269 18779 21327 18785
rect 19521 18751 19579 18757
rect 19521 18717 19533 18751
rect 19567 18717 19579 18751
rect 19521 18711 19579 18717
rect 20714 18708 20720 18760
rect 20772 18748 20778 18760
rect 21361 18751 21419 18757
rect 21361 18748 21373 18751
rect 20772 18720 21373 18748
rect 20772 18708 20778 18720
rect 21361 18717 21373 18720
rect 21407 18717 21419 18751
rect 21361 18711 21419 18717
rect 21450 18708 21456 18760
rect 21508 18748 21514 18760
rect 22296 18748 22324 18788
rect 22462 18776 22468 18788
rect 22520 18776 22526 18828
rect 25225 18819 25283 18825
rect 25225 18785 25237 18819
rect 25271 18785 25283 18819
rect 25225 18779 25283 18785
rect 25317 18819 25375 18825
rect 25317 18785 25329 18819
rect 25363 18816 25375 18819
rect 25498 18816 25504 18828
rect 25363 18788 25504 18816
rect 25363 18785 25375 18788
rect 25317 18779 25375 18785
rect 22646 18748 22652 18760
rect 21508 18720 21553 18748
rect 22296 18720 22652 18748
rect 21508 18708 21514 18720
rect 22646 18708 22652 18720
rect 22704 18708 22710 18760
rect 24765 18683 24823 18689
rect 24765 18649 24777 18683
rect 24811 18680 24823 18683
rect 25240 18680 25268 18779
rect 25498 18776 25504 18788
rect 25556 18776 25562 18828
rect 25961 18819 26019 18825
rect 25961 18785 25973 18819
rect 26007 18816 26019 18819
rect 26510 18816 26516 18828
rect 26007 18788 26516 18816
rect 26007 18785 26019 18788
rect 25961 18779 26019 18785
rect 26510 18776 26516 18788
rect 26568 18816 26574 18828
rect 26881 18819 26939 18825
rect 26881 18816 26893 18819
rect 26568 18788 26893 18816
rect 26568 18776 26574 18788
rect 26881 18785 26893 18788
rect 26927 18785 26939 18819
rect 26881 18779 26939 18785
rect 25406 18748 25412 18760
rect 25367 18720 25412 18748
rect 25406 18708 25412 18720
rect 25464 18708 25470 18760
rect 25866 18708 25872 18760
rect 25924 18748 25930 18760
rect 27065 18751 27123 18757
rect 27065 18748 27077 18751
rect 25924 18720 27077 18748
rect 25924 18708 25930 18720
rect 27065 18717 27077 18720
rect 27111 18717 27123 18751
rect 27065 18711 27123 18717
rect 26513 18683 26571 18689
rect 26513 18680 26525 18683
rect 24811 18652 26525 18680
rect 24811 18649 24823 18652
rect 24765 18643 24823 18649
rect 26513 18649 26525 18652
rect 26559 18649 26571 18683
rect 26513 18643 26571 18649
rect 1854 18612 1860 18624
rect 1815 18584 1860 18612
rect 1854 18572 1860 18584
rect 1912 18572 1918 18624
rect 3421 18615 3479 18621
rect 3421 18581 3433 18615
rect 3467 18612 3479 18615
rect 3878 18612 3884 18624
rect 3467 18584 3884 18612
rect 3467 18581 3479 18584
rect 3421 18575 3479 18581
rect 3878 18572 3884 18584
rect 3936 18572 3942 18624
rect 6917 18615 6975 18621
rect 6917 18581 6929 18615
rect 6963 18612 6975 18615
rect 7098 18612 7104 18624
rect 6963 18584 7104 18612
rect 6963 18581 6975 18584
rect 6917 18575 6975 18581
rect 7098 18572 7104 18584
rect 7156 18572 7162 18624
rect 8570 18612 8576 18624
rect 8531 18584 8576 18612
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 8941 18615 8999 18621
rect 8941 18581 8953 18615
rect 8987 18612 8999 18615
rect 9030 18612 9036 18624
rect 8987 18584 9036 18612
rect 8987 18581 8999 18584
rect 8941 18575 8999 18581
rect 9030 18572 9036 18584
rect 9088 18572 9094 18624
rect 10778 18612 10784 18624
rect 10739 18584 10784 18612
rect 10778 18572 10784 18584
rect 10836 18572 10842 18624
rect 14918 18572 14924 18624
rect 14976 18612 14982 18624
rect 15013 18615 15071 18621
rect 15013 18612 15025 18615
rect 14976 18584 15025 18612
rect 14976 18572 14982 18584
rect 15013 18581 15025 18584
rect 15059 18581 15071 18615
rect 17862 18612 17868 18624
rect 17823 18584 17868 18612
rect 15013 18575 15071 18581
rect 17862 18572 17868 18584
rect 17920 18572 17926 18624
rect 19978 18612 19984 18624
rect 19939 18584 19984 18612
rect 19978 18572 19984 18584
rect 20036 18572 20042 18624
rect 22005 18615 22063 18621
rect 22005 18581 22017 18615
rect 22051 18612 22063 18615
rect 22094 18612 22100 18624
rect 22051 18584 22100 18612
rect 22051 18581 22063 18584
rect 22005 18575 22063 18581
rect 22094 18572 22100 18584
rect 22152 18572 22158 18624
rect 27338 18572 27344 18624
rect 27396 18612 27402 18624
rect 27525 18615 27583 18621
rect 27525 18612 27537 18615
rect 27396 18584 27537 18612
rect 27396 18572 27402 18584
rect 27525 18581 27537 18584
rect 27571 18581 27583 18615
rect 27525 18575 27583 18581
rect 1104 18522 28888 18544
rect 1104 18470 5982 18522
rect 6034 18470 6046 18522
rect 6098 18470 6110 18522
rect 6162 18470 6174 18522
rect 6226 18470 15982 18522
rect 16034 18470 16046 18522
rect 16098 18470 16110 18522
rect 16162 18470 16174 18522
rect 16226 18470 25982 18522
rect 26034 18470 26046 18522
rect 26098 18470 26110 18522
rect 26162 18470 26174 18522
rect 26226 18470 28888 18522
rect 1104 18448 28888 18470
rect 3329 18411 3387 18417
rect 3329 18377 3341 18411
rect 3375 18408 3387 18411
rect 3970 18408 3976 18420
rect 3375 18380 3976 18408
rect 3375 18377 3387 18380
rect 3329 18371 3387 18377
rect 3970 18368 3976 18380
rect 4028 18368 4034 18420
rect 4893 18411 4951 18417
rect 4893 18377 4905 18411
rect 4939 18408 4951 18411
rect 5442 18408 5448 18420
rect 4939 18380 5448 18408
rect 4939 18377 4951 18380
rect 4893 18371 4951 18377
rect 5442 18368 5448 18380
rect 5500 18368 5506 18420
rect 7834 18408 7840 18420
rect 7795 18380 7840 18408
rect 7834 18368 7840 18380
rect 7892 18368 7898 18420
rect 10226 18368 10232 18420
rect 10284 18408 10290 18420
rect 10781 18411 10839 18417
rect 10781 18408 10793 18411
rect 10284 18380 10793 18408
rect 10284 18368 10290 18380
rect 10781 18377 10793 18380
rect 10827 18377 10839 18411
rect 10781 18371 10839 18377
rect 11882 18368 11888 18420
rect 11940 18408 11946 18420
rect 12437 18411 12495 18417
rect 12437 18408 12449 18411
rect 11940 18380 12449 18408
rect 11940 18368 11946 18380
rect 12437 18377 12449 18380
rect 12483 18377 12495 18411
rect 12437 18371 12495 18377
rect 17678 18368 17684 18420
rect 17736 18408 17742 18420
rect 18049 18411 18107 18417
rect 18049 18408 18061 18411
rect 17736 18380 18061 18408
rect 17736 18368 17742 18380
rect 18049 18377 18061 18380
rect 18095 18377 18107 18411
rect 19610 18408 19616 18420
rect 19571 18380 19616 18408
rect 18049 18371 18107 18377
rect 19610 18368 19616 18380
rect 19668 18368 19674 18420
rect 24029 18411 24087 18417
rect 24029 18377 24041 18411
rect 24075 18408 24087 18411
rect 25498 18408 25504 18420
rect 24075 18380 25504 18408
rect 24075 18377 24087 18380
rect 24029 18371 24087 18377
rect 25498 18368 25504 18380
rect 25556 18408 25562 18420
rect 26973 18411 27031 18417
rect 26973 18408 26985 18411
rect 25556 18380 26985 18408
rect 25556 18368 25562 18380
rect 26973 18377 26985 18380
rect 27019 18377 27031 18411
rect 26973 18371 27031 18377
rect 6825 18343 6883 18349
rect 6825 18309 6837 18343
rect 6871 18340 6883 18343
rect 7558 18340 7564 18352
rect 6871 18312 7564 18340
rect 6871 18309 6883 18312
rect 6825 18303 6883 18309
rect 7558 18300 7564 18312
rect 7616 18300 7622 18352
rect 9861 18343 9919 18349
rect 9861 18309 9873 18343
rect 9907 18340 9919 18343
rect 10318 18340 10324 18352
rect 9907 18312 10324 18340
rect 9907 18309 9919 18312
rect 9861 18303 9919 18309
rect 10318 18300 10324 18312
rect 10376 18300 10382 18352
rect 10594 18340 10600 18352
rect 10555 18312 10600 18340
rect 10594 18300 10600 18312
rect 10652 18300 10658 18352
rect 16758 18300 16764 18352
rect 16816 18340 16822 18352
rect 16945 18343 17003 18349
rect 16945 18340 16957 18343
rect 16816 18312 16957 18340
rect 16816 18300 16822 18312
rect 16945 18309 16957 18312
rect 16991 18340 17003 18343
rect 17865 18343 17923 18349
rect 17865 18340 17877 18343
rect 16991 18312 17877 18340
rect 16991 18309 17003 18312
rect 16945 18303 17003 18309
rect 17865 18309 17877 18312
rect 17911 18340 17923 18343
rect 17911 18312 18644 18340
rect 17911 18309 17923 18312
rect 17865 18303 17923 18309
rect 18616 18284 18644 18312
rect 19978 18300 19984 18352
rect 20036 18340 20042 18352
rect 25866 18340 25872 18352
rect 20036 18312 20116 18340
rect 25827 18312 25872 18340
rect 20036 18300 20042 18312
rect 3878 18272 3884 18284
rect 3839 18244 3884 18272
rect 3878 18232 3884 18244
rect 3936 18272 3942 18284
rect 4154 18272 4160 18284
rect 3936 18244 4160 18272
rect 3936 18232 3942 18244
rect 4154 18232 4160 18244
rect 4212 18232 4218 18284
rect 4338 18232 4344 18284
rect 4396 18272 4402 18284
rect 5537 18275 5595 18281
rect 5537 18272 5549 18275
rect 4396 18244 5549 18272
rect 4396 18232 4402 18244
rect 5537 18241 5549 18244
rect 5583 18272 5595 18275
rect 5905 18275 5963 18281
rect 5905 18272 5917 18275
rect 5583 18244 5917 18272
rect 5583 18241 5595 18244
rect 5537 18235 5595 18241
rect 5905 18241 5917 18244
rect 5951 18241 5963 18275
rect 5905 18235 5963 18241
rect 7282 18232 7288 18284
rect 7340 18272 7346 18284
rect 7377 18275 7435 18281
rect 7377 18272 7389 18275
rect 7340 18244 7389 18272
rect 7340 18232 7346 18244
rect 7377 18241 7389 18244
rect 7423 18241 7435 18275
rect 9030 18272 9036 18284
rect 8991 18244 9036 18272
rect 7377 18235 7435 18241
rect 9030 18232 9036 18244
rect 9088 18232 9094 18284
rect 10229 18275 10287 18281
rect 10229 18241 10241 18275
rect 10275 18272 10287 18275
rect 11422 18272 11428 18284
rect 10275 18244 11428 18272
rect 10275 18241 10287 18244
rect 10229 18235 10287 18241
rect 11422 18232 11428 18244
rect 11480 18232 11486 18284
rect 11885 18275 11943 18281
rect 11885 18241 11897 18275
rect 11931 18272 11943 18275
rect 12526 18272 12532 18284
rect 11931 18244 12532 18272
rect 11931 18241 11943 18244
rect 11885 18235 11943 18241
rect 12526 18232 12532 18244
rect 12584 18272 12590 18284
rect 13078 18272 13084 18284
rect 12584 18244 12940 18272
rect 12991 18244 13084 18272
rect 12584 18232 12590 18244
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18173 1455 18207
rect 3694 18204 3700 18216
rect 3655 18176 3700 18204
rect 1397 18167 1455 18173
rect 1412 18136 1440 18167
rect 3694 18164 3700 18176
rect 3752 18164 3758 18216
rect 9582 18204 9588 18216
rect 4172 18176 9588 18204
rect 2041 18139 2099 18145
rect 2041 18136 2053 18139
rect 1412 18108 2053 18136
rect 2041 18105 2053 18108
rect 2087 18136 2099 18139
rect 4172 18136 4200 18176
rect 9582 18164 9588 18176
rect 9640 18164 9646 18216
rect 10594 18164 10600 18216
rect 10652 18204 10658 18216
rect 11146 18204 11152 18216
rect 10652 18176 11152 18204
rect 10652 18164 10658 18176
rect 11146 18164 11152 18176
rect 11204 18164 11210 18216
rect 12805 18207 12863 18213
rect 12805 18204 12817 18207
rect 12176 18176 12817 18204
rect 5258 18136 5264 18148
rect 2087 18108 4200 18136
rect 4356 18108 5264 18136
rect 2087 18105 2099 18108
rect 2041 18099 2099 18105
rect 1581 18071 1639 18077
rect 1581 18037 1593 18071
rect 1627 18068 1639 18071
rect 1670 18068 1676 18080
rect 1627 18040 1676 18068
rect 1627 18037 1639 18040
rect 1581 18031 1639 18037
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 2409 18071 2467 18077
rect 2409 18037 2421 18071
rect 2455 18068 2467 18071
rect 2498 18068 2504 18080
rect 2455 18040 2504 18068
rect 2455 18037 2467 18040
rect 2409 18031 2467 18037
rect 2498 18028 2504 18040
rect 2556 18028 2562 18080
rect 2682 18028 2688 18080
rect 2740 18068 2746 18080
rect 2777 18071 2835 18077
rect 2777 18068 2789 18071
rect 2740 18040 2789 18068
rect 2740 18028 2746 18040
rect 2777 18037 2789 18040
rect 2823 18037 2835 18071
rect 2777 18031 2835 18037
rect 3237 18071 3295 18077
rect 3237 18037 3249 18071
rect 3283 18068 3295 18071
rect 3602 18068 3608 18080
rect 3283 18040 3608 18068
rect 3283 18037 3295 18040
rect 3237 18031 3295 18037
rect 3602 18028 3608 18040
rect 3660 18068 3666 18080
rect 3789 18071 3847 18077
rect 3789 18068 3801 18071
rect 3660 18040 3801 18068
rect 3660 18028 3666 18040
rect 3789 18037 3801 18040
rect 3835 18037 3847 18071
rect 3789 18031 3847 18037
rect 4246 18028 4252 18080
rect 4304 18068 4310 18080
rect 4356 18077 4384 18108
rect 5258 18096 5264 18108
rect 5316 18096 5322 18148
rect 7098 18096 7104 18148
rect 7156 18136 7162 18148
rect 7285 18139 7343 18145
rect 7285 18136 7297 18139
rect 7156 18108 7297 18136
rect 7156 18096 7162 18108
rect 7285 18105 7297 18108
rect 7331 18105 7343 18139
rect 8938 18136 8944 18148
rect 7285 18099 7343 18105
rect 8312 18108 8944 18136
rect 4341 18071 4399 18077
rect 4341 18068 4353 18071
rect 4304 18040 4353 18068
rect 4304 18028 4310 18040
rect 4341 18037 4353 18040
rect 4387 18037 4399 18071
rect 4341 18031 4399 18037
rect 4801 18071 4859 18077
rect 4801 18037 4813 18071
rect 4847 18068 4859 18071
rect 4982 18068 4988 18080
rect 4847 18040 4988 18068
rect 4847 18037 4859 18040
rect 4801 18031 4859 18037
rect 4982 18028 4988 18040
rect 5040 18068 5046 18080
rect 5353 18071 5411 18077
rect 5353 18068 5365 18071
rect 5040 18040 5365 18068
rect 5040 18028 5046 18040
rect 5353 18037 5365 18040
rect 5399 18037 5411 18071
rect 5353 18031 5411 18037
rect 5442 18028 5448 18080
rect 5500 18068 5506 18080
rect 6549 18071 6607 18077
rect 6549 18068 6561 18071
rect 5500 18040 6561 18068
rect 5500 18028 5506 18040
rect 6549 18037 6561 18040
rect 6595 18068 6607 18071
rect 7190 18068 7196 18080
rect 6595 18040 7196 18068
rect 6595 18037 6607 18040
rect 6549 18031 6607 18037
rect 7190 18028 7196 18040
rect 7248 18028 7254 18080
rect 7926 18028 7932 18080
rect 7984 18068 7990 18080
rect 8312 18077 8340 18108
rect 8938 18096 8944 18108
rect 8996 18096 9002 18148
rect 10686 18096 10692 18148
rect 10744 18136 10750 18148
rect 12176 18145 12204 18176
rect 12805 18173 12817 18176
rect 12851 18173 12863 18207
rect 12912 18204 12940 18244
rect 13078 18232 13084 18244
rect 13136 18272 13142 18284
rect 13449 18275 13507 18281
rect 13449 18272 13461 18275
rect 13136 18244 13461 18272
rect 13136 18232 13142 18244
rect 13449 18241 13461 18244
rect 13495 18241 13507 18275
rect 13449 18235 13507 18241
rect 17497 18275 17555 18281
rect 17497 18241 17509 18275
rect 17543 18272 17555 18275
rect 18138 18272 18144 18284
rect 17543 18244 18144 18272
rect 17543 18241 17555 18244
rect 17497 18235 17555 18241
rect 18138 18232 18144 18244
rect 18196 18272 18202 18284
rect 18509 18275 18567 18281
rect 18509 18272 18521 18275
rect 18196 18244 18521 18272
rect 18196 18232 18202 18244
rect 18509 18241 18521 18244
rect 18555 18241 18567 18275
rect 18509 18235 18567 18241
rect 18598 18232 18604 18284
rect 18656 18272 18662 18284
rect 20088 18281 20116 18312
rect 25866 18300 25872 18312
rect 25924 18340 25930 18352
rect 26513 18343 26571 18349
rect 26513 18340 26525 18343
rect 25924 18312 26525 18340
rect 25924 18300 25930 18312
rect 26513 18309 26525 18312
rect 26559 18340 26571 18343
rect 27985 18343 28043 18349
rect 27985 18340 27997 18343
rect 26559 18312 27997 18340
rect 26559 18309 26571 18312
rect 26513 18303 26571 18309
rect 20073 18275 20131 18281
rect 18656 18244 18701 18272
rect 18656 18232 18662 18244
rect 20073 18241 20085 18275
rect 20119 18241 20131 18275
rect 20073 18235 20131 18241
rect 20162 18232 20168 18284
rect 20220 18272 20226 18284
rect 20220 18244 20265 18272
rect 20220 18232 20226 18244
rect 21634 18232 21640 18284
rect 21692 18272 21698 18284
rect 22094 18272 22100 18284
rect 21692 18244 22100 18272
rect 21692 18232 21698 18244
rect 22094 18232 22100 18244
rect 22152 18232 22158 18284
rect 27540 18281 27568 18312
rect 27985 18309 27997 18312
rect 28031 18309 28043 18343
rect 27985 18303 28043 18309
rect 27525 18275 27583 18281
rect 27525 18241 27537 18275
rect 27571 18241 27583 18275
rect 27525 18235 27583 18241
rect 14185 18207 14243 18213
rect 14185 18204 14197 18207
rect 12912 18176 14197 18204
rect 12805 18167 12863 18173
rect 14185 18173 14197 18176
rect 14231 18204 14243 18207
rect 14231 18176 14596 18204
rect 14231 18173 14243 18176
rect 14185 18167 14243 18173
rect 12161 18139 12219 18145
rect 12161 18136 12173 18139
rect 10744 18108 12173 18136
rect 10744 18096 10750 18108
rect 12161 18105 12173 18108
rect 12207 18105 12219 18139
rect 12161 18099 12219 18105
rect 13906 18096 13912 18148
rect 13964 18136 13970 18148
rect 14430 18139 14488 18145
rect 14430 18136 14442 18139
rect 13964 18108 14442 18136
rect 13964 18096 13970 18108
rect 14430 18105 14442 18108
rect 14476 18105 14488 18139
rect 14430 18099 14488 18105
rect 8297 18071 8355 18077
rect 8297 18068 8309 18071
rect 7984 18040 8309 18068
rect 7984 18028 7990 18040
rect 8297 18037 8309 18040
rect 8343 18037 8355 18071
rect 8478 18068 8484 18080
rect 8439 18040 8484 18068
rect 8297 18031 8355 18037
rect 8478 18028 8484 18040
rect 8536 18028 8542 18080
rect 8570 18028 8576 18080
rect 8628 18068 8634 18080
rect 8849 18071 8907 18077
rect 8849 18068 8861 18071
rect 8628 18040 8861 18068
rect 8628 18028 8634 18040
rect 8849 18037 8861 18040
rect 8895 18037 8907 18071
rect 8849 18031 8907 18037
rect 10778 18028 10784 18080
rect 10836 18068 10842 18080
rect 11241 18071 11299 18077
rect 11241 18068 11253 18071
rect 10836 18040 11253 18068
rect 10836 18028 10842 18040
rect 11241 18037 11253 18040
rect 11287 18037 11299 18071
rect 11241 18031 11299 18037
rect 12897 18071 12955 18077
rect 12897 18037 12909 18071
rect 12943 18068 12955 18071
rect 12986 18068 12992 18080
rect 12943 18040 12992 18068
rect 12943 18037 12955 18040
rect 12897 18031 12955 18037
rect 12986 18028 12992 18040
rect 13044 18028 13050 18080
rect 14093 18071 14151 18077
rect 14093 18037 14105 18071
rect 14139 18068 14151 18071
rect 14568 18068 14596 18176
rect 18230 18164 18236 18216
rect 18288 18204 18294 18216
rect 18417 18207 18475 18213
rect 18417 18204 18429 18207
rect 18288 18176 18429 18204
rect 18288 18164 18294 18176
rect 18417 18173 18429 18176
rect 18463 18173 18475 18207
rect 18417 18167 18475 18173
rect 18874 18164 18880 18216
rect 18932 18204 18938 18216
rect 19981 18207 20039 18213
rect 19981 18204 19993 18207
rect 18932 18176 19993 18204
rect 18932 18164 18938 18176
rect 19981 18173 19993 18176
rect 20027 18204 20039 18207
rect 20254 18204 20260 18216
rect 20027 18176 20260 18204
rect 20027 18173 20039 18176
rect 19981 18167 20039 18173
rect 20254 18164 20260 18176
rect 20312 18164 20318 18216
rect 21453 18207 21511 18213
rect 21453 18173 21465 18207
rect 21499 18204 21511 18207
rect 21913 18207 21971 18213
rect 21913 18204 21925 18207
rect 21499 18176 21925 18204
rect 21499 18173 21511 18176
rect 21453 18167 21511 18173
rect 21913 18173 21925 18176
rect 21959 18204 21971 18207
rect 22002 18204 22008 18216
rect 21959 18176 22008 18204
rect 21959 18173 21971 18176
rect 21913 18167 21971 18173
rect 22002 18164 22008 18176
rect 22060 18164 22066 18216
rect 24489 18207 24547 18213
rect 24489 18204 24501 18207
rect 24320 18176 24501 18204
rect 19058 18136 19064 18148
rect 19019 18108 19064 18136
rect 19058 18096 19064 18108
rect 19116 18096 19122 18148
rect 20346 18096 20352 18148
rect 20404 18136 20410 18148
rect 21266 18136 21272 18148
rect 20404 18108 21272 18136
rect 20404 18096 20410 18108
rect 21266 18096 21272 18108
rect 21324 18096 21330 18148
rect 22094 18096 22100 18148
rect 22152 18136 22158 18148
rect 22462 18136 22468 18148
rect 22152 18108 22468 18136
rect 22152 18096 22158 18108
rect 22462 18096 22468 18108
rect 22520 18136 22526 18148
rect 22925 18139 22983 18145
rect 22925 18136 22937 18139
rect 22520 18108 22937 18136
rect 22520 18096 22526 18108
rect 22925 18105 22937 18108
rect 22971 18105 22983 18139
rect 22925 18099 22983 18105
rect 24320 18080 24348 18176
rect 24489 18173 24501 18176
rect 24535 18173 24547 18207
rect 24489 18167 24547 18173
rect 24670 18096 24676 18148
rect 24728 18145 24734 18148
rect 24728 18139 24792 18145
rect 24728 18105 24746 18139
rect 24780 18105 24792 18139
rect 24728 18099 24792 18105
rect 24728 18096 24734 18099
rect 15286 18068 15292 18080
rect 14139 18040 15292 18068
rect 14139 18037 14151 18040
rect 14093 18031 14151 18037
rect 15286 18028 15292 18040
rect 15344 18028 15350 18080
rect 15562 18068 15568 18080
rect 15523 18040 15568 18068
rect 15562 18028 15568 18040
rect 15620 18028 15626 18080
rect 15838 18028 15844 18080
rect 15896 18068 15902 18080
rect 16482 18068 16488 18080
rect 15896 18040 16488 18068
rect 15896 18028 15902 18040
rect 16482 18028 16488 18040
rect 16540 18028 16546 18080
rect 19426 18068 19432 18080
rect 19387 18040 19432 18068
rect 19426 18028 19432 18040
rect 19484 18028 19490 18080
rect 20714 18028 20720 18080
rect 20772 18068 20778 18080
rect 20901 18071 20959 18077
rect 20901 18068 20913 18071
rect 20772 18040 20913 18068
rect 20772 18028 20778 18040
rect 20901 18037 20913 18040
rect 20947 18037 20959 18071
rect 21542 18068 21548 18080
rect 21503 18040 21548 18068
rect 20901 18031 20959 18037
rect 21542 18028 21548 18040
rect 21600 18028 21606 18080
rect 21910 18028 21916 18080
rect 21968 18068 21974 18080
rect 22005 18071 22063 18077
rect 22005 18068 22017 18071
rect 21968 18040 22017 18068
rect 21968 18028 21974 18040
rect 22005 18037 22017 18040
rect 22051 18037 22063 18071
rect 22646 18068 22652 18080
rect 22607 18040 22652 18068
rect 22005 18031 22063 18037
rect 22646 18028 22652 18040
rect 22704 18028 22710 18080
rect 24302 18068 24308 18080
rect 24263 18040 24308 18068
rect 24302 18028 24308 18040
rect 24360 18028 24366 18080
rect 26234 18028 26240 18080
rect 26292 18068 26298 18080
rect 27338 18068 27344 18080
rect 26292 18040 27344 18068
rect 26292 18028 26298 18040
rect 27338 18028 27344 18040
rect 27396 18028 27402 18080
rect 27433 18071 27491 18077
rect 27433 18037 27445 18071
rect 27479 18068 27491 18071
rect 27522 18068 27528 18080
rect 27479 18040 27528 18068
rect 27479 18037 27491 18040
rect 27433 18031 27491 18037
rect 27522 18028 27528 18040
rect 27580 18028 27586 18080
rect 1104 17978 28888 18000
rect 1104 17926 10982 17978
rect 11034 17926 11046 17978
rect 11098 17926 11110 17978
rect 11162 17926 11174 17978
rect 11226 17926 20982 17978
rect 21034 17926 21046 17978
rect 21098 17926 21110 17978
rect 21162 17926 21174 17978
rect 21226 17926 28888 17978
rect 1104 17904 28888 17926
rect 1765 17867 1823 17873
rect 1765 17833 1777 17867
rect 1811 17864 1823 17867
rect 2222 17864 2228 17876
rect 1811 17836 2228 17864
rect 1811 17833 1823 17836
rect 1765 17827 1823 17833
rect 2222 17824 2228 17836
rect 2280 17824 2286 17876
rect 3421 17867 3479 17873
rect 3421 17833 3433 17867
rect 3467 17864 3479 17867
rect 3694 17864 3700 17876
rect 3467 17836 3700 17864
rect 3467 17833 3479 17836
rect 3421 17827 3479 17833
rect 3694 17824 3700 17836
rect 3752 17824 3758 17876
rect 4338 17864 4344 17876
rect 4299 17836 4344 17864
rect 4338 17824 4344 17836
rect 4396 17824 4402 17876
rect 4706 17864 4712 17876
rect 4667 17836 4712 17864
rect 4706 17824 4712 17836
rect 4764 17824 4770 17876
rect 5534 17824 5540 17876
rect 5592 17864 5598 17876
rect 6365 17867 6423 17873
rect 6365 17864 6377 17867
rect 5592 17836 6377 17864
rect 5592 17824 5598 17836
rect 6365 17833 6377 17836
rect 6411 17864 6423 17867
rect 6822 17864 6828 17876
rect 6411 17836 6828 17864
rect 6411 17833 6423 17836
rect 6365 17827 6423 17833
rect 6822 17824 6828 17836
rect 6880 17824 6886 17876
rect 7558 17824 7564 17876
rect 7616 17864 7622 17876
rect 7653 17867 7711 17873
rect 7653 17864 7665 17867
rect 7616 17836 7665 17864
rect 7616 17824 7622 17836
rect 7653 17833 7665 17836
rect 7699 17833 7711 17867
rect 7653 17827 7711 17833
rect 8021 17867 8079 17873
rect 8021 17833 8033 17867
rect 8067 17864 8079 17867
rect 8202 17864 8208 17876
rect 8067 17836 8208 17864
rect 8067 17833 8079 17836
rect 8021 17827 8079 17833
rect 8202 17824 8208 17836
rect 8260 17824 8266 17876
rect 8478 17824 8484 17876
rect 8536 17864 8542 17876
rect 9398 17864 9404 17876
rect 8536 17836 9404 17864
rect 8536 17824 8542 17836
rect 9398 17824 9404 17836
rect 9456 17824 9462 17876
rect 11422 17824 11428 17876
rect 11480 17864 11486 17876
rect 11609 17867 11667 17873
rect 11609 17864 11621 17867
rect 11480 17836 11621 17864
rect 11480 17824 11486 17836
rect 11609 17833 11621 17836
rect 11655 17833 11667 17867
rect 12158 17864 12164 17876
rect 12119 17836 12164 17864
rect 11609 17827 11667 17833
rect 4154 17756 4160 17808
rect 4212 17796 4218 17808
rect 5230 17799 5288 17805
rect 5230 17796 5242 17799
rect 4212 17768 5242 17796
rect 4212 17756 4218 17768
rect 5230 17765 5242 17768
rect 5276 17796 5288 17799
rect 5350 17796 5356 17808
rect 5276 17768 5356 17796
rect 5276 17765 5288 17768
rect 5230 17759 5288 17765
rect 5350 17756 5356 17768
rect 5408 17796 5414 17808
rect 6917 17799 6975 17805
rect 6917 17796 6929 17799
rect 5408 17768 6929 17796
rect 5408 17756 5414 17768
rect 6917 17765 6929 17768
rect 6963 17796 6975 17799
rect 7282 17796 7288 17808
rect 6963 17768 7288 17796
rect 6963 17765 6975 17768
rect 6917 17759 6975 17765
rect 7282 17756 7288 17768
rect 7340 17756 7346 17808
rect 8386 17796 8392 17808
rect 8299 17768 8392 17796
rect 8386 17756 8392 17768
rect 8444 17796 8450 17808
rect 10778 17796 10784 17808
rect 8444 17768 10784 17796
rect 8444 17756 8450 17768
rect 10778 17756 10784 17768
rect 10836 17756 10842 17808
rect 11624 17796 11652 17827
rect 12158 17824 12164 17836
rect 12216 17824 12222 17876
rect 13633 17867 13691 17873
rect 13633 17833 13645 17867
rect 13679 17864 13691 17867
rect 13722 17864 13728 17876
rect 13679 17836 13728 17864
rect 13679 17833 13691 17836
rect 13633 17827 13691 17833
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 17221 17867 17279 17873
rect 17221 17833 17233 17867
rect 17267 17833 17279 17867
rect 17221 17827 17279 17833
rect 19705 17867 19763 17873
rect 19705 17833 19717 17867
rect 19751 17864 19763 17867
rect 20070 17864 20076 17876
rect 19751 17836 20076 17864
rect 19751 17833 19763 17836
rect 19705 17827 19763 17833
rect 13078 17796 13084 17808
rect 11624 17768 13084 17796
rect 13078 17756 13084 17768
rect 13136 17756 13142 17808
rect 13814 17756 13820 17808
rect 13872 17796 13878 17808
rect 14093 17799 14151 17805
rect 14093 17796 14105 17799
rect 13872 17768 14105 17796
rect 13872 17756 13878 17768
rect 14093 17765 14105 17768
rect 14139 17765 14151 17799
rect 17236 17796 17264 17827
rect 20070 17824 20076 17836
rect 20128 17824 20134 17876
rect 20254 17864 20260 17876
rect 20215 17836 20260 17864
rect 20254 17824 20260 17836
rect 20312 17824 20318 17876
rect 20901 17867 20959 17873
rect 20901 17833 20913 17867
rect 20947 17864 20959 17867
rect 22094 17864 22100 17876
rect 20947 17836 22100 17864
rect 20947 17833 20959 17836
rect 20901 17827 20959 17833
rect 22094 17824 22100 17836
rect 22152 17824 22158 17876
rect 24949 17867 25007 17873
rect 24949 17833 24961 17867
rect 24995 17864 25007 17867
rect 25406 17864 25412 17876
rect 24995 17836 25412 17864
rect 24995 17833 25007 17836
rect 24949 17827 25007 17833
rect 25406 17824 25412 17836
rect 25464 17864 25470 17876
rect 26145 17867 26203 17873
rect 26145 17864 26157 17867
rect 25464 17836 26157 17864
rect 25464 17824 25470 17836
rect 26145 17833 26157 17836
rect 26191 17864 26203 17867
rect 26326 17864 26332 17876
rect 26191 17836 26332 17864
rect 26191 17833 26203 17836
rect 26145 17827 26203 17833
rect 26326 17824 26332 17836
rect 26384 17824 26390 17876
rect 26510 17864 26516 17876
rect 26471 17836 26516 17864
rect 26510 17824 26516 17836
rect 26568 17824 26574 17876
rect 18233 17799 18291 17805
rect 18233 17796 18245 17799
rect 17236 17768 18245 17796
rect 14093 17759 14151 17765
rect 18233 17765 18245 17768
rect 18279 17796 18291 17799
rect 18592 17799 18650 17805
rect 18592 17796 18604 17799
rect 18279 17768 18604 17796
rect 18279 17765 18291 17768
rect 18233 17759 18291 17765
rect 18592 17765 18604 17768
rect 18638 17796 18650 17799
rect 19794 17796 19800 17808
rect 18638 17768 19800 17796
rect 18638 17765 18650 17768
rect 18592 17759 18650 17765
rect 19794 17756 19800 17768
rect 19852 17796 19858 17808
rect 20717 17799 20775 17805
rect 20717 17796 20729 17799
rect 19852 17768 20729 17796
rect 19852 17756 19858 17768
rect 20717 17765 20729 17768
rect 20763 17796 20775 17799
rect 21450 17796 21456 17808
rect 20763 17768 21456 17796
rect 20763 17765 20775 17768
rect 20717 17759 20775 17765
rect 21450 17756 21456 17768
rect 21508 17756 21514 17808
rect 22462 17756 22468 17808
rect 22520 17796 22526 17808
rect 22710 17799 22768 17805
rect 22710 17796 22722 17799
rect 22520 17768 22722 17796
rect 22520 17756 22526 17768
rect 22710 17765 22722 17768
rect 22756 17765 22768 17799
rect 22710 17759 22768 17765
rect 25590 17756 25596 17808
rect 25648 17796 25654 17808
rect 26973 17799 27031 17805
rect 26973 17796 26985 17799
rect 25648 17768 26985 17796
rect 25648 17756 25654 17768
rect 26973 17765 26985 17768
rect 27019 17765 27031 17799
rect 26973 17759 27031 17765
rect 2130 17728 2136 17740
rect 2091 17700 2136 17728
rect 2130 17688 2136 17700
rect 2188 17728 2194 17740
rect 2682 17728 2688 17740
rect 2188 17700 2688 17728
rect 2188 17688 2194 17700
rect 2682 17688 2688 17700
rect 2740 17688 2746 17740
rect 4706 17688 4712 17740
rect 4764 17728 4770 17740
rect 4985 17731 5043 17737
rect 4985 17728 4997 17731
rect 4764 17700 4997 17728
rect 4764 17688 4770 17700
rect 4985 17697 4997 17700
rect 5031 17697 5043 17731
rect 4985 17691 5043 17697
rect 7377 17731 7435 17737
rect 7377 17697 7389 17731
rect 7423 17728 7435 17731
rect 7650 17728 7656 17740
rect 7423 17700 7656 17728
rect 7423 17697 7435 17700
rect 7377 17691 7435 17697
rect 7650 17688 7656 17700
rect 7708 17688 7714 17740
rect 8202 17688 8208 17740
rect 8260 17728 8266 17740
rect 9582 17728 9588 17740
rect 8260 17700 9588 17728
rect 8260 17688 8266 17700
rect 9582 17688 9588 17700
rect 9640 17728 9646 17740
rect 9677 17731 9735 17737
rect 9677 17728 9689 17731
rect 9640 17700 9689 17728
rect 9640 17688 9646 17700
rect 9677 17697 9689 17700
rect 9723 17697 9735 17731
rect 9677 17691 9735 17697
rect 9766 17688 9772 17740
rect 9824 17728 9830 17740
rect 9933 17731 9991 17737
rect 9933 17728 9945 17731
rect 9824 17700 9945 17728
rect 9824 17688 9830 17700
rect 9933 17697 9945 17700
rect 9979 17697 9991 17731
rect 13998 17728 14004 17740
rect 13959 17700 14004 17728
rect 9933 17691 9991 17697
rect 13998 17688 14004 17700
rect 14056 17688 14062 17740
rect 16097 17731 16155 17737
rect 16097 17728 16109 17731
rect 14200 17700 16109 17728
rect 14200 17672 14228 17700
rect 16097 17697 16109 17700
rect 16143 17728 16155 17731
rect 16390 17728 16396 17740
rect 16143 17700 16396 17728
rect 16143 17697 16155 17700
rect 16097 17691 16155 17697
rect 16390 17688 16396 17700
rect 16448 17688 16454 17740
rect 21266 17728 21272 17740
rect 21227 17700 21272 17728
rect 21266 17688 21272 17700
rect 21324 17688 21330 17740
rect 25409 17731 25467 17737
rect 25409 17697 25421 17731
rect 25455 17728 25467 17731
rect 25682 17728 25688 17740
rect 25455 17700 25688 17728
rect 25455 17697 25467 17700
rect 25409 17691 25467 17697
rect 25682 17688 25688 17700
rect 25740 17728 25746 17740
rect 26881 17731 26939 17737
rect 26881 17728 26893 17731
rect 25740 17700 26893 17728
rect 25740 17688 25746 17700
rect 26881 17697 26893 17700
rect 26927 17697 26939 17731
rect 26881 17691 26939 17697
rect 1854 17620 1860 17672
rect 1912 17660 1918 17672
rect 2225 17663 2283 17669
rect 2225 17660 2237 17663
rect 1912 17632 2237 17660
rect 1912 17620 1918 17632
rect 2225 17629 2237 17632
rect 2271 17629 2283 17663
rect 2225 17623 2283 17629
rect 2317 17663 2375 17669
rect 2317 17629 2329 17663
rect 2363 17660 2375 17663
rect 3142 17660 3148 17672
rect 2363 17632 3148 17660
rect 2363 17629 2375 17632
rect 2317 17623 2375 17629
rect 1673 17595 1731 17601
rect 1673 17561 1685 17595
rect 1719 17592 1731 17595
rect 2332 17592 2360 17623
rect 3142 17620 3148 17632
rect 3200 17620 3206 17672
rect 7466 17620 7472 17672
rect 7524 17660 7530 17672
rect 8481 17663 8539 17669
rect 8481 17660 8493 17663
rect 7524 17632 8493 17660
rect 7524 17620 7530 17632
rect 8481 17629 8493 17632
rect 8527 17629 8539 17663
rect 8662 17660 8668 17672
rect 8623 17632 8668 17660
rect 8481 17623 8539 17629
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 11514 17620 11520 17672
rect 11572 17660 11578 17672
rect 12710 17660 12716 17672
rect 11572 17632 12716 17660
rect 11572 17620 11578 17632
rect 12710 17620 12716 17632
rect 12768 17620 12774 17672
rect 14182 17660 14188 17672
rect 14143 17632 14188 17660
rect 14182 17620 14188 17632
rect 14240 17620 14246 17672
rect 15286 17620 15292 17672
rect 15344 17660 15350 17672
rect 15838 17660 15844 17672
rect 15344 17632 15844 17660
rect 15344 17620 15350 17632
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 17862 17620 17868 17672
rect 17920 17660 17926 17672
rect 18325 17663 18383 17669
rect 18325 17660 18337 17663
rect 17920 17632 18337 17660
rect 17920 17620 17926 17632
rect 18325 17629 18337 17632
rect 18371 17629 18383 17663
rect 21358 17660 21364 17672
rect 21319 17632 21364 17660
rect 18325 17623 18383 17629
rect 21358 17620 21364 17632
rect 21416 17620 21422 17672
rect 21450 17620 21456 17672
rect 21508 17660 21514 17672
rect 21508 17632 21553 17660
rect 21508 17620 21514 17632
rect 22370 17620 22376 17672
rect 22428 17660 22434 17672
rect 22465 17663 22523 17669
rect 22465 17660 22477 17663
rect 22428 17632 22477 17660
rect 22428 17620 22434 17632
rect 22465 17629 22477 17632
rect 22511 17629 22523 17663
rect 22465 17623 22523 17629
rect 24854 17620 24860 17672
rect 24912 17660 24918 17672
rect 26142 17660 26148 17672
rect 24912 17632 26148 17660
rect 24912 17620 24918 17632
rect 26142 17620 26148 17632
rect 26200 17620 26206 17672
rect 27157 17663 27215 17669
rect 27157 17629 27169 17663
rect 27203 17660 27215 17663
rect 27430 17660 27436 17672
rect 27203 17632 27436 17660
rect 27203 17629 27215 17632
rect 27157 17623 27215 17629
rect 27430 17620 27436 17632
rect 27488 17620 27494 17672
rect 1719 17564 2360 17592
rect 1719 17561 1731 17564
rect 1673 17555 1731 17561
rect 11238 17552 11244 17604
rect 11296 17592 11302 17604
rect 11977 17595 12035 17601
rect 11977 17592 11989 17595
rect 11296 17564 11989 17592
rect 11296 17552 11302 17564
rect 11977 17561 11989 17564
rect 12023 17561 12035 17595
rect 11977 17555 12035 17561
rect 19334 17552 19340 17604
rect 19392 17592 19398 17604
rect 22094 17592 22100 17604
rect 19392 17564 22100 17592
rect 19392 17552 19398 17564
rect 22094 17552 22100 17564
rect 22152 17552 22158 17604
rect 2774 17484 2780 17536
rect 2832 17524 2838 17536
rect 11057 17527 11115 17533
rect 2832 17496 2877 17524
rect 2832 17484 2838 17496
rect 11057 17493 11069 17527
rect 11103 17524 11115 17527
rect 11514 17524 11520 17536
rect 11103 17496 11520 17524
rect 11103 17493 11115 17496
rect 11057 17487 11115 17493
rect 11514 17484 11520 17496
rect 11572 17484 11578 17536
rect 12986 17524 12992 17536
rect 12947 17496 12992 17524
rect 12986 17484 12992 17496
rect 13044 17484 13050 17536
rect 21910 17524 21916 17536
rect 21871 17496 21916 17524
rect 21910 17484 21916 17496
rect 21968 17484 21974 17536
rect 23845 17527 23903 17533
rect 23845 17493 23857 17527
rect 23891 17524 23903 17527
rect 24118 17524 24124 17536
rect 23891 17496 24124 17524
rect 23891 17493 23903 17496
rect 23845 17487 23903 17493
rect 24118 17484 24124 17496
rect 24176 17484 24182 17536
rect 24581 17527 24639 17533
rect 24581 17493 24593 17527
rect 24627 17524 24639 17527
rect 24670 17524 24676 17536
rect 24627 17496 24676 17524
rect 24627 17493 24639 17496
rect 24581 17487 24639 17493
rect 24670 17484 24676 17496
rect 24728 17484 24734 17536
rect 25314 17524 25320 17536
rect 25275 17496 25320 17524
rect 25314 17484 25320 17496
rect 25372 17484 25378 17536
rect 27614 17524 27620 17536
rect 27575 17496 27620 17524
rect 27614 17484 27620 17496
rect 27672 17484 27678 17536
rect 1104 17434 28888 17456
rect 1104 17382 5982 17434
rect 6034 17382 6046 17434
rect 6098 17382 6110 17434
rect 6162 17382 6174 17434
rect 6226 17382 15982 17434
rect 16034 17382 16046 17434
rect 16098 17382 16110 17434
rect 16162 17382 16174 17434
rect 16226 17382 25982 17434
rect 26034 17382 26046 17434
rect 26098 17382 26110 17434
rect 26162 17382 26174 17434
rect 26226 17382 28888 17434
rect 1104 17360 28888 17382
rect 3142 17320 3148 17332
rect 3103 17292 3148 17320
rect 3142 17280 3148 17292
rect 3200 17280 3206 17332
rect 5350 17280 5356 17332
rect 5408 17320 5414 17332
rect 5629 17323 5687 17329
rect 5629 17320 5641 17323
rect 5408 17292 5641 17320
rect 5408 17280 5414 17292
rect 5629 17289 5641 17292
rect 5675 17320 5687 17323
rect 6181 17323 6239 17329
rect 6181 17320 6193 17323
rect 5675 17292 6193 17320
rect 5675 17289 5687 17292
rect 5629 17283 5687 17289
rect 6181 17289 6193 17292
rect 6227 17289 6239 17323
rect 6638 17320 6644 17332
rect 6599 17292 6644 17320
rect 6181 17283 6239 17289
rect 6638 17280 6644 17292
rect 6696 17280 6702 17332
rect 7837 17323 7895 17329
rect 7837 17289 7849 17323
rect 7883 17320 7895 17323
rect 8662 17320 8668 17332
rect 7883 17292 8668 17320
rect 7883 17289 7895 17292
rect 7837 17283 7895 17289
rect 8662 17280 8668 17292
rect 8720 17320 8726 17332
rect 9677 17323 9735 17329
rect 9677 17320 9689 17323
rect 8720 17292 9689 17320
rect 8720 17280 8726 17292
rect 9677 17289 9689 17292
rect 9723 17320 9735 17323
rect 9766 17320 9772 17332
rect 9723 17292 9772 17320
rect 9723 17289 9735 17292
rect 9677 17283 9735 17289
rect 9766 17280 9772 17292
rect 9824 17320 9830 17332
rect 10597 17323 10655 17329
rect 10597 17320 10609 17323
rect 9824 17292 10609 17320
rect 9824 17280 9830 17292
rect 10597 17289 10609 17292
rect 10643 17289 10655 17323
rect 10778 17320 10784 17332
rect 10739 17292 10784 17320
rect 10597 17283 10655 17289
rect 10778 17280 10784 17292
rect 10836 17280 10842 17332
rect 11790 17320 11796 17332
rect 11751 17292 11796 17320
rect 11790 17280 11796 17292
rect 11848 17280 11854 17332
rect 12437 17323 12495 17329
rect 12437 17289 12449 17323
rect 12483 17320 12495 17323
rect 12986 17320 12992 17332
rect 12483 17292 12992 17320
rect 12483 17289 12495 17292
rect 12437 17283 12495 17289
rect 12986 17280 12992 17292
rect 13044 17280 13050 17332
rect 13725 17323 13783 17329
rect 13725 17289 13737 17323
rect 13771 17320 13783 17323
rect 14182 17320 14188 17332
rect 13771 17292 14188 17320
rect 13771 17289 13783 17292
rect 13725 17283 13783 17289
rect 14182 17280 14188 17292
rect 14240 17280 14246 17332
rect 16390 17320 16396 17332
rect 16351 17292 16396 17320
rect 16390 17280 16396 17292
rect 16448 17320 16454 17332
rect 16945 17323 17003 17329
rect 16945 17320 16957 17323
rect 16448 17292 16957 17320
rect 16448 17280 16454 17292
rect 16945 17289 16957 17292
rect 16991 17289 17003 17323
rect 18322 17320 18328 17332
rect 18283 17292 18328 17320
rect 16945 17283 17003 17289
rect 18322 17280 18328 17292
rect 18380 17280 18386 17332
rect 19794 17320 19800 17332
rect 19755 17292 19800 17320
rect 19794 17280 19800 17292
rect 19852 17280 19858 17332
rect 20625 17323 20683 17329
rect 20625 17289 20637 17323
rect 20671 17320 20683 17323
rect 21450 17320 21456 17332
rect 20671 17292 21456 17320
rect 20671 17289 20683 17292
rect 20625 17283 20683 17289
rect 21450 17280 21456 17292
rect 21508 17320 21514 17332
rect 22462 17320 22468 17332
rect 21508 17292 22468 17320
rect 21508 17280 21514 17292
rect 22462 17280 22468 17292
rect 22520 17280 22526 17332
rect 25682 17320 25688 17332
rect 25643 17292 25688 17320
rect 25682 17280 25688 17292
rect 25740 17280 25746 17332
rect 27430 17320 27436 17332
rect 25792 17292 27436 17320
rect 9582 17212 9588 17264
rect 9640 17252 9646 17264
rect 10229 17255 10287 17261
rect 10229 17252 10241 17255
rect 9640 17224 10241 17252
rect 9640 17212 9646 17224
rect 10229 17221 10241 17224
rect 10275 17221 10287 17255
rect 10229 17215 10287 17221
rect 13740 17224 15056 17252
rect 11330 17184 11336 17196
rect 11291 17156 11336 17184
rect 11330 17144 11336 17156
rect 11388 17144 11394 17196
rect 12710 17144 12716 17196
rect 12768 17184 12774 17196
rect 12989 17187 13047 17193
rect 12989 17184 13001 17187
rect 12768 17156 13001 17184
rect 12768 17144 12774 17156
rect 12989 17153 13001 17156
rect 13035 17153 13047 17187
rect 12989 17147 13047 17153
rect 1486 17076 1492 17128
rect 1544 17116 1550 17128
rect 1673 17119 1731 17125
rect 1673 17116 1685 17119
rect 1544 17088 1685 17116
rect 1544 17076 1550 17088
rect 1673 17085 1685 17088
rect 1719 17116 1731 17119
rect 1765 17119 1823 17125
rect 1765 17116 1777 17119
rect 1719 17088 1777 17116
rect 1719 17085 1731 17088
rect 1673 17079 1731 17085
rect 1765 17085 1777 17088
rect 1811 17085 1823 17119
rect 1765 17079 1823 17085
rect 2032 17119 2090 17125
rect 2032 17085 2044 17119
rect 2078 17116 2090 17119
rect 2406 17116 2412 17128
rect 2078 17088 2412 17116
rect 2078 17085 2090 17088
rect 2032 17079 2090 17085
rect 2406 17076 2412 17088
rect 2464 17116 2470 17128
rect 2774 17116 2780 17128
rect 2464 17088 2780 17116
rect 2464 17076 2470 17088
rect 2774 17076 2780 17088
rect 2832 17076 2838 17128
rect 4249 17119 4307 17125
rect 4249 17085 4261 17119
rect 4295 17085 4307 17119
rect 4249 17079 4307 17085
rect 4157 17051 4215 17057
rect 4157 17017 4169 17051
rect 4203 17048 4215 17051
rect 4264 17048 4292 17079
rect 4338 17076 4344 17128
rect 4396 17116 4402 17128
rect 4505 17119 4563 17125
rect 4505 17116 4517 17119
rect 4396 17088 4517 17116
rect 4396 17076 4402 17088
rect 4505 17085 4517 17088
rect 4551 17085 4563 17119
rect 4505 17079 4563 17085
rect 8202 17076 8208 17128
rect 8260 17116 8266 17128
rect 8297 17119 8355 17125
rect 8297 17116 8309 17119
rect 8260 17088 8309 17116
rect 8260 17076 8266 17088
rect 8297 17085 8309 17088
rect 8343 17085 8355 17119
rect 11146 17116 11152 17128
rect 11107 17088 11152 17116
rect 8297 17079 8355 17085
rect 11146 17076 11152 17088
rect 11204 17076 11210 17128
rect 11790 17076 11796 17128
rect 11848 17116 11854 17128
rect 12805 17119 12863 17125
rect 12805 17116 12817 17119
rect 11848 17088 12817 17116
rect 11848 17076 11854 17088
rect 12805 17085 12817 17088
rect 12851 17116 12863 17119
rect 12851 17088 13032 17116
rect 12851 17085 12863 17088
rect 12805 17079 12863 17085
rect 13004 17060 13032 17088
rect 4706 17048 4712 17060
rect 4203 17020 4712 17048
rect 4203 17017 4215 17020
rect 4157 17011 4215 17017
rect 4706 17008 4712 17020
rect 4764 17008 4770 17060
rect 7101 17051 7159 17057
rect 7101 17017 7113 17051
rect 7147 17048 7159 17051
rect 7466 17048 7472 17060
rect 7147 17020 7472 17048
rect 7147 17017 7159 17020
rect 7101 17011 7159 17017
rect 7466 17008 7472 17020
rect 7524 17008 7530 17060
rect 8564 17051 8622 17057
rect 8564 17048 8576 17051
rect 8036 17020 8576 17048
rect 1854 16940 1860 16992
rect 1912 16980 1918 16992
rect 2774 16980 2780 16992
rect 1912 16952 2780 16980
rect 1912 16940 1918 16952
rect 2774 16940 2780 16952
rect 2832 16940 2838 16992
rect 3694 16980 3700 16992
rect 3655 16952 3700 16980
rect 3694 16940 3700 16952
rect 3752 16940 3758 16992
rect 7377 16983 7435 16989
rect 7377 16949 7389 16983
rect 7423 16980 7435 16983
rect 8036 16980 8064 17020
rect 8564 17017 8576 17020
rect 8610 17048 8622 17051
rect 9490 17048 9496 17060
rect 8610 17020 9496 17048
rect 8610 17017 8622 17020
rect 8564 17011 8622 17017
rect 9490 17008 9496 17020
rect 9548 17008 9554 17060
rect 11238 17048 11244 17060
rect 11199 17020 11244 17048
rect 11238 17008 11244 17020
rect 11296 17008 11302 17060
rect 12986 17008 12992 17060
rect 13044 17008 13050 17060
rect 8202 16980 8208 16992
rect 7423 16952 8064 16980
rect 8163 16952 8208 16980
rect 7423 16949 7435 16952
rect 7377 16943 7435 16949
rect 8202 16940 8208 16952
rect 8260 16940 8266 16992
rect 12250 16980 12256 16992
rect 12211 16952 12256 16980
rect 12250 16940 12256 16952
rect 12308 16980 12314 16992
rect 12897 16983 12955 16989
rect 12897 16980 12909 16983
rect 12308 16952 12909 16980
rect 12308 16940 12314 16952
rect 12897 16949 12909 16952
rect 12943 16980 12955 16983
rect 13740 16980 13768 17224
rect 14001 17187 14059 17193
rect 14001 17153 14013 17187
rect 14047 17184 14059 17187
rect 14918 17184 14924 17196
rect 14047 17156 14924 17184
rect 14047 17153 14059 17156
rect 14001 17147 14059 17153
rect 14918 17144 14924 17156
rect 14976 17144 14982 17196
rect 15028 17184 15056 17224
rect 18969 17187 19027 17193
rect 15028 17156 15148 17184
rect 15013 17119 15071 17125
rect 15013 17085 15025 17119
rect 15059 17085 15071 17119
rect 15120 17116 15148 17156
rect 18969 17153 18981 17187
rect 19015 17184 19027 17187
rect 19058 17184 19064 17196
rect 19015 17156 19064 17184
rect 19015 17153 19027 17156
rect 18969 17147 19027 17153
rect 19058 17144 19064 17156
rect 19116 17184 19122 17196
rect 19812 17184 19840 17280
rect 24670 17212 24676 17264
rect 24728 17252 24734 17264
rect 25041 17255 25099 17261
rect 25041 17252 25053 17255
rect 24728 17224 25053 17252
rect 24728 17212 24734 17224
rect 25041 17221 25053 17224
rect 25087 17252 25099 17255
rect 25792 17252 25820 17292
rect 27430 17280 27436 17292
rect 27488 17320 27494 17332
rect 28077 17323 28135 17329
rect 28077 17320 28089 17323
rect 27488 17292 28089 17320
rect 27488 17280 27494 17292
rect 28077 17289 28089 17292
rect 28123 17289 28135 17323
rect 28077 17283 28135 17289
rect 25087 17224 25820 17252
rect 25087 17221 25099 17224
rect 25041 17215 25099 17221
rect 19116 17156 19840 17184
rect 19116 17144 19122 17156
rect 25590 17144 25596 17196
rect 25648 17184 25654 17196
rect 25961 17187 26019 17193
rect 25961 17184 25973 17187
rect 25648 17156 25973 17184
rect 25648 17144 25654 17156
rect 25961 17153 25973 17156
rect 26007 17153 26019 17187
rect 25961 17147 26019 17153
rect 17773 17119 17831 17125
rect 17773 17116 17785 17119
rect 15120 17088 17785 17116
rect 15013 17079 15071 17085
rect 17773 17085 17785 17088
rect 17819 17116 17831 17119
rect 18598 17116 18604 17128
rect 17819 17088 18604 17116
rect 17819 17085 17831 17088
rect 17773 17079 17831 17085
rect 12943 16952 13768 16980
rect 12943 16949 12955 16952
rect 12897 16943 12955 16949
rect 13814 16940 13820 16992
rect 13872 16980 13878 16992
rect 14461 16983 14519 16989
rect 14461 16980 14473 16983
rect 13872 16952 14473 16980
rect 13872 16940 13878 16952
rect 14461 16949 14473 16952
rect 14507 16949 14519 16983
rect 14461 16943 14519 16949
rect 14921 16983 14979 16989
rect 14921 16949 14933 16983
rect 14967 16980 14979 16983
rect 15028 16980 15056 17079
rect 18598 17076 18604 17088
rect 18656 17116 18662 17128
rect 18785 17119 18843 17125
rect 18785 17116 18797 17119
rect 18656 17088 18797 17116
rect 18656 17076 18662 17088
rect 18785 17085 18797 17088
rect 18831 17085 18843 17119
rect 18785 17079 18843 17085
rect 20806 17076 20812 17128
rect 20864 17116 20870 17128
rect 21085 17119 21143 17125
rect 21085 17116 21097 17119
rect 20864 17088 21097 17116
rect 20864 17076 20870 17088
rect 21085 17085 21097 17088
rect 21131 17116 21143 17119
rect 22370 17116 22376 17128
rect 21131 17088 22376 17116
rect 21131 17085 21143 17088
rect 21085 17079 21143 17085
rect 22370 17076 22376 17088
rect 22428 17116 22434 17128
rect 23017 17119 23075 17125
rect 23017 17116 23029 17119
rect 22428 17088 23029 17116
rect 22428 17076 22434 17088
rect 23017 17085 23029 17088
rect 23063 17116 23075 17119
rect 23385 17119 23443 17125
rect 23385 17116 23397 17119
rect 23063 17088 23397 17116
rect 23063 17085 23075 17088
rect 23017 17079 23075 17085
rect 23385 17085 23397 17088
rect 23431 17116 23443 17119
rect 23661 17119 23719 17125
rect 23661 17116 23673 17119
rect 23431 17088 23673 17116
rect 23431 17085 23443 17088
rect 23385 17079 23443 17085
rect 23661 17085 23673 17088
rect 23707 17116 23719 17119
rect 24302 17116 24308 17128
rect 23707 17088 24308 17116
rect 23707 17085 23719 17088
rect 23661 17079 23719 17085
rect 24302 17076 24308 17088
rect 24360 17076 24366 17128
rect 26145 17119 26203 17125
rect 26145 17085 26157 17119
rect 26191 17116 26203 17119
rect 26234 17116 26240 17128
rect 26191 17088 26240 17116
rect 26191 17085 26203 17088
rect 26145 17079 26203 17085
rect 26234 17076 26240 17088
rect 26292 17076 26298 17128
rect 15280 17051 15338 17057
rect 15280 17017 15292 17051
rect 15326 17048 15338 17051
rect 15470 17048 15476 17060
rect 15326 17020 15476 17048
rect 15326 17017 15338 17020
rect 15280 17011 15338 17017
rect 15470 17008 15476 17020
rect 15528 17008 15534 17060
rect 20257 17051 20315 17057
rect 20257 17017 20269 17051
rect 20303 17048 20315 17051
rect 21352 17051 21410 17057
rect 21352 17048 21364 17051
rect 20303 17020 21364 17048
rect 20303 17017 20315 17020
rect 20257 17011 20315 17017
rect 21352 17017 21364 17020
rect 21398 17048 21410 17051
rect 21910 17048 21916 17060
rect 21398 17020 21916 17048
rect 21398 17017 21410 17020
rect 21352 17011 21410 17017
rect 21910 17008 21916 17020
rect 21968 17008 21974 17060
rect 23928 17051 23986 17057
rect 23928 17017 23940 17051
rect 23974 17048 23986 17051
rect 24118 17048 24124 17060
rect 23974 17020 24124 17048
rect 23974 17017 23986 17020
rect 23928 17011 23986 17017
rect 24118 17008 24124 17020
rect 24176 17008 24182 17060
rect 26326 17008 26332 17060
rect 26384 17057 26390 17060
rect 26384 17051 26448 17057
rect 26384 17017 26402 17051
rect 26436 17017 26448 17051
rect 26384 17011 26448 17017
rect 26384 17008 26390 17011
rect 15194 16980 15200 16992
rect 14967 16952 15200 16980
rect 14967 16949 14979 16952
rect 14921 16943 14979 16949
rect 15194 16940 15200 16952
rect 15252 16940 15258 16992
rect 17494 16980 17500 16992
rect 17407 16952 17500 16980
rect 17494 16940 17500 16952
rect 17552 16980 17558 16992
rect 18690 16980 18696 16992
rect 17552 16952 18696 16980
rect 17552 16940 17558 16952
rect 18690 16940 18696 16952
rect 18748 16940 18754 16992
rect 19429 16983 19487 16989
rect 19429 16949 19441 16983
rect 19475 16980 19487 16983
rect 19886 16980 19892 16992
rect 19475 16952 19892 16980
rect 19475 16949 19487 16952
rect 19429 16943 19487 16949
rect 19886 16940 19892 16952
rect 19944 16980 19950 16992
rect 20806 16980 20812 16992
rect 19944 16952 20812 16980
rect 19944 16940 19950 16952
rect 20806 16940 20812 16952
rect 20864 16980 20870 16992
rect 20901 16983 20959 16989
rect 20901 16980 20913 16983
rect 20864 16952 20913 16980
rect 20864 16940 20870 16952
rect 20901 16949 20913 16952
rect 20947 16949 20959 16983
rect 22462 16980 22468 16992
rect 22423 16952 22468 16980
rect 20901 16943 20959 16949
rect 22462 16940 22468 16952
rect 22520 16940 22526 16992
rect 27522 16980 27528 16992
rect 27483 16952 27528 16980
rect 27522 16940 27528 16952
rect 27580 16940 27586 16992
rect 1104 16890 28888 16912
rect 1104 16838 10982 16890
rect 11034 16838 11046 16890
rect 11098 16838 11110 16890
rect 11162 16838 11174 16890
rect 11226 16838 20982 16890
rect 21034 16838 21046 16890
rect 21098 16838 21110 16890
rect 21162 16838 21174 16890
rect 21226 16838 28888 16890
rect 1104 16816 28888 16838
rect 1673 16779 1731 16785
rect 1673 16745 1685 16779
rect 1719 16776 1731 16779
rect 2130 16776 2136 16788
rect 1719 16748 2136 16776
rect 1719 16745 1731 16748
rect 1673 16739 1731 16745
rect 2130 16736 2136 16748
rect 2188 16736 2194 16788
rect 2222 16736 2228 16788
rect 2280 16776 2286 16788
rect 3694 16776 3700 16788
rect 2280 16748 3700 16776
rect 2280 16736 2286 16748
rect 3694 16736 3700 16748
rect 3752 16736 3758 16788
rect 4706 16736 4712 16788
rect 4764 16776 4770 16788
rect 4985 16779 5043 16785
rect 4985 16776 4997 16779
rect 4764 16748 4997 16776
rect 4764 16736 4770 16748
rect 4985 16745 4997 16748
rect 5031 16745 5043 16779
rect 4985 16739 5043 16745
rect 7929 16779 7987 16785
rect 7929 16745 7941 16779
rect 7975 16776 7987 16779
rect 8478 16776 8484 16788
rect 7975 16748 8484 16776
rect 7975 16745 7987 16748
rect 7929 16739 7987 16745
rect 3142 16668 3148 16720
rect 3200 16708 3206 16720
rect 3329 16711 3387 16717
rect 3329 16708 3341 16711
rect 3200 16680 3341 16708
rect 3200 16668 3206 16680
rect 3329 16677 3341 16680
rect 3375 16708 3387 16711
rect 3418 16708 3424 16720
rect 3375 16680 3424 16708
rect 3375 16677 3387 16680
rect 3329 16671 3387 16677
rect 3418 16668 3424 16680
rect 3476 16668 3482 16720
rect 2038 16640 2044 16652
rect 1999 16612 2044 16640
rect 2038 16600 2044 16612
rect 2096 16600 2102 16652
rect 5000 16640 5028 16739
rect 8478 16736 8484 16748
rect 8536 16776 8542 16788
rect 9677 16779 9735 16785
rect 9677 16776 9689 16779
rect 8536 16748 9689 16776
rect 8536 16736 8542 16748
rect 9677 16745 9689 16748
rect 9723 16745 9735 16779
rect 9677 16739 9735 16745
rect 11241 16779 11299 16785
rect 11241 16745 11253 16779
rect 11287 16776 11299 16779
rect 11330 16776 11336 16788
rect 11287 16748 11336 16776
rect 11287 16745 11299 16748
rect 11241 16739 11299 16745
rect 11330 16736 11336 16748
rect 11388 16736 11394 16788
rect 12805 16779 12863 16785
rect 12805 16745 12817 16779
rect 12851 16776 12863 16779
rect 13078 16776 13084 16788
rect 12851 16748 13084 16776
rect 12851 16745 12863 16748
rect 12805 16739 12863 16745
rect 13078 16736 13084 16748
rect 13136 16736 13142 16788
rect 13725 16779 13783 16785
rect 13725 16745 13737 16779
rect 13771 16776 13783 16779
rect 13814 16776 13820 16788
rect 13771 16748 13820 16776
rect 13771 16745 13783 16748
rect 13725 16739 13783 16745
rect 13814 16736 13820 16748
rect 13872 16736 13878 16788
rect 15289 16779 15347 16785
rect 15289 16745 15301 16779
rect 15335 16776 15347 16779
rect 17218 16776 17224 16788
rect 15335 16748 17224 16776
rect 15335 16745 15347 16748
rect 15289 16739 15347 16745
rect 17218 16736 17224 16748
rect 17276 16776 17282 16788
rect 17313 16779 17371 16785
rect 17313 16776 17325 16779
rect 17276 16748 17325 16776
rect 17276 16736 17282 16748
rect 17313 16745 17325 16748
rect 17359 16745 17371 16779
rect 18414 16776 18420 16788
rect 18375 16748 18420 16776
rect 17313 16739 17371 16745
rect 18414 16736 18420 16748
rect 18472 16736 18478 16788
rect 20717 16779 20775 16785
rect 20717 16745 20729 16779
rect 20763 16776 20775 16779
rect 21358 16776 21364 16788
rect 20763 16748 21364 16776
rect 20763 16745 20775 16748
rect 20717 16739 20775 16745
rect 21358 16736 21364 16748
rect 21416 16736 21422 16788
rect 22462 16736 22468 16788
rect 22520 16776 22526 16788
rect 23017 16779 23075 16785
rect 23017 16776 23029 16779
rect 22520 16748 23029 16776
rect 22520 16736 22526 16748
rect 23017 16745 23029 16748
rect 23063 16745 23075 16779
rect 24670 16776 24676 16788
rect 24631 16748 24676 16776
rect 23017 16739 23075 16745
rect 24670 16736 24676 16748
rect 24728 16736 24734 16788
rect 24854 16776 24860 16788
rect 24815 16748 24860 16776
rect 24854 16736 24860 16748
rect 24912 16736 24918 16788
rect 25314 16776 25320 16788
rect 25275 16748 25320 16776
rect 25314 16736 25320 16748
rect 25372 16776 25378 16788
rect 26513 16779 26571 16785
rect 26513 16776 26525 16779
rect 25372 16748 26525 16776
rect 25372 16736 25378 16748
rect 26513 16745 26525 16748
rect 26559 16745 26571 16779
rect 26513 16739 26571 16745
rect 5626 16717 5632 16720
rect 5620 16708 5632 16717
rect 5587 16680 5632 16708
rect 5620 16671 5632 16680
rect 5626 16668 5632 16671
rect 5684 16668 5690 16720
rect 8294 16668 8300 16720
rect 8352 16708 8358 16720
rect 8389 16711 8447 16717
rect 8389 16708 8401 16711
rect 8352 16680 8401 16708
rect 8352 16668 8358 16680
rect 8389 16677 8401 16680
rect 8435 16677 8447 16711
rect 8389 16671 8447 16677
rect 9125 16711 9183 16717
rect 9125 16677 9137 16711
rect 9171 16708 9183 16711
rect 10137 16711 10195 16717
rect 10137 16708 10149 16711
rect 9171 16680 10149 16708
rect 9171 16677 9183 16680
rect 9125 16671 9183 16677
rect 10137 16677 10149 16680
rect 10183 16708 10195 16711
rect 10778 16708 10784 16720
rect 10183 16680 10784 16708
rect 10183 16677 10195 16680
rect 10137 16671 10195 16677
rect 10778 16668 10784 16680
rect 10836 16668 10842 16720
rect 15749 16711 15807 16717
rect 15749 16677 15761 16711
rect 15795 16708 15807 16711
rect 16574 16708 16580 16720
rect 15795 16680 16580 16708
rect 15795 16677 15807 16680
rect 15749 16671 15807 16677
rect 16574 16668 16580 16680
rect 16632 16668 16638 16720
rect 20349 16711 20407 16717
rect 20349 16677 20361 16711
rect 20395 16708 20407 16711
rect 21174 16708 21180 16720
rect 20395 16680 21180 16708
rect 20395 16677 20407 16680
rect 20349 16671 20407 16677
rect 21174 16668 21180 16680
rect 21232 16668 21238 16720
rect 25222 16708 25228 16720
rect 25183 16680 25228 16708
rect 25222 16668 25228 16680
rect 25280 16668 25286 16720
rect 5350 16640 5356 16652
rect 5000 16612 5356 16640
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 7558 16640 7564 16652
rect 7519 16612 7564 16640
rect 7558 16600 7564 16612
rect 7616 16600 7622 16652
rect 8018 16600 8024 16652
rect 8076 16600 8082 16652
rect 8481 16643 8539 16649
rect 8481 16609 8493 16643
rect 8527 16640 8539 16643
rect 8754 16640 8760 16652
rect 8527 16612 8760 16640
rect 8527 16609 8539 16612
rect 8481 16603 8539 16609
rect 8754 16600 8760 16612
rect 8812 16600 8818 16652
rect 9493 16643 9551 16649
rect 9493 16609 9505 16643
rect 9539 16640 9551 16643
rect 9582 16640 9588 16652
rect 9539 16612 9588 16640
rect 9539 16609 9551 16612
rect 9493 16603 9551 16609
rect 9582 16600 9588 16612
rect 9640 16600 9646 16652
rect 10045 16643 10103 16649
rect 10045 16609 10057 16643
rect 10091 16640 10103 16643
rect 10410 16640 10416 16652
rect 10091 16612 10416 16640
rect 10091 16609 10103 16612
rect 10045 16603 10103 16609
rect 10410 16600 10416 16612
rect 10468 16600 10474 16652
rect 11514 16600 11520 16652
rect 11572 16640 11578 16652
rect 11681 16643 11739 16649
rect 11681 16640 11693 16643
rect 11572 16612 11693 16640
rect 11572 16600 11578 16612
rect 11681 16609 11693 16612
rect 11727 16609 11739 16643
rect 11681 16603 11739 16609
rect 13814 16600 13820 16652
rect 13872 16640 13878 16652
rect 15013 16643 15071 16649
rect 15013 16640 15025 16643
rect 13872 16612 15025 16640
rect 13872 16600 13878 16612
rect 15013 16609 15025 16612
rect 15059 16640 15071 16643
rect 15470 16640 15476 16652
rect 15059 16612 15476 16640
rect 15059 16609 15071 16612
rect 15013 16603 15071 16609
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 15654 16600 15660 16652
rect 15712 16640 15718 16652
rect 16298 16640 16304 16652
rect 15712 16612 16304 16640
rect 15712 16600 15718 16612
rect 16298 16600 16304 16612
rect 16356 16600 16362 16652
rect 16666 16640 16672 16652
rect 16627 16612 16672 16640
rect 16666 16600 16672 16612
rect 16724 16640 16730 16652
rect 17221 16643 17279 16649
rect 17221 16640 17233 16643
rect 16724 16612 17233 16640
rect 16724 16600 16730 16612
rect 17221 16609 17233 16612
rect 17267 16609 17279 16643
rect 18782 16640 18788 16652
rect 18743 16612 18788 16640
rect 17221 16603 17279 16609
rect 18782 16600 18788 16612
rect 18840 16600 18846 16652
rect 21352 16643 21410 16649
rect 21352 16609 21364 16643
rect 21398 16640 21410 16643
rect 21634 16640 21640 16652
rect 21398 16612 21640 16640
rect 21398 16609 21410 16612
rect 21352 16603 21410 16609
rect 21634 16600 21640 16612
rect 21692 16600 21698 16652
rect 23566 16640 23572 16652
rect 23527 16612 23572 16640
rect 23566 16600 23572 16612
rect 23624 16600 23630 16652
rect 26878 16640 26884 16652
rect 26839 16612 26884 16640
rect 26878 16600 26884 16612
rect 26936 16600 26942 16652
rect 26970 16600 26976 16652
rect 27028 16640 27034 16652
rect 27028 16612 27073 16640
rect 27028 16600 27034 16612
rect 2130 16532 2136 16584
rect 2188 16572 2194 16584
rect 2317 16575 2375 16581
rect 2188 16544 2233 16572
rect 2188 16532 2194 16544
rect 2317 16541 2329 16575
rect 2363 16541 2375 16575
rect 2317 16535 2375 16541
rect 2332 16504 2360 16535
rect 2866 16532 2872 16584
rect 2924 16572 2930 16584
rect 4065 16575 4123 16581
rect 4065 16572 4077 16575
rect 2924 16544 4077 16572
rect 2924 16532 2930 16544
rect 4065 16541 4077 16544
rect 4111 16541 4123 16575
rect 4065 16535 4123 16541
rect 2406 16504 2412 16516
rect 2332 16476 2412 16504
rect 2406 16464 2412 16476
rect 2464 16504 2470 16516
rect 8036 16513 8064 16600
rect 8573 16575 8631 16581
rect 8573 16541 8585 16575
rect 8619 16572 8631 16575
rect 9030 16572 9036 16584
rect 8619 16544 9036 16572
rect 8619 16541 8631 16544
rect 8573 16535 8631 16541
rect 9030 16532 9036 16544
rect 9088 16572 9094 16584
rect 10226 16572 10232 16584
rect 9088 16544 10232 16572
rect 9088 16532 9094 16544
rect 10226 16532 10232 16544
rect 10284 16532 10290 16584
rect 11422 16572 11428 16584
rect 11383 16544 11428 16572
rect 11422 16532 11428 16544
rect 11480 16532 11486 16584
rect 14277 16575 14335 16581
rect 14277 16541 14289 16575
rect 14323 16572 14335 16575
rect 14458 16572 14464 16584
rect 14323 16544 14464 16572
rect 14323 16541 14335 16544
rect 14277 16535 14335 16541
rect 14458 16532 14464 16544
rect 14516 16572 14522 16584
rect 15102 16572 15108 16584
rect 14516 16544 15108 16572
rect 14516 16532 14522 16544
rect 15102 16532 15108 16544
rect 15160 16572 15166 16584
rect 15841 16575 15899 16581
rect 15841 16572 15853 16575
rect 15160 16544 15853 16572
rect 15160 16532 15166 16544
rect 15841 16541 15853 16544
rect 15887 16541 15899 16575
rect 17402 16572 17408 16584
rect 17363 16544 17408 16572
rect 15841 16535 15899 16541
rect 17402 16532 17408 16544
rect 17460 16532 17466 16584
rect 17586 16532 17592 16584
rect 17644 16572 17650 16584
rect 18877 16575 18935 16581
rect 18877 16572 18889 16575
rect 17644 16544 18889 16572
rect 17644 16532 17650 16544
rect 18877 16541 18889 16544
rect 18923 16541 18935 16575
rect 19058 16572 19064 16584
rect 19019 16544 19064 16572
rect 18877 16535 18935 16541
rect 19058 16532 19064 16544
rect 19116 16532 19122 16584
rect 20806 16532 20812 16584
rect 20864 16572 20870 16584
rect 21085 16575 21143 16581
rect 21085 16572 21097 16575
rect 20864 16544 21097 16572
rect 20864 16532 20870 16544
rect 21085 16541 21097 16544
rect 21131 16541 21143 16575
rect 21085 16535 21143 16541
rect 24670 16532 24676 16584
rect 24728 16572 24734 16584
rect 25409 16575 25467 16581
rect 25409 16572 25421 16575
rect 24728 16544 25421 16572
rect 24728 16532 24734 16544
rect 25409 16541 25421 16544
rect 25455 16541 25467 16575
rect 25409 16535 25467 16541
rect 25866 16532 25872 16584
rect 25924 16572 25930 16584
rect 27065 16575 27123 16581
rect 27065 16572 27077 16575
rect 25924 16544 27077 16572
rect 25924 16532 25930 16544
rect 27065 16541 27077 16544
rect 27111 16541 27123 16575
rect 27065 16535 27123 16541
rect 8021 16507 8079 16513
rect 2464 16476 3740 16504
rect 2464 16464 2470 16476
rect 3712 16448 3740 16476
rect 8021 16473 8033 16507
rect 8067 16473 8079 16507
rect 16850 16504 16856 16516
rect 16811 16476 16856 16504
rect 8021 16467 8079 16473
rect 16850 16464 16856 16476
rect 16908 16464 16914 16516
rect 24118 16504 24124 16516
rect 24031 16476 24124 16504
rect 24118 16464 24124 16476
rect 24176 16504 24182 16516
rect 25884 16504 25912 16532
rect 24176 16476 25912 16504
rect 24176 16464 24182 16476
rect 2682 16436 2688 16448
rect 2643 16408 2688 16436
rect 2682 16396 2688 16408
rect 2740 16396 2746 16448
rect 3694 16436 3700 16448
rect 3655 16408 3700 16436
rect 3694 16396 3700 16408
rect 3752 16396 3758 16448
rect 4522 16436 4528 16448
rect 4483 16408 4528 16436
rect 4522 16396 4528 16408
rect 4580 16396 4586 16448
rect 6362 16396 6368 16448
rect 6420 16436 6426 16448
rect 6733 16439 6791 16445
rect 6733 16436 6745 16439
rect 6420 16408 6745 16436
rect 6420 16396 6426 16408
rect 6733 16405 6745 16408
rect 6779 16405 6791 16439
rect 6733 16399 6791 16405
rect 10873 16439 10931 16445
rect 10873 16405 10885 16439
rect 10919 16436 10931 16439
rect 11054 16436 11060 16448
rect 10919 16408 11060 16436
rect 10919 16405 10931 16408
rect 10873 16399 10931 16405
rect 11054 16396 11060 16408
rect 11112 16396 11118 16448
rect 16393 16439 16451 16445
rect 16393 16405 16405 16439
rect 16439 16436 16451 16439
rect 17862 16436 17868 16448
rect 16439 16408 17868 16436
rect 16439 16405 16451 16408
rect 16393 16399 16451 16405
rect 17862 16396 17868 16408
rect 17920 16396 17926 16448
rect 18138 16436 18144 16448
rect 18099 16408 18144 16436
rect 18138 16396 18144 16408
rect 18196 16396 18202 16448
rect 22465 16439 22523 16445
rect 22465 16405 22477 16439
rect 22511 16436 22523 16439
rect 22554 16436 22560 16448
rect 22511 16408 22560 16436
rect 22511 16405 22523 16408
rect 22465 16399 22523 16405
rect 22554 16396 22560 16408
rect 22612 16396 22618 16448
rect 23474 16436 23480 16448
rect 23435 16408 23480 16436
rect 23474 16396 23480 16408
rect 23532 16396 23538 16448
rect 26237 16439 26295 16445
rect 26237 16405 26249 16439
rect 26283 16436 26295 16439
rect 26326 16436 26332 16448
rect 26283 16408 26332 16436
rect 26283 16405 26295 16408
rect 26237 16399 26295 16405
rect 26326 16396 26332 16408
rect 26384 16396 26390 16448
rect 1104 16346 28888 16368
rect 1104 16294 5982 16346
rect 6034 16294 6046 16346
rect 6098 16294 6110 16346
rect 6162 16294 6174 16346
rect 6226 16294 15982 16346
rect 16034 16294 16046 16346
rect 16098 16294 16110 16346
rect 16162 16294 16174 16346
rect 16226 16294 25982 16346
rect 26034 16294 26046 16346
rect 26098 16294 26110 16346
rect 26162 16294 26174 16346
rect 26226 16294 28888 16346
rect 1104 16272 28888 16294
rect 2866 16232 2872 16244
rect 2827 16204 2872 16232
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 4338 16192 4344 16244
rect 4396 16232 4402 16244
rect 4709 16235 4767 16241
rect 4709 16232 4721 16235
rect 4396 16204 4721 16232
rect 4396 16192 4402 16204
rect 4709 16201 4721 16204
rect 4755 16201 4767 16235
rect 5350 16232 5356 16244
rect 5311 16204 5356 16232
rect 4709 16195 4767 16201
rect 5350 16192 5356 16204
rect 5408 16192 5414 16244
rect 5626 16192 5632 16244
rect 5684 16232 5690 16244
rect 5721 16235 5779 16241
rect 5721 16232 5733 16235
rect 5684 16204 5733 16232
rect 5684 16192 5690 16204
rect 5721 16201 5733 16204
rect 5767 16201 5779 16235
rect 5721 16195 5779 16201
rect 8113 16235 8171 16241
rect 8113 16201 8125 16235
rect 8159 16232 8171 16235
rect 8202 16232 8208 16244
rect 8159 16204 8208 16232
rect 8159 16201 8171 16204
rect 8113 16195 8171 16201
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 9490 16192 9496 16244
rect 9548 16232 9554 16244
rect 9585 16235 9643 16241
rect 9585 16232 9597 16235
rect 9548 16204 9597 16232
rect 9548 16192 9554 16204
rect 9585 16201 9597 16204
rect 9631 16201 9643 16235
rect 10778 16232 10784 16244
rect 10739 16204 10784 16232
rect 9585 16195 9643 16201
rect 10778 16192 10784 16204
rect 10836 16192 10842 16244
rect 11790 16232 11796 16244
rect 11751 16204 11796 16232
rect 11790 16192 11796 16204
rect 11848 16192 11854 16244
rect 12434 16192 12440 16244
rect 12492 16232 12498 16244
rect 12492 16204 12537 16232
rect 12492 16192 12498 16204
rect 13078 16192 13084 16244
rect 13136 16232 13142 16244
rect 13449 16235 13507 16241
rect 13449 16232 13461 16235
rect 13136 16204 13461 16232
rect 13136 16192 13142 16204
rect 13449 16201 13461 16204
rect 13495 16201 13507 16235
rect 13449 16195 13507 16201
rect 15470 16192 15476 16244
rect 15528 16232 15534 16244
rect 15565 16235 15623 16241
rect 15565 16232 15577 16235
rect 15528 16204 15577 16232
rect 15528 16192 15534 16204
rect 15565 16201 15577 16204
rect 15611 16232 15623 16235
rect 17221 16235 17279 16241
rect 17221 16232 17233 16235
rect 15611 16204 17233 16232
rect 15611 16201 15623 16204
rect 15565 16195 15623 16201
rect 17221 16201 17233 16204
rect 17267 16232 17279 16235
rect 17402 16232 17408 16244
rect 17267 16204 17408 16232
rect 17267 16201 17279 16204
rect 17221 16195 17279 16201
rect 17402 16192 17408 16204
rect 17460 16192 17466 16244
rect 21266 16192 21272 16244
rect 21324 16232 21330 16244
rect 21361 16235 21419 16241
rect 21361 16232 21373 16235
rect 21324 16204 21373 16232
rect 21324 16192 21330 16204
rect 21361 16201 21373 16204
rect 21407 16201 21419 16235
rect 24578 16232 24584 16244
rect 24539 16204 24584 16232
rect 21361 16195 21419 16201
rect 24578 16192 24584 16204
rect 24636 16192 24642 16244
rect 25222 16192 25228 16244
rect 25280 16232 25286 16244
rect 25593 16235 25651 16241
rect 25593 16232 25605 16235
rect 25280 16204 25605 16232
rect 25280 16192 25286 16204
rect 25593 16201 25605 16204
rect 25639 16232 25651 16235
rect 25682 16232 25688 16244
rect 25639 16204 25688 16232
rect 25639 16201 25651 16204
rect 25593 16195 25651 16201
rect 25682 16192 25688 16204
rect 25740 16192 25746 16244
rect 28074 16232 28080 16244
rect 28035 16204 28080 16232
rect 28074 16192 28080 16204
rect 28132 16192 28138 16244
rect 2409 16099 2467 16105
rect 2409 16065 2421 16099
rect 2455 16096 2467 16099
rect 2682 16096 2688 16108
rect 2455 16068 2688 16096
rect 2455 16065 2467 16068
rect 2409 16059 2467 16065
rect 2682 16056 2688 16068
rect 2740 16056 2746 16108
rect 7377 16099 7435 16105
rect 7377 16065 7389 16099
rect 7423 16096 7435 16099
rect 7423 16068 8340 16096
rect 7423 16065 7435 16068
rect 7377 16059 7435 16065
rect 1486 15988 1492 16040
rect 1544 16028 1550 16040
rect 3145 16031 3203 16037
rect 3145 16028 3157 16031
rect 1544 16000 3157 16028
rect 1544 15988 1550 16000
rect 3145 15997 3157 16000
rect 3191 16028 3203 16031
rect 3329 16031 3387 16037
rect 3329 16028 3341 16031
rect 3191 16000 3341 16028
rect 3191 15997 3203 16000
rect 3145 15991 3203 15997
rect 3329 15997 3341 16000
rect 3375 15997 3387 16031
rect 3329 15991 3387 15997
rect 3418 15988 3424 16040
rect 3476 16028 3482 16040
rect 3585 16031 3643 16037
rect 3585 16028 3597 16031
rect 3476 16000 3597 16028
rect 3476 15988 3482 16000
rect 3585 15997 3597 16000
rect 3631 15997 3643 16031
rect 3585 15991 3643 15997
rect 5442 15988 5448 16040
rect 5500 16028 5506 16040
rect 8110 16028 8116 16040
rect 5500 16000 8116 16028
rect 5500 15988 5506 16000
rect 8110 15988 8116 16000
rect 8168 16028 8174 16040
rect 8205 16031 8263 16037
rect 8205 16028 8217 16031
rect 8168 16000 8217 16028
rect 8168 15988 8174 16000
rect 8205 15997 8217 16000
rect 8251 15997 8263 16031
rect 8205 15991 8263 15997
rect 1578 15920 1584 15972
rect 1636 15960 1642 15972
rect 1673 15963 1731 15969
rect 1673 15960 1685 15963
rect 1636 15932 1685 15960
rect 1636 15920 1642 15932
rect 1673 15929 1685 15932
rect 1719 15960 1731 15963
rect 2133 15963 2191 15969
rect 2133 15960 2145 15963
rect 1719 15932 2145 15960
rect 1719 15929 1731 15932
rect 1673 15923 1731 15929
rect 2133 15929 2145 15932
rect 2179 15960 2191 15963
rect 4246 15960 4252 15972
rect 2179 15932 4252 15960
rect 2179 15929 2191 15932
rect 2133 15923 2191 15929
rect 4246 15920 4252 15932
rect 4304 15920 4310 15972
rect 8312 15960 8340 16068
rect 11054 16056 11060 16108
rect 11112 16096 11118 16108
rect 11330 16096 11336 16108
rect 11112 16068 11336 16096
rect 11112 16056 11118 16068
rect 11330 16056 11336 16068
rect 11388 16056 11394 16108
rect 12253 16099 12311 16105
rect 12253 16065 12265 16099
rect 12299 16096 12311 16099
rect 12342 16096 12348 16108
rect 12299 16068 12348 16096
rect 12299 16065 12311 16068
rect 12253 16059 12311 16065
rect 12342 16056 12348 16068
rect 12400 16056 12406 16108
rect 13096 16105 13124 16192
rect 16209 16167 16267 16173
rect 16209 16133 16221 16167
rect 16255 16164 16267 16167
rect 16298 16164 16304 16176
rect 16255 16136 16304 16164
rect 16255 16133 16267 16136
rect 16209 16127 16267 16133
rect 16298 16124 16304 16136
rect 16356 16124 16362 16176
rect 20809 16167 20867 16173
rect 20809 16133 20821 16167
rect 20855 16164 20867 16167
rect 21634 16164 21640 16176
rect 20855 16136 21640 16164
rect 20855 16133 20867 16136
rect 20809 16127 20867 16133
rect 21634 16124 21640 16136
rect 21692 16124 21698 16176
rect 21910 16124 21916 16176
rect 21968 16164 21974 16176
rect 24489 16167 24547 16173
rect 21968 16136 22048 16164
rect 21968 16124 21974 16136
rect 13081 16099 13139 16105
rect 13081 16065 13093 16099
rect 13127 16065 13139 16099
rect 13081 16059 13139 16065
rect 21542 16056 21548 16108
rect 21600 16056 21606 16108
rect 22020 16105 22048 16136
rect 24489 16133 24501 16167
rect 24535 16164 24547 16167
rect 24670 16164 24676 16176
rect 24535 16136 24676 16164
rect 24535 16133 24547 16136
rect 24489 16127 24547 16133
rect 24670 16124 24676 16136
rect 24728 16164 24734 16176
rect 25958 16164 25964 16176
rect 24728 16136 25176 16164
rect 25919 16136 25964 16164
rect 24728 16124 24734 16136
rect 25148 16105 25176 16136
rect 25958 16124 25964 16136
rect 26016 16124 26022 16176
rect 22005 16099 22063 16105
rect 22005 16065 22017 16099
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 25133 16099 25191 16105
rect 25133 16065 25145 16099
rect 25179 16065 25191 16099
rect 25133 16059 25191 16065
rect 10594 15988 10600 16040
rect 10652 16028 10658 16040
rect 11606 16028 11612 16040
rect 10652 16000 11612 16028
rect 10652 15988 10658 16000
rect 11606 15988 11612 16000
rect 11664 15988 11670 16040
rect 14458 16037 14464 16040
rect 14185 16031 14243 16037
rect 14185 15997 14197 16031
rect 14231 15997 14243 16031
rect 14452 16028 14464 16037
rect 14419 16000 14464 16028
rect 14185 15991 14243 15997
rect 14452 15991 14464 16000
rect 8386 15960 8392 15972
rect 8312 15932 8392 15960
rect 8386 15920 8392 15932
rect 8444 15969 8450 15972
rect 8444 15963 8508 15969
rect 8444 15929 8462 15963
rect 8496 15929 8508 15963
rect 8444 15923 8508 15929
rect 10689 15963 10747 15969
rect 10689 15929 10701 15963
rect 10735 15960 10747 15963
rect 10735 15932 11284 15960
rect 10735 15929 10747 15932
rect 10689 15923 10747 15929
rect 8444 15920 8450 15923
rect 1762 15892 1768 15904
rect 1723 15864 1768 15892
rect 1762 15852 1768 15864
rect 1820 15852 1826 15904
rect 2225 15895 2283 15901
rect 2225 15861 2237 15895
rect 2271 15892 2283 15895
rect 2498 15892 2504 15904
rect 2271 15864 2504 15892
rect 2271 15861 2283 15864
rect 2225 15855 2283 15861
rect 2498 15852 2504 15864
rect 2556 15852 2562 15904
rect 6086 15892 6092 15904
rect 6047 15864 6092 15892
rect 6086 15852 6092 15864
rect 6144 15852 6150 15904
rect 7745 15895 7803 15901
rect 7745 15861 7757 15895
rect 7791 15892 7803 15895
rect 8754 15892 8760 15904
rect 7791 15864 8760 15892
rect 7791 15861 7803 15864
rect 7745 15855 7803 15861
rect 8754 15852 8760 15864
rect 8812 15852 8818 15904
rect 10229 15895 10287 15901
rect 10229 15861 10241 15895
rect 10275 15892 10287 15895
rect 10410 15892 10416 15904
rect 10275 15864 10416 15892
rect 10275 15861 10287 15864
rect 10229 15855 10287 15861
rect 10410 15852 10416 15864
rect 10468 15852 10474 15904
rect 10778 15852 10784 15904
rect 10836 15892 10842 15904
rect 11256 15901 11284 15932
rect 11790 15920 11796 15972
rect 11848 15960 11854 15972
rect 11848 15932 12296 15960
rect 11848 15920 11854 15932
rect 11149 15895 11207 15901
rect 11149 15892 11161 15895
rect 10836 15864 11161 15892
rect 10836 15852 10842 15864
rect 11149 15861 11161 15864
rect 11195 15861 11207 15895
rect 11149 15855 11207 15861
rect 11241 15895 11299 15901
rect 11241 15861 11253 15895
rect 11287 15892 11299 15895
rect 11606 15892 11612 15904
rect 11287 15864 11612 15892
rect 11287 15861 11299 15864
rect 11241 15855 11299 15861
rect 11606 15852 11612 15864
rect 11664 15852 11670 15904
rect 12268 15892 12296 15932
rect 12342 15920 12348 15972
rect 12400 15960 12406 15972
rect 12805 15963 12863 15969
rect 12805 15960 12817 15963
rect 12400 15932 12817 15960
rect 12400 15920 12406 15932
rect 12805 15929 12817 15932
rect 12851 15929 12863 15963
rect 12805 15923 12863 15929
rect 13078 15920 13084 15972
rect 13136 15960 13142 15972
rect 14093 15963 14151 15969
rect 14093 15960 14105 15963
rect 13136 15932 14105 15960
rect 13136 15920 13142 15932
rect 14093 15929 14105 15932
rect 14139 15960 14151 15963
rect 14200 15960 14228 15991
rect 14458 15988 14464 15991
rect 14516 15988 14522 16040
rect 17862 15988 17868 16040
rect 17920 16028 17926 16040
rect 18049 16031 18107 16037
rect 18049 16028 18061 16031
rect 17920 16000 18061 16028
rect 17920 15988 17926 16000
rect 18049 15997 18061 16000
rect 18095 15997 18107 16031
rect 18049 15991 18107 15997
rect 18138 15988 18144 16040
rect 18196 16028 18202 16040
rect 18305 16031 18363 16037
rect 18305 16028 18317 16031
rect 18196 16000 18317 16028
rect 18196 15988 18202 16000
rect 18305 15997 18317 16000
rect 18351 15997 18363 16031
rect 21560 16028 21588 16056
rect 21821 16031 21879 16037
rect 21821 16028 21833 16031
rect 21560 16000 21833 16028
rect 18305 15991 18363 15997
rect 21821 15997 21833 16000
rect 21867 16028 21879 16031
rect 22741 16031 22799 16037
rect 22741 16028 22753 16031
rect 21867 16000 22753 16028
rect 21867 15997 21879 16000
rect 21821 15991 21879 15997
rect 22741 15997 22753 16000
rect 22787 15997 22799 16031
rect 22741 15991 22799 15997
rect 23474 15988 23480 16040
rect 23532 16028 23538 16040
rect 24762 16028 24768 16040
rect 23532 16000 24768 16028
rect 23532 15988 23538 16000
rect 24762 15988 24768 16000
rect 24820 16028 24826 16040
rect 24949 16031 25007 16037
rect 24949 16028 24961 16031
rect 24820 16000 24961 16028
rect 24820 15988 24826 16000
rect 24949 15997 24961 16000
rect 24995 15997 25007 16031
rect 26142 16028 26148 16040
rect 26103 16000 26148 16028
rect 24949 15991 25007 15997
rect 26142 15988 26148 16000
rect 26200 15988 26206 16040
rect 26418 16037 26424 16040
rect 26412 16028 26424 16037
rect 26331 16000 26424 16028
rect 26412 15991 26424 16000
rect 26476 16028 26482 16040
rect 27522 16028 27528 16040
rect 26476 16000 27528 16028
rect 26418 15988 26424 15991
rect 26476 15988 26482 16000
rect 27522 15988 27528 16000
rect 27580 15988 27586 16040
rect 15286 15960 15292 15972
rect 14139 15932 15292 15960
rect 14139 15929 14151 15932
rect 14093 15923 14151 15929
rect 15286 15920 15292 15932
rect 15344 15920 15350 15972
rect 16482 15920 16488 15972
rect 16540 15960 16546 15972
rect 16853 15963 16911 15969
rect 16853 15960 16865 15963
rect 16540 15932 16865 15960
rect 16540 15920 16546 15932
rect 16853 15929 16865 15932
rect 16899 15929 16911 15963
rect 16853 15923 16911 15929
rect 21729 15963 21787 15969
rect 21729 15929 21741 15963
rect 21775 15960 21787 15963
rect 22186 15960 22192 15972
rect 21775 15932 22192 15960
rect 21775 15929 21787 15932
rect 21729 15923 21787 15929
rect 22186 15920 22192 15932
rect 22244 15960 22250 15972
rect 23109 15963 23167 15969
rect 23109 15960 23121 15963
rect 22244 15932 23121 15960
rect 22244 15920 22250 15932
rect 23109 15929 23121 15932
rect 23155 15929 23167 15963
rect 23109 15923 23167 15929
rect 23198 15920 23204 15972
rect 23256 15960 23262 15972
rect 24121 15963 24179 15969
rect 24121 15960 24133 15963
rect 23256 15932 24133 15960
rect 23256 15920 23262 15932
rect 24121 15929 24133 15932
rect 24167 15960 24179 15963
rect 25041 15963 25099 15969
rect 25041 15960 25053 15963
rect 24167 15932 25053 15960
rect 24167 15929 24179 15932
rect 24121 15923 24179 15929
rect 25041 15929 25053 15932
rect 25087 15929 25099 15963
rect 25041 15923 25099 15929
rect 12894 15892 12900 15904
rect 12268 15864 12900 15892
rect 12894 15852 12900 15864
rect 12952 15852 12958 15904
rect 16574 15892 16580 15904
rect 16535 15864 16580 15892
rect 16574 15852 16580 15864
rect 16632 15852 16638 15904
rect 17586 15852 17592 15904
rect 17644 15892 17650 15904
rect 17773 15895 17831 15901
rect 17773 15892 17785 15895
rect 17644 15864 17785 15892
rect 17644 15852 17650 15864
rect 17773 15861 17785 15864
rect 17819 15861 17831 15895
rect 17773 15855 17831 15861
rect 18506 15852 18512 15904
rect 18564 15892 18570 15904
rect 19429 15895 19487 15901
rect 19429 15892 19441 15895
rect 18564 15864 19441 15892
rect 18564 15852 18570 15864
rect 19429 15861 19441 15864
rect 19475 15861 19487 15895
rect 19978 15892 19984 15904
rect 19939 15864 19984 15892
rect 19429 15855 19487 15861
rect 19978 15852 19984 15864
rect 20036 15852 20042 15904
rect 20806 15852 20812 15904
rect 20864 15892 20870 15904
rect 21085 15895 21143 15901
rect 21085 15892 21097 15895
rect 20864 15864 21097 15892
rect 20864 15852 20870 15864
rect 21085 15861 21097 15864
rect 21131 15861 21143 15895
rect 21085 15855 21143 15861
rect 21910 15852 21916 15904
rect 21968 15892 21974 15904
rect 22373 15895 22431 15901
rect 22373 15892 22385 15895
rect 21968 15864 22385 15892
rect 21968 15852 21974 15864
rect 22373 15861 22385 15864
rect 22419 15892 22431 15895
rect 22554 15892 22560 15904
rect 22419 15864 22560 15892
rect 22419 15861 22431 15864
rect 22373 15855 22431 15861
rect 22554 15852 22560 15864
rect 22612 15852 22618 15904
rect 27338 15852 27344 15904
rect 27396 15892 27402 15904
rect 27525 15895 27583 15901
rect 27525 15892 27537 15895
rect 27396 15864 27537 15892
rect 27396 15852 27402 15864
rect 27525 15861 27537 15864
rect 27571 15861 27583 15895
rect 27525 15855 27583 15861
rect 1104 15802 28888 15824
rect 1104 15750 10982 15802
rect 11034 15750 11046 15802
rect 11098 15750 11110 15802
rect 11162 15750 11174 15802
rect 11226 15750 20982 15802
rect 21034 15750 21046 15802
rect 21098 15750 21110 15802
rect 21162 15750 21174 15802
rect 21226 15750 28888 15802
rect 1104 15728 28888 15750
rect 2774 15648 2780 15700
rect 2832 15688 2838 15700
rect 4065 15691 4123 15697
rect 4065 15688 4077 15691
rect 2832 15660 4077 15688
rect 2832 15648 2838 15660
rect 4065 15657 4077 15660
rect 4111 15657 4123 15691
rect 4522 15688 4528 15700
rect 4483 15660 4528 15688
rect 4065 15651 4123 15657
rect 4522 15648 4528 15660
rect 4580 15648 4586 15700
rect 8110 15648 8116 15700
rect 8168 15688 8174 15700
rect 8205 15691 8263 15697
rect 8205 15688 8217 15691
rect 8168 15660 8217 15688
rect 8168 15648 8174 15660
rect 8205 15657 8217 15660
rect 8251 15688 8263 15691
rect 8294 15688 8300 15700
rect 8251 15660 8300 15688
rect 8251 15657 8263 15660
rect 8205 15651 8263 15657
rect 8294 15648 8300 15660
rect 8352 15648 8358 15700
rect 8570 15688 8576 15700
rect 8531 15660 8576 15688
rect 8570 15648 8576 15660
rect 8628 15648 8634 15700
rect 9674 15688 9680 15700
rect 9635 15660 9680 15688
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 10226 15688 10232 15700
rect 9784 15660 10232 15688
rect 7929 15623 7987 15629
rect 7929 15589 7941 15623
rect 7975 15620 7987 15623
rect 8386 15620 8392 15632
rect 7975 15592 8392 15620
rect 7975 15589 7987 15592
rect 7929 15583 7987 15589
rect 8386 15580 8392 15592
rect 8444 15620 8450 15632
rect 9125 15623 9183 15629
rect 9125 15620 9137 15623
rect 8444 15592 9137 15620
rect 8444 15580 8450 15592
rect 9125 15589 9137 15592
rect 9171 15620 9183 15623
rect 9493 15623 9551 15629
rect 9493 15620 9505 15623
rect 9171 15592 9505 15620
rect 9171 15589 9183 15592
rect 9125 15583 9183 15589
rect 9493 15589 9505 15592
rect 9539 15620 9551 15623
rect 9784 15620 9812 15660
rect 10226 15648 10232 15660
rect 10284 15688 10290 15700
rect 13173 15691 13231 15697
rect 13173 15688 13185 15691
rect 10284 15660 13185 15688
rect 10284 15648 10290 15660
rect 13173 15657 13185 15660
rect 13219 15657 13231 15691
rect 14458 15688 14464 15700
rect 14419 15660 14464 15688
rect 13173 15651 13231 15657
rect 14458 15648 14464 15660
rect 14516 15648 14522 15700
rect 17218 15688 17224 15700
rect 17179 15660 17224 15688
rect 17218 15648 17224 15660
rect 17276 15648 17282 15700
rect 17773 15691 17831 15697
rect 17773 15657 17785 15691
rect 17819 15688 17831 15691
rect 19058 15688 19064 15700
rect 17819 15660 19064 15688
rect 17819 15657 17831 15660
rect 17773 15651 17831 15657
rect 19058 15648 19064 15660
rect 19116 15648 19122 15700
rect 21085 15691 21143 15697
rect 21085 15657 21097 15691
rect 21131 15688 21143 15691
rect 21358 15688 21364 15700
rect 21131 15660 21364 15688
rect 21131 15657 21143 15660
rect 21085 15651 21143 15657
rect 21358 15648 21364 15660
rect 21416 15648 21422 15700
rect 21634 15648 21640 15700
rect 21692 15688 21698 15700
rect 22097 15691 22155 15697
rect 22097 15688 22109 15691
rect 21692 15660 22109 15688
rect 21692 15648 21698 15660
rect 22097 15657 22109 15660
rect 22143 15657 22155 15691
rect 23198 15688 23204 15700
rect 23159 15660 23204 15688
rect 22097 15651 22155 15657
rect 23198 15648 23204 15660
rect 23256 15648 23262 15700
rect 24762 15688 24768 15700
rect 24723 15660 24768 15688
rect 24762 15648 24768 15660
rect 24820 15648 24826 15700
rect 25866 15688 25872 15700
rect 25827 15660 25872 15688
rect 25866 15648 25872 15660
rect 25924 15648 25930 15700
rect 27522 15688 27528 15700
rect 27483 15660 27528 15688
rect 27522 15648 27528 15660
rect 27580 15648 27586 15700
rect 9539 15592 9812 15620
rect 9539 15589 9551 15592
rect 9493 15583 9551 15589
rect 11330 15580 11336 15632
rect 11388 15620 11394 15632
rect 12038 15623 12096 15629
rect 12038 15620 12050 15623
rect 11388 15592 12050 15620
rect 11388 15580 11394 15592
rect 12038 15589 12050 15592
rect 12084 15620 12096 15623
rect 12158 15620 12164 15632
rect 12084 15592 12164 15620
rect 12084 15589 12096 15592
rect 12038 15583 12096 15589
rect 12158 15580 12164 15592
rect 12216 15580 12222 15632
rect 15562 15629 15568 15632
rect 15556 15620 15568 15629
rect 15523 15592 15568 15620
rect 15556 15583 15568 15592
rect 15562 15580 15568 15583
rect 15620 15580 15626 15632
rect 1486 15552 1492 15564
rect 1447 15524 1492 15552
rect 1486 15512 1492 15524
rect 1544 15512 1550 15564
rect 1756 15555 1814 15561
rect 1756 15521 1768 15555
rect 1802 15552 1814 15555
rect 2590 15552 2596 15564
rect 1802 15524 2596 15552
rect 1802 15521 1814 15524
rect 1756 15515 1814 15521
rect 2590 15512 2596 15524
rect 2648 15512 2654 15564
rect 4430 15552 4436 15564
rect 4391 15524 4436 15552
rect 4430 15512 4436 15524
rect 4488 15512 4494 15564
rect 5261 15555 5319 15561
rect 5261 15521 5273 15555
rect 5307 15552 5319 15555
rect 5988 15555 6046 15561
rect 5988 15552 6000 15555
rect 5307 15524 6000 15552
rect 5307 15521 5319 15524
rect 5261 15515 5319 15521
rect 5988 15521 6000 15524
rect 6034 15552 6046 15555
rect 6362 15552 6368 15564
rect 6034 15524 6368 15552
rect 6034 15521 6046 15524
rect 5988 15515 6046 15521
rect 6362 15512 6368 15524
rect 6420 15512 6426 15564
rect 9674 15512 9680 15564
rect 9732 15552 9738 15564
rect 10045 15555 10103 15561
rect 10045 15552 10057 15555
rect 9732 15524 10057 15552
rect 9732 15512 9738 15524
rect 10045 15521 10057 15524
rect 10091 15521 10103 15555
rect 10045 15515 10103 15521
rect 17402 15512 17408 15564
rect 17460 15552 17466 15564
rect 18506 15561 18512 15564
rect 18489 15555 18512 15561
rect 18489 15552 18501 15555
rect 17460 15524 18501 15552
rect 17460 15512 17466 15524
rect 18489 15521 18501 15524
rect 18564 15552 18570 15564
rect 18564 15524 18637 15552
rect 18489 15515 18512 15521
rect 18506 15512 18512 15515
rect 18564 15512 18570 15524
rect 20622 15512 20628 15564
rect 20680 15552 20686 15564
rect 21453 15555 21511 15561
rect 21453 15552 21465 15555
rect 20680 15524 21465 15552
rect 20680 15512 20686 15524
rect 21453 15521 21465 15524
rect 21499 15521 21511 15555
rect 23566 15552 23572 15564
rect 23527 15524 23572 15552
rect 21453 15515 21511 15521
rect 23566 15512 23572 15524
rect 23624 15512 23630 15564
rect 24670 15552 24676 15564
rect 24583 15524 24676 15552
rect 24670 15512 24676 15524
rect 24728 15552 24734 15564
rect 25133 15555 25191 15561
rect 25133 15552 25145 15555
rect 24728 15524 25145 15552
rect 24728 15512 24734 15524
rect 25133 15521 25145 15524
rect 25179 15552 25191 15555
rect 25590 15552 25596 15564
rect 25179 15524 25596 15552
rect 25179 15521 25191 15524
rect 25133 15515 25191 15521
rect 25590 15512 25596 15524
rect 25648 15512 25654 15564
rect 26881 15555 26939 15561
rect 26881 15521 26893 15555
rect 26927 15552 26939 15555
rect 27430 15552 27436 15564
rect 26927 15524 27436 15552
rect 26927 15521 26939 15524
rect 26881 15515 26939 15521
rect 27430 15512 27436 15524
rect 27488 15512 27494 15564
rect 3694 15484 3700 15496
rect 2884 15456 3700 15484
rect 2884 15425 2912 15456
rect 3694 15444 3700 15456
rect 3752 15484 3758 15496
rect 4614 15484 4620 15496
rect 3752 15456 4620 15484
rect 3752 15444 3758 15456
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 5442 15444 5448 15496
rect 5500 15484 5506 15496
rect 5721 15487 5779 15493
rect 5721 15484 5733 15487
rect 5500 15456 5733 15484
rect 5500 15444 5506 15456
rect 5721 15453 5733 15456
rect 5767 15453 5779 15487
rect 5721 15447 5779 15453
rect 9766 15444 9772 15496
rect 9824 15484 9830 15496
rect 10137 15487 10195 15493
rect 10137 15484 10149 15487
rect 9824 15456 10149 15484
rect 9824 15444 9830 15456
rect 10137 15453 10149 15456
rect 10183 15453 10195 15487
rect 10318 15484 10324 15496
rect 10279 15456 10324 15484
rect 10137 15447 10195 15453
rect 10318 15444 10324 15456
rect 10376 15444 10382 15496
rect 11422 15444 11428 15496
rect 11480 15484 11486 15496
rect 11517 15487 11575 15493
rect 11517 15484 11529 15487
rect 11480 15456 11529 15484
rect 11480 15444 11486 15456
rect 11517 15453 11529 15456
rect 11563 15484 11575 15487
rect 11790 15484 11796 15496
rect 11563 15456 11796 15484
rect 11563 15453 11575 15456
rect 11517 15447 11575 15453
rect 11790 15444 11796 15456
rect 11848 15444 11854 15496
rect 15286 15484 15292 15496
rect 15247 15456 15292 15484
rect 15286 15444 15292 15456
rect 15344 15444 15350 15496
rect 18233 15487 18291 15493
rect 18233 15484 18245 15487
rect 18064 15456 18245 15484
rect 2869 15419 2927 15425
rect 2869 15385 2881 15419
rect 2915 15385 2927 15419
rect 2869 15379 2927 15385
rect 3513 15351 3571 15357
rect 3513 15317 3525 15351
rect 3559 15348 3571 15351
rect 3878 15348 3884 15360
rect 3559 15320 3884 15348
rect 3559 15317 3571 15320
rect 3513 15311 3571 15317
rect 3878 15308 3884 15320
rect 3936 15308 3942 15360
rect 5626 15348 5632 15360
rect 5587 15320 5632 15348
rect 5626 15308 5632 15320
rect 5684 15348 5690 15360
rect 7101 15351 7159 15357
rect 7101 15348 7113 15351
rect 5684 15320 7113 15348
rect 5684 15308 5690 15320
rect 7101 15317 7113 15320
rect 7147 15317 7159 15351
rect 10778 15348 10784 15360
rect 10739 15320 10784 15348
rect 7101 15311 7159 15317
rect 10778 15308 10784 15320
rect 10836 15308 10842 15360
rect 13817 15351 13875 15357
rect 13817 15317 13829 15351
rect 13863 15348 13875 15351
rect 14090 15348 14096 15360
rect 13863 15320 14096 15348
rect 13863 15317 13875 15320
rect 13817 15311 13875 15317
rect 14090 15308 14096 15320
rect 14148 15308 14154 15360
rect 16482 15308 16488 15360
rect 16540 15348 16546 15360
rect 16669 15351 16727 15357
rect 16669 15348 16681 15351
rect 16540 15320 16681 15348
rect 16540 15308 16546 15320
rect 16669 15317 16681 15320
rect 16715 15317 16727 15351
rect 16669 15311 16727 15317
rect 17862 15308 17868 15360
rect 17920 15348 17926 15360
rect 18064 15357 18092 15456
rect 18233 15453 18245 15456
rect 18279 15453 18291 15487
rect 18233 15447 18291 15453
rect 21545 15487 21603 15493
rect 21545 15453 21557 15487
rect 21591 15453 21603 15487
rect 21545 15447 21603 15453
rect 21729 15487 21787 15493
rect 21729 15453 21741 15487
rect 21775 15484 21787 15487
rect 21910 15484 21916 15496
rect 21775 15456 21916 15484
rect 21775 15453 21787 15456
rect 21729 15447 21787 15453
rect 18049 15351 18107 15357
rect 18049 15348 18061 15351
rect 17920 15320 18061 15348
rect 17920 15308 17926 15320
rect 18049 15317 18061 15320
rect 18095 15317 18107 15351
rect 18049 15311 18107 15317
rect 18230 15308 18236 15360
rect 18288 15348 18294 15360
rect 19613 15351 19671 15357
rect 19613 15348 19625 15351
rect 18288 15320 19625 15348
rect 18288 15308 18294 15320
rect 19613 15317 19625 15320
rect 19659 15317 19671 15351
rect 19613 15311 19671 15317
rect 20257 15351 20315 15357
rect 20257 15317 20269 15351
rect 20303 15348 20315 15351
rect 20530 15348 20536 15360
rect 20303 15320 20536 15348
rect 20303 15317 20315 15320
rect 20257 15311 20315 15317
rect 20530 15308 20536 15320
rect 20588 15308 20594 15360
rect 20714 15348 20720 15360
rect 20675 15320 20720 15348
rect 20714 15308 20720 15320
rect 20772 15348 20778 15360
rect 21560 15348 21588 15447
rect 21910 15444 21916 15456
rect 21968 15444 21974 15496
rect 23658 15484 23664 15496
rect 23619 15456 23664 15484
rect 23658 15444 23664 15456
rect 23716 15444 23722 15496
rect 23845 15487 23903 15493
rect 23845 15453 23857 15487
rect 23891 15453 23903 15487
rect 25222 15484 25228 15496
rect 25183 15456 25228 15484
rect 23845 15447 23903 15453
rect 23474 15376 23480 15428
rect 23532 15416 23538 15428
rect 23860 15416 23888 15447
rect 25222 15444 25228 15456
rect 25280 15444 25286 15496
rect 25409 15487 25467 15493
rect 25409 15453 25421 15487
rect 25455 15484 25467 15487
rect 25866 15484 25872 15496
rect 25455 15456 25872 15484
rect 25455 15453 25467 15456
rect 25409 15447 25467 15453
rect 25314 15416 25320 15428
rect 23532 15388 25320 15416
rect 23532 15376 23538 15388
rect 25314 15376 25320 15388
rect 25372 15416 25378 15428
rect 25424 15416 25452 15447
rect 25866 15444 25872 15456
rect 25924 15444 25930 15496
rect 26142 15484 26148 15496
rect 26055 15456 26148 15484
rect 25372 15388 25452 15416
rect 25372 15376 25378 15388
rect 24302 15348 24308 15360
rect 20772 15320 21588 15348
rect 24263 15320 24308 15348
rect 20772 15308 20778 15320
rect 24302 15308 24308 15320
rect 24360 15348 24366 15360
rect 26068 15348 26096 15456
rect 26142 15444 26148 15456
rect 26200 15444 26206 15496
rect 26602 15444 26608 15496
rect 26660 15484 26666 15496
rect 26973 15487 27031 15493
rect 26973 15484 26985 15487
rect 26660 15456 26985 15484
rect 26660 15444 26666 15456
rect 26973 15453 26985 15456
rect 27019 15453 27031 15487
rect 26973 15447 27031 15453
rect 27157 15487 27215 15493
rect 27157 15453 27169 15487
rect 27203 15484 27215 15487
rect 27522 15484 27528 15496
rect 27203 15456 27528 15484
rect 27203 15453 27215 15456
rect 27157 15447 27215 15453
rect 27522 15444 27528 15456
rect 27580 15444 27586 15496
rect 26510 15348 26516 15360
rect 24360 15320 26096 15348
rect 26471 15320 26516 15348
rect 24360 15308 24366 15320
rect 26510 15308 26516 15320
rect 26568 15308 26574 15360
rect 1104 15258 28888 15280
rect 1104 15206 5982 15258
rect 6034 15206 6046 15258
rect 6098 15206 6110 15258
rect 6162 15206 6174 15258
rect 6226 15206 15982 15258
rect 16034 15206 16046 15258
rect 16098 15206 16110 15258
rect 16162 15206 16174 15258
rect 16226 15206 25982 15258
rect 26034 15206 26046 15258
rect 26098 15206 26110 15258
rect 26162 15206 26174 15258
rect 26226 15206 28888 15258
rect 1104 15184 28888 15206
rect 1949 15147 2007 15153
rect 1949 15113 1961 15147
rect 1995 15144 2007 15147
rect 2038 15144 2044 15156
rect 1995 15116 2044 15144
rect 1995 15113 2007 15116
rect 1949 15107 2007 15113
rect 2038 15104 2044 15116
rect 2096 15104 2102 15156
rect 5442 15104 5448 15156
rect 5500 15144 5506 15156
rect 6181 15147 6239 15153
rect 6181 15144 6193 15147
rect 5500 15116 6193 15144
rect 5500 15104 5506 15116
rect 6181 15113 6193 15116
rect 6227 15113 6239 15147
rect 6181 15107 6239 15113
rect 7558 15104 7564 15156
rect 7616 15144 7622 15156
rect 7837 15147 7895 15153
rect 7837 15144 7849 15147
rect 7616 15116 7849 15144
rect 7616 15104 7622 15116
rect 7837 15113 7849 15116
rect 7883 15113 7895 15147
rect 7837 15107 7895 15113
rect 8941 15147 8999 15153
rect 8941 15113 8953 15147
rect 8987 15144 8999 15147
rect 9766 15144 9772 15156
rect 8987 15116 9772 15144
rect 8987 15113 8999 15116
rect 8941 15107 8999 15113
rect 9766 15104 9772 15116
rect 9824 15104 9830 15156
rect 11514 15144 11520 15156
rect 11475 15116 11520 15144
rect 11514 15104 11520 15116
rect 11572 15104 11578 15156
rect 12158 15144 12164 15156
rect 12119 15116 12164 15144
rect 12158 15104 12164 15116
rect 12216 15104 12222 15156
rect 14090 15104 14096 15156
rect 14148 15144 14154 15156
rect 16025 15147 16083 15153
rect 16025 15144 16037 15147
rect 14148 15116 16037 15144
rect 14148 15104 14154 15116
rect 16025 15113 16037 15116
rect 16071 15113 16083 15147
rect 16025 15107 16083 15113
rect 20073 15147 20131 15153
rect 20073 15113 20085 15147
rect 20119 15144 20131 15147
rect 20622 15144 20628 15156
rect 20119 15116 20628 15144
rect 20119 15113 20131 15116
rect 20073 15107 20131 15113
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 21637 15147 21695 15153
rect 21637 15113 21649 15147
rect 21683 15144 21695 15147
rect 22186 15144 22192 15156
rect 21683 15116 22192 15144
rect 21683 15113 21695 15116
rect 21637 15107 21695 15113
rect 22186 15104 22192 15116
rect 22244 15104 22250 15156
rect 3510 15076 3516 15088
rect 3471 15048 3516 15076
rect 3510 15036 3516 15048
rect 3568 15036 3574 15088
rect 7650 15076 7656 15088
rect 7611 15048 7656 15076
rect 7650 15036 7656 15048
rect 7708 15036 7714 15088
rect 8294 15036 8300 15088
rect 8352 15076 8358 15088
rect 9214 15076 9220 15088
rect 8352 15048 9220 15076
rect 8352 15036 8358 15048
rect 9214 15036 9220 15048
rect 9272 15076 9278 15088
rect 12897 15079 12955 15085
rect 9272 15048 9444 15076
rect 9272 15036 9278 15048
rect 2590 15008 2596 15020
rect 2551 14980 2596 15008
rect 2590 14968 2596 14980
rect 2648 15008 2654 15020
rect 3878 15008 3884 15020
rect 2648 14980 3884 15008
rect 2648 14968 2654 14980
rect 3878 14968 3884 14980
rect 3936 15008 3942 15020
rect 4065 15011 4123 15017
rect 4065 15008 4077 15011
rect 3936 14980 4077 15008
rect 3936 14968 3942 14980
rect 4065 14977 4077 14980
rect 4111 15008 4123 15011
rect 4525 15011 4583 15017
rect 4525 15008 4537 15011
rect 4111 14980 4537 15008
rect 4111 14977 4123 14980
rect 4065 14971 4123 14977
rect 4525 14977 4537 14980
rect 4571 14977 4583 15011
rect 4525 14971 4583 14977
rect 5813 15011 5871 15017
rect 5813 14977 5825 15011
rect 5859 15008 5871 15011
rect 6362 15008 6368 15020
rect 5859 14980 6368 15008
rect 5859 14977 5871 14980
rect 5813 14971 5871 14977
rect 6362 14968 6368 14980
rect 6420 14968 6426 15020
rect 7282 15008 7288 15020
rect 7243 14980 7288 15008
rect 7282 14968 7288 14980
rect 7340 14968 7346 15020
rect 1857 14943 1915 14949
rect 1857 14909 1869 14943
rect 1903 14940 1915 14943
rect 1946 14940 1952 14952
rect 1903 14912 1952 14940
rect 1903 14909 1915 14912
rect 1857 14903 1915 14909
rect 1946 14900 1952 14912
rect 2004 14900 2010 14952
rect 2317 14943 2375 14949
rect 2317 14909 2329 14943
rect 2363 14940 2375 14943
rect 2682 14940 2688 14952
rect 2363 14912 2688 14940
rect 2363 14909 2375 14912
rect 2317 14903 2375 14909
rect 2682 14900 2688 14912
rect 2740 14900 2746 14952
rect 4246 14900 4252 14952
rect 4304 14940 4310 14952
rect 5077 14943 5135 14949
rect 5077 14940 5089 14943
rect 4304 14912 5089 14940
rect 4304 14900 4310 14912
rect 5077 14909 5089 14912
rect 5123 14940 5135 14943
rect 5123 14912 5488 14940
rect 5123 14909 5135 14912
rect 5077 14903 5135 14909
rect 1964 14872 1992 14900
rect 2409 14875 2467 14881
rect 2409 14872 2421 14875
rect 1964 14844 2421 14872
rect 2409 14841 2421 14844
rect 2455 14841 2467 14875
rect 2409 14835 2467 14841
rect 5460 14816 5488 14912
rect 7190 14900 7196 14952
rect 7248 14940 7254 14952
rect 7668 14940 7696 15036
rect 8386 15008 8392 15020
rect 8347 14980 8392 15008
rect 8386 14968 8392 14980
rect 8444 14968 8450 15020
rect 9416 15017 9444 15048
rect 12897 15045 12909 15079
rect 12943 15076 12955 15079
rect 13909 15079 13967 15085
rect 13909 15076 13921 15079
rect 12943 15048 13921 15076
rect 12943 15045 12955 15048
rect 12897 15039 12955 15045
rect 13909 15045 13921 15048
rect 13955 15076 13967 15079
rect 13955 15048 14964 15076
rect 13955 15045 13967 15048
rect 13909 15039 13967 15045
rect 9401 15011 9459 15017
rect 9401 14977 9413 15011
rect 9447 14977 9459 15011
rect 9401 14971 9459 14977
rect 11790 14968 11796 15020
rect 11848 15008 11854 15020
rect 11885 15011 11943 15017
rect 11885 15008 11897 15011
rect 11848 14980 11897 15008
rect 11848 14968 11854 14980
rect 11885 14977 11897 14980
rect 11931 15008 11943 15011
rect 13078 15008 13084 15020
rect 11931 14980 13084 15008
rect 11931 14977 11943 14980
rect 11885 14971 11943 14977
rect 13078 14968 13084 14980
rect 13136 14968 13142 15020
rect 13538 15008 13544 15020
rect 13499 14980 13544 15008
rect 13538 14968 13544 14980
rect 13596 14968 13602 15020
rect 14274 15008 14280 15020
rect 14235 14980 14280 15008
rect 14274 14968 14280 14980
rect 14332 15008 14338 15020
rect 14936 15017 14964 15048
rect 15562 15036 15568 15088
rect 15620 15076 15626 15088
rect 15838 15076 15844 15088
rect 15620 15048 15844 15076
rect 15620 15036 15626 15048
rect 15838 15036 15844 15048
rect 15896 15036 15902 15088
rect 17586 15036 17592 15088
rect 17644 15076 17650 15088
rect 17644 15048 24256 15076
rect 17644 15036 17650 15048
rect 14921 15011 14979 15017
rect 14332 14980 14872 15008
rect 14332 14968 14338 14980
rect 14844 14952 14872 14980
rect 14921 14977 14933 15011
rect 14967 14977 14979 15011
rect 15102 15008 15108 15020
rect 15063 14980 15108 15008
rect 14921 14971 14979 14977
rect 15102 14968 15108 14980
rect 15160 15008 15166 15020
rect 16482 15008 16488 15020
rect 15160 14980 16488 15008
rect 15160 14968 15166 14980
rect 16482 14968 16488 14980
rect 16540 15008 16546 15020
rect 16577 15011 16635 15017
rect 16577 15008 16589 15011
rect 16540 14980 16589 15008
rect 16540 14968 16546 14980
rect 16577 14977 16589 14980
rect 16623 14977 16635 15011
rect 19150 15008 19156 15020
rect 19111 14980 19156 15008
rect 16577 14971 16635 14977
rect 19150 14968 19156 14980
rect 19208 14968 19214 15020
rect 19613 15011 19671 15017
rect 19613 14977 19625 15011
rect 19659 15008 19671 15011
rect 20717 15011 20775 15017
rect 20717 15008 20729 15011
rect 19659 14980 20729 15008
rect 19659 14977 19671 14980
rect 19613 14971 19671 14977
rect 20717 14977 20729 14980
rect 20763 15008 20775 15011
rect 21634 15008 21640 15020
rect 20763 14980 21640 15008
rect 20763 14977 20775 14980
rect 20717 14971 20775 14977
rect 21634 14968 21640 14980
rect 21692 15008 21698 15020
rect 22189 15011 22247 15017
rect 22189 15008 22201 15011
rect 21692 14980 22201 15008
rect 21692 14968 21698 14980
rect 22189 14977 22201 14980
rect 22235 15008 22247 15011
rect 22830 15008 22836 15020
rect 22235 14980 22836 15008
rect 22235 14977 22247 14980
rect 22189 14971 22247 14977
rect 22830 14968 22836 14980
rect 22888 14968 22894 15020
rect 23198 15008 23204 15020
rect 23159 14980 23204 15008
rect 23198 14968 23204 14980
rect 23256 14968 23262 15020
rect 8205 14943 8263 14949
rect 8205 14940 8217 14943
rect 7248 14912 8217 14940
rect 7248 14900 7254 14912
rect 8205 14909 8217 14912
rect 8251 14909 8263 14943
rect 13262 14940 13268 14952
rect 13223 14912 13268 14940
rect 8205 14903 8263 14909
rect 13262 14900 13268 14912
rect 13320 14900 13326 14952
rect 14826 14940 14832 14952
rect 14739 14912 14832 14940
rect 14826 14900 14832 14912
rect 14884 14900 14890 14952
rect 15286 14900 15292 14952
rect 15344 14940 15350 14952
rect 15565 14943 15623 14949
rect 15565 14940 15577 14943
rect 15344 14912 15577 14940
rect 15344 14900 15350 14912
rect 15565 14909 15577 14912
rect 15611 14940 15623 14943
rect 17862 14940 17868 14952
rect 15611 14912 17868 14940
rect 15611 14909 15623 14912
rect 15565 14903 15623 14909
rect 17862 14900 17868 14912
rect 17920 14900 17926 14952
rect 21177 14943 21235 14949
rect 21177 14909 21189 14943
rect 21223 14940 21235 14943
rect 22002 14940 22008 14952
rect 21223 14912 22008 14940
rect 21223 14909 21235 14912
rect 21177 14903 21235 14909
rect 22002 14900 22008 14912
rect 22060 14900 22066 14952
rect 5537 14875 5595 14881
rect 5537 14841 5549 14875
rect 5583 14872 5595 14875
rect 5902 14872 5908 14884
rect 5583 14844 5908 14872
rect 5583 14841 5595 14844
rect 5537 14835 5595 14841
rect 5902 14832 5908 14844
rect 5960 14872 5966 14884
rect 5960 14844 7880 14872
rect 5960 14832 5966 14844
rect 7852 14816 7880 14844
rect 9490 14832 9496 14884
rect 9548 14872 9554 14884
rect 9646 14875 9704 14881
rect 9646 14872 9658 14875
rect 9548 14844 9658 14872
rect 9548 14832 9554 14844
rect 9646 14841 9658 14844
rect 9692 14841 9704 14875
rect 13357 14875 13415 14881
rect 13357 14872 13369 14875
rect 9646 14835 9704 14841
rect 12912 14844 13369 14872
rect 12912 14816 12940 14844
rect 13357 14841 13369 14844
rect 13403 14841 13415 14875
rect 13357 14835 13415 14841
rect 13998 14832 14004 14884
rect 14056 14872 14062 14884
rect 16393 14875 16451 14881
rect 14056 14844 14504 14872
rect 14056 14832 14062 14844
rect 2958 14804 2964 14816
rect 2919 14776 2964 14804
rect 2958 14764 2964 14776
rect 3016 14764 3022 14816
rect 3421 14807 3479 14813
rect 3421 14773 3433 14807
rect 3467 14804 3479 14807
rect 3786 14804 3792 14816
rect 3467 14776 3792 14804
rect 3467 14773 3479 14776
rect 3421 14767 3479 14773
rect 3786 14764 3792 14776
rect 3844 14804 3850 14816
rect 3881 14807 3939 14813
rect 3881 14804 3893 14807
rect 3844 14776 3893 14804
rect 3844 14764 3850 14776
rect 3881 14773 3893 14776
rect 3927 14773 3939 14807
rect 3881 14767 3939 14773
rect 3970 14764 3976 14816
rect 4028 14804 4034 14816
rect 4798 14804 4804 14816
rect 4028 14776 4804 14804
rect 4028 14764 4034 14776
rect 4798 14764 4804 14776
rect 4856 14764 4862 14816
rect 5166 14804 5172 14816
rect 5127 14776 5172 14804
rect 5166 14764 5172 14776
rect 5224 14764 5230 14816
rect 5442 14764 5448 14816
rect 5500 14804 5506 14816
rect 5629 14807 5687 14813
rect 5629 14804 5641 14807
rect 5500 14776 5641 14804
rect 5500 14764 5506 14776
rect 5629 14773 5641 14776
rect 5675 14773 5687 14807
rect 5629 14767 5687 14773
rect 6362 14764 6368 14816
rect 6420 14804 6426 14816
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 6420 14776 6561 14804
rect 6420 14764 6426 14776
rect 6549 14773 6561 14776
rect 6595 14773 6607 14807
rect 6549 14767 6607 14773
rect 6638 14764 6644 14816
rect 6696 14804 6702 14816
rect 6825 14807 6883 14813
rect 6825 14804 6837 14807
rect 6696 14776 6837 14804
rect 6696 14764 6702 14776
rect 6825 14773 6837 14776
rect 6871 14773 6883 14807
rect 6825 14767 6883 14773
rect 7834 14764 7840 14816
rect 7892 14804 7898 14816
rect 8297 14807 8355 14813
rect 8297 14804 8309 14807
rect 7892 14776 8309 14804
rect 7892 14764 7898 14776
rect 8297 14773 8309 14776
rect 8343 14773 8355 14807
rect 8297 14767 8355 14773
rect 10781 14807 10839 14813
rect 10781 14773 10793 14807
rect 10827 14804 10839 14807
rect 11330 14804 11336 14816
rect 10827 14776 11336 14804
rect 10827 14773 10839 14776
rect 10781 14767 10839 14773
rect 11330 14764 11336 14776
rect 11388 14764 11394 14816
rect 12805 14807 12863 14813
rect 12805 14773 12817 14807
rect 12851 14804 12863 14807
rect 12894 14804 12900 14816
rect 12851 14776 12900 14804
rect 12851 14773 12863 14776
rect 12805 14767 12863 14773
rect 12894 14764 12900 14776
rect 12952 14764 12958 14816
rect 14476 14813 14504 14844
rect 16393 14841 16405 14875
rect 16439 14872 16451 14875
rect 16666 14872 16672 14884
rect 16439 14844 16672 14872
rect 16439 14841 16451 14844
rect 16393 14835 16451 14841
rect 16666 14832 16672 14844
rect 16724 14832 16730 14884
rect 18417 14875 18475 14881
rect 18417 14841 18429 14875
rect 18463 14872 18475 14875
rect 18598 14872 18604 14884
rect 18463 14844 18604 14872
rect 18463 14841 18475 14844
rect 18417 14835 18475 14841
rect 18598 14832 18604 14844
rect 18656 14872 18662 14884
rect 18877 14875 18935 14881
rect 18877 14872 18889 14875
rect 18656 14844 18889 14872
rect 18656 14832 18662 14844
rect 18877 14841 18889 14844
rect 18923 14841 18935 14875
rect 23566 14872 23572 14884
rect 18877 14835 18935 14841
rect 22940 14844 23572 14872
rect 22940 14816 22968 14844
rect 23566 14832 23572 14844
rect 23624 14832 23630 14884
rect 14461 14807 14519 14813
rect 14461 14773 14473 14807
rect 14507 14773 14519 14807
rect 14461 14767 14519 14773
rect 16482 14764 16488 14816
rect 16540 14804 16546 14816
rect 17037 14807 17095 14813
rect 17037 14804 17049 14807
rect 16540 14776 17049 14804
rect 16540 14764 16546 14776
rect 17037 14773 17049 14776
rect 17083 14773 17095 14807
rect 17402 14804 17408 14816
rect 17363 14776 17408 14804
rect 17037 14767 17095 14773
rect 17402 14764 17408 14776
rect 17460 14764 17466 14816
rect 17862 14804 17868 14816
rect 17823 14776 17868 14804
rect 17862 14764 17868 14776
rect 17920 14764 17926 14816
rect 18506 14804 18512 14816
rect 18467 14776 18512 14804
rect 18506 14764 18512 14776
rect 18564 14764 18570 14816
rect 18966 14804 18972 14816
rect 18927 14776 18972 14804
rect 18966 14764 18972 14776
rect 19024 14764 19030 14816
rect 19886 14804 19892 14816
rect 19847 14776 19892 14804
rect 19886 14764 19892 14776
rect 19944 14804 19950 14816
rect 20438 14804 20444 14816
rect 19944 14776 20444 14804
rect 19944 14764 19950 14776
rect 20438 14764 20444 14776
rect 20496 14764 20502 14816
rect 20530 14764 20536 14816
rect 20588 14804 20594 14816
rect 20588 14776 20633 14804
rect 20588 14764 20594 14776
rect 21266 14764 21272 14816
rect 21324 14804 21330 14816
rect 21453 14807 21511 14813
rect 21453 14804 21465 14807
rect 21324 14776 21465 14804
rect 21324 14764 21330 14776
rect 21453 14773 21465 14776
rect 21499 14804 21511 14807
rect 21726 14804 21732 14816
rect 21499 14776 21732 14804
rect 21499 14773 21511 14776
rect 21453 14767 21511 14773
rect 21726 14764 21732 14776
rect 21784 14804 21790 14816
rect 22097 14807 22155 14813
rect 22097 14804 22109 14807
rect 21784 14776 22109 14804
rect 21784 14764 21790 14776
rect 22097 14773 22109 14776
rect 22143 14773 22155 14807
rect 22922 14804 22928 14816
rect 22883 14776 22928 14804
rect 22097 14767 22155 14773
rect 22922 14764 22928 14776
rect 22980 14764 22986 14816
rect 24228 14813 24256 15048
rect 27338 15008 27344 15020
rect 27299 14980 27344 15008
rect 27338 14968 27344 14980
rect 27396 14968 27402 15020
rect 24302 14900 24308 14952
rect 24360 14940 24366 14952
rect 24360 14912 24405 14940
rect 24360 14900 24366 14912
rect 26510 14900 26516 14952
rect 26568 14940 26574 14952
rect 27249 14943 27307 14949
rect 27249 14940 27261 14943
rect 26568 14912 27261 14940
rect 26568 14900 26574 14912
rect 27249 14909 27261 14912
rect 27295 14909 27307 14943
rect 27249 14903 27307 14909
rect 24394 14832 24400 14884
rect 24452 14872 24458 14884
rect 24550 14875 24608 14881
rect 24550 14872 24562 14875
rect 24452 14844 24562 14872
rect 24452 14832 24458 14844
rect 24550 14841 24562 14844
rect 24596 14841 24608 14875
rect 24550 14835 24608 14841
rect 27614 14832 27620 14884
rect 27672 14872 27678 14884
rect 28169 14875 28227 14881
rect 28169 14872 28181 14875
rect 27672 14844 28181 14872
rect 27672 14832 27678 14844
rect 28169 14841 28181 14844
rect 28215 14841 28227 14875
rect 28169 14835 28227 14841
rect 24213 14807 24271 14813
rect 24213 14773 24225 14807
rect 24259 14804 24271 14807
rect 25130 14804 25136 14816
rect 24259 14776 25136 14804
rect 24259 14773 24271 14776
rect 24213 14767 24271 14773
rect 25130 14764 25136 14776
rect 25188 14764 25194 14816
rect 25682 14804 25688 14816
rect 25643 14776 25688 14804
rect 25682 14764 25688 14776
rect 25740 14764 25746 14816
rect 26602 14804 26608 14816
rect 26563 14776 26608 14804
rect 26602 14764 26608 14776
rect 26660 14764 26666 14816
rect 26786 14804 26792 14816
rect 26747 14776 26792 14804
rect 26786 14764 26792 14776
rect 26844 14764 26850 14816
rect 27157 14807 27215 14813
rect 27157 14773 27169 14807
rect 27203 14804 27215 14807
rect 27338 14804 27344 14816
rect 27203 14776 27344 14804
rect 27203 14773 27215 14776
rect 27157 14767 27215 14773
rect 27338 14764 27344 14776
rect 27396 14804 27402 14816
rect 27801 14807 27859 14813
rect 27801 14804 27813 14807
rect 27396 14776 27813 14804
rect 27396 14764 27402 14776
rect 27801 14773 27813 14776
rect 27847 14773 27859 14807
rect 27801 14767 27859 14773
rect 1104 14714 28888 14736
rect 1104 14662 10982 14714
rect 11034 14662 11046 14714
rect 11098 14662 11110 14714
rect 11162 14662 11174 14714
rect 11226 14662 20982 14714
rect 21034 14662 21046 14714
rect 21098 14662 21110 14714
rect 21162 14662 21174 14714
rect 21226 14662 28888 14714
rect 1104 14640 28888 14662
rect 1949 14603 2007 14609
rect 1949 14569 1961 14603
rect 1995 14600 2007 14603
rect 2130 14600 2136 14612
rect 1995 14572 2136 14600
rect 1995 14569 2007 14572
rect 1949 14563 2007 14569
rect 2130 14560 2136 14572
rect 2188 14560 2194 14612
rect 2774 14600 2780 14612
rect 2332 14572 2780 14600
rect 2038 14424 2044 14476
rect 2096 14464 2102 14476
rect 2332 14473 2360 14572
rect 2774 14560 2780 14572
rect 2832 14560 2838 14612
rect 2958 14600 2964 14612
rect 2919 14572 2964 14600
rect 2958 14560 2964 14572
rect 3016 14560 3022 14612
rect 3605 14603 3663 14609
rect 3605 14569 3617 14603
rect 3651 14600 3663 14603
rect 3970 14600 3976 14612
rect 3651 14572 3976 14600
rect 3651 14569 3663 14572
rect 3605 14563 3663 14569
rect 3970 14560 3976 14572
rect 4028 14560 4034 14612
rect 4614 14600 4620 14612
rect 4575 14572 4620 14600
rect 4614 14560 4620 14572
rect 4672 14560 4678 14612
rect 4798 14560 4804 14612
rect 4856 14600 4862 14612
rect 5261 14603 5319 14609
rect 5261 14600 5273 14603
rect 4856 14572 5273 14600
rect 4856 14560 4862 14572
rect 5261 14569 5273 14572
rect 5307 14600 5319 14603
rect 5902 14600 5908 14612
rect 5307 14572 5908 14600
rect 5307 14569 5319 14572
rect 5261 14563 5319 14569
rect 5902 14560 5908 14572
rect 5960 14560 5966 14612
rect 7558 14560 7564 14612
rect 7616 14600 7622 14612
rect 8389 14603 8447 14609
rect 8389 14600 8401 14603
rect 7616 14572 8401 14600
rect 7616 14560 7622 14572
rect 8389 14569 8401 14572
rect 8435 14569 8447 14603
rect 8389 14563 8447 14569
rect 8478 14560 8484 14612
rect 8536 14600 8542 14612
rect 8536 14572 8581 14600
rect 8536 14560 8542 14572
rect 12158 14560 12164 14612
rect 12216 14600 12222 14612
rect 12437 14603 12495 14609
rect 12437 14600 12449 14603
rect 12216 14572 12449 14600
rect 12216 14560 12222 14572
rect 12437 14569 12449 14572
rect 12483 14569 12495 14603
rect 12437 14563 12495 14569
rect 13081 14603 13139 14609
rect 13081 14569 13093 14603
rect 13127 14600 13139 14603
rect 13262 14600 13268 14612
rect 13127 14572 13268 14600
rect 13127 14569 13139 14572
rect 13081 14563 13139 14569
rect 13262 14560 13268 14572
rect 13320 14560 13326 14612
rect 13633 14603 13691 14609
rect 13633 14569 13645 14603
rect 13679 14600 13691 14603
rect 13722 14600 13728 14612
rect 13679 14572 13728 14600
rect 13679 14569 13691 14572
rect 13633 14563 13691 14569
rect 13722 14560 13728 14572
rect 13780 14560 13786 14612
rect 14090 14600 14096 14612
rect 14051 14572 14096 14600
rect 14090 14560 14096 14572
rect 14148 14560 14154 14612
rect 15289 14603 15347 14609
rect 15289 14569 15301 14603
rect 15335 14600 15347 14603
rect 16482 14600 16488 14612
rect 15335 14572 16488 14600
rect 15335 14569 15347 14572
rect 15289 14563 15347 14569
rect 16482 14560 16488 14572
rect 16540 14560 16546 14612
rect 17126 14600 17132 14612
rect 17087 14572 17132 14600
rect 17126 14560 17132 14572
rect 17184 14560 17190 14612
rect 18230 14600 18236 14612
rect 18191 14572 18236 14600
rect 18230 14560 18236 14572
rect 18288 14560 18294 14612
rect 18506 14560 18512 14612
rect 18564 14600 18570 14612
rect 19613 14603 19671 14609
rect 19613 14600 19625 14603
rect 18564 14572 19625 14600
rect 18564 14560 18570 14572
rect 19613 14569 19625 14572
rect 19659 14600 19671 14603
rect 20254 14600 20260 14612
rect 19659 14572 20260 14600
rect 19659 14569 19671 14572
rect 19613 14563 19671 14569
rect 20254 14560 20260 14572
rect 20312 14560 20318 14612
rect 20349 14603 20407 14609
rect 20349 14569 20361 14603
rect 20395 14600 20407 14603
rect 20622 14600 20628 14612
rect 20395 14572 20628 14600
rect 20395 14569 20407 14572
rect 20349 14563 20407 14569
rect 20622 14560 20628 14572
rect 20680 14560 20686 14612
rect 20717 14603 20775 14609
rect 20717 14569 20729 14603
rect 20763 14600 20775 14603
rect 21910 14600 21916 14612
rect 20763 14572 21916 14600
rect 20763 14569 20775 14572
rect 20717 14563 20775 14569
rect 21910 14560 21916 14572
rect 21968 14560 21974 14612
rect 22830 14600 22836 14612
rect 22791 14572 22836 14600
rect 22830 14560 22836 14572
rect 22888 14560 22894 14612
rect 23474 14600 23480 14612
rect 23435 14572 23480 14600
rect 23474 14560 23480 14572
rect 23532 14560 23538 14612
rect 23750 14600 23756 14612
rect 23711 14572 23756 14600
rect 23750 14560 23756 14572
rect 23808 14560 23814 14612
rect 25961 14603 26019 14609
rect 25961 14569 25973 14603
rect 26007 14600 26019 14603
rect 26510 14600 26516 14612
rect 26007 14572 26516 14600
rect 26007 14569 26019 14572
rect 25961 14563 26019 14569
rect 26510 14560 26516 14572
rect 26568 14560 26574 14612
rect 27246 14560 27252 14612
rect 27304 14600 27310 14612
rect 27525 14603 27583 14609
rect 27525 14600 27537 14603
rect 27304 14572 27537 14600
rect 27304 14560 27310 14572
rect 27525 14569 27537 14572
rect 27571 14569 27583 14603
rect 27525 14563 27583 14569
rect 5626 14492 5632 14544
rect 5684 14541 5690 14544
rect 5684 14535 5748 14541
rect 5684 14501 5702 14535
rect 5736 14501 5748 14535
rect 16390 14532 16396 14544
rect 16351 14504 16396 14532
rect 5684 14495 5748 14501
rect 5684 14492 5690 14495
rect 16390 14492 16396 14504
rect 16448 14492 16454 14544
rect 18969 14535 19027 14541
rect 18969 14501 18981 14535
rect 19015 14532 19027 14535
rect 19150 14532 19156 14544
rect 19015 14504 19156 14532
rect 19015 14501 19027 14504
rect 18969 14495 19027 14501
rect 19150 14492 19156 14504
rect 19208 14492 19214 14544
rect 26329 14535 26387 14541
rect 26329 14501 26341 14535
rect 26375 14532 26387 14535
rect 26418 14532 26424 14544
rect 26375 14504 26424 14532
rect 26375 14501 26387 14504
rect 26329 14495 26387 14501
rect 26418 14492 26424 14504
rect 26476 14492 26482 14544
rect 2317 14467 2375 14473
rect 2317 14464 2329 14467
rect 2096 14436 2329 14464
rect 2096 14424 2102 14436
rect 2317 14433 2329 14436
rect 2363 14433 2375 14467
rect 4065 14467 4123 14473
rect 4065 14464 4077 14467
rect 2317 14427 2375 14433
rect 2424 14436 4077 14464
rect 2424 14408 2452 14436
rect 4065 14433 4077 14436
rect 4111 14464 4123 14467
rect 4706 14464 4712 14476
rect 4111 14436 4712 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 4706 14424 4712 14436
rect 4764 14424 4770 14476
rect 5445 14467 5503 14473
rect 5445 14433 5457 14467
rect 5491 14464 5503 14467
rect 5534 14464 5540 14476
rect 5491 14436 5540 14464
rect 5491 14433 5503 14436
rect 5445 14427 5503 14433
rect 5534 14424 5540 14436
rect 5592 14424 5598 14476
rect 9214 14424 9220 14476
rect 9272 14464 9278 14476
rect 9953 14467 10011 14473
rect 9272 14436 9536 14464
rect 9272 14424 9278 14436
rect 2406 14396 2412 14408
rect 2367 14368 2412 14396
rect 2406 14356 2412 14368
rect 2464 14356 2470 14408
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14396 2651 14399
rect 3878 14396 3884 14408
rect 2639 14368 3884 14396
rect 2639 14365 2651 14368
rect 2593 14359 2651 14365
rect 3878 14356 3884 14368
rect 3936 14356 3942 14408
rect 8294 14356 8300 14408
rect 8352 14396 8358 14408
rect 8665 14399 8723 14405
rect 8665 14396 8677 14399
rect 8352 14368 8677 14396
rect 8352 14356 8358 14368
rect 8665 14365 8677 14368
rect 8711 14396 8723 14399
rect 9398 14396 9404 14408
rect 8711 14368 9404 14396
rect 8711 14365 8723 14368
rect 8665 14359 8723 14365
rect 9398 14356 9404 14368
rect 9456 14356 9462 14408
rect 9508 14396 9536 14436
rect 9953 14433 9965 14467
rect 9999 14464 10011 14467
rect 10318 14464 10324 14476
rect 9999 14436 10324 14464
rect 9999 14433 10011 14436
rect 9953 14427 10011 14433
rect 10318 14424 10324 14436
rect 10376 14464 10382 14476
rect 11330 14473 11336 14476
rect 11324 14464 11336 14473
rect 10376 14436 11336 14464
rect 10376 14424 10382 14436
rect 11324 14427 11336 14436
rect 11330 14424 11336 14427
rect 11388 14424 11394 14476
rect 13998 14464 14004 14476
rect 13959 14436 14004 14464
rect 13998 14424 14004 14436
rect 14056 14424 14062 14476
rect 15654 14464 15660 14476
rect 15615 14436 15660 14464
rect 15654 14424 15660 14436
rect 15712 14424 15718 14476
rect 15749 14467 15807 14473
rect 15749 14433 15761 14467
rect 15795 14464 15807 14467
rect 16298 14464 16304 14476
rect 15795 14436 16304 14464
rect 15795 14433 15807 14436
rect 15749 14427 15807 14433
rect 16298 14424 16304 14436
rect 16356 14424 16362 14476
rect 16482 14424 16488 14476
rect 16540 14464 16546 14476
rect 17497 14467 17555 14473
rect 17497 14464 17509 14467
rect 16540 14436 17509 14464
rect 16540 14424 16546 14436
rect 17497 14433 17509 14436
rect 17543 14433 17555 14467
rect 17497 14427 17555 14433
rect 19334 14424 19340 14476
rect 19392 14464 19398 14476
rect 19702 14464 19708 14476
rect 19392 14436 19708 14464
rect 19392 14424 19398 14436
rect 19702 14424 19708 14436
rect 19760 14424 19766 14476
rect 21720 14467 21778 14473
rect 21720 14433 21732 14467
rect 21766 14464 21778 14467
rect 22186 14464 22192 14476
rect 21766 14436 22192 14464
rect 21766 14433 21778 14436
rect 21720 14427 21778 14433
rect 22186 14424 22192 14436
rect 22244 14424 22250 14476
rect 23474 14424 23480 14476
rect 23532 14464 23538 14476
rect 24193 14467 24251 14473
rect 24193 14464 24205 14467
rect 23532 14436 24205 14464
rect 23532 14424 23538 14436
rect 24193 14433 24205 14436
rect 24239 14433 24251 14467
rect 26878 14464 26884 14476
rect 26839 14436 26884 14464
rect 24193 14427 24251 14433
rect 26878 14424 26884 14436
rect 26936 14424 26942 14476
rect 11057 14399 11115 14405
rect 11057 14396 11069 14399
rect 9508 14368 11069 14396
rect 11057 14365 11069 14368
rect 11103 14365 11115 14399
rect 11057 14359 11115 14365
rect 1670 14328 1676 14340
rect 1583 14300 1676 14328
rect 1670 14288 1676 14300
rect 1728 14328 1734 14340
rect 2682 14328 2688 14340
rect 1728 14300 2688 14328
rect 1728 14288 1734 14300
rect 2682 14288 2688 14300
rect 2740 14288 2746 14340
rect 6730 14288 6736 14340
rect 6788 14328 6794 14340
rect 7377 14331 7435 14337
rect 7377 14328 7389 14331
rect 6788 14300 7389 14328
rect 6788 14288 6794 14300
rect 7377 14297 7389 14300
rect 7423 14297 7435 14331
rect 7377 14291 7435 14297
rect 7466 14288 7472 14340
rect 7524 14328 7530 14340
rect 8021 14331 8079 14337
rect 8021 14328 8033 14331
rect 7524 14300 8033 14328
rect 7524 14288 7530 14300
rect 8021 14297 8033 14300
rect 8067 14297 8079 14331
rect 8021 14291 8079 14297
rect 1486 14220 1492 14272
rect 1544 14260 1550 14272
rect 2590 14260 2596 14272
rect 1544 14232 2596 14260
rect 1544 14220 1550 14232
rect 2590 14220 2596 14232
rect 2648 14260 2654 14272
rect 2958 14260 2964 14272
rect 2648 14232 2964 14260
rect 2648 14220 2654 14232
rect 2958 14220 2964 14232
rect 3016 14220 3022 14272
rect 4246 14260 4252 14272
rect 4207 14232 4252 14260
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 6822 14260 6828 14272
rect 6783 14232 6828 14260
rect 6822 14220 6828 14232
rect 6880 14220 6886 14272
rect 7834 14260 7840 14272
rect 7795 14232 7840 14260
rect 7834 14220 7840 14232
rect 7892 14220 7898 14272
rect 9122 14260 9128 14272
rect 9083 14232 9128 14260
rect 9122 14220 9128 14232
rect 9180 14220 9186 14272
rect 9490 14260 9496 14272
rect 9451 14232 9496 14260
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 10318 14260 10324 14272
rect 10279 14232 10324 14260
rect 10318 14220 10324 14232
rect 10376 14220 10382 14272
rect 10870 14260 10876 14272
rect 10831 14232 10876 14260
rect 10870 14220 10876 14232
rect 10928 14220 10934 14272
rect 11072 14260 11100 14359
rect 13814 14356 13820 14408
rect 13872 14396 13878 14408
rect 14185 14399 14243 14405
rect 14185 14396 14197 14399
rect 13872 14368 14197 14396
rect 13872 14356 13878 14368
rect 14185 14365 14197 14368
rect 14231 14365 14243 14399
rect 15838 14396 15844 14408
rect 15799 14368 15844 14396
rect 14185 14359 14243 14365
rect 15838 14356 15844 14368
rect 15896 14356 15902 14408
rect 16758 14356 16764 14408
rect 16816 14396 16822 14408
rect 17589 14399 17647 14405
rect 17589 14396 17601 14399
rect 16816 14368 17601 14396
rect 16816 14356 16822 14368
rect 17589 14365 17601 14368
rect 17635 14365 17647 14399
rect 17770 14396 17776 14408
rect 17731 14368 17776 14396
rect 17589 14359 17647 14365
rect 17770 14356 17776 14368
rect 17828 14356 17834 14408
rect 19889 14399 19947 14405
rect 19889 14365 19901 14399
rect 19935 14396 19947 14399
rect 20070 14396 20076 14408
rect 19935 14368 20076 14396
rect 19935 14365 19947 14368
rect 19889 14359 19947 14365
rect 20070 14356 20076 14368
rect 20128 14356 20134 14408
rect 20806 14356 20812 14408
rect 20864 14396 20870 14408
rect 21453 14399 21511 14405
rect 21453 14396 21465 14399
rect 20864 14368 21465 14396
rect 20864 14356 20870 14368
rect 13449 14331 13507 14337
rect 13449 14297 13461 14331
rect 13495 14328 13507 14331
rect 13538 14328 13544 14340
rect 13495 14300 13544 14328
rect 13495 14297 13507 14300
rect 13449 14291 13507 14297
rect 13538 14288 13544 14300
rect 13596 14328 13602 14340
rect 15013 14331 15071 14337
rect 15013 14328 15025 14331
rect 13596 14300 15025 14328
rect 13596 14288 13602 14300
rect 15013 14297 15025 14300
rect 15059 14328 15071 14331
rect 15856 14328 15884 14356
rect 15059 14300 15884 14328
rect 15059 14297 15071 14300
rect 15013 14291 15071 14297
rect 21100 14272 21128 14368
rect 21453 14365 21465 14368
rect 21499 14365 21511 14399
rect 21453 14359 21511 14365
rect 23842 14356 23848 14408
rect 23900 14396 23906 14408
rect 23937 14399 23995 14405
rect 23937 14396 23949 14399
rect 23900 14368 23949 14396
rect 23900 14356 23906 14368
rect 23937 14365 23949 14368
rect 23983 14365 23995 14399
rect 26970 14396 26976 14408
rect 26931 14368 26976 14396
rect 23937 14359 23995 14365
rect 11422 14260 11428 14272
rect 11072 14232 11428 14260
rect 11422 14220 11428 14232
rect 11480 14220 11486 14272
rect 16666 14260 16672 14272
rect 16627 14232 16672 14260
rect 16666 14220 16672 14232
rect 16724 14220 16730 14272
rect 18506 14260 18512 14272
rect 18467 14232 18512 14260
rect 18506 14220 18512 14232
rect 18564 14260 18570 14272
rect 18966 14260 18972 14272
rect 18564 14232 18972 14260
rect 18564 14220 18570 14232
rect 18966 14220 18972 14232
rect 19024 14220 19030 14272
rect 19242 14260 19248 14272
rect 19203 14232 19248 14260
rect 19242 14220 19248 14232
rect 19300 14220 19306 14272
rect 21082 14260 21088 14272
rect 21043 14232 21088 14260
rect 21082 14220 21088 14232
rect 21140 14220 21146 14272
rect 23952 14260 23980 14359
rect 26970 14356 26976 14368
rect 27028 14356 27034 14408
rect 27065 14399 27123 14405
rect 27065 14365 27077 14399
rect 27111 14365 27123 14399
rect 27065 14359 27123 14365
rect 27080 14328 27108 14359
rect 27706 14328 27712 14340
rect 25884 14300 27712 14328
rect 25884 14272 25912 14300
rect 27706 14288 27712 14300
rect 27764 14288 27770 14340
rect 24302 14260 24308 14272
rect 23952 14232 24308 14260
rect 24302 14220 24308 14232
rect 24360 14220 24366 14272
rect 25317 14263 25375 14269
rect 25317 14229 25329 14263
rect 25363 14260 25375 14263
rect 25866 14260 25872 14272
rect 25363 14232 25872 14260
rect 25363 14229 25375 14232
rect 25317 14223 25375 14229
rect 25866 14220 25872 14232
rect 25924 14220 25930 14272
rect 26326 14220 26332 14272
rect 26384 14260 26390 14272
rect 26513 14263 26571 14269
rect 26513 14260 26525 14263
rect 26384 14232 26525 14260
rect 26384 14220 26390 14232
rect 26513 14229 26525 14232
rect 26559 14229 26571 14263
rect 26513 14223 26571 14229
rect 26878 14220 26884 14272
rect 26936 14260 26942 14272
rect 27154 14260 27160 14272
rect 26936 14232 27160 14260
rect 26936 14220 26942 14232
rect 27154 14220 27160 14232
rect 27212 14220 27218 14272
rect 1104 14170 28888 14192
rect 1104 14118 5982 14170
rect 6034 14118 6046 14170
rect 6098 14118 6110 14170
rect 6162 14118 6174 14170
rect 6226 14118 15982 14170
rect 16034 14118 16046 14170
rect 16098 14118 16110 14170
rect 16162 14118 16174 14170
rect 16226 14118 25982 14170
rect 26034 14118 26046 14170
rect 26098 14118 26110 14170
rect 26162 14118 26174 14170
rect 26226 14118 28888 14170
rect 1104 14096 28888 14118
rect 2038 14056 2044 14068
rect 1999 14028 2044 14056
rect 2038 14016 2044 14028
rect 2096 14016 2102 14068
rect 2406 14056 2412 14068
rect 2367 14028 2412 14056
rect 2406 14016 2412 14028
rect 2464 14016 2470 14068
rect 4617 14059 4675 14065
rect 4617 14025 4629 14059
rect 4663 14056 4675 14059
rect 4706 14056 4712 14068
rect 4663 14028 4712 14056
rect 4663 14025 4675 14028
rect 4617 14019 4675 14025
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 5258 14016 5264 14068
rect 5316 14056 5322 14068
rect 5534 14056 5540 14068
rect 5316 14028 5540 14056
rect 5316 14016 5322 14028
rect 5534 14016 5540 14028
rect 5592 14056 5598 14068
rect 6181 14059 6239 14065
rect 6181 14056 6193 14059
rect 5592 14028 6193 14056
rect 5592 14016 5598 14028
rect 6181 14025 6193 14028
rect 6227 14056 6239 14059
rect 6365 14059 6423 14065
rect 6365 14056 6377 14059
rect 6227 14028 6377 14056
rect 6227 14025 6239 14028
rect 6181 14019 6239 14025
rect 6365 14025 6377 14028
rect 6411 14025 6423 14059
rect 6546 14056 6552 14068
rect 6507 14028 6552 14056
rect 6365 14019 6423 14025
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 8294 14056 8300 14068
rect 8255 14028 8300 14056
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 9217 14059 9275 14065
rect 9217 14025 9229 14059
rect 9263 14056 9275 14059
rect 9582 14056 9588 14068
rect 9263 14028 9588 14056
rect 9263 14025 9275 14028
rect 9217 14019 9275 14025
rect 9582 14016 9588 14028
rect 9640 14016 9646 14068
rect 10318 14016 10324 14068
rect 10376 14056 10382 14068
rect 10781 14059 10839 14065
rect 10781 14056 10793 14059
rect 10376 14028 10793 14056
rect 10376 14016 10382 14028
rect 10781 14025 10793 14028
rect 10827 14025 10839 14059
rect 14734 14056 14740 14068
rect 14695 14028 14740 14056
rect 10781 14019 10839 14025
rect 14734 14016 14740 14028
rect 14792 14016 14798 14068
rect 16482 14056 16488 14068
rect 16443 14028 16488 14056
rect 16482 14016 16488 14028
rect 16540 14016 16546 14068
rect 20070 14056 20076 14068
rect 20031 14028 20076 14056
rect 20070 14016 20076 14028
rect 20128 14016 20134 14068
rect 21358 14016 21364 14068
rect 21416 14056 21422 14068
rect 22002 14056 22008 14068
rect 21416 14028 22008 14056
rect 21416 14016 21422 14028
rect 22002 14016 22008 14028
rect 22060 14016 22066 14068
rect 23474 14056 23480 14068
rect 23435 14028 23480 14056
rect 23474 14016 23480 14028
rect 23532 14016 23538 14068
rect 24210 14056 24216 14068
rect 24171 14028 24216 14056
rect 24210 14016 24216 14028
rect 24268 14016 24274 14068
rect 25314 14056 25320 14068
rect 25275 14028 25320 14056
rect 25314 14016 25320 14028
rect 25372 14016 25378 14068
rect 27706 14056 27712 14068
rect 27667 14028 27712 14056
rect 27706 14016 27712 14028
rect 27764 14016 27770 14068
rect 1581 13991 1639 13997
rect 1581 13957 1593 13991
rect 1627 13988 1639 13991
rect 1854 13988 1860 14000
rect 1627 13960 1860 13988
rect 1627 13957 1639 13960
rect 1581 13951 1639 13957
rect 1854 13948 1860 13960
rect 1912 13948 1918 14000
rect 5169 13991 5227 13997
rect 5169 13957 5181 13991
rect 5215 13988 5227 13991
rect 5215 13960 5488 13988
rect 5215 13957 5227 13960
rect 5169 13951 5227 13957
rect 2590 13920 2596 13932
rect 2551 13892 2596 13920
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 1670 13852 1676 13864
rect 1443 13824 1676 13852
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 1670 13812 1676 13824
rect 1728 13812 1734 13864
rect 2866 13793 2872 13796
rect 2860 13784 2872 13793
rect 2827 13756 2872 13784
rect 2860 13747 2872 13756
rect 2866 13744 2872 13747
rect 2924 13744 2930 13796
rect 5460 13784 5488 13960
rect 6270 13948 6276 14000
rect 6328 13988 6334 14000
rect 6825 13991 6883 13997
rect 6825 13988 6837 13991
rect 6328 13960 6837 13988
rect 6328 13948 6334 13960
rect 6825 13957 6837 13960
rect 6871 13957 6883 13991
rect 10594 13988 10600 14000
rect 10555 13960 10600 13988
rect 6825 13951 6883 13957
rect 10594 13948 10600 13960
rect 10652 13948 10658 14000
rect 13814 13988 13820 14000
rect 13775 13960 13820 13988
rect 13814 13948 13820 13960
rect 13872 13948 13878 14000
rect 14921 13991 14979 13997
rect 14921 13957 14933 13991
rect 14967 13988 14979 13991
rect 16666 13988 16672 14000
rect 14967 13960 16672 13988
rect 14967 13957 14979 13960
rect 14921 13951 14979 13957
rect 16666 13948 16672 13960
rect 16724 13948 16730 14000
rect 19426 13988 19432 14000
rect 19387 13960 19432 13988
rect 19426 13948 19432 13960
rect 19484 13948 19490 14000
rect 26970 13948 26976 14000
rect 27028 13988 27034 14000
rect 28077 13991 28135 13997
rect 28077 13988 28089 13991
rect 27028 13960 28089 13988
rect 27028 13948 27034 13960
rect 28077 13957 28089 13960
rect 28123 13957 28135 13991
rect 28077 13951 28135 13957
rect 5813 13923 5871 13929
rect 5813 13889 5825 13923
rect 5859 13920 5871 13923
rect 6362 13920 6368 13932
rect 5859 13892 6368 13920
rect 5859 13889 5871 13892
rect 5813 13883 5871 13889
rect 6362 13880 6368 13892
rect 6420 13920 6426 13932
rect 7469 13923 7527 13929
rect 7469 13920 7481 13923
rect 6420 13892 7481 13920
rect 6420 13880 6426 13892
rect 7469 13889 7481 13892
rect 7515 13920 7527 13923
rect 7837 13923 7895 13929
rect 7837 13920 7849 13923
rect 7515 13892 7849 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 7837 13889 7849 13892
rect 7883 13889 7895 13923
rect 7837 13883 7895 13889
rect 9033 13923 9091 13929
rect 9033 13889 9045 13923
rect 9079 13920 9091 13923
rect 9490 13920 9496 13932
rect 9079 13892 9496 13920
rect 9079 13889 9091 13892
rect 9033 13883 9091 13889
rect 9490 13880 9496 13892
rect 9548 13920 9554 13932
rect 9861 13923 9919 13929
rect 9861 13920 9873 13923
rect 9548 13892 9873 13920
rect 9548 13880 9554 13892
rect 9861 13889 9873 13892
rect 9907 13920 9919 13923
rect 10410 13920 10416 13932
rect 9907 13892 10416 13920
rect 9907 13889 9919 13892
rect 9861 13883 9919 13889
rect 10410 13880 10416 13892
rect 10468 13880 10474 13932
rect 5534 13812 5540 13864
rect 5592 13852 5598 13864
rect 5592 13824 5637 13852
rect 5592 13812 5598 13824
rect 6546 13812 6552 13864
rect 6604 13852 6610 13864
rect 7285 13855 7343 13861
rect 7285 13852 7297 13855
rect 6604 13824 7297 13852
rect 6604 13812 6610 13824
rect 7285 13821 7297 13824
rect 7331 13821 7343 13855
rect 7285 13815 7343 13821
rect 5718 13784 5724 13796
rect 5460 13756 5724 13784
rect 5718 13744 5724 13756
rect 5776 13784 5782 13796
rect 6730 13784 6736 13796
rect 5776 13756 6736 13784
rect 5776 13744 5782 13756
rect 6730 13744 6736 13756
rect 6788 13744 6794 13796
rect 3878 13676 3884 13728
rect 3936 13716 3942 13728
rect 3973 13719 4031 13725
rect 3973 13716 3985 13719
rect 3936 13688 3985 13716
rect 3936 13676 3942 13688
rect 3973 13685 3985 13688
rect 4019 13685 4031 13719
rect 3973 13679 4031 13685
rect 4522 13676 4528 13728
rect 4580 13716 4586 13728
rect 5077 13719 5135 13725
rect 5077 13716 5089 13719
rect 4580 13688 5089 13716
rect 4580 13676 4586 13688
rect 5077 13685 5089 13688
rect 5123 13716 5135 13719
rect 5629 13719 5687 13725
rect 5629 13716 5641 13719
rect 5123 13688 5641 13716
rect 5123 13685 5135 13688
rect 5077 13679 5135 13685
rect 5629 13685 5641 13688
rect 5675 13716 5687 13719
rect 5902 13716 5908 13728
rect 5675 13688 5908 13716
rect 5675 13685 5687 13688
rect 5629 13679 5687 13685
rect 5902 13676 5908 13688
rect 5960 13676 5966 13728
rect 6365 13719 6423 13725
rect 6365 13685 6377 13719
rect 6411 13716 6423 13719
rect 7006 13716 7012 13728
rect 6411 13688 7012 13716
rect 6411 13685 6423 13688
rect 6365 13679 6423 13685
rect 7006 13676 7012 13688
rect 7064 13676 7070 13728
rect 7098 13676 7104 13728
rect 7156 13716 7162 13728
rect 7193 13719 7251 13725
rect 7193 13716 7205 13719
rect 7156 13688 7205 13716
rect 7156 13676 7162 13688
rect 7193 13685 7205 13688
rect 7239 13685 7251 13719
rect 7300 13716 7328 13815
rect 8202 13812 8208 13864
rect 8260 13852 8266 13864
rect 8573 13855 8631 13861
rect 8573 13852 8585 13855
rect 8260 13824 8585 13852
rect 8260 13812 8266 13824
rect 8573 13821 8585 13824
rect 8619 13821 8631 13855
rect 8573 13815 8631 13821
rect 9122 13812 9128 13864
rect 9180 13852 9186 13864
rect 10318 13852 10324 13864
rect 9180 13824 9536 13852
rect 9180 13812 9186 13824
rect 8570 13716 8576 13728
rect 7300 13688 8576 13716
rect 7193 13679 7251 13685
rect 8570 13676 8576 13688
rect 8628 13676 8634 13728
rect 9508 13716 9536 13824
rect 9600 13824 10324 13852
rect 9600 13793 9628 13824
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 10612 13852 10640 13948
rect 10870 13880 10876 13932
rect 10928 13920 10934 13932
rect 11333 13923 11391 13929
rect 11333 13920 11345 13923
rect 10928 13892 11345 13920
rect 10928 13880 10934 13892
rect 11333 13889 11345 13892
rect 11379 13920 11391 13923
rect 11422 13920 11428 13932
rect 11379 13892 11428 13920
rect 11379 13889 11391 13892
rect 11333 13883 11391 13889
rect 11422 13880 11428 13892
rect 11480 13880 11486 13932
rect 14461 13923 14519 13929
rect 14461 13889 14473 13923
rect 14507 13920 14519 13923
rect 15565 13923 15623 13929
rect 15565 13920 15577 13923
rect 14507 13892 15577 13920
rect 14507 13889 14519 13892
rect 14461 13883 14519 13889
rect 15565 13889 15577 13892
rect 15611 13920 15623 13923
rect 15838 13920 15844 13932
rect 15611 13892 15844 13920
rect 15611 13889 15623 13892
rect 15565 13883 15623 13889
rect 15838 13880 15844 13892
rect 15896 13880 15902 13932
rect 20625 13923 20683 13929
rect 20625 13889 20637 13923
rect 20671 13920 20683 13923
rect 20671 13892 21220 13920
rect 20671 13889 20683 13892
rect 20625 13883 20683 13889
rect 11241 13855 11299 13861
rect 11241 13852 11253 13855
rect 10612 13824 11253 13852
rect 11241 13821 11253 13824
rect 11287 13821 11299 13855
rect 11882 13852 11888 13864
rect 11795 13824 11888 13852
rect 11241 13815 11299 13821
rect 11882 13812 11888 13824
rect 11940 13852 11946 13864
rect 12253 13855 12311 13861
rect 12253 13852 12265 13855
rect 11940 13824 12265 13852
rect 11940 13812 11946 13824
rect 12253 13821 12265 13824
rect 12299 13852 12311 13855
rect 12437 13855 12495 13861
rect 12437 13852 12449 13855
rect 12299 13824 12449 13852
rect 12299 13821 12311 13824
rect 12253 13815 12311 13821
rect 12437 13821 12449 13824
rect 12483 13852 12495 13855
rect 13078 13852 13084 13864
rect 12483 13824 13084 13852
rect 12483 13821 12495 13824
rect 12437 13815 12495 13821
rect 13078 13812 13084 13824
rect 13136 13812 13142 13864
rect 14734 13812 14740 13864
rect 14792 13852 14798 13864
rect 15381 13855 15439 13861
rect 15381 13852 15393 13855
rect 14792 13824 15393 13852
rect 14792 13812 14798 13824
rect 15381 13821 15393 13824
rect 15427 13852 15439 13855
rect 15746 13852 15752 13864
rect 15427 13824 15752 13852
rect 15427 13821 15439 13824
rect 15381 13815 15439 13821
rect 15746 13812 15752 13824
rect 15804 13812 15810 13864
rect 16022 13852 16028 13864
rect 15983 13824 16028 13852
rect 16022 13812 16028 13824
rect 16080 13852 16086 13864
rect 16298 13852 16304 13864
rect 16080 13824 16304 13852
rect 16080 13812 16086 13824
rect 16298 13812 16304 13824
rect 16356 13812 16362 13864
rect 16390 13812 16396 13864
rect 16448 13852 16454 13864
rect 16758 13852 16764 13864
rect 16448 13824 16764 13852
rect 16448 13812 16454 13824
rect 16758 13812 16764 13824
rect 16816 13812 16822 13864
rect 17497 13855 17555 13861
rect 17497 13821 17509 13855
rect 17543 13852 17555 13855
rect 17770 13852 17776 13864
rect 17543 13824 17776 13852
rect 17543 13821 17555 13824
rect 17497 13815 17555 13821
rect 17770 13812 17776 13824
rect 17828 13812 17834 13864
rect 18049 13855 18107 13861
rect 18049 13821 18061 13855
rect 18095 13821 18107 13855
rect 21082 13852 21088 13864
rect 18049 13815 18107 13821
rect 20916 13824 21088 13852
rect 9585 13787 9643 13793
rect 9585 13753 9597 13787
rect 9631 13753 9643 13787
rect 9585 13747 9643 13753
rect 9677 13787 9735 13793
rect 9677 13753 9689 13787
rect 9723 13784 9735 13787
rect 11514 13784 11520 13796
rect 9723 13756 11520 13784
rect 9723 13753 9735 13756
rect 9677 13747 9735 13753
rect 9692 13716 9720 13747
rect 11514 13744 11520 13756
rect 11572 13744 11578 13796
rect 12710 13793 12716 13796
rect 12704 13784 12716 13793
rect 12671 13756 12716 13784
rect 12704 13747 12716 13756
rect 12710 13744 12716 13747
rect 12768 13744 12774 13796
rect 14182 13744 14188 13796
rect 14240 13784 14246 13796
rect 17402 13784 17408 13796
rect 14240 13756 17408 13784
rect 14240 13744 14246 13756
rect 17402 13744 17408 13756
rect 17460 13744 17466 13796
rect 17862 13784 17868 13796
rect 17775 13756 17868 13784
rect 10226 13716 10232 13728
rect 9508 13688 9720 13716
rect 10187 13688 10232 13716
rect 10226 13676 10232 13688
rect 10284 13676 10290 13728
rect 10870 13676 10876 13728
rect 10928 13716 10934 13728
rect 11149 13719 11207 13725
rect 11149 13716 11161 13719
rect 10928 13688 11161 13716
rect 10928 13676 10934 13688
rect 11149 13685 11161 13688
rect 11195 13685 11207 13719
rect 11149 13679 11207 13685
rect 14918 13676 14924 13728
rect 14976 13716 14982 13728
rect 15289 13719 15347 13725
rect 15289 13716 15301 13719
rect 14976 13688 15301 13716
rect 14976 13676 14982 13688
rect 15289 13685 15301 13688
rect 15335 13716 15347 13719
rect 15562 13716 15568 13728
rect 15335 13688 15568 13716
rect 15335 13685 15347 13688
rect 15289 13679 15347 13685
rect 15562 13676 15568 13688
rect 15620 13676 15626 13728
rect 16574 13676 16580 13728
rect 16632 13716 16638 13728
rect 16945 13719 17003 13725
rect 16945 13716 16957 13719
rect 16632 13688 16957 13716
rect 16632 13676 16638 13688
rect 16945 13685 16957 13688
rect 16991 13685 17003 13719
rect 16945 13679 17003 13685
rect 17126 13676 17132 13728
rect 17184 13716 17190 13728
rect 17788 13725 17816 13756
rect 17862 13744 17868 13756
rect 17920 13784 17926 13796
rect 18064 13784 18092 13815
rect 17920 13756 18092 13784
rect 17920 13744 17926 13756
rect 18230 13744 18236 13796
rect 18288 13793 18294 13796
rect 18288 13787 18352 13793
rect 18288 13753 18306 13787
rect 18340 13753 18352 13787
rect 18288 13747 18352 13753
rect 18288 13744 18294 13747
rect 17773 13719 17831 13725
rect 17773 13716 17785 13719
rect 17184 13688 17785 13716
rect 17184 13676 17190 13688
rect 17773 13685 17785 13688
rect 17819 13685 17831 13719
rect 17773 13679 17831 13685
rect 20806 13676 20812 13728
rect 20864 13716 20870 13728
rect 20916 13725 20944 13824
rect 21082 13812 21088 13824
rect 21140 13812 21146 13864
rect 21192 13852 21220 13892
rect 23474 13880 23480 13932
rect 23532 13920 23538 13932
rect 24765 13923 24823 13929
rect 24765 13920 24777 13923
rect 23532 13892 24777 13920
rect 23532 13880 23538 13892
rect 24765 13889 24777 13892
rect 24811 13920 24823 13923
rect 25682 13920 25688 13932
rect 24811 13892 25688 13920
rect 24811 13889 24823 13892
rect 24765 13883 24823 13889
rect 25682 13880 25688 13892
rect 25740 13880 25746 13932
rect 21341 13855 21399 13861
rect 21341 13852 21353 13855
rect 21192 13824 21353 13852
rect 21341 13821 21353 13824
rect 21387 13852 21399 13855
rect 23109 13855 23167 13861
rect 21387 13824 22140 13852
rect 21387 13821 21399 13824
rect 21341 13815 21399 13821
rect 22112 13796 22140 13824
rect 23109 13821 23121 13855
rect 23155 13852 23167 13855
rect 24670 13852 24676 13864
rect 23155 13824 24676 13852
rect 23155 13821 23167 13824
rect 23109 13815 23167 13821
rect 24670 13812 24676 13824
rect 24728 13812 24734 13864
rect 25777 13855 25835 13861
rect 25777 13821 25789 13855
rect 25823 13821 25835 13855
rect 25777 13815 25835 13821
rect 22094 13744 22100 13796
rect 22152 13744 22158 13796
rect 25593 13787 25651 13793
rect 25593 13784 25605 13787
rect 23952 13756 25605 13784
rect 20901 13719 20959 13725
rect 20901 13716 20913 13719
rect 20864 13688 20913 13716
rect 20864 13676 20870 13688
rect 20901 13685 20913 13688
rect 20947 13685 20959 13719
rect 20901 13679 20959 13685
rect 22186 13676 22192 13728
rect 22244 13716 22250 13728
rect 22465 13719 22523 13725
rect 22465 13716 22477 13719
rect 22244 13688 22477 13716
rect 22244 13676 22250 13688
rect 22465 13685 22477 13688
rect 22511 13685 22523 13719
rect 22465 13679 22523 13685
rect 23842 13676 23848 13728
rect 23900 13716 23906 13728
rect 23952 13725 23980 13756
rect 25593 13753 25605 13756
rect 25639 13784 25651 13787
rect 25792 13784 25820 13815
rect 25866 13812 25872 13864
rect 25924 13852 25930 13864
rect 26033 13855 26091 13861
rect 26033 13852 26045 13855
rect 25924 13824 26045 13852
rect 25924 13812 25930 13824
rect 26033 13821 26045 13824
rect 26079 13821 26091 13855
rect 26033 13815 26091 13821
rect 25639 13756 25820 13784
rect 25639 13753 25651 13756
rect 25593 13747 25651 13753
rect 23937 13719 23995 13725
rect 23937 13716 23949 13719
rect 23900 13688 23949 13716
rect 23900 13676 23906 13688
rect 23937 13685 23949 13688
rect 23983 13685 23995 13719
rect 24578 13716 24584 13728
rect 24539 13688 24584 13716
rect 23937 13679 23995 13685
rect 24578 13676 24584 13688
rect 24636 13676 24642 13728
rect 27154 13716 27160 13728
rect 27115 13688 27160 13716
rect 27154 13676 27160 13688
rect 27212 13676 27218 13728
rect 1104 13626 28888 13648
rect 1104 13574 10982 13626
rect 11034 13574 11046 13626
rect 11098 13574 11110 13626
rect 11162 13574 11174 13626
rect 11226 13574 20982 13626
rect 21034 13574 21046 13626
rect 21098 13574 21110 13626
rect 21162 13574 21174 13626
rect 21226 13574 28888 13626
rect 1104 13552 28888 13574
rect 2498 13472 2504 13524
rect 2556 13512 2562 13524
rect 4065 13515 4123 13521
rect 4065 13512 4077 13515
rect 2556 13484 4077 13512
rect 2556 13472 2562 13484
rect 4065 13481 4077 13484
rect 4111 13481 4123 13515
rect 4522 13512 4528 13524
rect 4483 13484 4528 13512
rect 4065 13475 4123 13481
rect 4522 13472 4528 13484
rect 4580 13472 4586 13524
rect 6273 13515 6331 13521
rect 6273 13481 6285 13515
rect 6319 13512 6331 13515
rect 6362 13512 6368 13524
rect 6319 13484 6368 13512
rect 6319 13481 6331 13484
rect 6273 13475 6331 13481
rect 6362 13472 6368 13484
rect 6420 13472 6426 13524
rect 6914 13512 6920 13524
rect 6472 13484 6920 13512
rect 3878 13444 3884 13456
rect 3839 13416 3884 13444
rect 3878 13404 3884 13416
rect 3936 13404 3942 13456
rect 6472 13444 6500 13484
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 9677 13515 9735 13521
rect 9677 13481 9689 13515
rect 9723 13512 9735 13515
rect 9766 13512 9772 13524
rect 9723 13484 9772 13512
rect 9723 13481 9735 13484
rect 9677 13475 9735 13481
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 10042 13512 10048 13524
rect 9955 13484 10048 13512
rect 10042 13472 10048 13484
rect 10100 13512 10106 13524
rect 10226 13512 10232 13524
rect 10100 13484 10232 13512
rect 10100 13472 10106 13484
rect 10226 13472 10232 13484
rect 10284 13472 10290 13524
rect 11241 13515 11299 13521
rect 11241 13481 11253 13515
rect 11287 13512 11299 13515
rect 11330 13512 11336 13524
rect 11287 13484 11336 13512
rect 11287 13481 11299 13484
rect 11241 13475 11299 13481
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 11514 13512 11520 13524
rect 11475 13484 11520 13512
rect 11514 13472 11520 13484
rect 11572 13472 11578 13524
rect 11790 13472 11796 13524
rect 11848 13512 11854 13524
rect 11885 13515 11943 13521
rect 11885 13512 11897 13515
rect 11848 13484 11897 13512
rect 11848 13472 11854 13484
rect 11885 13481 11897 13484
rect 11931 13481 11943 13515
rect 11885 13475 11943 13481
rect 13541 13515 13599 13521
rect 13541 13481 13553 13515
rect 13587 13512 13599 13515
rect 13722 13512 13728 13524
rect 13587 13484 13728 13512
rect 13587 13481 13599 13484
rect 13541 13475 13599 13481
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 14090 13512 14096 13524
rect 14051 13484 14096 13512
rect 14090 13472 14096 13484
rect 14148 13472 14154 13524
rect 16666 13472 16672 13524
rect 16724 13512 16730 13524
rect 18230 13512 18236 13524
rect 16724 13484 18236 13512
rect 16724 13472 16730 13484
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 19153 13515 19211 13521
rect 19153 13481 19165 13515
rect 19199 13512 19211 13515
rect 19242 13512 19248 13524
rect 19199 13484 19248 13512
rect 19199 13481 19211 13484
rect 19153 13475 19211 13481
rect 19242 13472 19248 13484
rect 19300 13472 19306 13524
rect 20254 13512 20260 13524
rect 20215 13484 20260 13512
rect 20254 13472 20260 13484
rect 20312 13472 20318 13524
rect 20714 13472 20720 13524
rect 20772 13512 20778 13524
rect 21177 13515 21235 13521
rect 21177 13512 21189 13515
rect 20772 13484 21189 13512
rect 20772 13472 20778 13484
rect 21177 13481 21189 13484
rect 21223 13481 21235 13515
rect 22738 13512 22744 13524
rect 22699 13484 22744 13512
rect 21177 13475 21235 13481
rect 22738 13472 22744 13484
rect 22796 13472 22802 13524
rect 23109 13515 23167 13521
rect 23109 13481 23121 13515
rect 23155 13512 23167 13515
rect 23198 13512 23204 13524
rect 23155 13484 23204 13512
rect 23155 13481 23167 13484
rect 23109 13475 23167 13481
rect 23198 13472 23204 13484
rect 23256 13472 23262 13524
rect 23474 13472 23480 13524
rect 23532 13512 23538 13524
rect 24121 13515 24179 13521
rect 24121 13512 24133 13515
rect 23532 13484 24133 13512
rect 23532 13472 23538 13484
rect 24121 13481 24133 13484
rect 24167 13481 24179 13515
rect 24121 13475 24179 13481
rect 24486 13472 24492 13524
rect 24544 13512 24550 13524
rect 24765 13515 24823 13521
rect 24765 13512 24777 13515
rect 24544 13484 24777 13512
rect 24544 13472 24550 13484
rect 24765 13481 24777 13484
rect 24811 13481 24823 13515
rect 25866 13512 25872 13524
rect 25827 13484 25872 13512
rect 24765 13475 24823 13481
rect 25866 13472 25872 13484
rect 25924 13472 25930 13524
rect 27614 13512 27620 13524
rect 27575 13484 27620 13512
rect 27614 13472 27620 13484
rect 27672 13472 27678 13524
rect 5644 13416 6500 13444
rect 1486 13376 1492 13388
rect 1447 13348 1492 13376
rect 1486 13336 1492 13348
rect 1544 13336 1550 13388
rect 1756 13379 1814 13385
rect 1756 13345 1768 13379
rect 1802 13376 1814 13379
rect 2314 13376 2320 13388
rect 1802 13348 2320 13376
rect 1802 13345 1814 13348
rect 1756 13339 1814 13345
rect 2314 13336 2320 13348
rect 2372 13336 2378 13388
rect 4433 13379 4491 13385
rect 4433 13345 4445 13379
rect 4479 13376 4491 13379
rect 4614 13376 4620 13388
rect 4479 13348 4620 13376
rect 4479 13345 4491 13348
rect 4433 13339 4491 13345
rect 4614 13336 4620 13348
rect 4672 13376 4678 13388
rect 5644 13385 5672 13416
rect 6822 13404 6828 13456
rect 6880 13444 6886 13456
rect 7374 13453 7380 13456
rect 7368 13444 7380 13453
rect 6880 13416 7380 13444
rect 6880 13404 6886 13416
rect 7368 13407 7380 13416
rect 7374 13404 7380 13407
rect 7432 13404 7438 13456
rect 14918 13444 14924 13456
rect 14879 13416 14924 13444
rect 14918 13404 14924 13416
rect 14976 13404 14982 13456
rect 19610 13444 19616 13456
rect 19571 13416 19616 13444
rect 19610 13404 19616 13416
rect 19668 13404 19674 13456
rect 20898 13404 20904 13456
rect 20956 13444 20962 13456
rect 21358 13444 21364 13456
rect 20956 13416 21364 13444
rect 20956 13404 20962 13416
rect 21358 13404 21364 13416
rect 21416 13404 21422 13456
rect 22649 13447 22707 13453
rect 22649 13413 22661 13447
rect 22695 13444 22707 13447
rect 24578 13444 24584 13456
rect 22695 13416 24584 13444
rect 22695 13413 22707 13416
rect 22649 13407 22707 13413
rect 24578 13404 24584 13416
rect 24636 13404 24642 13456
rect 5629 13379 5687 13385
rect 4672 13348 5304 13376
rect 4672 13336 4678 13348
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13308 4767 13311
rect 4798 13308 4804 13320
rect 4755 13280 4804 13308
rect 4755 13277 4767 13280
rect 4709 13271 4767 13277
rect 2866 13240 2872 13252
rect 2779 13212 2872 13240
rect 2866 13200 2872 13212
rect 2924 13240 2930 13252
rect 3513 13243 3571 13249
rect 3513 13240 3525 13243
rect 2924 13212 3525 13240
rect 2924 13200 2930 13212
rect 3513 13209 3525 13212
rect 3559 13240 3571 13243
rect 4724 13240 4752 13271
rect 4798 13268 4804 13280
rect 4856 13268 4862 13320
rect 5276 13317 5304 13348
rect 5629 13345 5641 13379
rect 5675 13345 5687 13379
rect 5629 13339 5687 13345
rect 5810 13336 5816 13388
rect 5868 13376 5874 13388
rect 6362 13376 6368 13388
rect 5868 13348 6368 13376
rect 5868 13336 5874 13348
rect 6362 13336 6368 13348
rect 6420 13336 6426 13388
rect 7006 13336 7012 13388
rect 7064 13376 7070 13388
rect 7101 13379 7159 13385
rect 7101 13376 7113 13379
rect 7064 13348 7113 13376
rect 7064 13336 7070 13348
rect 7101 13345 7113 13348
rect 7147 13345 7159 13379
rect 9033 13379 9091 13385
rect 9033 13376 9045 13379
rect 7101 13339 7159 13345
rect 7208 13348 9045 13376
rect 5261 13311 5319 13317
rect 5261 13277 5273 13311
rect 5307 13308 5319 13311
rect 5534 13308 5540 13320
rect 5307 13280 5540 13308
rect 5307 13277 5319 13280
rect 5261 13271 5319 13277
rect 5534 13268 5540 13280
rect 5592 13308 5598 13320
rect 6822 13308 6828 13320
rect 5592 13280 6828 13308
rect 5592 13268 5598 13280
rect 6822 13268 6828 13280
rect 6880 13268 6886 13320
rect 7208 13308 7236 13348
rect 9033 13345 9045 13348
rect 9079 13345 9091 13379
rect 9033 13339 9091 13345
rect 9493 13379 9551 13385
rect 9493 13345 9505 13379
rect 9539 13376 9551 13379
rect 10137 13379 10195 13385
rect 10137 13376 10149 13379
rect 9539 13348 10149 13376
rect 9539 13345 9551 13348
rect 9493 13339 9551 13345
rect 10137 13345 10149 13348
rect 10183 13376 10195 13379
rect 11330 13376 11336 13388
rect 10183 13348 11336 13376
rect 10183 13345 10195 13348
rect 10137 13339 10195 13345
rect 11330 13336 11336 13348
rect 11388 13336 11394 13388
rect 11422 13336 11428 13388
rect 11480 13376 11486 13388
rect 11790 13376 11796 13388
rect 11480 13348 11796 13376
rect 11480 13336 11486 13348
rect 11790 13336 11796 13348
rect 11848 13376 11854 13388
rect 11848 13348 12112 13376
rect 11848 13336 11854 13348
rect 6932 13280 7236 13308
rect 10321 13311 10379 13317
rect 3559 13212 4752 13240
rect 3559 13209 3571 13212
rect 3513 13203 3571 13209
rect 5166 13200 5172 13252
rect 5224 13240 5230 13252
rect 6932 13240 6960 13280
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 10410 13308 10416 13320
rect 10367 13280 10416 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 10410 13268 10416 13280
rect 10468 13268 10474 13320
rect 11974 13308 11980 13320
rect 11935 13280 11980 13308
rect 11974 13268 11980 13280
rect 12032 13268 12038 13320
rect 12084 13317 12112 13348
rect 13906 13336 13912 13388
rect 13964 13376 13970 13388
rect 14001 13379 14059 13385
rect 14001 13376 14013 13379
rect 13964 13348 14013 13376
rect 13964 13336 13970 13348
rect 14001 13345 14013 13348
rect 14047 13376 14059 13379
rect 15473 13379 15531 13385
rect 15473 13376 15485 13379
rect 14047 13348 15485 13376
rect 14047 13345 14059 13348
rect 14001 13339 14059 13345
rect 15473 13345 15485 13348
rect 15519 13376 15531 13379
rect 15654 13376 15660 13388
rect 15519 13348 15660 13376
rect 15519 13345 15531 13348
rect 15473 13339 15531 13345
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 16752 13379 16810 13385
rect 16752 13345 16764 13379
rect 16798 13376 16810 13379
rect 17494 13376 17500 13388
rect 16798 13348 17500 13376
rect 16798 13345 16810 13348
rect 16752 13339 16810 13345
rect 17494 13336 17500 13348
rect 17552 13336 17558 13388
rect 21545 13379 21603 13385
rect 21545 13376 21557 13379
rect 20732 13348 21557 13376
rect 12069 13311 12127 13317
rect 12069 13277 12081 13311
rect 12115 13277 12127 13311
rect 14182 13308 14188 13320
rect 14143 13280 14188 13308
rect 12069 13271 12127 13277
rect 5224 13212 6960 13240
rect 12084 13240 12112 13271
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 16485 13311 16543 13317
rect 16485 13277 16497 13311
rect 16531 13277 16543 13311
rect 19702 13308 19708 13320
rect 19663 13280 19708 13308
rect 16485 13271 16543 13277
rect 12710 13240 12716 13252
rect 12084 13212 12716 13240
rect 5224 13200 5230 13212
rect 12710 13200 12716 13212
rect 12768 13240 12774 13252
rect 12897 13243 12955 13249
rect 12897 13240 12909 13243
rect 12768 13212 12909 13240
rect 12768 13200 12774 13212
rect 12897 13209 12909 13212
rect 12943 13209 12955 13243
rect 12897 13203 12955 13209
rect 5810 13172 5816 13184
rect 5771 13144 5816 13172
rect 5810 13132 5816 13144
rect 5868 13132 5874 13184
rect 6917 13175 6975 13181
rect 6917 13141 6929 13175
rect 6963 13172 6975 13175
rect 7098 13172 7104 13184
rect 6963 13144 7104 13172
rect 6963 13141 6975 13144
rect 6917 13135 6975 13141
rect 7098 13132 7104 13144
rect 7156 13172 7162 13184
rect 8018 13172 8024 13184
rect 7156 13144 8024 13172
rect 7156 13132 7162 13144
rect 8018 13132 8024 13144
rect 8076 13132 8082 13184
rect 8481 13175 8539 13181
rect 8481 13141 8493 13175
rect 8527 13172 8539 13175
rect 8846 13172 8852 13184
rect 8527 13144 8852 13172
rect 8527 13141 8539 13144
rect 8481 13135 8539 13141
rect 8846 13132 8852 13144
rect 8904 13132 8910 13184
rect 10873 13175 10931 13181
rect 10873 13141 10885 13175
rect 10919 13172 10931 13175
rect 10962 13172 10968 13184
rect 10919 13144 10968 13172
rect 10919 13141 10931 13144
rect 10873 13135 10931 13141
rect 10962 13132 10968 13144
rect 11020 13132 11026 13184
rect 12618 13172 12624 13184
rect 12579 13144 12624 13172
rect 12618 13132 12624 13144
rect 12676 13132 12682 13184
rect 13630 13172 13636 13184
rect 13591 13144 13636 13172
rect 13630 13132 13636 13144
rect 13688 13132 13694 13184
rect 15102 13132 15108 13184
rect 15160 13172 15166 13184
rect 15378 13172 15384 13184
rect 15160 13144 15384 13172
rect 15160 13132 15166 13144
rect 15378 13132 15384 13144
rect 15436 13132 15442 13184
rect 15838 13132 15844 13184
rect 15896 13172 15902 13184
rect 15933 13175 15991 13181
rect 15933 13172 15945 13175
rect 15896 13144 15945 13172
rect 15896 13132 15902 13144
rect 15933 13141 15945 13144
rect 15979 13141 15991 13175
rect 16298 13172 16304 13184
rect 16259 13144 16304 13172
rect 15933 13135 15991 13141
rect 16298 13132 16304 13144
rect 16356 13132 16362 13184
rect 16500 13172 16528 13271
rect 19702 13268 19708 13280
rect 19760 13268 19766 13320
rect 19794 13268 19800 13320
rect 19852 13308 19858 13320
rect 19852 13280 19897 13308
rect 19852 13268 19858 13280
rect 20732 13249 20760 13348
rect 21545 13345 21557 13348
rect 21591 13345 21603 13379
rect 23750 13376 23756 13388
rect 23711 13348 23756 13376
rect 21545 13339 21603 13345
rect 23750 13336 23756 13348
rect 23808 13336 23814 13388
rect 24670 13376 24676 13388
rect 24631 13348 24676 13376
rect 24670 13336 24676 13348
rect 24728 13336 24734 13388
rect 25682 13336 25688 13388
rect 25740 13376 25746 13388
rect 26881 13379 26939 13385
rect 26881 13376 26893 13379
rect 25740 13348 26893 13376
rect 25740 13336 25746 13348
rect 26881 13345 26893 13348
rect 26927 13376 26939 13379
rect 27522 13376 27528 13388
rect 26927 13348 27528 13376
rect 26927 13345 26939 13348
rect 26881 13339 26939 13345
rect 27522 13336 27528 13348
rect 27580 13336 27586 13388
rect 21634 13308 21640 13320
rect 21595 13280 21640 13308
rect 21634 13268 21640 13280
rect 21692 13268 21698 13320
rect 21726 13268 21732 13320
rect 21784 13308 21790 13320
rect 21821 13311 21879 13317
rect 21821 13308 21833 13311
rect 21784 13280 21833 13308
rect 21784 13268 21790 13280
rect 21821 13277 21833 13280
rect 21867 13277 21879 13311
rect 23198 13308 23204 13320
rect 23159 13280 23204 13308
rect 21821 13271 21879 13277
rect 23198 13268 23204 13280
rect 23256 13268 23262 13320
rect 23293 13311 23351 13317
rect 23293 13277 23305 13311
rect 23339 13277 23351 13311
rect 23293 13271 23351 13277
rect 24949 13311 25007 13317
rect 24949 13277 24961 13311
rect 24995 13308 25007 13311
rect 25314 13308 25320 13320
rect 24995 13280 25320 13308
rect 24995 13277 25007 13280
rect 24949 13271 25007 13277
rect 19245 13243 19303 13249
rect 19245 13209 19257 13243
rect 19291 13240 19303 13243
rect 20717 13243 20775 13249
rect 20717 13240 20729 13243
rect 19291 13212 20729 13240
rect 19291 13209 19303 13212
rect 19245 13203 19303 13209
rect 20717 13209 20729 13212
rect 20763 13209 20775 13243
rect 23308 13240 23336 13271
rect 25314 13268 25320 13280
rect 25372 13268 25378 13320
rect 25866 13268 25872 13320
rect 25924 13308 25930 13320
rect 26970 13308 26976 13320
rect 25924 13280 26976 13308
rect 25924 13268 25930 13280
rect 26970 13268 26976 13280
rect 27028 13268 27034 13320
rect 27154 13308 27160 13320
rect 27115 13280 27160 13308
rect 27154 13268 27160 13280
rect 27212 13268 27218 13320
rect 20717 13203 20775 13209
rect 22204 13212 23336 13240
rect 22204 13184 22232 13212
rect 23382 13200 23388 13252
rect 23440 13240 23446 13252
rect 25590 13240 25596 13252
rect 23440 13212 25596 13240
rect 23440 13200 23446 13212
rect 25590 13200 25596 13212
rect 25648 13200 25654 13252
rect 26237 13243 26295 13249
rect 26237 13209 26249 13243
rect 26283 13240 26295 13243
rect 26418 13240 26424 13252
rect 26283 13212 26424 13240
rect 26283 13209 26295 13212
rect 26237 13203 26295 13209
rect 26418 13200 26424 13212
rect 26476 13240 26482 13252
rect 27172 13240 27200 13268
rect 26476 13212 27200 13240
rect 26476 13200 26482 13212
rect 17126 13172 17132 13184
rect 16500 13144 17132 13172
rect 17126 13132 17132 13144
rect 17184 13132 17190 13184
rect 17770 13132 17776 13184
rect 17828 13172 17834 13184
rect 17865 13175 17923 13181
rect 17865 13172 17877 13175
rect 17828 13144 17877 13172
rect 17828 13132 17834 13144
rect 17865 13141 17877 13144
rect 17911 13141 17923 13175
rect 17865 13135 17923 13141
rect 18322 13132 18328 13184
rect 18380 13172 18386 13184
rect 18417 13175 18475 13181
rect 18417 13172 18429 13175
rect 18380 13144 18429 13172
rect 18380 13132 18386 13144
rect 18417 13141 18429 13144
rect 18463 13141 18475 13175
rect 22186 13172 22192 13184
rect 22147 13144 22192 13172
rect 18417 13135 18475 13141
rect 22186 13132 22192 13144
rect 22244 13132 22250 13184
rect 24302 13172 24308 13184
rect 24263 13144 24308 13172
rect 24302 13132 24308 13144
rect 24360 13132 24366 13184
rect 25314 13172 25320 13184
rect 25275 13144 25320 13172
rect 25314 13132 25320 13144
rect 25372 13132 25378 13184
rect 26326 13132 26332 13184
rect 26384 13172 26390 13184
rect 26513 13175 26571 13181
rect 26513 13172 26525 13175
rect 26384 13144 26525 13172
rect 26384 13132 26390 13144
rect 26513 13141 26525 13144
rect 26559 13141 26571 13175
rect 26513 13135 26571 13141
rect 1104 13082 28888 13104
rect 1104 13030 5982 13082
rect 6034 13030 6046 13082
rect 6098 13030 6110 13082
rect 6162 13030 6174 13082
rect 6226 13030 15982 13082
rect 16034 13030 16046 13082
rect 16098 13030 16110 13082
rect 16162 13030 16174 13082
rect 16226 13030 25982 13082
rect 26034 13030 26046 13082
rect 26098 13030 26110 13082
rect 26162 13030 26174 13082
rect 26226 13030 28888 13082
rect 1104 13008 28888 13030
rect 566 12928 572 12980
rect 624 12968 630 12980
rect 4525 12971 4583 12977
rect 624 12940 2636 12968
rect 624 12928 630 12940
rect 2608 12900 2636 12940
rect 4525 12937 4537 12971
rect 4571 12968 4583 12971
rect 4614 12968 4620 12980
rect 4571 12940 4620 12968
rect 4571 12937 4583 12940
rect 4525 12931 4583 12937
rect 4614 12928 4620 12940
rect 4672 12928 4678 12980
rect 4798 12968 4804 12980
rect 4759 12940 4804 12968
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 5534 12928 5540 12980
rect 5592 12968 5598 12980
rect 6457 12971 6515 12977
rect 6457 12968 6469 12971
rect 5592 12940 6469 12968
rect 5592 12928 5598 12940
rect 6457 12937 6469 12940
rect 6503 12968 6515 12971
rect 6549 12971 6607 12977
rect 6549 12968 6561 12971
rect 6503 12940 6561 12968
rect 6503 12937 6515 12940
rect 6457 12931 6515 12937
rect 6549 12937 6561 12940
rect 6595 12937 6607 12971
rect 6549 12931 6607 12937
rect 7006 12928 7012 12980
rect 7064 12968 7070 12980
rect 8573 12971 8631 12977
rect 8573 12968 8585 12971
rect 7064 12940 8585 12968
rect 7064 12928 7070 12940
rect 8573 12937 8585 12940
rect 8619 12937 8631 12971
rect 8573 12931 8631 12937
rect 11241 12971 11299 12977
rect 11241 12937 11253 12971
rect 11287 12968 11299 12971
rect 11514 12968 11520 12980
rect 11287 12940 11520 12968
rect 11287 12937 11299 12940
rect 11241 12931 11299 12937
rect 3050 12900 3056 12912
rect 2608 12872 3056 12900
rect 3050 12860 3056 12872
rect 3108 12900 3114 12912
rect 4982 12900 4988 12912
rect 3108 12872 4988 12900
rect 3108 12860 3114 12872
rect 4982 12860 4988 12872
rect 5040 12900 5046 12912
rect 6178 12900 6184 12912
rect 5040 12872 6184 12900
rect 5040 12860 5046 12872
rect 6178 12860 6184 12872
rect 6236 12860 6242 12912
rect 6273 12903 6331 12909
rect 6273 12869 6285 12903
rect 6319 12900 6331 12903
rect 6914 12900 6920 12912
rect 6319 12872 6920 12900
rect 6319 12869 6331 12872
rect 6273 12863 6331 12869
rect 6914 12860 6920 12872
rect 6972 12860 6978 12912
rect 1486 12792 1492 12844
rect 1544 12832 1550 12844
rect 1673 12835 1731 12841
rect 1673 12832 1685 12835
rect 1544 12804 1685 12832
rect 1544 12792 1550 12804
rect 1673 12801 1685 12804
rect 1719 12801 1731 12835
rect 1673 12795 1731 12801
rect 1688 12764 1716 12795
rect 4062 12792 4068 12844
rect 4120 12832 4126 12844
rect 4157 12835 4215 12841
rect 4157 12832 4169 12835
rect 4120 12804 4169 12832
rect 4120 12792 4126 12804
rect 4157 12801 4169 12804
rect 4203 12832 4215 12835
rect 4522 12832 4528 12844
rect 4203 12804 4528 12832
rect 4203 12801 4215 12804
rect 4157 12795 4215 12801
rect 4522 12792 4528 12804
rect 4580 12792 4586 12844
rect 5626 12792 5632 12844
rect 5684 12832 5690 12844
rect 5721 12835 5779 12841
rect 5721 12832 5733 12835
rect 5684 12804 5733 12832
rect 5684 12792 5690 12804
rect 5721 12801 5733 12804
rect 5767 12832 5779 12835
rect 6546 12832 6552 12844
rect 5767 12804 6552 12832
rect 5767 12801 5779 12804
rect 5721 12795 5779 12801
rect 6546 12792 6552 12804
rect 6604 12832 6610 12844
rect 7653 12835 7711 12841
rect 7653 12832 7665 12835
rect 6604 12804 7665 12832
rect 6604 12792 6610 12804
rect 7653 12801 7665 12804
rect 7699 12801 7711 12835
rect 8588 12832 8616 12931
rect 11514 12928 11520 12940
rect 11572 12968 11578 12980
rect 11974 12968 11980 12980
rect 11572 12940 11980 12968
rect 11572 12928 11578 12940
rect 11974 12928 11980 12940
rect 12032 12928 12038 12980
rect 13725 12971 13783 12977
rect 13725 12937 13737 12971
rect 13771 12968 13783 12971
rect 14090 12968 14096 12980
rect 13771 12940 14096 12968
rect 13771 12937 13783 12940
rect 13725 12931 13783 12937
rect 14090 12928 14096 12940
rect 14148 12928 14154 12980
rect 14829 12971 14887 12977
rect 14829 12937 14841 12971
rect 14875 12968 14887 12971
rect 15838 12968 15844 12980
rect 14875 12940 15844 12968
rect 14875 12937 14887 12940
rect 14829 12931 14887 12937
rect 15838 12928 15844 12940
rect 15896 12968 15902 12980
rect 17494 12968 17500 12980
rect 15896 12940 16804 12968
rect 17455 12940 17500 12968
rect 15896 12928 15902 12940
rect 10137 12903 10195 12909
rect 10137 12869 10149 12903
rect 10183 12900 10195 12903
rect 10870 12900 10876 12912
rect 10183 12872 10876 12900
rect 10183 12869 10195 12872
rect 10137 12863 10195 12869
rect 10870 12860 10876 12872
rect 10928 12860 10934 12912
rect 11698 12860 11704 12912
rect 11756 12900 11762 12912
rect 11793 12903 11851 12909
rect 11793 12900 11805 12903
rect 11756 12872 11805 12900
rect 11756 12860 11762 12872
rect 11793 12869 11805 12872
rect 11839 12900 11851 12903
rect 12158 12900 12164 12912
rect 11839 12872 12020 12900
rect 12119 12872 12164 12900
rect 11839 12869 11851 12872
rect 11793 12863 11851 12869
rect 11992 12844 12020 12872
rect 12158 12860 12164 12872
rect 12216 12860 12222 12912
rect 14734 12900 14740 12912
rect 14647 12872 14740 12900
rect 14734 12860 14740 12872
rect 14792 12900 14798 12912
rect 15102 12900 15108 12912
rect 14792 12872 15108 12900
rect 14792 12860 14798 12872
rect 15102 12860 15108 12872
rect 15160 12900 15166 12912
rect 16393 12903 16451 12909
rect 15160 12872 15332 12900
rect 15160 12860 15166 12872
rect 8757 12835 8815 12841
rect 8757 12832 8769 12835
rect 8588 12804 8769 12832
rect 7653 12795 7711 12801
rect 8757 12801 8769 12804
rect 8803 12801 8815 12835
rect 8757 12795 8815 12801
rect 10962 12792 10968 12844
rect 11020 12832 11026 12844
rect 11333 12835 11391 12841
rect 11333 12832 11345 12835
rect 11020 12804 11345 12832
rect 11020 12792 11026 12804
rect 11333 12801 11345 12804
rect 11379 12801 11391 12835
rect 11333 12795 11391 12801
rect 11974 12792 11980 12844
rect 12032 12792 12038 12844
rect 2222 12764 2228 12776
rect 1688 12736 2228 12764
rect 2222 12724 2228 12736
rect 2280 12724 2286 12776
rect 5166 12724 5172 12776
rect 5224 12764 5230 12776
rect 5537 12767 5595 12773
rect 5537 12764 5549 12767
rect 5224 12736 5549 12764
rect 5224 12724 5230 12736
rect 5537 12733 5549 12736
rect 5583 12733 5595 12767
rect 7558 12764 7564 12776
rect 7519 12736 7564 12764
rect 5537 12727 5595 12733
rect 7558 12724 7564 12736
rect 7616 12764 7622 12776
rect 8113 12767 8171 12773
rect 8113 12764 8125 12767
rect 7616 12736 8125 12764
rect 7616 12724 7622 12736
rect 8113 12733 8125 12736
rect 8159 12733 8171 12767
rect 8113 12727 8171 12733
rect 8846 12724 8852 12776
rect 8904 12764 8910 12776
rect 9013 12767 9071 12773
rect 9013 12764 9025 12767
rect 8904 12736 9025 12764
rect 8904 12724 8910 12736
rect 9013 12733 9025 12736
rect 9059 12733 9071 12767
rect 12176 12764 12204 12860
rect 12342 12792 12348 12844
rect 12400 12832 12406 12844
rect 12618 12832 12624 12844
rect 12400 12804 12624 12832
rect 12400 12792 12406 12804
rect 12618 12792 12624 12804
rect 12676 12832 12682 12844
rect 15304 12841 15332 12872
rect 16393 12869 16405 12903
rect 16439 12900 16451 12903
rect 16482 12900 16488 12912
rect 16439 12872 16488 12900
rect 16439 12869 16451 12872
rect 16393 12863 16451 12869
rect 16482 12860 16488 12872
rect 16540 12860 16546 12912
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 12676 12804 13001 12832
rect 12676 12792 12682 12804
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 15289 12835 15347 12841
rect 15289 12801 15301 12835
rect 15335 12801 15347 12835
rect 15289 12795 15347 12801
rect 15378 12792 15384 12844
rect 15436 12832 15442 12844
rect 15473 12835 15531 12841
rect 15473 12832 15485 12835
rect 15436 12804 15485 12832
rect 15436 12792 15442 12804
rect 15473 12801 15485 12804
rect 15519 12832 15531 12835
rect 15933 12835 15991 12841
rect 15933 12832 15945 12835
rect 15519 12804 15945 12832
rect 15519 12801 15531 12804
rect 15473 12795 15531 12801
rect 15933 12801 15945 12804
rect 15979 12832 15991 12835
rect 16666 12832 16672 12844
rect 15979 12804 16672 12832
rect 15979 12801 15991 12804
rect 15933 12795 15991 12801
rect 16666 12792 16672 12804
rect 16724 12792 16730 12844
rect 12897 12767 12955 12773
rect 12897 12764 12909 12767
rect 12176 12736 12909 12764
rect 9013 12727 9071 12733
rect 12897 12733 12909 12736
rect 12943 12733 12955 12767
rect 12897 12727 12955 12733
rect 13906 12724 13912 12776
rect 13964 12764 13970 12776
rect 14001 12767 14059 12773
rect 14001 12764 14013 12767
rect 13964 12736 14013 12764
rect 13964 12724 13970 12736
rect 14001 12733 14013 12736
rect 14047 12733 14059 12767
rect 14001 12727 14059 12733
rect 15102 12724 15108 12776
rect 15160 12764 15166 12776
rect 15197 12767 15255 12773
rect 15197 12764 15209 12767
rect 15160 12736 15209 12764
rect 15160 12724 15166 12736
rect 15197 12733 15209 12736
rect 15243 12764 15255 12767
rect 16574 12764 16580 12776
rect 15243 12736 16580 12764
rect 15243 12733 15255 12736
rect 15197 12727 15255 12733
rect 16574 12724 16580 12736
rect 16632 12724 16638 12776
rect 16776 12773 16804 12940
rect 17494 12928 17500 12940
rect 17552 12928 17558 12980
rect 19702 12928 19708 12980
rect 19760 12968 19766 12980
rect 19981 12971 20039 12977
rect 19981 12968 19993 12971
rect 19760 12940 19993 12968
rect 19760 12928 19766 12940
rect 19981 12937 19993 12940
rect 20027 12937 20039 12971
rect 19981 12931 20039 12937
rect 21910 12928 21916 12980
rect 21968 12968 21974 12980
rect 22094 12968 22100 12980
rect 21968 12940 22100 12968
rect 21968 12928 21974 12940
rect 22094 12928 22100 12940
rect 22152 12968 22158 12980
rect 22373 12971 22431 12977
rect 22373 12968 22385 12971
rect 22152 12940 22385 12968
rect 22152 12928 22158 12940
rect 22373 12937 22385 12940
rect 22419 12937 22431 12971
rect 23014 12968 23020 12980
rect 22927 12940 23020 12968
rect 22373 12931 22431 12937
rect 23014 12928 23020 12940
rect 23072 12968 23078 12980
rect 23198 12968 23204 12980
rect 23072 12940 23204 12968
rect 23072 12928 23078 12940
rect 23198 12928 23204 12940
rect 23256 12928 23262 12980
rect 24486 12928 24492 12980
rect 24544 12968 24550 12980
rect 24857 12971 24915 12977
rect 24857 12968 24869 12971
rect 24544 12940 24869 12968
rect 24544 12928 24550 12940
rect 24857 12937 24869 12940
rect 24903 12937 24915 12971
rect 25682 12968 25688 12980
rect 25643 12940 25688 12968
rect 24857 12931 24915 12937
rect 25682 12928 25688 12940
rect 25740 12928 25746 12980
rect 27154 12928 27160 12980
rect 27212 12968 27218 12980
rect 28077 12971 28135 12977
rect 28077 12968 28089 12971
rect 27212 12940 28089 12968
rect 27212 12928 27218 12940
rect 28077 12937 28089 12940
rect 28123 12937 28135 12971
rect 28077 12931 28135 12937
rect 17034 12832 17040 12844
rect 16947 12804 17040 12832
rect 17034 12792 17040 12804
rect 17092 12832 17098 12844
rect 17512 12832 17540 12928
rect 19429 12903 19487 12909
rect 19429 12869 19441 12903
rect 19475 12900 19487 12903
rect 20070 12900 20076 12912
rect 19475 12872 20076 12900
rect 19475 12869 19487 12872
rect 19429 12863 19487 12869
rect 20070 12860 20076 12872
rect 20128 12860 20134 12912
rect 23750 12860 23756 12912
rect 23808 12900 23814 12912
rect 23808 12872 24256 12900
rect 23808 12860 23814 12872
rect 17092 12804 17540 12832
rect 17092 12792 17098 12804
rect 23198 12792 23204 12844
rect 23256 12832 23262 12844
rect 24228 12841 24256 12872
rect 24762 12860 24768 12912
rect 24820 12900 24826 12912
rect 25866 12900 25872 12912
rect 24820 12872 25872 12900
rect 24820 12860 24826 12872
rect 25866 12860 25872 12872
rect 25924 12900 25930 12912
rect 25961 12903 26019 12909
rect 25961 12900 25973 12903
rect 25924 12872 25973 12900
rect 25924 12860 25930 12872
rect 25961 12869 25973 12872
rect 26007 12869 26019 12903
rect 25961 12863 26019 12869
rect 23477 12835 23535 12841
rect 23477 12832 23489 12835
rect 23256 12804 23489 12832
rect 23256 12792 23262 12804
rect 23477 12801 23489 12804
rect 23523 12832 23535 12835
rect 24213 12835 24271 12841
rect 23523 12804 24164 12832
rect 23523 12801 23535 12804
rect 23477 12795 23535 12801
rect 16761 12767 16819 12773
rect 16761 12733 16773 12767
rect 16807 12733 16819 12767
rect 16761 12727 16819 12733
rect 17126 12724 17132 12776
rect 17184 12764 17190 12776
rect 18322 12773 18328 12776
rect 17865 12767 17923 12773
rect 17865 12764 17877 12767
rect 17184 12736 17877 12764
rect 17184 12724 17190 12736
rect 17865 12733 17877 12736
rect 17911 12764 17923 12767
rect 18049 12767 18107 12773
rect 18049 12764 18061 12767
rect 17911 12736 18061 12764
rect 17911 12733 17923 12736
rect 17865 12727 17923 12733
rect 18049 12733 18061 12736
rect 18095 12733 18107 12767
rect 18316 12764 18328 12773
rect 18283 12736 18328 12764
rect 18049 12727 18107 12733
rect 18316 12727 18328 12736
rect 1940 12699 1998 12705
rect 1940 12665 1952 12699
rect 1986 12696 1998 12699
rect 5629 12699 5687 12705
rect 1986 12668 3464 12696
rect 1986 12665 1998 12668
rect 1940 12659 1998 12665
rect 3436 12640 3464 12668
rect 5629 12665 5641 12699
rect 5675 12696 5687 12699
rect 5718 12696 5724 12708
rect 5675 12668 5724 12696
rect 5675 12665 5687 12668
rect 5629 12659 5687 12665
rect 5718 12656 5724 12668
rect 5776 12656 5782 12708
rect 6457 12699 6515 12705
rect 6457 12665 6469 12699
rect 6503 12696 6515 12699
rect 7466 12696 7472 12708
rect 6503 12668 7472 12696
rect 6503 12665 6515 12668
rect 6457 12659 6515 12665
rect 7466 12656 7472 12668
rect 7524 12656 7530 12708
rect 16114 12656 16120 12708
rect 16172 12696 16178 12708
rect 16853 12699 16911 12705
rect 16853 12696 16865 12699
rect 16172 12668 16865 12696
rect 16172 12656 16178 12668
rect 16853 12665 16865 12668
rect 16899 12665 16911 12699
rect 18064 12696 18092 12727
rect 18322 12724 18328 12727
rect 18380 12724 18386 12776
rect 20714 12764 20720 12776
rect 20627 12736 20720 12764
rect 20714 12724 20720 12736
rect 20772 12764 20778 12776
rect 20993 12767 21051 12773
rect 20993 12764 21005 12767
rect 20772 12736 21005 12764
rect 20772 12724 20778 12736
rect 20993 12733 21005 12736
rect 21039 12733 21051 12767
rect 20993 12727 21051 12733
rect 23106 12724 23112 12776
rect 23164 12764 23170 12776
rect 23290 12764 23296 12776
rect 23164 12736 23296 12764
rect 23164 12724 23170 12736
rect 23290 12724 23296 12736
rect 23348 12724 23354 12776
rect 24136 12773 24164 12804
rect 24213 12801 24225 12835
rect 24259 12801 24271 12835
rect 24394 12832 24400 12844
rect 24355 12804 24400 12832
rect 24213 12795 24271 12801
rect 24394 12792 24400 12804
rect 24452 12792 24458 12844
rect 27246 12792 27252 12844
rect 27304 12832 27310 12844
rect 27304 12804 27568 12832
rect 27304 12792 27310 12804
rect 27540 12776 27568 12804
rect 24121 12767 24179 12773
rect 24121 12733 24133 12767
rect 24167 12733 24179 12767
rect 26142 12764 26148 12776
rect 26103 12736 26148 12764
rect 24121 12727 24179 12733
rect 26142 12724 26148 12736
rect 26200 12724 26206 12776
rect 26418 12773 26424 12776
rect 26412 12764 26424 12773
rect 26379 12736 26424 12764
rect 26412 12727 26424 12736
rect 26418 12724 26424 12727
rect 26476 12724 26482 12776
rect 27522 12724 27528 12776
rect 27580 12724 27586 12776
rect 19242 12696 19248 12708
rect 18064 12668 19248 12696
rect 16853 12659 16911 12665
rect 19242 12656 19248 12668
rect 19300 12656 19306 12708
rect 19886 12656 19892 12708
rect 19944 12696 19950 12708
rect 20441 12699 20499 12705
rect 20441 12696 20453 12699
rect 19944 12668 20453 12696
rect 19944 12656 19950 12668
rect 20441 12665 20453 12668
rect 20487 12696 20499 12699
rect 21238 12699 21296 12705
rect 21238 12696 21250 12699
rect 20487 12668 21250 12696
rect 20487 12665 20499 12668
rect 20441 12659 20499 12665
rect 21238 12665 21250 12668
rect 21284 12665 21296 12699
rect 21238 12659 21296 12665
rect 23474 12656 23480 12708
rect 23532 12696 23538 12708
rect 24670 12696 24676 12708
rect 23532 12668 24676 12696
rect 23532 12656 23538 12668
rect 24670 12656 24676 12668
rect 24728 12696 24734 12708
rect 25133 12699 25191 12705
rect 25133 12696 25145 12699
rect 24728 12668 25145 12696
rect 24728 12656 24734 12668
rect 25133 12665 25145 12668
rect 25179 12665 25191 12699
rect 25133 12659 25191 12665
rect 26970 12656 26976 12708
rect 27028 12696 27034 12708
rect 27246 12696 27252 12708
rect 27028 12668 27252 12696
rect 27028 12656 27034 12668
rect 27246 12656 27252 12668
rect 27304 12656 27310 12708
rect 2314 12588 2320 12640
rect 2372 12628 2378 12640
rect 2498 12628 2504 12640
rect 2372 12600 2504 12628
rect 2372 12588 2378 12600
rect 2498 12588 2504 12600
rect 2556 12628 2562 12640
rect 3053 12631 3111 12637
rect 3053 12628 3065 12631
rect 2556 12600 3065 12628
rect 2556 12588 2562 12600
rect 3053 12597 3065 12600
rect 3099 12597 3111 12631
rect 3053 12591 3111 12597
rect 3418 12588 3424 12640
rect 3476 12628 3482 12640
rect 3605 12631 3663 12637
rect 3605 12628 3617 12631
rect 3476 12600 3617 12628
rect 3476 12588 3482 12600
rect 3605 12597 3617 12600
rect 3651 12597 3663 12631
rect 5166 12628 5172 12640
rect 5127 12600 5172 12628
rect 3605 12591 3663 12597
rect 5166 12588 5172 12600
rect 5224 12588 5230 12640
rect 7101 12631 7159 12637
rect 7101 12597 7113 12631
rect 7147 12628 7159 12631
rect 7282 12628 7288 12640
rect 7147 12600 7288 12628
rect 7147 12597 7159 12600
rect 7101 12591 7159 12597
rect 7282 12588 7288 12600
rect 7340 12588 7346 12640
rect 10778 12628 10784 12640
rect 10739 12600 10784 12628
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 12492 12600 12537 12628
rect 12492 12588 12498 12600
rect 12710 12588 12716 12640
rect 12768 12628 12774 12640
rect 12805 12631 12863 12637
rect 12805 12628 12817 12631
rect 12768 12600 12817 12628
rect 12768 12588 12774 12600
rect 12805 12597 12817 12600
rect 12851 12628 12863 12631
rect 12986 12628 12992 12640
rect 12851 12600 12992 12628
rect 12851 12597 12863 12600
rect 12805 12591 12863 12597
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 16301 12631 16359 12637
rect 16301 12597 16313 12631
rect 16347 12628 16359 12631
rect 17126 12628 17132 12640
rect 16347 12600 17132 12628
rect 16347 12597 16359 12600
rect 16301 12591 16359 12597
rect 17126 12588 17132 12600
rect 17184 12588 17190 12640
rect 19334 12588 19340 12640
rect 19392 12628 19398 12640
rect 20717 12631 20775 12637
rect 20717 12628 20729 12631
rect 19392 12600 20729 12628
rect 19392 12588 19398 12600
rect 20717 12597 20729 12600
rect 20763 12628 20775 12631
rect 20809 12631 20867 12637
rect 20809 12628 20821 12631
rect 20763 12600 20821 12628
rect 20763 12597 20775 12600
rect 20717 12591 20775 12597
rect 20809 12597 20821 12600
rect 20855 12597 20867 12631
rect 23750 12628 23756 12640
rect 23711 12600 23756 12628
rect 20809 12591 20867 12597
rect 23750 12588 23756 12600
rect 23808 12588 23814 12640
rect 27154 12588 27160 12640
rect 27212 12628 27218 12640
rect 27525 12631 27583 12637
rect 27525 12628 27537 12631
rect 27212 12600 27537 12628
rect 27212 12588 27218 12600
rect 27525 12597 27537 12600
rect 27571 12597 27583 12631
rect 27525 12591 27583 12597
rect 1104 12538 28888 12560
rect 1104 12486 10982 12538
rect 11034 12486 11046 12538
rect 11098 12486 11110 12538
rect 11162 12486 11174 12538
rect 11226 12486 20982 12538
rect 21034 12486 21046 12538
rect 21098 12486 21110 12538
rect 21162 12486 21174 12538
rect 21226 12486 28888 12538
rect 1104 12464 28888 12486
rect 1949 12427 2007 12433
rect 1949 12393 1961 12427
rect 1995 12424 2007 12427
rect 2222 12424 2228 12436
rect 1995 12396 2228 12424
rect 1995 12393 2007 12396
rect 1949 12387 2007 12393
rect 2222 12384 2228 12396
rect 2280 12384 2286 12436
rect 3694 12384 3700 12436
rect 3752 12424 3758 12436
rect 5810 12424 5816 12436
rect 3752 12396 5816 12424
rect 3752 12384 3758 12396
rect 5810 12384 5816 12396
rect 5868 12384 5874 12436
rect 7006 12424 7012 12436
rect 6967 12396 7012 12424
rect 7006 12384 7012 12396
rect 7064 12384 7070 12436
rect 7098 12384 7104 12436
rect 7156 12424 7162 12436
rect 8202 12424 8208 12436
rect 7156 12396 8208 12424
rect 7156 12384 7162 12396
rect 8202 12384 8208 12396
rect 8260 12384 8266 12436
rect 8846 12424 8852 12436
rect 8807 12396 8852 12424
rect 8846 12384 8852 12396
rect 8904 12384 8910 12436
rect 9953 12427 10011 12433
rect 9953 12393 9965 12427
rect 9999 12424 10011 12427
rect 10410 12424 10416 12436
rect 9999 12396 10416 12424
rect 9999 12393 10011 12396
rect 9953 12387 10011 12393
rect 10410 12384 10416 12396
rect 10468 12384 10474 12436
rect 10778 12384 10784 12436
rect 10836 12424 10842 12436
rect 11790 12424 11796 12436
rect 10836 12396 11796 12424
rect 10836 12384 10842 12396
rect 11790 12384 11796 12396
rect 11848 12424 11854 12436
rect 11977 12427 12035 12433
rect 11977 12424 11989 12427
rect 11848 12396 11989 12424
rect 11848 12384 11854 12396
rect 11977 12393 11989 12396
rect 12023 12393 12035 12427
rect 11977 12387 12035 12393
rect 12621 12427 12679 12433
rect 12621 12393 12633 12427
rect 12667 12424 12679 12427
rect 12710 12424 12716 12436
rect 12667 12396 12716 12424
rect 12667 12393 12679 12396
rect 12621 12387 12679 12393
rect 12710 12384 12716 12396
rect 12768 12384 12774 12436
rect 13998 12424 14004 12436
rect 13959 12396 14004 12424
rect 13998 12384 14004 12396
rect 14056 12384 14062 12436
rect 14921 12427 14979 12433
rect 14921 12393 14933 12427
rect 14967 12424 14979 12427
rect 15102 12424 15108 12436
rect 14967 12396 15108 12424
rect 14967 12393 14979 12396
rect 14921 12387 14979 12393
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 15565 12427 15623 12433
rect 15565 12393 15577 12427
rect 15611 12393 15623 12427
rect 15565 12387 15623 12393
rect 5166 12316 5172 12368
rect 5224 12356 5230 12368
rect 5718 12356 5724 12368
rect 5224 12328 5724 12356
rect 5224 12316 5230 12328
rect 5718 12316 5724 12328
rect 5776 12356 5782 12368
rect 10870 12365 10876 12368
rect 9125 12359 9183 12365
rect 9125 12356 9137 12359
rect 5776 12328 9137 12356
rect 5776 12316 5782 12328
rect 9125 12325 9137 12328
rect 9171 12325 9183 12359
rect 10864 12356 10876 12365
rect 10783 12328 10876 12356
rect 9125 12319 9183 12325
rect 10864 12319 10876 12328
rect 10928 12356 10934 12368
rect 11422 12356 11428 12368
rect 10928 12328 11428 12356
rect 10870 12316 10876 12319
rect 10928 12316 10934 12328
rect 11422 12316 11428 12328
rect 11480 12356 11486 12368
rect 12342 12356 12348 12368
rect 11480 12328 12348 12356
rect 11480 12316 11486 12328
rect 12342 12316 12348 12328
rect 12400 12316 12406 12368
rect 13725 12359 13783 12365
rect 13725 12325 13737 12359
rect 13771 12356 13783 12359
rect 14182 12356 14188 12368
rect 13771 12328 14188 12356
rect 13771 12325 13783 12328
rect 13725 12319 13783 12325
rect 14182 12316 14188 12328
rect 14240 12316 14246 12368
rect 15580 12356 15608 12387
rect 15838 12384 15844 12436
rect 15896 12424 15902 12436
rect 16025 12427 16083 12433
rect 16025 12424 16037 12427
rect 15896 12396 16037 12424
rect 15896 12384 15902 12396
rect 16025 12393 16037 12396
rect 16071 12393 16083 12427
rect 16025 12387 16083 12393
rect 16669 12427 16727 12433
rect 16669 12393 16681 12427
rect 16715 12424 16727 12427
rect 17034 12424 17040 12436
rect 16715 12396 17040 12424
rect 16715 12393 16727 12396
rect 16669 12387 16727 12393
rect 17034 12384 17040 12396
rect 17092 12384 17098 12436
rect 18322 12384 18328 12436
rect 18380 12424 18386 12436
rect 18509 12427 18567 12433
rect 18509 12424 18521 12427
rect 18380 12396 18521 12424
rect 18380 12384 18386 12396
rect 18509 12393 18521 12396
rect 18555 12393 18567 12427
rect 18509 12387 18567 12393
rect 19337 12427 19395 12433
rect 19337 12393 19349 12427
rect 19383 12424 19395 12427
rect 19610 12424 19616 12436
rect 19383 12396 19616 12424
rect 19383 12393 19395 12396
rect 19337 12387 19395 12393
rect 19610 12384 19616 12396
rect 19668 12384 19674 12436
rect 19705 12427 19763 12433
rect 19705 12393 19717 12427
rect 19751 12424 19763 12427
rect 19794 12424 19800 12436
rect 19751 12396 19800 12424
rect 19751 12393 19763 12396
rect 19705 12387 19763 12393
rect 19794 12384 19800 12396
rect 19852 12384 19858 12436
rect 21269 12427 21327 12433
rect 21269 12393 21281 12427
rect 21315 12424 21327 12427
rect 21726 12424 21732 12436
rect 21315 12396 21732 12424
rect 21315 12393 21327 12396
rect 21269 12387 21327 12393
rect 21726 12384 21732 12396
rect 21784 12384 21790 12436
rect 21821 12427 21879 12433
rect 21821 12393 21833 12427
rect 21867 12424 21879 12427
rect 22738 12424 22744 12436
rect 21867 12396 22744 12424
rect 21867 12393 21879 12396
rect 21821 12387 21879 12393
rect 22738 12384 22744 12396
rect 22796 12384 22802 12436
rect 22833 12427 22891 12433
rect 22833 12393 22845 12427
rect 22879 12424 22891 12427
rect 23106 12424 23112 12436
rect 22879 12396 23112 12424
rect 22879 12393 22891 12396
rect 22833 12387 22891 12393
rect 23106 12384 23112 12396
rect 23164 12384 23170 12436
rect 26510 12384 26516 12436
rect 26568 12424 26574 12436
rect 26970 12424 26976 12436
rect 26568 12396 26976 12424
rect 26568 12384 26574 12396
rect 26970 12384 26976 12396
rect 27028 12384 27034 12436
rect 16114 12356 16120 12368
rect 15580 12328 16120 12356
rect 16114 12316 16120 12328
rect 16172 12356 16178 12368
rect 16298 12356 16304 12368
rect 16172 12328 16304 12356
rect 16172 12316 16178 12328
rect 16298 12316 16304 12328
rect 16356 12316 16362 12368
rect 2777 12291 2835 12297
rect 2777 12257 2789 12291
rect 2823 12257 2835 12291
rect 2777 12251 2835 12257
rect 1397 12223 1455 12229
rect 1397 12189 1409 12223
rect 1443 12220 1455 12223
rect 1670 12220 1676 12232
rect 1443 12192 1676 12220
rect 1443 12189 1455 12192
rect 1397 12183 1455 12189
rect 1670 12180 1676 12192
rect 1728 12180 1734 12232
rect 2406 12084 2412 12096
rect 2367 12056 2412 12084
rect 2406 12044 2412 12056
rect 2464 12044 2470 12096
rect 2792 12084 2820 12251
rect 2866 12248 2872 12300
rect 2924 12288 2930 12300
rect 3421 12291 3479 12297
rect 3421 12288 3433 12291
rect 2924 12260 3433 12288
rect 2924 12248 2930 12260
rect 3421 12257 3433 12260
rect 3467 12257 3479 12291
rect 3421 12251 3479 12257
rect 4065 12291 4123 12297
rect 4065 12257 4077 12291
rect 4111 12288 4123 12291
rect 4154 12288 4160 12300
rect 4111 12260 4160 12288
rect 4111 12257 4123 12260
rect 4065 12251 4123 12257
rect 4154 12248 4160 12260
rect 4212 12248 4218 12300
rect 5813 12291 5871 12297
rect 5813 12257 5825 12291
rect 5859 12288 5871 12291
rect 6362 12288 6368 12300
rect 5859 12260 6368 12288
rect 5859 12257 5871 12260
rect 5813 12251 5871 12257
rect 6362 12248 6368 12260
rect 6420 12248 6426 12300
rect 6638 12248 6644 12300
rect 6696 12288 6702 12300
rect 7469 12291 7527 12297
rect 7469 12288 7481 12291
rect 6696 12260 7481 12288
rect 6696 12248 6702 12260
rect 7469 12257 7481 12260
rect 7515 12257 7527 12291
rect 7469 12251 7527 12257
rect 7558 12248 7564 12300
rect 7616 12288 7622 12300
rect 15930 12288 15936 12300
rect 7616 12260 7661 12288
rect 15843 12260 15936 12288
rect 7616 12248 7622 12260
rect 15930 12248 15936 12260
rect 15988 12288 15994 12300
rect 16482 12288 16488 12300
rect 15988 12260 16488 12288
rect 15988 12248 15994 12260
rect 16482 12248 16488 12260
rect 16540 12248 16546 12300
rect 17126 12288 17132 12300
rect 17087 12260 17132 12288
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 17396 12291 17454 12297
rect 17396 12257 17408 12291
rect 17442 12288 17454 12291
rect 17770 12288 17776 12300
rect 17442 12260 17776 12288
rect 17442 12257 17454 12260
rect 17396 12251 17454 12257
rect 17770 12248 17776 12260
rect 17828 12248 17834 12300
rect 19812 12288 19840 12384
rect 21542 12316 21548 12368
rect 21600 12356 21606 12368
rect 21913 12359 21971 12365
rect 21913 12356 21925 12359
rect 21600 12328 21925 12356
rect 21600 12316 21606 12328
rect 21913 12325 21925 12328
rect 21959 12325 21971 12359
rect 23842 12356 23848 12368
rect 21913 12319 21971 12325
rect 23400 12328 23848 12356
rect 22186 12288 22192 12300
rect 19812 12260 22192 12288
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12220 3111 12223
rect 3510 12220 3516 12232
rect 3099 12192 3516 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 3510 12180 3516 12192
rect 3568 12180 3574 12232
rect 5902 12220 5908 12232
rect 5863 12192 5908 12220
rect 5902 12180 5908 12192
rect 5960 12180 5966 12232
rect 6089 12223 6147 12229
rect 6089 12189 6101 12223
rect 6135 12220 6147 12223
rect 6135 12192 6592 12220
rect 6135 12189 6147 12192
rect 6089 12183 6147 12189
rect 5074 12112 5080 12164
rect 5132 12152 5138 12164
rect 5261 12155 5319 12161
rect 5261 12152 5273 12155
rect 5132 12124 5273 12152
rect 5132 12112 5138 12124
rect 5261 12121 5273 12124
rect 5307 12152 5319 12155
rect 6104 12152 6132 12183
rect 6564 12164 6592 12192
rect 7650 12180 7656 12232
rect 7708 12220 7714 12232
rect 10594 12220 10600 12232
rect 7708 12192 7753 12220
rect 10555 12192 10600 12220
rect 7708 12180 7714 12192
rect 10594 12180 10600 12192
rect 10652 12180 10658 12232
rect 16209 12223 16267 12229
rect 16209 12189 16221 12223
rect 16255 12220 16267 12223
rect 16666 12220 16672 12232
rect 16255 12192 16672 12220
rect 16255 12189 16267 12192
rect 16209 12183 16267 12189
rect 16666 12180 16672 12192
rect 16724 12220 16730 12232
rect 16942 12220 16948 12232
rect 16724 12192 16948 12220
rect 16724 12180 16730 12192
rect 16942 12180 16948 12192
rect 17000 12180 17006 12232
rect 21928 12220 21956 12260
rect 22186 12248 22192 12260
rect 22244 12288 22250 12300
rect 23109 12291 23167 12297
rect 23109 12288 23121 12291
rect 22244 12260 23121 12288
rect 22244 12248 22250 12260
rect 23109 12257 23121 12260
rect 23155 12257 23167 12291
rect 23109 12251 23167 12257
rect 23400 12232 23428 12328
rect 23842 12316 23848 12328
rect 23900 12356 23906 12368
rect 26142 12356 26148 12368
rect 23900 12328 26148 12356
rect 23900 12316 23906 12328
rect 26142 12316 26148 12328
rect 26200 12316 26206 12368
rect 23474 12248 23480 12300
rect 23532 12288 23538 12300
rect 23641 12291 23699 12297
rect 23641 12288 23653 12291
rect 23532 12260 23653 12288
rect 23532 12248 23538 12260
rect 23641 12257 23653 12260
rect 23687 12288 23699 12291
rect 24394 12288 24400 12300
rect 23687 12260 24400 12288
rect 23687 12257 23699 12260
rect 23641 12251 23699 12257
rect 24394 12248 24400 12260
rect 24452 12288 24458 12300
rect 25314 12288 25320 12300
rect 24452 12260 25320 12288
rect 24452 12248 24458 12260
rect 25314 12248 25320 12260
rect 25372 12248 25378 12300
rect 25590 12248 25596 12300
rect 25648 12288 25654 12300
rect 26510 12288 26516 12300
rect 25648 12260 26516 12288
rect 25648 12248 25654 12260
rect 26510 12248 26516 12260
rect 26568 12288 26574 12300
rect 26881 12291 26939 12297
rect 26881 12288 26893 12291
rect 26568 12260 26893 12288
rect 26568 12248 26574 12260
rect 26881 12257 26893 12260
rect 26927 12257 26939 12291
rect 26881 12251 26939 12257
rect 22005 12223 22063 12229
rect 22005 12220 22017 12223
rect 21928 12192 22017 12220
rect 22005 12189 22017 12192
rect 22051 12189 22063 12223
rect 23382 12220 23388 12232
rect 23343 12192 23388 12220
rect 22005 12183 22063 12189
rect 23382 12180 23388 12192
rect 23440 12180 23446 12232
rect 27154 12220 27160 12232
rect 27115 12192 27160 12220
rect 27154 12180 27160 12192
rect 27212 12180 27218 12232
rect 5307 12124 6132 12152
rect 5307 12121 5319 12124
rect 5261 12115 5319 12121
rect 6546 12112 6552 12164
rect 6604 12152 6610 12164
rect 6641 12155 6699 12161
rect 6641 12152 6653 12155
rect 6604 12124 6653 12152
rect 6604 12112 6610 12124
rect 6641 12121 6653 12124
rect 6687 12152 6699 12155
rect 7668 12152 7696 12180
rect 6687 12124 7696 12152
rect 20717 12155 20775 12161
rect 6687 12121 6699 12124
rect 6641 12115 6699 12121
rect 20717 12121 20729 12155
rect 20763 12152 20775 12155
rect 21453 12155 21511 12161
rect 21453 12152 21465 12155
rect 20763 12124 21465 12152
rect 20763 12121 20775 12124
rect 20717 12115 20775 12121
rect 21453 12121 21465 12124
rect 21499 12152 21511 12155
rect 21634 12152 21640 12164
rect 21499 12124 21640 12152
rect 21499 12121 21511 12124
rect 21453 12115 21511 12121
rect 21634 12112 21640 12124
rect 21692 12112 21698 12164
rect 3878 12084 3884 12096
rect 2792 12056 3884 12084
rect 3878 12044 3884 12056
rect 3936 12044 3942 12096
rect 4246 12084 4252 12096
rect 4207 12056 4252 12084
rect 4246 12044 4252 12056
rect 4304 12044 4310 12096
rect 4614 12084 4620 12096
rect 4575 12056 4620 12084
rect 4614 12044 4620 12056
rect 4672 12044 4678 12096
rect 5445 12087 5503 12093
rect 5445 12053 5457 12087
rect 5491 12084 5503 12087
rect 5534 12084 5540 12096
rect 5491 12056 5540 12084
rect 5491 12053 5503 12056
rect 5445 12047 5503 12053
rect 5534 12044 5540 12056
rect 5592 12044 5598 12096
rect 8110 12084 8116 12096
rect 8071 12056 8116 12084
rect 8110 12044 8116 12056
rect 8168 12044 8174 12096
rect 10226 12084 10232 12096
rect 10187 12056 10232 12084
rect 10226 12044 10232 12056
rect 10284 12044 10290 12096
rect 20073 12087 20131 12093
rect 20073 12053 20085 12087
rect 20119 12084 20131 12087
rect 20162 12084 20168 12096
rect 20119 12056 20168 12084
rect 20119 12053 20131 12056
rect 20073 12047 20131 12053
rect 20162 12044 20168 12056
rect 20220 12044 20226 12096
rect 24765 12087 24823 12093
rect 24765 12053 24777 12087
rect 24811 12084 24823 12087
rect 24946 12084 24952 12096
rect 24811 12056 24952 12084
rect 24811 12053 24823 12056
rect 24765 12047 24823 12053
rect 24946 12044 24952 12056
rect 25004 12044 25010 12096
rect 25777 12087 25835 12093
rect 25777 12053 25789 12087
rect 25823 12084 25835 12087
rect 25866 12084 25872 12096
rect 25823 12056 25872 12084
rect 25823 12053 25835 12056
rect 25777 12047 25835 12053
rect 25866 12044 25872 12056
rect 25924 12084 25930 12096
rect 26513 12087 26571 12093
rect 26513 12084 26525 12087
rect 25924 12056 26525 12084
rect 25924 12044 25930 12056
rect 26513 12053 26525 12056
rect 26559 12053 26571 12087
rect 26513 12047 26571 12053
rect 1104 11994 28888 12016
rect 1104 11942 5982 11994
rect 6034 11942 6046 11994
rect 6098 11942 6110 11994
rect 6162 11942 6174 11994
rect 6226 11942 15982 11994
rect 16034 11942 16046 11994
rect 16098 11942 16110 11994
rect 16162 11942 16174 11994
rect 16226 11942 25982 11994
rect 26034 11942 26046 11994
rect 26098 11942 26110 11994
rect 26162 11942 26174 11994
rect 26226 11942 28888 11994
rect 1104 11920 28888 11942
rect 1673 11883 1731 11889
rect 1673 11849 1685 11883
rect 1719 11880 1731 11883
rect 2498 11880 2504 11892
rect 1719 11852 2504 11880
rect 1719 11849 1731 11852
rect 1673 11843 1731 11849
rect 2498 11840 2504 11852
rect 2556 11840 2562 11892
rect 4154 11880 4160 11892
rect 4115 11852 4160 11880
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 5074 11880 5080 11892
rect 5035 11852 5080 11880
rect 5074 11840 5080 11852
rect 5132 11840 5138 11892
rect 6273 11883 6331 11889
rect 6273 11849 6285 11883
rect 6319 11880 6331 11883
rect 6362 11880 6368 11892
rect 6319 11852 6368 11880
rect 6319 11849 6331 11852
rect 6273 11843 6331 11849
rect 6362 11840 6368 11852
rect 6420 11840 6426 11892
rect 6638 11880 6644 11892
rect 6599 11852 6644 11880
rect 6638 11840 6644 11852
rect 6696 11840 6702 11892
rect 7558 11840 7564 11892
rect 7616 11880 7622 11892
rect 7837 11883 7895 11889
rect 7837 11880 7849 11883
rect 7616 11852 7849 11880
rect 7616 11840 7622 11852
rect 7837 11849 7849 11852
rect 7883 11849 7895 11883
rect 7837 11843 7895 11849
rect 8389 11883 8447 11889
rect 8389 11849 8401 11883
rect 8435 11880 8447 11883
rect 9214 11880 9220 11892
rect 8435 11852 9220 11880
rect 8435 11849 8447 11852
rect 8389 11843 8447 11849
rect 9214 11840 9220 11852
rect 9272 11840 9278 11892
rect 9398 11880 9404 11892
rect 9359 11852 9404 11880
rect 9398 11840 9404 11852
rect 9456 11840 9462 11892
rect 10042 11880 10048 11892
rect 10003 11852 10048 11880
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 10594 11840 10600 11892
rect 10652 11880 10658 11892
rect 11149 11883 11207 11889
rect 11149 11880 11161 11883
rect 10652 11852 11161 11880
rect 10652 11840 10658 11852
rect 11149 11849 11161 11852
rect 11195 11880 11207 11883
rect 11882 11880 11888 11892
rect 11195 11852 11888 11880
rect 11195 11849 11207 11852
rect 11149 11843 11207 11849
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 15289 11883 15347 11889
rect 15289 11849 15301 11883
rect 15335 11880 15347 11883
rect 15378 11880 15384 11892
rect 15335 11852 15384 11880
rect 15335 11849 15347 11852
rect 15289 11843 15347 11849
rect 15378 11840 15384 11852
rect 15436 11840 15442 11892
rect 15838 11840 15844 11892
rect 15896 11880 15902 11892
rect 15933 11883 15991 11889
rect 15933 11880 15945 11883
rect 15896 11852 15945 11880
rect 15896 11840 15902 11852
rect 15933 11849 15945 11852
rect 15979 11849 15991 11883
rect 16390 11880 16396 11892
rect 16351 11852 16396 11880
rect 15933 11843 15991 11849
rect 16390 11840 16396 11852
rect 16448 11840 16454 11892
rect 17126 11840 17132 11892
rect 17184 11880 17190 11892
rect 17405 11883 17463 11889
rect 17405 11880 17417 11883
rect 17184 11852 17417 11880
rect 17184 11840 17190 11852
rect 17405 11849 17417 11852
rect 17451 11849 17463 11883
rect 17770 11880 17776 11892
rect 17731 11852 17776 11880
rect 17405 11843 17463 11849
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 19886 11840 19892 11892
rect 19944 11880 19950 11892
rect 21361 11883 21419 11889
rect 21361 11880 21373 11883
rect 19944 11852 21373 11880
rect 19944 11840 19950 11852
rect 21361 11849 21373 11852
rect 21407 11849 21419 11883
rect 21361 11843 21419 11849
rect 21542 11840 21548 11892
rect 21600 11880 21606 11892
rect 21913 11883 21971 11889
rect 21913 11880 21925 11883
rect 21600 11852 21925 11880
rect 21600 11840 21606 11852
rect 21913 11849 21925 11852
rect 21959 11849 21971 11883
rect 21913 11843 21971 11849
rect 23109 11883 23167 11889
rect 23109 11849 23121 11883
rect 23155 11880 23167 11883
rect 23198 11880 23204 11892
rect 23155 11852 23204 11880
rect 23155 11849 23167 11852
rect 23109 11843 23167 11849
rect 9950 11812 9956 11824
rect 9911 11784 9956 11812
rect 9950 11772 9956 11784
rect 10008 11812 10014 11824
rect 11422 11812 11428 11824
rect 10008 11784 10456 11812
rect 11383 11784 11428 11812
rect 10008 11772 10014 11784
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11744 4767 11747
rect 5721 11747 5779 11753
rect 5721 11744 5733 11747
rect 4755 11716 5733 11744
rect 4755 11713 4767 11716
rect 4709 11707 4767 11713
rect 5721 11713 5733 11716
rect 5767 11744 5779 11747
rect 7374 11744 7380 11756
rect 5767 11716 7380 11744
rect 5767 11713 5779 11716
rect 5721 11707 5779 11713
rect 7374 11704 7380 11716
rect 7432 11744 7438 11756
rect 7558 11744 7564 11756
rect 7432 11716 7564 11744
rect 7432 11704 7438 11716
rect 7558 11704 7564 11716
rect 7616 11744 7622 11756
rect 8110 11744 8116 11756
rect 7616 11716 8116 11744
rect 7616 11704 7622 11716
rect 8110 11704 8116 11716
rect 8168 11704 8174 11756
rect 8297 11747 8355 11753
rect 8297 11713 8309 11747
rect 8343 11744 8355 11747
rect 8846 11744 8852 11756
rect 8343 11716 8852 11744
rect 8343 11713 8355 11716
rect 8297 11707 8355 11713
rect 8846 11704 8852 11716
rect 8904 11744 8910 11756
rect 8941 11747 8999 11753
rect 8941 11744 8953 11747
rect 8904 11716 8953 11744
rect 8904 11704 8910 11716
rect 8941 11713 8953 11716
rect 8987 11713 8999 11747
rect 8941 11707 8999 11713
rect 2041 11679 2099 11685
rect 2041 11645 2053 11679
rect 2087 11676 2099 11679
rect 2133 11679 2191 11685
rect 2133 11676 2145 11679
rect 2087 11648 2145 11676
rect 2087 11645 2099 11648
rect 2041 11639 2099 11645
rect 2133 11645 2145 11648
rect 2179 11676 2191 11679
rect 2222 11676 2228 11688
rect 2179 11648 2228 11676
rect 2179 11645 2191 11648
rect 2133 11639 2191 11645
rect 2222 11636 2228 11648
rect 2280 11676 2286 11688
rect 2280 11648 4660 11676
rect 2280 11636 2286 11648
rect 2378 11611 2436 11617
rect 2378 11608 2390 11611
rect 2240 11580 2390 11608
rect 2240 11552 2268 11580
rect 2378 11577 2390 11580
rect 2424 11577 2436 11611
rect 4632 11608 4660 11648
rect 7098 11636 7104 11688
rect 7156 11676 7162 11688
rect 7193 11679 7251 11685
rect 7193 11676 7205 11679
rect 7156 11648 7205 11676
rect 7156 11636 7162 11648
rect 7193 11645 7205 11648
rect 7239 11645 7251 11679
rect 7193 11639 7251 11645
rect 7282 11636 7288 11688
rect 7340 11676 7346 11688
rect 10428 11685 10456 11784
rect 11422 11772 11428 11784
rect 11480 11772 11486 11824
rect 20990 11772 20996 11824
rect 21048 11812 21054 11824
rect 22373 11815 22431 11821
rect 22373 11812 22385 11815
rect 21048 11784 22385 11812
rect 21048 11772 21054 11784
rect 21376 11756 21404 11784
rect 22373 11781 22385 11784
rect 22419 11812 22431 11815
rect 22738 11812 22744 11824
rect 22419 11784 22744 11812
rect 22419 11781 22431 11784
rect 22373 11775 22431 11781
rect 22738 11772 22744 11784
rect 22796 11772 22802 11824
rect 10594 11744 10600 11756
rect 10555 11716 10600 11744
rect 10594 11704 10600 11716
rect 10652 11744 10658 11756
rect 10778 11744 10784 11756
rect 10652 11716 10784 11744
rect 10652 11704 10658 11716
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 17034 11744 17040 11756
rect 16995 11716 17040 11744
rect 17034 11704 17040 11716
rect 17092 11704 17098 11756
rect 18325 11747 18383 11753
rect 18325 11713 18337 11747
rect 18371 11744 18383 11747
rect 19061 11747 19119 11753
rect 19061 11744 19073 11747
rect 18371 11716 19073 11744
rect 18371 11713 18383 11716
rect 18325 11707 18383 11713
rect 19061 11713 19073 11716
rect 19107 11744 19119 11747
rect 19794 11744 19800 11756
rect 19107 11716 19800 11744
rect 19107 11713 19119 11716
rect 19061 11707 19119 11713
rect 19794 11704 19800 11716
rect 19852 11704 19858 11756
rect 21358 11704 21364 11756
rect 21416 11704 21422 11756
rect 10413 11679 10471 11685
rect 7340 11648 7385 11676
rect 7340 11636 7346 11648
rect 10413 11645 10425 11679
rect 10459 11645 10471 11679
rect 10413 11639 10471 11645
rect 19334 11636 19340 11688
rect 19392 11676 19398 11688
rect 19981 11679 20039 11685
rect 19981 11676 19993 11679
rect 19392 11648 19993 11676
rect 19392 11636 19398 11648
rect 4798 11608 4804 11620
rect 4632 11580 4804 11608
rect 2378 11571 2436 11577
rect 4798 11568 4804 11580
rect 4856 11608 4862 11620
rect 5258 11608 5264 11620
rect 4856 11580 5264 11608
rect 4856 11568 4862 11580
rect 5258 11568 5264 11580
rect 5316 11568 5322 11620
rect 5629 11611 5687 11617
rect 5629 11577 5641 11611
rect 5675 11608 5687 11611
rect 5718 11608 5724 11620
rect 5675 11580 5724 11608
rect 5675 11577 5687 11580
rect 5629 11571 5687 11577
rect 5718 11568 5724 11580
rect 5776 11568 5782 11620
rect 8757 11611 8815 11617
rect 8757 11608 8769 11611
rect 6840 11580 8769 11608
rect 2222 11500 2228 11552
rect 2280 11500 2286 11552
rect 3418 11500 3424 11552
rect 3476 11540 3482 11552
rect 3513 11543 3571 11549
rect 3513 11540 3525 11543
rect 3476 11512 3525 11540
rect 3476 11500 3482 11512
rect 3513 11509 3525 11512
rect 3559 11509 3571 11543
rect 5166 11540 5172 11552
rect 5127 11512 5172 11540
rect 3513 11503 3571 11509
rect 5166 11500 5172 11512
rect 5224 11500 5230 11552
rect 5534 11540 5540 11552
rect 5495 11512 5540 11540
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 6840 11549 6868 11580
rect 8757 11577 8769 11580
rect 8803 11608 8815 11611
rect 9214 11608 9220 11620
rect 8803 11580 9220 11608
rect 8803 11577 8815 11580
rect 8757 11571 8815 11577
rect 9214 11568 9220 11580
rect 9272 11568 9278 11620
rect 11790 11608 11796 11620
rect 11751 11580 11796 11608
rect 11790 11568 11796 11580
rect 11848 11568 11854 11620
rect 15657 11611 15715 11617
rect 15657 11577 15669 11611
rect 15703 11608 15715 11611
rect 16482 11608 16488 11620
rect 15703 11580 16488 11608
rect 15703 11577 15715 11580
rect 15657 11571 15715 11577
rect 16482 11568 16488 11580
rect 16540 11568 16546 11620
rect 18785 11611 18843 11617
rect 18785 11577 18797 11611
rect 18831 11608 18843 11611
rect 19242 11608 19248 11620
rect 18831 11580 19248 11608
rect 18831 11577 18843 11580
rect 18785 11571 18843 11577
rect 19242 11568 19248 11580
rect 19300 11608 19306 11620
rect 19429 11611 19487 11617
rect 19429 11608 19441 11611
rect 19300 11580 19441 11608
rect 19300 11568 19306 11580
rect 19429 11577 19441 11580
rect 19475 11577 19487 11611
rect 19429 11571 19487 11577
rect 6825 11543 6883 11549
rect 6825 11509 6837 11543
rect 6871 11509 6883 11543
rect 8846 11540 8852 11552
rect 8807 11512 8852 11540
rect 6825 11503 6883 11509
rect 8846 11500 8852 11512
rect 8904 11500 8910 11552
rect 10502 11540 10508 11552
rect 10463 11512 10508 11540
rect 10502 11500 10508 11512
rect 10560 11500 10566 11552
rect 15746 11500 15752 11552
rect 15804 11540 15810 11552
rect 16761 11543 16819 11549
rect 16761 11540 16773 11543
rect 15804 11512 16773 11540
rect 15804 11500 15810 11512
rect 16761 11509 16773 11512
rect 16807 11509 16819 11543
rect 16761 11503 16819 11509
rect 16850 11500 16856 11552
rect 16908 11540 16914 11552
rect 18414 11540 18420 11552
rect 16908 11512 16953 11540
rect 18375 11512 18420 11540
rect 16908 11500 16914 11512
rect 18414 11500 18420 11512
rect 18472 11500 18478 11552
rect 18874 11540 18880 11552
rect 18835 11512 18880 11540
rect 18874 11500 18880 11512
rect 18932 11500 18938 11552
rect 19702 11500 19708 11552
rect 19760 11540 19766 11552
rect 19812 11549 19840 11648
rect 19981 11645 19993 11648
rect 20027 11676 20039 11679
rect 22465 11679 22523 11685
rect 20027 11648 22416 11676
rect 20027 11645 20039 11648
rect 19981 11639 20039 11645
rect 20162 11568 20168 11620
rect 20220 11617 20226 11620
rect 20220 11611 20284 11617
rect 20220 11577 20238 11611
rect 20272 11577 20284 11611
rect 22388 11608 22416 11648
rect 22465 11645 22477 11679
rect 22511 11676 22523 11679
rect 23124 11676 23152 11843
rect 23198 11840 23204 11852
rect 23256 11840 23262 11892
rect 24026 11880 24032 11892
rect 23987 11852 24032 11880
rect 24026 11840 24032 11852
rect 24084 11840 24090 11892
rect 26510 11840 26516 11892
rect 26568 11880 26574 11892
rect 26605 11883 26663 11889
rect 26605 11880 26617 11883
rect 26568 11852 26617 11880
rect 26568 11840 26574 11852
rect 26605 11849 26617 11852
rect 26651 11849 26663 11883
rect 26970 11880 26976 11892
rect 26931 11852 26976 11880
rect 26605 11843 26663 11849
rect 24670 11812 24676 11824
rect 24504 11784 24676 11812
rect 24504 11753 24532 11784
rect 24670 11772 24676 11784
rect 24728 11812 24734 11824
rect 25593 11815 25651 11821
rect 25593 11812 25605 11815
rect 24728 11784 25605 11812
rect 24728 11772 24734 11784
rect 25593 11781 25605 11784
rect 25639 11781 25651 11815
rect 26620 11812 26648 11843
rect 26970 11840 26976 11852
rect 27028 11840 27034 11892
rect 27154 11840 27160 11892
rect 27212 11880 27218 11892
rect 28077 11883 28135 11889
rect 28077 11880 28089 11883
rect 27212 11852 28089 11880
rect 27212 11840 27218 11852
rect 28077 11849 28089 11852
rect 28123 11849 28135 11883
rect 28077 11843 28135 11849
rect 27062 11812 27068 11824
rect 26620 11784 27068 11812
rect 25593 11775 25651 11781
rect 27062 11772 27068 11784
rect 27120 11772 27126 11824
rect 24489 11747 24547 11753
rect 24489 11713 24501 11747
rect 24535 11713 24547 11747
rect 24489 11707 24547 11713
rect 24581 11747 24639 11753
rect 24581 11713 24593 11747
rect 24627 11713 24639 11747
rect 24581 11707 24639 11713
rect 24596 11676 24624 11707
rect 24946 11704 24952 11756
rect 25004 11744 25010 11756
rect 25501 11747 25559 11753
rect 25501 11744 25513 11747
rect 25004 11716 25513 11744
rect 25004 11704 25010 11716
rect 25501 11713 25513 11716
rect 25547 11744 25559 11747
rect 26145 11747 26203 11753
rect 26145 11744 26157 11747
rect 25547 11716 26157 11744
rect 25547 11713 25559 11716
rect 25501 11707 25559 11713
rect 26145 11713 26157 11716
rect 26191 11713 26203 11747
rect 26145 11707 26203 11713
rect 24762 11676 24768 11688
rect 22511 11648 23152 11676
rect 23860 11648 24768 11676
rect 22511 11645 22523 11648
rect 22465 11639 22523 11645
rect 23382 11608 23388 11620
rect 22388 11580 23388 11608
rect 20220 11571 20284 11577
rect 20220 11568 20226 11571
rect 23382 11568 23388 11580
rect 23440 11568 23446 11620
rect 23860 11552 23888 11648
rect 24762 11636 24768 11648
rect 24820 11636 24826 11688
rect 25866 11636 25872 11688
rect 25924 11676 25930 11688
rect 25961 11679 26019 11685
rect 25961 11676 25973 11679
rect 25924 11648 25973 11676
rect 25924 11636 25930 11648
rect 25961 11645 25973 11648
rect 26007 11645 26019 11679
rect 25961 11639 26019 11645
rect 26970 11636 26976 11688
rect 27028 11676 27034 11688
rect 27157 11679 27215 11685
rect 27157 11676 27169 11679
rect 27028 11648 27169 11676
rect 27028 11636 27034 11648
rect 27157 11645 27169 11648
rect 27203 11676 27215 11679
rect 27709 11679 27767 11685
rect 27709 11676 27721 11679
rect 27203 11648 27721 11676
rect 27203 11645 27215 11648
rect 27157 11639 27215 11645
rect 27709 11645 27721 11648
rect 27755 11645 27767 11679
rect 27709 11639 27767 11645
rect 25133 11611 25191 11617
rect 25133 11577 25145 11611
rect 25179 11608 25191 11611
rect 26053 11611 26111 11617
rect 26053 11608 26065 11611
rect 25179 11580 26065 11608
rect 25179 11577 25191 11580
rect 25133 11571 25191 11577
rect 26053 11577 26065 11580
rect 26099 11608 26111 11611
rect 26510 11608 26516 11620
rect 26099 11580 26516 11608
rect 26099 11577 26111 11580
rect 26053 11571 26111 11577
rect 26510 11568 26516 11580
rect 26568 11568 26574 11620
rect 19797 11543 19855 11549
rect 19797 11540 19809 11543
rect 19760 11512 19809 11540
rect 19760 11500 19766 11512
rect 19797 11509 19809 11512
rect 19843 11509 19855 11543
rect 22646 11540 22652 11552
rect 22607 11512 22652 11540
rect 19797 11503 19855 11509
rect 22646 11500 22652 11512
rect 22704 11500 22710 11552
rect 23842 11540 23848 11552
rect 23803 11512 23848 11540
rect 23842 11500 23848 11512
rect 23900 11500 23906 11552
rect 24397 11543 24455 11549
rect 24397 11509 24409 11543
rect 24443 11540 24455 11543
rect 24946 11540 24952 11552
rect 24443 11512 24952 11540
rect 24443 11509 24455 11512
rect 24397 11503 24455 11509
rect 24946 11500 24952 11512
rect 25004 11500 25010 11552
rect 27338 11540 27344 11552
rect 27299 11512 27344 11540
rect 27338 11500 27344 11512
rect 27396 11500 27402 11552
rect 1104 11450 28888 11472
rect 1104 11398 10982 11450
rect 11034 11398 11046 11450
rect 11098 11398 11110 11450
rect 11162 11398 11174 11450
rect 11226 11398 20982 11450
rect 21034 11398 21046 11450
rect 21098 11398 21110 11450
rect 21162 11398 21174 11450
rect 21226 11398 28888 11450
rect 1104 11376 28888 11398
rect 2409 11339 2467 11345
rect 2409 11305 2421 11339
rect 2455 11336 2467 11339
rect 2866 11336 2872 11348
rect 2455 11308 2872 11336
rect 2455 11305 2467 11308
rect 2409 11299 2467 11305
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 3510 11336 3516 11348
rect 3423 11308 3516 11336
rect 3510 11296 3516 11308
rect 3568 11336 3574 11348
rect 6825 11339 6883 11345
rect 6825 11336 6837 11339
rect 3568 11308 6837 11336
rect 3568 11296 3574 11308
rect 6825 11305 6837 11308
rect 6871 11305 6883 11339
rect 6825 11299 6883 11305
rect 7469 11339 7527 11345
rect 7469 11305 7481 11339
rect 7515 11336 7527 11339
rect 7650 11336 7656 11348
rect 7515 11308 7656 11336
rect 7515 11305 7527 11308
rect 7469 11299 7527 11305
rect 7650 11296 7656 11308
rect 7708 11296 7714 11348
rect 8386 11336 8392 11348
rect 8347 11308 8392 11336
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 9306 11336 9312 11348
rect 9267 11308 9312 11336
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 10229 11339 10287 11345
rect 10229 11305 10241 11339
rect 10275 11305 10287 11339
rect 10229 11299 10287 11305
rect 1394 11228 1400 11280
rect 1452 11268 1458 11280
rect 1673 11271 1731 11277
rect 1673 11268 1685 11271
rect 1452 11240 1685 11268
rect 1452 11228 1458 11240
rect 1673 11237 1685 11240
rect 1719 11268 1731 11271
rect 2590 11268 2596 11280
rect 1719 11240 2596 11268
rect 1719 11237 1731 11240
rect 1673 11231 1731 11237
rect 2590 11228 2596 11240
rect 2648 11228 2654 11280
rect 2774 11228 2780 11280
rect 2832 11268 2838 11280
rect 3326 11268 3332 11280
rect 2832 11240 3332 11268
rect 2832 11228 2838 11240
rect 3326 11228 3332 11240
rect 3384 11228 3390 11280
rect 5442 11228 5448 11280
rect 5500 11268 5506 11280
rect 6270 11268 6276 11280
rect 5500 11240 6276 11268
rect 5500 11228 5506 11240
rect 6270 11228 6276 11240
rect 6328 11228 6334 11280
rect 7558 11228 7564 11280
rect 7616 11268 7622 11280
rect 7745 11271 7803 11277
rect 7745 11268 7757 11271
rect 7616 11240 7757 11268
rect 7616 11228 7622 11240
rect 7745 11237 7757 11240
rect 7791 11237 7803 11271
rect 10244 11268 10272 11299
rect 10502 11296 10508 11348
rect 10560 11336 10566 11348
rect 11241 11339 11299 11345
rect 11241 11336 11253 11339
rect 10560 11308 11253 11336
rect 10560 11296 10566 11308
rect 11241 11305 11253 11308
rect 11287 11305 11299 11339
rect 11241 11299 11299 11305
rect 11330 11296 11336 11348
rect 11388 11336 11394 11348
rect 11793 11339 11851 11345
rect 11793 11336 11805 11339
rect 11388 11308 11805 11336
rect 11388 11296 11394 11308
rect 11793 11305 11805 11308
rect 11839 11305 11851 11339
rect 11793 11299 11851 11305
rect 12253 11339 12311 11345
rect 12253 11305 12265 11339
rect 12299 11336 12311 11339
rect 12342 11336 12348 11348
rect 12299 11308 12348 11336
rect 12299 11305 12311 11308
rect 12253 11299 12311 11305
rect 12342 11296 12348 11308
rect 12400 11296 12406 11348
rect 16025 11339 16083 11345
rect 16025 11305 16037 11339
rect 16071 11336 16083 11339
rect 16117 11339 16175 11345
rect 16117 11336 16129 11339
rect 16071 11308 16129 11336
rect 16071 11305 16083 11308
rect 16025 11299 16083 11305
rect 16117 11305 16129 11308
rect 16163 11336 16175 11339
rect 16850 11336 16856 11348
rect 16163 11308 16856 11336
rect 16163 11305 16175 11308
rect 16117 11299 16175 11305
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 16942 11296 16948 11348
rect 17000 11336 17006 11348
rect 17129 11339 17187 11345
rect 17129 11336 17141 11339
rect 17000 11308 17141 11336
rect 17000 11296 17006 11308
rect 17129 11305 17141 11308
rect 17175 11305 17187 11339
rect 17129 11299 17187 11305
rect 17681 11339 17739 11345
rect 17681 11305 17693 11339
rect 17727 11336 17739 11339
rect 18785 11339 18843 11345
rect 18785 11336 18797 11339
rect 17727 11308 18797 11336
rect 17727 11305 17739 11308
rect 17681 11299 17739 11305
rect 18785 11305 18797 11308
rect 18831 11336 18843 11339
rect 18874 11336 18880 11348
rect 18831 11308 18880 11336
rect 18831 11305 18843 11308
rect 18785 11299 18843 11305
rect 18874 11296 18880 11308
rect 18932 11296 18938 11348
rect 19245 11339 19303 11345
rect 19245 11305 19257 11339
rect 19291 11336 19303 11339
rect 21269 11339 21327 11345
rect 21269 11336 21281 11339
rect 19291 11308 21281 11336
rect 19291 11305 19303 11308
rect 19245 11299 19303 11305
rect 21269 11305 21281 11308
rect 21315 11336 21327 11339
rect 22186 11336 22192 11348
rect 21315 11308 22192 11336
rect 21315 11305 21327 11308
rect 21269 11299 21327 11305
rect 22186 11296 22192 11308
rect 22244 11296 22250 11348
rect 23474 11336 23480 11348
rect 23435 11308 23480 11336
rect 23474 11296 23480 11308
rect 23532 11296 23538 11348
rect 23569 11339 23627 11345
rect 23569 11305 23581 11339
rect 23615 11305 23627 11339
rect 23569 11299 23627 11305
rect 12161 11271 12219 11277
rect 12161 11268 12173 11271
rect 10244 11240 12173 11268
rect 7745 11231 7803 11237
rect 12161 11237 12173 11240
rect 12207 11268 12219 11271
rect 12526 11268 12532 11280
rect 12207 11240 12532 11268
rect 12207 11237 12219 11240
rect 12161 11231 12219 11237
rect 12526 11228 12532 11240
rect 12584 11228 12590 11280
rect 16298 11228 16304 11280
rect 16356 11268 16362 11280
rect 16485 11271 16543 11277
rect 16485 11268 16497 11271
rect 16356 11240 16497 11268
rect 16356 11228 16362 11240
rect 16485 11237 16497 11240
rect 16531 11237 16543 11271
rect 16485 11231 16543 11237
rect 19153 11271 19211 11277
rect 19153 11237 19165 11271
rect 19199 11268 19211 11271
rect 19199 11240 19748 11268
rect 19199 11237 19211 11240
rect 19153 11231 19211 11237
rect 4062 11200 4068 11212
rect 4023 11172 4068 11200
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 5718 11209 5724 11212
rect 5712 11200 5724 11209
rect 5679 11172 5724 11200
rect 5712 11163 5724 11172
rect 5718 11160 5724 11163
rect 5776 11160 5782 11212
rect 8294 11200 8300 11212
rect 8255 11172 8300 11200
rect 8294 11160 8300 11172
rect 8352 11200 8358 11212
rect 8941 11203 8999 11209
rect 8941 11200 8953 11203
rect 8352 11172 8953 11200
rect 8352 11160 8358 11172
rect 8941 11169 8953 11172
rect 8987 11169 8999 11203
rect 8941 11163 8999 11169
rect 10410 11160 10416 11212
rect 10468 11200 10474 11212
rect 10597 11203 10655 11209
rect 10597 11200 10609 11203
rect 10468 11172 10609 11200
rect 10468 11160 10474 11172
rect 10597 11169 10609 11172
rect 10643 11169 10655 11203
rect 10597 11163 10655 11169
rect 15470 11160 15476 11212
rect 15528 11200 15534 11212
rect 16577 11203 16635 11209
rect 16577 11200 16589 11203
rect 15528 11172 16589 11200
rect 15528 11160 15534 11172
rect 16577 11169 16589 11172
rect 16623 11169 16635 11203
rect 16577 11163 16635 11169
rect 17678 11160 17684 11212
rect 17736 11200 17742 11212
rect 19720 11209 19748 11240
rect 20806 11228 20812 11280
rect 20864 11268 20870 11280
rect 21361 11271 21419 11277
rect 21361 11268 21373 11271
rect 20864 11240 21373 11268
rect 20864 11228 20870 11240
rect 21361 11237 21373 11240
rect 21407 11268 21419 11271
rect 22002 11268 22008 11280
rect 21407 11240 22008 11268
rect 21407 11237 21419 11240
rect 21361 11231 21419 11237
rect 22002 11228 22008 11240
rect 22060 11228 22066 11280
rect 23584 11268 23612 11299
rect 23750 11296 23756 11348
rect 23808 11336 23814 11348
rect 24029 11339 24087 11345
rect 24029 11336 24041 11339
rect 23808 11308 24041 11336
rect 23808 11296 23814 11308
rect 24029 11305 24041 11308
rect 24075 11305 24087 11339
rect 24670 11336 24676 11348
rect 24631 11308 24676 11336
rect 24029 11299 24087 11305
rect 24670 11296 24676 11308
rect 24728 11296 24734 11348
rect 24946 11336 24952 11348
rect 24907 11308 24952 11336
rect 24946 11296 24952 11308
rect 25004 11296 25010 11348
rect 26326 11336 26332 11348
rect 26287 11308 26332 11336
rect 26326 11296 26332 11308
rect 26384 11296 26390 11348
rect 26510 11336 26516 11348
rect 26471 11308 26516 11336
rect 26510 11296 26516 11308
rect 26568 11296 26574 11348
rect 24964 11268 24992 11296
rect 23584 11240 24992 11268
rect 26344 11268 26372 11296
rect 26973 11271 27031 11277
rect 26973 11268 26985 11271
rect 26344 11240 26985 11268
rect 26973 11237 26985 11240
rect 27019 11237 27031 11271
rect 26973 11231 27031 11237
rect 18049 11203 18107 11209
rect 18049 11200 18061 11203
rect 17736 11172 18061 11200
rect 17736 11160 17742 11172
rect 18049 11169 18061 11172
rect 18095 11169 18107 11203
rect 18049 11163 18107 11169
rect 19613 11203 19671 11209
rect 19613 11169 19625 11203
rect 19659 11169 19671 11203
rect 19613 11163 19671 11169
rect 19705 11203 19763 11209
rect 19705 11169 19717 11203
rect 19751 11200 19763 11203
rect 19751 11172 19932 11200
rect 19751 11169 19763 11172
rect 19705 11163 19763 11169
rect 2866 11132 2872 11144
rect 2827 11104 2872 11132
rect 2866 11092 2872 11104
rect 2924 11092 2930 11144
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11101 3019 11135
rect 5445 11135 5503 11141
rect 5445 11132 5457 11135
rect 2961 11095 3019 11101
rect 4816 11104 5457 11132
rect 2222 10996 2228 11008
rect 2183 10968 2228 10996
rect 2222 10956 2228 10968
rect 2280 10956 2286 11008
rect 2314 10956 2320 11008
rect 2372 10996 2378 11008
rect 2976 10996 3004 11095
rect 3881 11067 3939 11073
rect 3881 11033 3893 11067
rect 3927 11064 3939 11067
rect 3927 11036 4016 11064
rect 3927 11033 3939 11036
rect 3881 11027 3939 11033
rect 2372 10968 3004 10996
rect 3988 10996 4016 11036
rect 4062 11024 4068 11076
rect 4120 11064 4126 11076
rect 4249 11067 4307 11073
rect 4249 11064 4261 11067
rect 4120 11036 4261 11064
rect 4120 11024 4126 11036
rect 4249 11033 4261 11036
rect 4295 11033 4307 11067
rect 4249 11027 4307 11033
rect 4816 11008 4844 11104
rect 5445 11101 5457 11104
rect 5491 11101 5503 11135
rect 5445 11095 5503 11101
rect 8481 11135 8539 11141
rect 8481 11101 8493 11135
rect 8527 11101 8539 11135
rect 10686 11132 10692 11144
rect 10647 11104 10692 11132
rect 8481 11095 8539 11101
rect 7926 11064 7932 11076
rect 7887 11036 7932 11064
rect 7926 11024 7932 11036
rect 7984 11024 7990 11076
rect 8294 11024 8300 11076
rect 8352 11064 8358 11076
rect 8496 11064 8524 11095
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 10870 11132 10876 11144
rect 10831 11104 10876 11132
rect 10870 11092 10876 11104
rect 10928 11092 10934 11144
rect 12345 11135 12403 11141
rect 12345 11101 12357 11135
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 16761 11135 16819 11141
rect 16761 11101 16773 11135
rect 16807 11132 16819 11135
rect 16942 11132 16948 11144
rect 16807 11104 16948 11132
rect 16807 11101 16819 11104
rect 16761 11095 16819 11101
rect 8352 11036 8524 11064
rect 10137 11067 10195 11073
rect 8352 11024 8358 11036
rect 10137 11033 10149 11067
rect 10183 11064 10195 11067
rect 10594 11064 10600 11076
rect 10183 11036 10600 11064
rect 10183 11033 10195 11036
rect 10137 11027 10195 11033
rect 10594 11024 10600 11036
rect 10652 11064 10658 11076
rect 11790 11064 11796 11076
rect 10652 11036 11796 11064
rect 10652 11024 10658 11036
rect 11790 11024 11796 11036
rect 11848 11064 11854 11076
rect 12360 11064 12388 11095
rect 16942 11092 16948 11104
rect 17000 11092 17006 11144
rect 17589 11135 17647 11141
rect 17589 11101 17601 11135
rect 17635 11132 17647 11135
rect 17954 11132 17960 11144
rect 17635 11104 17960 11132
rect 17635 11101 17647 11104
rect 17589 11095 17647 11101
rect 17954 11092 17960 11104
rect 18012 11132 18018 11144
rect 18141 11135 18199 11141
rect 18141 11132 18153 11135
rect 18012 11104 18153 11132
rect 18012 11092 18018 11104
rect 18141 11101 18153 11104
rect 18187 11101 18199 11135
rect 18141 11095 18199 11101
rect 18233 11135 18291 11141
rect 18233 11101 18245 11135
rect 18279 11101 18291 11135
rect 18233 11095 18291 11101
rect 11848 11036 12388 11064
rect 11848 11024 11854 11036
rect 18248 11008 18276 11095
rect 19628 11064 19656 11163
rect 19794 11132 19800 11144
rect 19755 11104 19800 11132
rect 19794 11092 19800 11104
rect 19852 11092 19858 11144
rect 19904 11132 19932 11172
rect 23290 11160 23296 11212
rect 23348 11200 23354 11212
rect 23937 11203 23995 11209
rect 23937 11200 23949 11203
rect 23348 11172 23949 11200
rect 23348 11160 23354 11172
rect 23937 11169 23949 11172
rect 23983 11200 23995 11203
rect 24302 11200 24308 11212
rect 23983 11172 24308 11200
rect 23983 11169 23995 11172
rect 23937 11163 23995 11169
rect 24302 11160 24308 11172
rect 24360 11160 24366 11212
rect 25130 11160 25136 11212
rect 25188 11200 25194 11212
rect 25317 11203 25375 11209
rect 25317 11200 25329 11203
rect 25188 11172 25329 11200
rect 25188 11160 25194 11172
rect 25317 11169 25329 11172
rect 25363 11200 25375 11203
rect 26881 11203 26939 11209
rect 26881 11200 26893 11203
rect 25363 11172 26893 11200
rect 25363 11169 25375 11172
rect 25317 11163 25375 11169
rect 26881 11169 26893 11172
rect 26927 11169 26939 11203
rect 26881 11163 26939 11169
rect 20806 11132 20812 11144
rect 19904 11104 20812 11132
rect 20806 11092 20812 11104
rect 20864 11092 20870 11144
rect 21545 11135 21603 11141
rect 21545 11101 21557 11135
rect 21591 11132 21603 11135
rect 21910 11132 21916 11144
rect 21591 11104 21916 11132
rect 21591 11101 21603 11104
rect 21545 11095 21603 11101
rect 21910 11092 21916 11104
rect 21968 11092 21974 11144
rect 22094 11092 22100 11144
rect 22152 11132 22158 11144
rect 22465 11135 22523 11141
rect 22465 11132 22477 11135
rect 22152 11104 22477 11132
rect 22152 11092 22158 11104
rect 22465 11101 22477 11104
rect 22511 11101 22523 11135
rect 24210 11132 24216 11144
rect 24123 11104 24216 11132
rect 22465 11095 22523 11101
rect 24210 11092 24216 11104
rect 24268 11132 24274 11144
rect 24854 11132 24860 11144
rect 24268 11104 24860 11132
rect 24268 11092 24274 11104
rect 24854 11092 24860 11104
rect 24912 11092 24918 11144
rect 27065 11135 27123 11141
rect 27065 11132 27077 11135
rect 25332 11104 27077 11132
rect 25332 11076 25360 11104
rect 27065 11101 27077 11104
rect 27111 11132 27123 11135
rect 27154 11132 27160 11144
rect 27111 11104 27160 11132
rect 27111 11101 27123 11104
rect 27065 11095 27123 11101
rect 27154 11092 27160 11104
rect 27212 11092 27218 11144
rect 20349 11067 20407 11073
rect 20349 11064 20361 11067
rect 19628 11036 20361 11064
rect 20349 11033 20361 11036
rect 20395 11064 20407 11067
rect 20622 11064 20628 11076
rect 20395 11036 20628 11064
rect 20395 11033 20407 11036
rect 20349 11027 20407 11033
rect 20622 11024 20628 11036
rect 20680 11024 20686 11076
rect 20901 11067 20959 11073
rect 20901 11033 20913 11067
rect 20947 11064 20959 11067
rect 21818 11064 21824 11076
rect 20947 11036 21824 11064
rect 20947 11033 20959 11036
rect 20901 11027 20959 11033
rect 21818 11024 21824 11036
rect 21876 11024 21882 11076
rect 22005 11067 22063 11073
rect 22005 11033 22017 11067
rect 22051 11064 22063 11067
rect 22278 11064 22284 11076
rect 22051 11036 22284 11064
rect 22051 11033 22063 11036
rect 22005 11027 22063 11033
rect 22278 11024 22284 11036
rect 22336 11024 22342 11076
rect 25314 11024 25320 11076
rect 25372 11024 25378 11076
rect 25406 11024 25412 11076
rect 25464 11064 25470 11076
rect 25501 11067 25559 11073
rect 25501 11064 25513 11067
rect 25464 11036 25513 11064
rect 25464 11024 25470 11036
rect 25501 11033 25513 11036
rect 25547 11033 25559 11067
rect 25501 11027 25559 11033
rect 4430 10996 4436 11008
rect 3988 10968 4436 10996
rect 2372 10956 2378 10968
rect 4430 10956 4436 10968
rect 4488 10956 4494 11008
rect 4709 10999 4767 11005
rect 4709 10965 4721 10999
rect 4755 10996 4767 10999
rect 4798 10996 4804 11008
rect 4755 10968 4804 10996
rect 4755 10965 4767 10968
rect 4709 10959 4767 10965
rect 4798 10956 4804 10968
rect 4856 10956 4862 11008
rect 4982 10996 4988 11008
rect 4943 10968 4988 10996
rect 4982 10956 4988 10968
rect 5040 10956 5046 11008
rect 15657 10999 15715 11005
rect 15657 10965 15669 10999
rect 15703 10996 15715 10999
rect 15746 10996 15752 11008
rect 15703 10968 15752 10996
rect 15703 10965 15715 10968
rect 15657 10959 15715 10965
rect 15746 10956 15752 10968
rect 15804 10956 15810 11008
rect 18230 10956 18236 11008
rect 18288 10956 18294 11008
rect 1104 10906 28888 10928
rect 1104 10854 5982 10906
rect 6034 10854 6046 10906
rect 6098 10854 6110 10906
rect 6162 10854 6174 10906
rect 6226 10854 15982 10906
rect 16034 10854 16046 10906
rect 16098 10854 16110 10906
rect 16162 10854 16174 10906
rect 16226 10854 25982 10906
rect 26034 10854 26046 10906
rect 26098 10854 26110 10906
rect 26162 10854 26174 10906
rect 26226 10854 28888 10906
rect 1104 10832 28888 10854
rect 2682 10792 2688 10804
rect 2643 10764 2688 10792
rect 2682 10752 2688 10764
rect 2740 10752 2746 10804
rect 3326 10752 3332 10804
rect 3384 10792 3390 10804
rect 3697 10795 3755 10801
rect 3697 10792 3709 10795
rect 3384 10764 3709 10792
rect 3384 10752 3390 10764
rect 3697 10761 3709 10764
rect 3743 10761 3755 10795
rect 4154 10792 4160 10804
rect 4067 10764 4160 10792
rect 3697 10755 3755 10761
rect 4154 10752 4160 10764
rect 4212 10792 4218 10804
rect 5350 10792 5356 10804
rect 4212 10764 5356 10792
rect 4212 10752 4218 10764
rect 5350 10752 5356 10764
rect 5408 10752 5414 10804
rect 6822 10792 6828 10804
rect 6783 10764 6828 10792
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 10229 10795 10287 10801
rect 10229 10761 10241 10795
rect 10275 10792 10287 10795
rect 10502 10792 10508 10804
rect 10275 10764 10508 10792
rect 10275 10761 10287 10764
rect 10229 10755 10287 10761
rect 10502 10752 10508 10764
rect 10560 10752 10566 10804
rect 10870 10752 10876 10804
rect 10928 10792 10934 10804
rect 11241 10795 11299 10801
rect 11241 10792 11253 10795
rect 10928 10764 11253 10792
rect 10928 10752 10934 10764
rect 11241 10761 11253 10764
rect 11287 10761 11299 10795
rect 11790 10792 11796 10804
rect 11751 10764 11796 10792
rect 11241 10755 11299 10761
rect 11790 10752 11796 10764
rect 11848 10752 11854 10804
rect 12253 10795 12311 10801
rect 12253 10761 12265 10795
rect 12299 10792 12311 10795
rect 12342 10792 12348 10804
rect 12299 10764 12348 10792
rect 12299 10761 12311 10764
rect 12253 10755 12311 10761
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 12526 10752 12532 10804
rect 12584 10792 12590 10804
rect 12621 10795 12679 10801
rect 12621 10792 12633 10795
rect 12584 10764 12633 10792
rect 12584 10752 12590 10764
rect 12621 10761 12633 10764
rect 12667 10761 12679 10795
rect 15378 10792 15384 10804
rect 15339 10764 15384 10792
rect 12621 10755 12679 10761
rect 15378 10752 15384 10764
rect 15436 10752 15442 10804
rect 15562 10752 15568 10804
rect 15620 10792 15626 10804
rect 15749 10795 15807 10801
rect 15749 10792 15761 10795
rect 15620 10764 15761 10792
rect 15620 10752 15626 10764
rect 15749 10761 15761 10764
rect 15795 10792 15807 10795
rect 16025 10795 16083 10801
rect 16025 10792 16037 10795
rect 15795 10764 16037 10792
rect 15795 10761 15807 10764
rect 15749 10755 15807 10761
rect 16025 10761 16037 10764
rect 16071 10761 16083 10795
rect 16025 10755 16083 10761
rect 16209 10795 16267 10801
rect 16209 10761 16221 10795
rect 16255 10792 16267 10795
rect 16298 10792 16304 10804
rect 16255 10764 16304 10792
rect 16255 10761 16267 10764
rect 16209 10755 16267 10761
rect 16298 10752 16304 10764
rect 16356 10752 16362 10804
rect 17954 10752 17960 10804
rect 18012 10792 18018 10804
rect 18049 10795 18107 10801
rect 18049 10792 18061 10795
rect 18012 10764 18061 10792
rect 18012 10752 18018 10764
rect 18049 10761 18061 10764
rect 18095 10761 18107 10795
rect 18049 10755 18107 10761
rect 19337 10795 19395 10801
rect 19337 10761 19349 10795
rect 19383 10792 19395 10795
rect 19794 10792 19800 10804
rect 19383 10764 19800 10792
rect 19383 10761 19395 10764
rect 19337 10755 19395 10761
rect 19794 10752 19800 10764
rect 19852 10752 19858 10804
rect 21821 10795 21879 10801
rect 21821 10761 21833 10795
rect 21867 10792 21879 10795
rect 21910 10792 21916 10804
rect 21867 10764 21916 10792
rect 21867 10761 21879 10764
rect 21821 10755 21879 10761
rect 21910 10752 21916 10764
rect 21968 10752 21974 10804
rect 22002 10752 22008 10804
rect 22060 10792 22066 10804
rect 22097 10795 22155 10801
rect 22097 10792 22109 10795
rect 22060 10764 22109 10792
rect 22060 10752 22066 10764
rect 22097 10761 22109 10764
rect 22143 10761 22155 10795
rect 22097 10755 22155 10761
rect 22186 10752 22192 10804
rect 22244 10792 22250 10804
rect 22465 10795 22523 10801
rect 22465 10792 22477 10795
rect 22244 10764 22477 10792
rect 22244 10752 22250 10764
rect 22465 10761 22477 10764
rect 22511 10761 22523 10795
rect 23382 10792 23388 10804
rect 23343 10764 23388 10792
rect 22465 10755 22523 10761
rect 23382 10752 23388 10764
rect 23440 10752 23446 10804
rect 24854 10752 24860 10804
rect 24912 10792 24918 10804
rect 25041 10795 25099 10801
rect 25041 10792 25053 10795
rect 24912 10764 25053 10792
rect 24912 10752 24918 10764
rect 25041 10761 25053 10764
rect 25087 10761 25099 10795
rect 25041 10755 25099 10761
rect 25130 10752 25136 10804
rect 25188 10792 25194 10804
rect 25593 10795 25651 10801
rect 25593 10792 25605 10795
rect 25188 10764 25605 10792
rect 25188 10752 25194 10764
rect 25593 10761 25605 10764
rect 25639 10792 25651 10795
rect 26237 10795 26295 10801
rect 26237 10792 26249 10795
rect 25639 10764 26249 10792
rect 25639 10761 25651 10764
rect 25593 10755 25651 10761
rect 26237 10761 26249 10764
rect 26283 10761 26295 10795
rect 26418 10792 26424 10804
rect 26379 10764 26424 10792
rect 26237 10755 26295 10761
rect 26418 10752 26424 10764
rect 26476 10752 26482 10804
rect 2225 10727 2283 10733
rect 2225 10693 2237 10727
rect 2271 10724 2283 10727
rect 2866 10724 2872 10736
rect 2271 10696 2872 10724
rect 2271 10693 2283 10696
rect 2225 10687 2283 10693
rect 2866 10684 2872 10696
rect 2924 10684 2930 10736
rect 9401 10727 9459 10733
rect 9401 10693 9413 10727
rect 9447 10724 9459 10727
rect 10888 10724 10916 10752
rect 9447 10696 10916 10724
rect 9447 10693 9459 10696
rect 9401 10687 9459 10693
rect 3329 10659 3387 10665
rect 3329 10656 3341 10659
rect 2240 10628 3341 10656
rect 2240 10600 2268 10628
rect 3329 10625 3341 10628
rect 3375 10656 3387 10659
rect 3510 10656 3516 10668
rect 3375 10628 3516 10656
rect 3375 10625 3387 10628
rect 3329 10619 3387 10625
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 5718 10616 5724 10668
rect 5776 10656 5782 10668
rect 7377 10659 7435 10665
rect 7377 10656 7389 10659
rect 5776 10628 7389 10656
rect 5776 10616 5782 10628
rect 7377 10625 7389 10628
rect 7423 10656 7435 10659
rect 7837 10659 7895 10665
rect 7837 10656 7849 10659
rect 7423 10628 7849 10656
rect 7423 10625 7435 10628
rect 7377 10619 7435 10625
rect 7837 10625 7849 10628
rect 7883 10625 7895 10659
rect 10045 10659 10103 10665
rect 10045 10656 10057 10659
rect 7837 10619 7895 10625
rect 8220 10628 10057 10656
rect 1394 10588 1400 10600
rect 1355 10560 1400 10588
rect 1394 10548 1400 10560
rect 1452 10548 1458 10600
rect 2222 10548 2228 10600
rect 2280 10548 2286 10600
rect 2593 10591 2651 10597
rect 2593 10557 2605 10591
rect 2639 10588 2651 10591
rect 3053 10591 3111 10597
rect 3053 10588 3065 10591
rect 2639 10560 3065 10588
rect 2639 10557 2651 10560
rect 2593 10551 2651 10557
rect 3053 10557 3065 10560
rect 3099 10588 3111 10591
rect 3142 10588 3148 10600
rect 3099 10560 3148 10588
rect 3099 10557 3111 10560
rect 3053 10551 3111 10557
rect 3142 10548 3148 10560
rect 3200 10548 3206 10600
rect 4246 10588 4252 10600
rect 4207 10560 4252 10588
rect 4246 10548 4252 10560
rect 4304 10548 4310 10600
rect 4522 10597 4528 10600
rect 4516 10588 4528 10597
rect 4435 10560 4528 10588
rect 4516 10551 4528 10560
rect 4580 10588 4586 10600
rect 4982 10588 4988 10600
rect 4580 10560 4988 10588
rect 4522 10548 4528 10551
rect 4580 10548 4586 10560
rect 4982 10548 4988 10560
rect 5040 10548 5046 10600
rect 6641 10591 6699 10597
rect 6641 10557 6653 10591
rect 6687 10588 6699 10591
rect 7285 10591 7343 10597
rect 7285 10588 7297 10591
rect 6687 10560 7297 10588
rect 6687 10557 6699 10560
rect 6641 10551 6699 10557
rect 7285 10557 7297 10560
rect 7331 10588 7343 10591
rect 8220 10588 8248 10628
rect 10045 10625 10057 10628
rect 10091 10656 10103 10659
rect 10686 10656 10692 10668
rect 10091 10628 10692 10656
rect 10091 10625 10103 10628
rect 10045 10619 10103 10625
rect 10686 10616 10692 10628
rect 10744 10616 10750 10668
rect 10888 10665 10916 10696
rect 15838 10684 15844 10736
rect 15896 10724 15902 10736
rect 16393 10727 16451 10733
rect 16393 10724 16405 10727
rect 15896 10696 16405 10724
rect 15896 10684 15902 10696
rect 16393 10693 16405 10696
rect 16439 10693 16451 10727
rect 16393 10687 16451 10693
rect 17865 10727 17923 10733
rect 17865 10693 17877 10727
rect 17911 10724 17923 10727
rect 18138 10724 18144 10736
rect 17911 10696 18144 10724
rect 17911 10693 17923 10696
rect 17865 10687 17923 10693
rect 18138 10684 18144 10696
rect 18196 10684 18202 10736
rect 27433 10727 27491 10733
rect 27433 10724 27445 10727
rect 26896 10696 27445 10724
rect 26896 10668 26924 10696
rect 27433 10693 27445 10696
rect 27479 10693 27491 10727
rect 27433 10687 27491 10693
rect 10873 10659 10931 10665
rect 10873 10625 10885 10659
rect 10919 10625 10931 10659
rect 16942 10656 16948 10668
rect 16903 10628 16948 10656
rect 10873 10619 10931 10625
rect 16942 10616 16948 10628
rect 17000 10616 17006 10668
rect 18322 10616 18328 10668
rect 18380 10656 18386 10668
rect 18601 10659 18659 10665
rect 18601 10656 18613 10659
rect 18380 10628 18613 10656
rect 18380 10616 18386 10628
rect 18601 10625 18613 10628
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 23109 10659 23167 10665
rect 23109 10625 23121 10659
rect 23155 10656 23167 10659
rect 26878 10656 26884 10668
rect 23155 10628 23796 10656
rect 26839 10628 26884 10656
rect 23155 10625 23167 10628
rect 23109 10619 23167 10625
rect 8386 10588 8392 10600
rect 7331 10560 8248 10588
rect 8299 10560 8392 10588
rect 7331 10557 7343 10560
rect 7285 10551 7343 10557
rect 8386 10548 8392 10560
rect 8444 10588 8450 10600
rect 9033 10591 9091 10597
rect 9033 10588 9045 10591
rect 8444 10560 9045 10588
rect 8444 10548 8450 10560
rect 9033 10557 9045 10560
rect 9079 10588 9091 10591
rect 10594 10588 10600 10600
rect 9079 10560 10600 10588
rect 9079 10557 9091 10560
rect 9033 10551 9091 10557
rect 10594 10548 10600 10560
rect 10652 10548 10658 10600
rect 10704 10588 10732 10616
rect 17405 10591 17463 10597
rect 17405 10588 17417 10591
rect 10704 10560 17417 10588
rect 17405 10557 17417 10560
rect 17451 10588 17463 10591
rect 17586 10588 17592 10600
rect 17451 10560 17592 10588
rect 17451 10557 17463 10560
rect 17405 10551 17463 10557
rect 17586 10548 17592 10560
rect 17644 10548 17650 10600
rect 18417 10591 18475 10597
rect 18417 10557 18429 10591
rect 18463 10588 18475 10591
rect 18690 10588 18696 10600
rect 18463 10560 18696 10588
rect 18463 10557 18475 10560
rect 18417 10551 18475 10557
rect 18690 10548 18696 10560
rect 18748 10548 18754 10600
rect 19702 10548 19708 10600
rect 19760 10588 19766 10600
rect 20070 10597 20076 10600
rect 19797 10591 19855 10597
rect 19797 10588 19809 10591
rect 19760 10560 19809 10588
rect 19760 10548 19766 10560
rect 19797 10557 19809 10560
rect 19843 10557 19855 10591
rect 20064 10588 20076 10597
rect 20031 10560 20076 10588
rect 19797 10551 19855 10557
rect 20064 10551 20076 10560
rect 20070 10548 20076 10551
rect 20128 10548 20134 10600
rect 23382 10548 23388 10600
rect 23440 10588 23446 10600
rect 23661 10591 23719 10597
rect 23661 10588 23673 10591
rect 23440 10560 23673 10588
rect 23440 10548 23446 10560
rect 23661 10557 23673 10560
rect 23707 10557 23719 10591
rect 23768 10588 23796 10628
rect 26878 10616 26884 10628
rect 26936 10616 26942 10668
rect 27065 10659 27123 10665
rect 27065 10625 27077 10659
rect 27111 10656 27123 10659
rect 27154 10656 27160 10668
rect 27111 10628 27160 10656
rect 27111 10625 27123 10628
rect 27065 10619 27123 10625
rect 27154 10616 27160 10628
rect 27212 10656 27218 10668
rect 27522 10656 27528 10668
rect 27212 10628 27528 10656
rect 27212 10616 27218 10628
rect 27522 10616 27528 10628
rect 27580 10656 27586 10668
rect 28169 10659 28227 10665
rect 28169 10656 28181 10659
rect 27580 10628 28181 10656
rect 27580 10616 27586 10628
rect 28169 10625 28181 10628
rect 28215 10625 28227 10659
rect 28169 10619 28227 10625
rect 23934 10597 23940 10600
rect 23928 10588 23940 10597
rect 23768 10560 23940 10588
rect 23661 10551 23719 10557
rect 23928 10551 23940 10560
rect 23992 10588 23998 10600
rect 24210 10588 24216 10600
rect 23992 10560 24216 10588
rect 2314 10480 2320 10532
rect 2372 10520 2378 10532
rect 5074 10520 5080 10532
rect 2372 10492 5080 10520
rect 2372 10480 2378 10492
rect 5074 10480 5080 10492
rect 5132 10520 5138 10532
rect 5718 10520 5724 10532
rect 5132 10492 5724 10520
rect 5132 10480 5138 10492
rect 1581 10455 1639 10461
rect 1581 10421 1593 10455
rect 1627 10452 1639 10455
rect 1854 10452 1860 10464
rect 1627 10424 1860 10452
rect 1627 10421 1639 10424
rect 1581 10415 1639 10421
rect 1854 10412 1860 10424
rect 1912 10412 1918 10464
rect 3142 10452 3148 10464
rect 3103 10424 3148 10452
rect 3142 10412 3148 10424
rect 3200 10412 3206 10464
rect 4246 10412 4252 10464
rect 4304 10452 4310 10464
rect 4798 10452 4804 10464
rect 4304 10424 4804 10452
rect 4304 10412 4310 10424
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 5644 10461 5672 10492
rect 5718 10480 5724 10492
rect 5776 10480 5782 10532
rect 7190 10520 7196 10532
rect 7103 10492 7196 10520
rect 7190 10480 7196 10492
rect 7248 10520 7254 10532
rect 9769 10523 9827 10529
rect 9769 10520 9781 10523
rect 7248 10492 9781 10520
rect 7248 10480 7254 10492
rect 9769 10489 9781 10492
rect 9815 10520 9827 10523
rect 10410 10520 10416 10532
rect 9815 10492 10416 10520
rect 9815 10489 9827 10492
rect 9769 10483 9827 10489
rect 10410 10480 10416 10492
rect 10468 10480 10474 10532
rect 16666 10480 16672 10532
rect 16724 10520 16730 10532
rect 16761 10523 16819 10529
rect 16761 10520 16773 10523
rect 16724 10492 16773 10520
rect 16724 10480 16730 10492
rect 16761 10489 16773 10492
rect 16807 10489 16819 10523
rect 16761 10483 16819 10489
rect 18138 10480 18144 10532
rect 18196 10520 18202 10532
rect 18509 10523 18567 10529
rect 18509 10520 18521 10523
rect 18196 10492 18521 10520
rect 18196 10480 18202 10492
rect 18509 10489 18521 10492
rect 18555 10489 18567 10523
rect 18509 10483 18567 10489
rect 19150 10480 19156 10532
rect 19208 10520 19214 10532
rect 23676 10520 23704 10551
rect 23934 10548 23940 10551
rect 23992 10548 23998 10560
rect 24210 10548 24216 10560
rect 24268 10548 24274 10600
rect 26786 10588 26792 10600
rect 26747 10560 26792 10588
rect 26786 10548 26792 10560
rect 26844 10588 26850 10600
rect 27801 10591 27859 10597
rect 27801 10588 27813 10591
rect 26844 10560 27813 10588
rect 26844 10548 26850 10560
rect 27801 10557 27813 10560
rect 27847 10557 27859 10591
rect 27801 10551 27859 10557
rect 24854 10520 24860 10532
rect 19208 10492 21220 10520
rect 23676 10492 24860 10520
rect 19208 10480 19214 10492
rect 5629 10455 5687 10461
rect 5629 10421 5641 10455
rect 5675 10421 5687 10455
rect 6178 10452 6184 10464
rect 6139 10424 6184 10452
rect 5629 10415 5687 10421
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 8294 10452 8300 10464
rect 8255 10424 8300 10452
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 8573 10455 8631 10461
rect 8573 10421 8585 10455
rect 8619 10452 8631 10455
rect 8662 10452 8668 10464
rect 8619 10424 8668 10452
rect 8619 10421 8631 10424
rect 8573 10415 8631 10421
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 10318 10412 10324 10464
rect 10376 10452 10382 10464
rect 10689 10455 10747 10461
rect 10689 10452 10701 10455
rect 10376 10424 10701 10452
rect 10376 10412 10382 10424
rect 10689 10421 10701 10424
rect 10735 10421 10747 10455
rect 10689 10415 10747 10421
rect 16025 10455 16083 10461
rect 16025 10421 16037 10455
rect 16071 10452 16083 10455
rect 16853 10455 16911 10461
rect 16853 10452 16865 10455
rect 16071 10424 16865 10452
rect 16071 10421 16083 10424
rect 16025 10415 16083 10421
rect 16853 10421 16865 10424
rect 16899 10421 16911 10455
rect 19702 10452 19708 10464
rect 19663 10424 19708 10452
rect 16853 10415 16911 10421
rect 19702 10412 19708 10424
rect 19760 10412 19766 10464
rect 21192 10461 21220 10492
rect 24854 10480 24860 10492
rect 24912 10480 24918 10532
rect 21177 10455 21235 10461
rect 21177 10421 21189 10455
rect 21223 10421 21235 10455
rect 21177 10415 21235 10421
rect 1104 10362 28888 10384
rect 1104 10310 10982 10362
rect 11034 10310 11046 10362
rect 11098 10310 11110 10362
rect 11162 10310 11174 10362
rect 11226 10310 20982 10362
rect 21034 10310 21046 10362
rect 21098 10310 21110 10362
rect 21162 10310 21174 10362
rect 21226 10310 28888 10362
rect 1104 10288 28888 10310
rect 1946 10248 1952 10260
rect 1907 10220 1952 10248
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 2314 10248 2320 10260
rect 2275 10220 2320 10248
rect 2314 10208 2320 10220
rect 2372 10208 2378 10260
rect 2406 10208 2412 10260
rect 2464 10248 2470 10260
rect 3510 10248 3516 10260
rect 2464 10220 3280 10248
rect 3471 10220 3516 10248
rect 2464 10208 2470 10220
rect 1397 10183 1455 10189
rect 1397 10149 1409 10183
rect 1443 10180 1455 10183
rect 2866 10180 2872 10192
rect 1443 10152 2872 10180
rect 1443 10149 1455 10152
rect 1397 10143 1455 10149
rect 2866 10140 2872 10152
rect 2924 10140 2930 10192
rect 3252 10189 3280 10220
rect 3510 10208 3516 10220
rect 3568 10208 3574 10260
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 4430 10248 4436 10260
rect 4120 10220 4436 10248
rect 4120 10208 4126 10220
rect 4430 10208 4436 10220
rect 4488 10208 4494 10260
rect 5074 10248 5080 10260
rect 5035 10220 5080 10248
rect 5074 10208 5080 10220
rect 5132 10248 5138 10260
rect 5445 10251 5503 10257
rect 5445 10248 5457 10251
rect 5132 10220 5457 10248
rect 5132 10208 5138 10220
rect 5445 10217 5457 10220
rect 5491 10217 5503 10251
rect 5626 10248 5632 10260
rect 5587 10220 5632 10248
rect 5445 10211 5503 10217
rect 3237 10183 3295 10189
rect 3237 10149 3249 10183
rect 3283 10180 3295 10183
rect 4522 10180 4528 10192
rect 3283 10152 4528 10180
rect 3283 10149 3295 10152
rect 3237 10143 3295 10149
rect 4522 10140 4528 10152
rect 4580 10140 4586 10192
rect 2777 10115 2835 10121
rect 2777 10081 2789 10115
rect 2823 10112 2835 10115
rect 3050 10112 3056 10124
rect 2823 10084 3056 10112
rect 2823 10081 2835 10084
rect 2777 10075 2835 10081
rect 3050 10072 3056 10084
rect 3108 10112 3114 10124
rect 3970 10112 3976 10124
rect 3108 10084 3976 10112
rect 3108 10072 3114 10084
rect 3970 10072 3976 10084
rect 4028 10072 4034 10124
rect 5460 10112 5488 10211
rect 5626 10208 5632 10220
rect 5684 10208 5690 10260
rect 5718 10208 5724 10260
rect 5776 10248 5782 10260
rect 5994 10248 6000 10260
rect 5776 10220 6000 10248
rect 5776 10208 5782 10220
rect 5994 10208 6000 10220
rect 6052 10208 6058 10260
rect 6546 10208 6552 10260
rect 6604 10248 6610 10260
rect 6917 10251 6975 10257
rect 6917 10248 6929 10251
rect 6604 10220 6929 10248
rect 6604 10208 6610 10220
rect 6917 10217 6929 10220
rect 6963 10248 6975 10251
rect 7190 10248 7196 10260
rect 6963 10220 7196 10248
rect 6963 10217 6975 10220
rect 6917 10211 6975 10217
rect 7190 10208 7196 10220
rect 7248 10208 7254 10260
rect 8478 10208 8484 10260
rect 8536 10248 8542 10260
rect 8941 10251 8999 10257
rect 8941 10248 8953 10251
rect 8536 10220 8953 10248
rect 8536 10208 8542 10220
rect 8941 10217 8953 10220
rect 8987 10217 8999 10251
rect 8941 10211 8999 10217
rect 9214 10208 9220 10260
rect 9272 10248 9278 10260
rect 9309 10251 9367 10257
rect 9309 10248 9321 10251
rect 9272 10220 9321 10248
rect 9272 10208 9278 10220
rect 9309 10217 9321 10220
rect 9355 10217 9367 10251
rect 10594 10248 10600 10260
rect 10555 10220 10600 10248
rect 9309 10211 9367 10217
rect 10594 10208 10600 10220
rect 10652 10208 10658 10260
rect 15470 10208 15476 10260
rect 15528 10248 15534 10260
rect 16025 10251 16083 10257
rect 16025 10248 16037 10251
rect 15528 10220 16037 10248
rect 15528 10208 15534 10220
rect 16025 10217 16037 10220
rect 16071 10217 16083 10251
rect 16025 10211 16083 10217
rect 16485 10251 16543 10257
rect 16485 10217 16497 10251
rect 16531 10248 16543 10251
rect 16666 10248 16672 10260
rect 16531 10220 16672 10248
rect 16531 10217 16543 10220
rect 16485 10211 16543 10217
rect 16666 10208 16672 10220
rect 16724 10208 16730 10260
rect 17126 10248 17132 10260
rect 17087 10220 17132 10248
rect 17126 10208 17132 10220
rect 17184 10208 17190 10260
rect 18322 10208 18328 10260
rect 18380 10248 18386 10260
rect 18417 10251 18475 10257
rect 18417 10248 18429 10251
rect 18380 10220 18429 10248
rect 18380 10208 18386 10220
rect 18417 10217 18429 10220
rect 18463 10217 18475 10251
rect 19242 10248 19248 10260
rect 19203 10220 19248 10248
rect 18417 10211 18475 10217
rect 19242 10208 19248 10220
rect 19300 10208 19306 10260
rect 20070 10208 20076 10260
rect 20128 10248 20134 10260
rect 20257 10251 20315 10257
rect 20257 10248 20269 10251
rect 20128 10220 20269 10248
rect 20128 10208 20134 10220
rect 20257 10217 20269 10220
rect 20303 10217 20315 10251
rect 20257 10211 20315 10217
rect 20622 10208 20628 10260
rect 20680 10248 20686 10260
rect 20901 10251 20959 10257
rect 20901 10248 20913 10251
rect 20680 10220 20913 10248
rect 20680 10208 20686 10220
rect 20901 10217 20913 10220
rect 20947 10217 20959 10251
rect 20901 10211 20959 10217
rect 21269 10251 21327 10257
rect 21269 10217 21281 10251
rect 21315 10248 21327 10251
rect 22002 10248 22008 10260
rect 21315 10220 22008 10248
rect 21315 10217 21327 10220
rect 21269 10211 21327 10217
rect 22002 10208 22008 10220
rect 22060 10208 22066 10260
rect 23750 10208 23756 10260
rect 23808 10248 23814 10260
rect 24029 10251 24087 10257
rect 24029 10248 24041 10251
rect 23808 10220 24041 10248
rect 23808 10208 23814 10220
rect 24029 10217 24041 10220
rect 24075 10217 24087 10251
rect 24394 10248 24400 10260
rect 24355 10220 24400 10248
rect 24029 10211 24087 10217
rect 24394 10208 24400 10220
rect 24452 10208 24458 10260
rect 25314 10208 25320 10260
rect 25372 10248 25378 10260
rect 26237 10251 26295 10257
rect 26237 10248 26249 10251
rect 25372 10220 26249 10248
rect 25372 10208 25378 10220
rect 26237 10217 26249 10220
rect 26283 10217 26295 10251
rect 26237 10211 26295 10217
rect 26513 10251 26571 10257
rect 26513 10217 26525 10251
rect 26559 10248 26571 10251
rect 26694 10248 26700 10260
rect 26559 10220 26700 10248
rect 26559 10217 26571 10220
rect 26513 10211 26571 10217
rect 26694 10208 26700 10220
rect 26752 10208 26758 10260
rect 26970 10248 26976 10260
rect 26931 10220 26976 10248
rect 26970 10208 26976 10220
rect 27028 10208 27034 10260
rect 6086 10180 6092 10192
rect 6047 10152 6092 10180
rect 6086 10140 6092 10152
rect 6144 10140 6150 10192
rect 6178 10140 6184 10192
rect 6236 10180 6242 10192
rect 18141 10183 18199 10189
rect 6236 10152 6500 10180
rect 6236 10140 6242 10152
rect 5460 10084 6224 10112
rect 2869 10047 2927 10053
rect 2869 10013 2881 10047
rect 2915 10013 2927 10047
rect 2869 10007 2927 10013
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10044 3019 10047
rect 3237 10047 3295 10053
rect 3237 10044 3249 10047
rect 3007 10016 3249 10044
rect 3007 10013 3019 10016
rect 2961 10007 3019 10013
rect 3237 10013 3249 10016
rect 3283 10013 3295 10047
rect 4525 10047 4583 10053
rect 4525 10044 4537 10047
rect 3237 10007 3295 10013
rect 3896 10016 4537 10044
rect 2130 9936 2136 9988
rect 2188 9976 2194 9988
rect 2409 9979 2467 9985
rect 2409 9976 2421 9979
rect 2188 9948 2421 9976
rect 2188 9936 2194 9948
rect 2409 9945 2421 9948
rect 2455 9945 2467 9979
rect 2884 9976 2912 10007
rect 3142 9976 3148 9988
rect 2884 9948 3148 9976
rect 2409 9939 2467 9945
rect 3142 9936 3148 9948
rect 3200 9936 3206 9988
rect 3896 9920 3924 10016
rect 4525 10013 4537 10016
rect 4571 10013 4583 10047
rect 4706 10044 4712 10056
rect 4667 10016 4712 10044
rect 4525 10007 4583 10013
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 6196 10053 6224 10084
rect 6472 10056 6500 10152
rect 18141 10149 18153 10183
rect 18187 10180 18199 10183
rect 18690 10180 18696 10192
rect 18187 10152 18696 10180
rect 18187 10149 18199 10152
rect 18141 10143 18199 10149
rect 18690 10140 18696 10152
rect 18748 10140 18754 10192
rect 19058 10140 19064 10192
rect 19116 10180 19122 10192
rect 19705 10183 19763 10189
rect 19705 10180 19717 10183
rect 19116 10152 19717 10180
rect 19116 10140 19122 10152
rect 19705 10149 19717 10152
rect 19751 10149 19763 10183
rect 19705 10143 19763 10149
rect 20346 10140 20352 10192
rect 20404 10180 20410 10192
rect 21174 10180 21180 10192
rect 20404 10152 21180 10180
rect 20404 10140 20410 10152
rect 21174 10140 21180 10152
rect 21232 10180 21238 10192
rect 21361 10183 21419 10189
rect 21361 10180 21373 10183
rect 21232 10152 21373 10180
rect 21232 10140 21238 10152
rect 21361 10149 21373 10152
rect 21407 10149 21419 10183
rect 21361 10143 21419 10149
rect 23109 10183 23167 10189
rect 23109 10149 23121 10183
rect 23155 10180 23167 10183
rect 23290 10180 23296 10192
rect 23155 10152 23296 10180
rect 23155 10149 23167 10152
rect 23109 10143 23167 10149
rect 23290 10140 23296 10152
rect 23348 10140 23354 10192
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 7561 10115 7619 10121
rect 7561 10112 7573 10115
rect 6972 10084 7573 10112
rect 6972 10072 6978 10084
rect 7561 10081 7573 10084
rect 7607 10112 7619 10115
rect 8573 10115 8631 10121
rect 8573 10112 8585 10115
rect 7607 10084 8585 10112
rect 7607 10081 7619 10084
rect 7561 10075 7619 10081
rect 8573 10081 8585 10084
rect 8619 10081 8631 10115
rect 8573 10075 8631 10081
rect 17037 10115 17095 10121
rect 17037 10081 17049 10115
rect 17083 10112 17095 10115
rect 17402 10112 17408 10124
rect 17083 10084 17408 10112
rect 17083 10081 17095 10084
rect 17037 10075 17095 10081
rect 17402 10072 17408 10084
rect 17460 10072 17466 10124
rect 19150 10112 19156 10124
rect 19111 10084 19156 10112
rect 19150 10072 19156 10084
rect 19208 10072 19214 10124
rect 19334 10072 19340 10124
rect 19392 10112 19398 10124
rect 19518 10112 19524 10124
rect 19392 10084 19524 10112
rect 19392 10072 19398 10084
rect 19518 10072 19524 10084
rect 19576 10112 19582 10124
rect 19613 10115 19671 10121
rect 19613 10112 19625 10115
rect 19576 10084 19625 10112
rect 19576 10072 19582 10084
rect 19613 10081 19625 10084
rect 19659 10081 19671 10115
rect 19613 10075 19671 10081
rect 23753 10115 23811 10121
rect 23753 10081 23765 10115
rect 23799 10112 23811 10115
rect 23934 10112 23940 10124
rect 23799 10084 23940 10112
rect 23799 10081 23811 10084
rect 23753 10075 23811 10081
rect 23934 10072 23940 10084
rect 23992 10072 23998 10124
rect 24118 10072 24124 10124
rect 24176 10112 24182 10124
rect 24213 10115 24271 10121
rect 24213 10112 24225 10115
rect 24176 10084 24225 10112
rect 24176 10072 24182 10084
rect 24213 10081 24225 10084
rect 24259 10081 24271 10115
rect 25314 10112 25320 10124
rect 25275 10084 25320 10112
rect 24213 10075 24271 10081
rect 25314 10072 25320 10084
rect 25372 10072 25378 10124
rect 26786 10072 26792 10124
rect 26844 10112 26850 10124
rect 26881 10115 26939 10121
rect 26881 10112 26893 10115
rect 26844 10084 26893 10112
rect 26844 10072 26850 10084
rect 26881 10081 26893 10084
rect 26927 10081 26939 10115
rect 26881 10075 26939 10081
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 6454 10004 6460 10056
rect 6512 10004 6518 10056
rect 6638 10004 6644 10056
rect 6696 10044 6702 10056
rect 7653 10047 7711 10053
rect 7653 10044 7665 10047
rect 6696 10016 7665 10044
rect 6696 10004 6702 10016
rect 7653 10013 7665 10016
rect 7699 10013 7711 10047
rect 7653 10007 7711 10013
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 8110 10044 8116 10056
rect 7883 10016 8116 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 3970 9936 3976 9988
rect 4028 9976 4034 9988
rect 4065 9979 4123 9985
rect 4065 9976 4077 9979
rect 4028 9948 4077 9976
rect 4028 9936 4034 9948
rect 4065 9945 4077 9948
rect 4111 9945 4123 9979
rect 7190 9976 7196 9988
rect 7151 9948 7196 9976
rect 4065 9939 4123 9945
rect 7190 9936 7196 9948
rect 7248 9936 7254 9988
rect 7668 9976 7696 10007
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 10318 10044 10324 10056
rect 10279 10016 10324 10044
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 17310 10044 17316 10056
rect 17271 10016 17316 10044
rect 17310 10004 17316 10016
rect 17368 10004 17374 10056
rect 17773 10047 17831 10053
rect 17773 10013 17785 10047
rect 17819 10044 17831 10047
rect 18230 10044 18236 10056
rect 17819 10016 18236 10044
rect 17819 10013 17831 10016
rect 17773 10007 17831 10013
rect 18230 10004 18236 10016
rect 18288 10044 18294 10056
rect 18966 10044 18972 10056
rect 18288 10016 18972 10044
rect 18288 10004 18294 10016
rect 18966 10004 18972 10016
rect 19024 10044 19030 10056
rect 19889 10047 19947 10053
rect 19889 10044 19901 10047
rect 19024 10016 19901 10044
rect 19024 10004 19030 10016
rect 19889 10013 19901 10016
rect 19935 10044 19947 10047
rect 20162 10044 20168 10056
rect 19935 10016 20168 10044
rect 19935 10013 19947 10016
rect 19889 10007 19947 10013
rect 20162 10004 20168 10016
rect 20220 10044 20226 10056
rect 21545 10047 21603 10053
rect 21545 10044 21557 10047
rect 20220 10016 21557 10044
rect 20220 10004 20226 10016
rect 21545 10013 21557 10016
rect 21591 10044 21603 10047
rect 21818 10044 21824 10056
rect 21591 10016 21824 10044
rect 21591 10013 21603 10016
rect 21545 10007 21603 10013
rect 21818 10004 21824 10016
rect 21876 10004 21882 10056
rect 23106 10004 23112 10056
rect 23164 10044 23170 10056
rect 23201 10047 23259 10053
rect 23201 10044 23213 10047
rect 23164 10016 23213 10044
rect 23164 10004 23170 10016
rect 23201 10013 23213 10016
rect 23247 10013 23259 10047
rect 27154 10044 27160 10056
rect 27115 10016 27160 10044
rect 23201 10007 23259 10013
rect 27154 10004 27160 10016
rect 27212 10004 27218 10056
rect 8205 9979 8263 9985
rect 8205 9976 8217 9979
rect 7668 9948 8217 9976
rect 8205 9945 8217 9948
rect 8251 9945 8263 9979
rect 8205 9939 8263 9945
rect 3878 9908 3884 9920
rect 3839 9880 3884 9908
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 16666 9908 16672 9920
rect 16627 9880 16672 9908
rect 16666 9868 16672 9880
rect 16724 9868 16730 9920
rect 25501 9911 25559 9917
rect 25501 9877 25513 9911
rect 25547 9908 25559 9911
rect 25590 9908 25596 9920
rect 25547 9880 25596 9908
rect 25547 9877 25559 9880
rect 25501 9871 25559 9877
rect 25590 9868 25596 9880
rect 25648 9868 25654 9920
rect 1104 9818 28888 9840
rect 1104 9766 5982 9818
rect 6034 9766 6046 9818
rect 6098 9766 6110 9818
rect 6162 9766 6174 9818
rect 6226 9766 15982 9818
rect 16034 9766 16046 9818
rect 16098 9766 16110 9818
rect 16162 9766 16174 9818
rect 16226 9766 25982 9818
rect 26034 9766 26046 9818
rect 26098 9766 26110 9818
rect 26162 9766 26174 9818
rect 26226 9766 28888 9818
rect 1104 9744 28888 9766
rect 2406 9664 2412 9716
rect 2464 9704 2470 9716
rect 3510 9704 3516 9716
rect 2464 9676 2728 9704
rect 2464 9664 2470 9676
rect 2700 9645 2728 9676
rect 3068 9676 3516 9704
rect 2685 9639 2743 9645
rect 2685 9605 2697 9639
rect 2731 9605 2743 9639
rect 2685 9599 2743 9605
rect 1946 9528 1952 9580
rect 2004 9568 2010 9580
rect 2041 9571 2099 9577
rect 2041 9568 2053 9571
rect 2004 9540 2053 9568
rect 2004 9528 2010 9540
rect 2041 9537 2053 9540
rect 2087 9537 2099 9571
rect 2222 9568 2228 9580
rect 2183 9540 2228 9568
rect 2041 9531 2099 9537
rect 2222 9528 2228 9540
rect 2280 9528 2286 9580
rect 2958 9528 2964 9580
rect 3016 9568 3022 9580
rect 3068 9568 3096 9676
rect 3510 9664 3516 9676
rect 3568 9664 3574 9716
rect 4522 9704 4528 9716
rect 4483 9676 4528 9704
rect 4522 9664 4528 9676
rect 4580 9664 4586 9716
rect 5718 9704 5724 9716
rect 5460 9676 5724 9704
rect 5169 9639 5227 9645
rect 5169 9605 5181 9639
rect 5215 9636 5227 9639
rect 5460 9636 5488 9676
rect 5718 9664 5724 9676
rect 5776 9664 5782 9716
rect 6273 9707 6331 9713
rect 6273 9673 6285 9707
rect 6319 9704 6331 9707
rect 6362 9704 6368 9716
rect 6319 9676 6368 9704
rect 6319 9673 6331 9676
rect 6273 9667 6331 9673
rect 6362 9664 6368 9676
rect 6420 9664 6426 9716
rect 17126 9704 17132 9716
rect 6840 9676 8156 9704
rect 5215 9608 5488 9636
rect 5215 9605 5227 9608
rect 5169 9599 5227 9605
rect 6086 9596 6092 9648
rect 6144 9636 6150 9648
rect 6840 9636 6868 9676
rect 8128 9648 8156 9676
rect 16592 9676 17132 9704
rect 6144 9608 6868 9636
rect 6144 9596 6150 9608
rect 8110 9596 8116 9648
rect 8168 9636 8174 9648
rect 8849 9639 8907 9645
rect 8849 9636 8861 9639
rect 8168 9608 8861 9636
rect 8168 9596 8174 9608
rect 8849 9605 8861 9608
rect 8895 9605 8907 9639
rect 8849 9599 8907 9605
rect 15746 9596 15752 9648
rect 15804 9636 15810 9648
rect 16301 9639 16359 9645
rect 16301 9636 16313 9639
rect 15804 9608 16313 9636
rect 15804 9596 15810 9608
rect 16301 9605 16313 9608
rect 16347 9636 16359 9639
rect 16592 9636 16620 9676
rect 17126 9664 17132 9676
rect 17184 9664 17190 9716
rect 19150 9664 19156 9716
rect 19208 9704 19214 9716
rect 19208 9676 19288 9704
rect 19208 9664 19214 9676
rect 16347 9608 16620 9636
rect 18877 9639 18935 9645
rect 16347 9605 16359 9608
rect 16301 9599 16359 9605
rect 18877 9605 18889 9639
rect 18923 9636 18935 9639
rect 19058 9636 19064 9648
rect 18923 9608 19064 9636
rect 18923 9605 18935 9608
rect 18877 9599 18935 9605
rect 19058 9596 19064 9608
rect 19116 9596 19122 9648
rect 19260 9636 19288 9676
rect 21174 9664 21180 9716
rect 21232 9704 21238 9716
rect 21269 9707 21327 9713
rect 21269 9704 21281 9707
rect 21232 9676 21281 9704
rect 21232 9664 21238 9676
rect 21269 9673 21281 9676
rect 21315 9673 21327 9707
rect 21269 9667 21327 9673
rect 21729 9707 21787 9713
rect 21729 9673 21741 9707
rect 21775 9704 21787 9707
rect 22002 9704 22008 9716
rect 21775 9676 22008 9704
rect 21775 9673 21787 9676
rect 21729 9667 21787 9673
rect 22002 9664 22008 9676
rect 22060 9664 22066 9716
rect 24118 9704 24124 9716
rect 24079 9676 24124 9704
rect 24118 9664 24124 9676
rect 24176 9664 24182 9716
rect 25225 9707 25283 9713
rect 25225 9673 25237 9707
rect 25271 9704 25283 9707
rect 25314 9704 25320 9716
rect 25271 9676 25320 9704
rect 25271 9673 25283 9676
rect 25225 9667 25283 9673
rect 25314 9664 25320 9676
rect 25372 9664 25378 9716
rect 26970 9664 26976 9716
rect 27028 9704 27034 9716
rect 27341 9707 27399 9713
rect 27341 9704 27353 9707
rect 27028 9676 27353 9704
rect 27028 9664 27034 9676
rect 27341 9673 27353 9676
rect 27387 9673 27399 9707
rect 27341 9667 27399 9673
rect 25498 9636 25504 9648
rect 19260 9608 19380 9636
rect 25459 9608 25504 9636
rect 3016 9540 3096 9568
rect 5537 9571 5595 9577
rect 3016 9528 3022 9540
rect 5537 9537 5549 9571
rect 5583 9568 5595 9571
rect 5810 9568 5816 9580
rect 5583 9540 5816 9568
rect 5583 9537 5595 9540
rect 5537 9531 5595 9537
rect 3053 9503 3111 9509
rect 3053 9469 3065 9503
rect 3099 9500 3111 9503
rect 3145 9503 3203 9509
rect 3145 9500 3157 9503
rect 3099 9472 3157 9500
rect 3099 9469 3111 9472
rect 3053 9463 3111 9469
rect 3145 9469 3157 9472
rect 3191 9500 3203 9503
rect 4798 9500 4804 9512
rect 3191 9472 4804 9500
rect 3191 9469 3203 9472
rect 3145 9463 3203 9469
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 5644 9509 5672 9540
rect 5810 9528 5816 9540
rect 5868 9528 5874 9580
rect 15930 9568 15936 9580
rect 15843 9540 15936 9568
rect 15930 9528 15936 9540
rect 15988 9568 15994 9580
rect 16850 9568 16856 9580
rect 15988 9540 16856 9568
rect 15988 9528 15994 9540
rect 16850 9528 16856 9540
rect 16908 9528 16914 9580
rect 17037 9571 17095 9577
rect 17037 9537 17049 9571
rect 17083 9568 17095 9571
rect 17310 9568 17316 9580
rect 17083 9540 17316 9568
rect 17083 9537 17095 9540
rect 17037 9531 17095 9537
rect 17310 9528 17316 9540
rect 17368 9568 17374 9580
rect 17770 9568 17776 9580
rect 17368 9540 17776 9568
rect 17368 9528 17374 9540
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 19352 9568 19380 9608
rect 25498 9596 25504 9608
rect 25556 9596 25562 9648
rect 26329 9639 26387 9645
rect 26329 9605 26341 9639
rect 26375 9636 26387 9639
rect 27246 9636 27252 9648
rect 26375 9608 27252 9636
rect 26375 9605 26387 9608
rect 26329 9599 26387 9605
rect 19352 9540 19472 9568
rect 5629 9503 5687 9509
rect 5629 9469 5641 9503
rect 5675 9500 5687 9503
rect 6917 9503 6975 9509
rect 6917 9500 6929 9503
rect 5675 9472 5709 9500
rect 6564 9472 6929 9500
rect 5675 9469 5687 9472
rect 5629 9463 5687 9469
rect 1486 9392 1492 9444
rect 1544 9432 1550 9444
rect 1670 9432 1676 9444
rect 1544 9404 1676 9432
rect 1544 9392 1550 9404
rect 1670 9392 1676 9404
rect 1728 9392 1734 9444
rect 1946 9432 1952 9444
rect 1907 9404 1952 9432
rect 1946 9392 1952 9404
rect 2004 9392 2010 9444
rect 3418 9441 3424 9444
rect 3412 9432 3424 9441
rect 3379 9404 3424 9432
rect 3412 9395 3424 9404
rect 3418 9392 3424 9395
rect 3476 9392 3482 9444
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 5810 9364 5816 9376
rect 5771 9336 5816 9364
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 6454 9324 6460 9376
rect 6512 9364 6518 9376
rect 6564 9373 6592 9472
rect 6917 9469 6929 9472
rect 6963 9469 6975 9503
rect 18506 9500 18512 9512
rect 18419 9472 18512 9500
rect 6917 9463 6975 9469
rect 18506 9460 18512 9472
rect 18564 9500 18570 9512
rect 19337 9503 19395 9509
rect 19337 9500 19349 9503
rect 18564 9472 19349 9500
rect 18564 9460 18570 9472
rect 19337 9469 19349 9472
rect 19383 9469 19395 9503
rect 19444 9500 19472 9540
rect 19593 9503 19651 9509
rect 19593 9500 19605 9503
rect 19444 9472 19605 9500
rect 19337 9463 19395 9469
rect 19593 9469 19605 9472
rect 19639 9500 19651 9503
rect 19886 9500 19892 9512
rect 19639 9472 19892 9500
rect 19639 9469 19651 9472
rect 19593 9463 19651 9469
rect 7098 9392 7104 9444
rect 7156 9441 7162 9444
rect 7156 9435 7220 9441
rect 7156 9401 7174 9435
rect 7208 9401 7220 9435
rect 7156 9395 7220 9401
rect 7156 9392 7162 9395
rect 15470 9392 15476 9444
rect 15528 9432 15534 9444
rect 15565 9435 15623 9441
rect 15565 9432 15577 9435
rect 15528 9404 15577 9432
rect 15528 9392 15534 9404
rect 15565 9401 15577 9404
rect 15611 9432 15623 9435
rect 16761 9435 16819 9441
rect 16761 9432 16773 9435
rect 15611 9404 16773 9432
rect 15611 9401 15623 9404
rect 15565 9395 15623 9401
rect 16761 9401 16773 9404
rect 16807 9401 16819 9435
rect 19352 9432 19380 9463
rect 19886 9460 19892 9472
rect 19944 9460 19950 9512
rect 24210 9500 24216 9512
rect 24171 9472 24216 9500
rect 24210 9460 24216 9472
rect 24268 9500 24274 9512
rect 24765 9503 24823 9509
rect 24765 9500 24777 9503
rect 24268 9472 24777 9500
rect 24268 9460 24274 9472
rect 24765 9469 24777 9472
rect 24811 9469 24823 9503
rect 24765 9463 24823 9469
rect 25222 9460 25228 9512
rect 25280 9500 25286 9512
rect 26436 9509 26464 9608
rect 27246 9596 27252 9608
rect 27304 9596 27310 9648
rect 25317 9503 25375 9509
rect 25317 9500 25329 9503
rect 25280 9472 25329 9500
rect 25280 9460 25286 9472
rect 25317 9469 25329 9472
rect 25363 9500 25375 9503
rect 25869 9503 25927 9509
rect 25869 9500 25881 9503
rect 25363 9472 25881 9500
rect 25363 9469 25375 9472
rect 25317 9463 25375 9469
rect 25869 9469 25881 9472
rect 25915 9469 25927 9503
rect 25869 9463 25927 9469
rect 26421 9503 26479 9509
rect 26421 9469 26433 9503
rect 26467 9469 26479 9503
rect 27522 9500 27528 9512
rect 27483 9472 27528 9500
rect 26421 9463 26479 9469
rect 19702 9432 19708 9444
rect 19352 9404 19708 9432
rect 16761 9395 16819 9401
rect 19702 9392 19708 9404
rect 19760 9392 19766 9444
rect 25884 9432 25912 9463
rect 27522 9460 27528 9472
rect 27580 9500 27586 9512
rect 28077 9503 28135 9509
rect 28077 9500 28089 9503
rect 27580 9472 28089 9500
rect 27580 9460 27586 9472
rect 28077 9469 28089 9472
rect 28123 9469 28135 9503
rect 28077 9463 28135 9469
rect 26786 9432 26792 9444
rect 25884 9404 26792 9432
rect 26786 9392 26792 9404
rect 26844 9432 26850 9444
rect 26973 9435 27031 9441
rect 26973 9432 26985 9435
rect 26844 9404 26985 9432
rect 26844 9392 26850 9404
rect 26973 9401 26985 9404
rect 27019 9401 27031 9435
rect 26973 9395 27031 9401
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 6512 9336 6561 9364
rect 6512 9324 6518 9336
rect 6549 9333 6561 9336
rect 6595 9333 6607 9367
rect 6549 9327 6607 9333
rect 7466 9324 7472 9376
rect 7524 9364 7530 9376
rect 8297 9367 8355 9373
rect 8297 9364 8309 9367
rect 7524 9336 8309 9364
rect 7524 9324 7530 9336
rect 8297 9333 8309 9336
rect 8343 9333 8355 9367
rect 16390 9364 16396 9376
rect 16351 9336 16396 9364
rect 8297 9327 8355 9333
rect 16390 9324 16396 9336
rect 16448 9324 16454 9376
rect 17402 9364 17408 9376
rect 17363 9336 17408 9364
rect 17402 9324 17408 9336
rect 17460 9324 17466 9376
rect 17770 9364 17776 9376
rect 17731 9336 17776 9364
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 19242 9364 19248 9376
rect 19203 9336 19248 9364
rect 19242 9324 19248 9336
rect 19300 9324 19306 9376
rect 20254 9324 20260 9376
rect 20312 9364 20318 9376
rect 20717 9367 20775 9373
rect 20717 9364 20729 9367
rect 20312 9336 20729 9364
rect 20312 9324 20318 9336
rect 20717 9333 20729 9336
rect 20763 9333 20775 9367
rect 20717 9327 20775 9333
rect 22094 9324 22100 9376
rect 22152 9364 22158 9376
rect 24394 9364 24400 9376
rect 22152 9336 22197 9364
rect 24355 9336 24400 9364
rect 22152 9324 22158 9336
rect 24394 9324 24400 9336
rect 24452 9324 24458 9376
rect 26605 9367 26663 9373
rect 26605 9333 26617 9367
rect 26651 9364 26663 9367
rect 26878 9364 26884 9376
rect 26651 9336 26884 9364
rect 26651 9333 26663 9336
rect 26605 9327 26663 9333
rect 26878 9324 26884 9336
rect 26936 9324 26942 9376
rect 27709 9367 27767 9373
rect 27709 9333 27721 9367
rect 27755 9364 27767 9367
rect 27798 9364 27804 9376
rect 27755 9336 27804 9364
rect 27755 9333 27767 9336
rect 27709 9327 27767 9333
rect 27798 9324 27804 9336
rect 27856 9324 27862 9376
rect 1104 9274 28888 9296
rect 1104 9222 10982 9274
rect 11034 9222 11046 9274
rect 11098 9222 11110 9274
rect 11162 9222 11174 9274
rect 11226 9222 20982 9274
rect 21034 9222 21046 9274
rect 21098 9222 21110 9274
rect 21162 9222 21174 9274
rect 21226 9222 28888 9274
rect 1104 9200 28888 9222
rect 1673 9163 1731 9169
rect 1673 9129 1685 9163
rect 1719 9160 1731 9163
rect 1946 9160 1952 9172
rect 1719 9132 1952 9160
rect 1719 9129 1731 9132
rect 1673 9123 1731 9129
rect 1946 9120 1952 9132
rect 2004 9120 2010 9172
rect 3237 9163 3295 9169
rect 3237 9129 3249 9163
rect 3283 9160 3295 9163
rect 3418 9160 3424 9172
rect 3283 9132 3424 9160
rect 3283 9129 3295 9132
rect 3237 9123 3295 9129
rect 3418 9120 3424 9132
rect 3476 9160 3482 9172
rect 4341 9163 4399 9169
rect 4341 9160 4353 9163
rect 3476 9132 4353 9160
rect 3476 9120 3482 9132
rect 4341 9129 4353 9132
rect 4387 9160 4399 9163
rect 4706 9160 4712 9172
rect 4387 9132 4712 9160
rect 4387 9129 4399 9132
rect 4341 9123 4399 9129
rect 4706 9120 4712 9132
rect 4764 9160 4770 9172
rect 6086 9160 6092 9172
rect 4764 9132 6092 9160
rect 4764 9120 4770 9132
rect 6086 9120 6092 9132
rect 6144 9120 6150 9172
rect 7006 9120 7012 9172
rect 7064 9160 7070 9172
rect 7374 9160 7380 9172
rect 7064 9132 7380 9160
rect 7064 9120 7070 9132
rect 7374 9120 7380 9132
rect 7432 9160 7438 9172
rect 7561 9163 7619 9169
rect 7561 9160 7573 9163
rect 7432 9132 7573 9160
rect 7432 9120 7438 9132
rect 7561 9129 7573 9132
rect 7607 9129 7619 9163
rect 7561 9123 7619 9129
rect 7653 9163 7711 9169
rect 7653 9129 7665 9163
rect 7699 9160 7711 9163
rect 7742 9160 7748 9172
rect 7699 9132 7748 9160
rect 7699 9129 7711 9132
rect 7653 9123 7711 9129
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 15470 9160 15476 9172
rect 15431 9132 15476 9160
rect 15470 9120 15476 9132
rect 15528 9120 15534 9172
rect 18966 9120 18972 9172
rect 19024 9160 19030 9172
rect 19061 9163 19119 9169
rect 19061 9160 19073 9163
rect 19024 9132 19073 9160
rect 19024 9120 19030 9132
rect 19061 9129 19073 9132
rect 19107 9129 19119 9163
rect 19061 9123 19119 9129
rect 20714 9120 20720 9172
rect 20772 9160 20778 9172
rect 21361 9163 21419 9169
rect 21361 9160 21373 9163
rect 20772 9132 21373 9160
rect 20772 9120 20778 9132
rect 21361 9129 21373 9132
rect 21407 9160 21419 9163
rect 21542 9160 21548 9172
rect 21407 9132 21548 9160
rect 21407 9129 21419 9132
rect 21361 9123 21419 9129
rect 21542 9120 21548 9132
rect 21600 9120 21606 9172
rect 27154 9160 27160 9172
rect 27115 9132 27160 9160
rect 27154 9120 27160 9132
rect 27212 9120 27218 9172
rect 1486 9052 1492 9104
rect 1544 9092 1550 9104
rect 2317 9095 2375 9101
rect 2317 9092 2329 9095
rect 1544 9064 2329 9092
rect 1544 9052 1550 9064
rect 2317 9061 2329 9064
rect 2363 9061 2375 9095
rect 2317 9055 2375 9061
rect 2409 9095 2467 9101
rect 2409 9061 2421 9095
rect 2455 9092 2467 9095
rect 2774 9092 2780 9104
rect 2455 9064 2780 9092
rect 2455 9061 2467 9064
rect 2409 9055 2467 9061
rect 2774 9052 2780 9064
rect 2832 9092 2838 9104
rect 4154 9092 4160 9104
rect 2832 9064 4160 9092
rect 2832 9052 2838 9064
rect 4154 9052 4160 9064
rect 4212 9052 4218 9104
rect 21269 9095 21327 9101
rect 21269 9061 21281 9095
rect 21315 9092 21327 9095
rect 21450 9092 21456 9104
rect 21315 9064 21456 9092
rect 21315 9061 21327 9064
rect 21269 9055 21327 9061
rect 21450 9052 21456 9064
rect 21508 9052 21514 9104
rect 3881 9027 3939 9033
rect 3881 8993 3893 9027
rect 3927 9024 3939 9027
rect 4976 9027 5034 9033
rect 4976 9024 4988 9027
rect 3927 8996 4988 9024
rect 3927 8993 3939 8996
rect 3881 8987 3939 8993
rect 4976 8993 4988 8996
rect 5022 9024 5034 9027
rect 5258 9024 5264 9036
rect 5022 8996 5264 9024
rect 5022 8993 5034 8996
rect 4976 8987 5034 8993
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 16393 9027 16451 9033
rect 16393 8993 16405 9027
rect 16439 9024 16451 9027
rect 16752 9027 16810 9033
rect 16752 9024 16764 9027
rect 16439 8996 16764 9024
rect 16439 8993 16451 8996
rect 16393 8987 16451 8993
rect 16752 8993 16764 8996
rect 16798 9024 16810 9027
rect 17770 9024 17776 9036
rect 16798 8996 17776 9024
rect 16798 8993 16810 8996
rect 16752 8987 16810 8993
rect 17770 8984 17776 8996
rect 17828 8984 17834 9036
rect 19518 8984 19524 9036
rect 19576 9024 19582 9036
rect 19613 9027 19671 9033
rect 19613 9024 19625 9027
rect 19576 8996 19625 9024
rect 19576 8984 19582 8996
rect 19613 8993 19625 8996
rect 19659 8993 19671 9027
rect 25314 9024 25320 9036
rect 25275 8996 25320 9024
rect 19613 8987 19671 8993
rect 25314 8984 25320 8996
rect 25372 8984 25378 9036
rect 26510 9024 26516 9036
rect 26471 8996 26516 9024
rect 26510 8984 26516 8996
rect 26568 8984 26574 9036
rect 2222 8916 2228 8968
rect 2280 8956 2286 8968
rect 2593 8959 2651 8965
rect 2593 8956 2605 8959
rect 2280 8928 2605 8956
rect 2280 8916 2286 8928
rect 2593 8925 2605 8928
rect 2639 8956 2651 8959
rect 2958 8956 2964 8968
rect 2639 8928 2964 8956
rect 2639 8925 2651 8928
rect 2593 8919 2651 8925
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 4706 8956 4712 8968
rect 4667 8928 4712 8956
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 7009 8959 7067 8965
rect 7009 8925 7021 8959
rect 7055 8956 7067 8959
rect 7098 8956 7104 8968
rect 7055 8928 7104 8956
rect 7055 8925 7067 8928
rect 7009 8919 7067 8925
rect 7098 8916 7104 8928
rect 7156 8956 7162 8968
rect 7837 8959 7895 8965
rect 7837 8956 7849 8959
rect 7156 8928 7849 8956
rect 7156 8916 7162 8928
rect 7837 8925 7849 8928
rect 7883 8956 7895 8959
rect 16482 8956 16488 8968
rect 7883 8928 8248 8956
rect 16443 8928 16488 8956
rect 7883 8925 7895 8928
rect 7837 8919 7895 8925
rect 6822 8848 6828 8900
rect 6880 8888 6886 8900
rect 7193 8891 7251 8897
rect 7193 8888 7205 8891
rect 6880 8860 7205 8888
rect 6880 8848 6886 8860
rect 7193 8857 7205 8860
rect 7239 8857 7251 8891
rect 7193 8851 7251 8857
rect 8220 8832 8248 8928
rect 16482 8916 16488 8928
rect 16540 8916 16546 8968
rect 19702 8956 19708 8968
rect 19663 8928 19708 8956
rect 19702 8916 19708 8928
rect 19760 8916 19766 8968
rect 19886 8956 19892 8968
rect 19847 8928 19892 8956
rect 19886 8916 19892 8928
rect 19944 8956 19950 8968
rect 21545 8959 21603 8965
rect 19944 8928 21404 8956
rect 19944 8916 19950 8928
rect 20806 8848 20812 8900
rect 20864 8888 20870 8900
rect 20901 8891 20959 8897
rect 20901 8888 20913 8891
rect 20864 8860 20913 8888
rect 20864 8848 20870 8860
rect 20901 8857 20913 8860
rect 20947 8857 20959 8891
rect 21376 8888 21404 8928
rect 21545 8925 21557 8959
rect 21591 8956 21603 8959
rect 21818 8956 21824 8968
rect 21591 8928 21824 8956
rect 21591 8925 21603 8928
rect 21545 8919 21603 8925
rect 21818 8916 21824 8928
rect 21876 8956 21882 8968
rect 22094 8956 22100 8968
rect 21876 8928 22100 8956
rect 21876 8916 21882 8928
rect 22094 8916 22100 8928
rect 22152 8916 22158 8968
rect 21726 8888 21732 8900
rect 21376 8860 21732 8888
rect 20901 8851 20959 8857
rect 21726 8848 21732 8860
rect 21784 8848 21790 8900
rect 1949 8823 2007 8829
rect 1949 8789 1961 8823
rect 1995 8820 2007 8823
rect 2130 8820 2136 8832
rect 1995 8792 2136 8820
rect 1995 8789 2007 8792
rect 1949 8783 2007 8789
rect 2130 8780 2136 8792
rect 2188 8780 2194 8832
rect 8202 8780 8208 8832
rect 8260 8820 8266 8832
rect 8389 8823 8447 8829
rect 8389 8820 8401 8823
rect 8260 8792 8401 8820
rect 8260 8780 8266 8792
rect 8389 8789 8401 8792
rect 8435 8789 8447 8823
rect 17862 8820 17868 8832
rect 17823 8792 17868 8820
rect 8389 8783 8447 8789
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 18782 8820 18788 8832
rect 18743 8792 18788 8820
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 19245 8823 19303 8829
rect 19245 8789 19257 8823
rect 19291 8820 19303 8823
rect 19334 8820 19340 8832
rect 19291 8792 19340 8820
rect 19291 8789 19303 8792
rect 19245 8783 19303 8789
rect 19334 8780 19340 8792
rect 19392 8780 19398 8832
rect 20070 8780 20076 8832
rect 20128 8820 20134 8832
rect 20257 8823 20315 8829
rect 20257 8820 20269 8823
rect 20128 8792 20269 8820
rect 20128 8780 20134 8792
rect 20257 8789 20269 8792
rect 20303 8789 20315 8823
rect 25498 8820 25504 8832
rect 25459 8792 25504 8820
rect 20257 8783 20315 8789
rect 25498 8780 25504 8792
rect 25556 8780 25562 8832
rect 25866 8780 25872 8832
rect 25924 8820 25930 8832
rect 26697 8823 26755 8829
rect 26697 8820 26709 8823
rect 25924 8792 26709 8820
rect 25924 8780 25930 8792
rect 26697 8789 26709 8792
rect 26743 8789 26755 8823
rect 26697 8783 26755 8789
rect 1104 8730 28888 8752
rect 1104 8678 5982 8730
rect 6034 8678 6046 8730
rect 6098 8678 6110 8730
rect 6162 8678 6174 8730
rect 6226 8678 15982 8730
rect 16034 8678 16046 8730
rect 16098 8678 16110 8730
rect 16162 8678 16174 8730
rect 16226 8678 25982 8730
rect 26034 8678 26046 8730
rect 26098 8678 26110 8730
rect 26162 8678 26174 8730
rect 26226 8678 28888 8730
rect 1104 8656 28888 8678
rect 1486 8576 1492 8628
rect 1544 8616 1550 8628
rect 1581 8619 1639 8625
rect 1581 8616 1593 8619
rect 1544 8588 1593 8616
rect 1544 8576 1550 8588
rect 1581 8585 1593 8588
rect 1627 8585 1639 8619
rect 1581 8579 1639 8585
rect 3789 8619 3847 8625
rect 3789 8585 3801 8619
rect 3835 8616 3847 8619
rect 4062 8616 4068 8628
rect 3835 8588 4068 8616
rect 3835 8585 3847 8588
rect 3789 8579 3847 8585
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 5997 8619 6055 8625
rect 5997 8585 6009 8619
rect 6043 8616 6055 8619
rect 6546 8616 6552 8628
rect 6043 8588 6552 8616
rect 6043 8585 6055 8588
rect 5997 8579 6055 8585
rect 2774 8508 2780 8560
rect 2832 8548 2838 8560
rect 5534 8548 5540 8560
rect 2832 8520 2877 8548
rect 5495 8520 5540 8548
rect 2832 8508 2838 8520
rect 5534 8508 5540 8520
rect 5592 8508 5598 8560
rect 1578 8440 1584 8492
rect 1636 8480 1642 8492
rect 1946 8480 1952 8492
rect 1636 8452 1952 8480
rect 1636 8440 1642 8452
rect 1946 8440 1952 8452
rect 2004 8480 2010 8492
rect 2225 8483 2283 8489
rect 2225 8480 2237 8483
rect 2004 8452 2237 8480
rect 2004 8440 2010 8452
rect 2225 8449 2237 8452
rect 2271 8449 2283 8483
rect 2225 8443 2283 8449
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8480 2467 8483
rect 2682 8480 2688 8492
rect 2455 8452 2688 8480
rect 2455 8449 2467 8452
rect 2409 8443 2467 8449
rect 2682 8440 2688 8452
rect 2740 8440 2746 8492
rect 3510 8440 3516 8492
rect 3568 8480 3574 8492
rect 3697 8483 3755 8489
rect 3697 8480 3709 8483
rect 3568 8452 3709 8480
rect 3568 8440 3574 8452
rect 3697 8449 3709 8452
rect 3743 8480 3755 8483
rect 4246 8480 4252 8492
rect 3743 8452 4252 8480
rect 3743 8449 3755 8452
rect 3697 8443 3755 8449
rect 4246 8440 4252 8452
rect 4304 8440 4310 8492
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8480 4491 8483
rect 5258 8480 5264 8492
rect 4479 8452 5264 8480
rect 4479 8449 4491 8452
rect 4433 8443 4491 8449
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 1670 8372 1676 8424
rect 1728 8412 1734 8424
rect 2958 8412 2964 8424
rect 1728 8384 2964 8412
rect 1728 8372 1734 8384
rect 2958 8372 2964 8384
rect 3016 8412 3022 8424
rect 3145 8415 3203 8421
rect 3145 8412 3157 8415
rect 3016 8384 3157 8412
rect 3016 8372 3022 8384
rect 3145 8381 3157 8384
rect 3191 8381 3203 8415
rect 3145 8375 3203 8381
rect 5353 8415 5411 8421
rect 5353 8381 5365 8415
rect 5399 8412 5411 8415
rect 6012 8412 6040 8579
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 6730 8576 6736 8628
rect 6788 8616 6794 8628
rect 6825 8619 6883 8625
rect 6825 8616 6837 8619
rect 6788 8588 6837 8616
rect 6788 8576 6794 8588
rect 6825 8585 6837 8588
rect 6871 8585 6883 8619
rect 6825 8579 6883 8585
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 7837 8619 7895 8625
rect 7837 8616 7849 8619
rect 7800 8588 7849 8616
rect 7800 8576 7806 8588
rect 7837 8585 7849 8588
rect 7883 8585 7895 8619
rect 7837 8579 7895 8585
rect 16301 8619 16359 8625
rect 16301 8585 16313 8619
rect 16347 8616 16359 8619
rect 16482 8616 16488 8628
rect 16347 8588 16488 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 16482 8576 16488 8588
rect 16540 8576 16546 8628
rect 20717 8619 20775 8625
rect 20717 8585 20729 8619
rect 20763 8616 20775 8619
rect 21450 8616 21456 8628
rect 20763 8588 21456 8616
rect 20763 8585 20775 8588
rect 20717 8579 20775 8585
rect 21450 8576 21456 8588
rect 21508 8576 21514 8628
rect 22094 8576 22100 8628
rect 22152 8616 22158 8628
rect 22189 8619 22247 8625
rect 22189 8616 22201 8619
rect 22152 8588 22201 8616
rect 22152 8576 22158 8588
rect 22189 8585 22201 8588
rect 22235 8585 22247 8619
rect 22189 8579 22247 8585
rect 25225 8619 25283 8625
rect 25225 8585 25237 8619
rect 25271 8616 25283 8619
rect 25314 8616 25320 8628
rect 25271 8588 25320 8616
rect 25271 8585 25283 8588
rect 25225 8579 25283 8585
rect 25314 8576 25320 8588
rect 25372 8576 25378 8628
rect 25774 8576 25780 8628
rect 25832 8616 25838 8628
rect 25869 8619 25927 8625
rect 25869 8616 25881 8619
rect 25832 8588 25881 8616
rect 25832 8576 25838 8588
rect 25869 8585 25881 8588
rect 25915 8585 25927 8619
rect 25869 8579 25927 8585
rect 26510 8576 26516 8628
rect 26568 8616 26574 8628
rect 27341 8619 27399 8625
rect 27341 8616 27353 8619
rect 26568 8588 27353 8616
rect 26568 8576 26574 8588
rect 27341 8585 27353 8588
rect 27387 8585 27399 8619
rect 27706 8616 27712 8628
rect 27667 8588 27712 8616
rect 27341 8579 27399 8585
rect 27706 8576 27712 8588
rect 27764 8576 27770 8628
rect 8389 8551 8447 8557
rect 8389 8548 8401 8551
rect 7300 8520 8401 8548
rect 7300 8489 7328 8520
rect 8389 8517 8401 8520
rect 8435 8548 8447 8551
rect 9401 8551 9459 8557
rect 9401 8548 9413 8551
rect 8435 8520 9413 8548
rect 8435 8517 8447 8520
rect 8389 8511 8447 8517
rect 9401 8517 9413 8520
rect 9447 8517 9459 8551
rect 9401 8511 9459 8517
rect 15933 8551 15991 8557
rect 15933 8517 15945 8551
rect 15979 8548 15991 8551
rect 21177 8551 21235 8557
rect 21177 8548 21189 8551
rect 15979 8520 17080 8548
rect 15979 8517 15991 8520
rect 15933 8511 15991 8517
rect 17052 8492 17080 8520
rect 20088 8520 21189 8548
rect 20088 8492 20116 8520
rect 21177 8517 21189 8520
rect 21223 8517 21235 8551
rect 21177 8511 21235 8517
rect 21634 8508 21640 8560
rect 21692 8548 21698 8560
rect 26234 8548 26240 8560
rect 21692 8520 26240 8548
rect 21692 8508 21698 8520
rect 26234 8508 26240 8520
rect 26292 8508 26298 8560
rect 26602 8548 26608 8560
rect 26563 8520 26608 8548
rect 26602 8508 26608 8520
rect 26660 8508 26666 8560
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 7466 8480 7472 8492
rect 7427 8452 7472 8480
rect 7285 8443 7343 8449
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 8202 8440 8208 8492
rect 8260 8480 8266 8492
rect 8941 8483 8999 8489
rect 8941 8480 8953 8483
rect 8260 8452 8953 8480
rect 8260 8440 8266 8452
rect 8941 8449 8953 8452
rect 8987 8449 8999 8483
rect 8941 8443 8999 8449
rect 15565 8483 15623 8489
rect 15565 8449 15577 8483
rect 15611 8480 15623 8483
rect 16666 8480 16672 8492
rect 15611 8452 16672 8480
rect 15611 8449 15623 8452
rect 15565 8443 15623 8449
rect 16666 8440 16672 8452
rect 16724 8480 16730 8492
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 16724 8452 16865 8480
rect 16724 8440 16730 8452
rect 16853 8449 16865 8452
rect 16899 8449 16911 8483
rect 17034 8480 17040 8492
rect 16995 8452 17040 8480
rect 16853 8443 16911 8449
rect 17034 8440 17040 8452
rect 17092 8480 17098 8492
rect 17773 8483 17831 8489
rect 17773 8480 17785 8483
rect 17092 8452 17785 8480
rect 17092 8440 17098 8452
rect 17773 8449 17785 8452
rect 17819 8480 17831 8483
rect 17862 8480 17868 8492
rect 17819 8452 17868 8480
rect 17819 8449 17831 8452
rect 17773 8443 17831 8449
rect 17862 8440 17868 8452
rect 17920 8480 17926 8492
rect 18601 8483 18659 8489
rect 18601 8480 18613 8483
rect 17920 8452 18613 8480
rect 17920 8440 17926 8452
rect 18601 8449 18613 8452
rect 18647 8449 18659 8483
rect 18601 8443 18659 8449
rect 19337 8483 19395 8489
rect 19337 8449 19349 8483
rect 19383 8480 19395 8483
rect 19702 8480 19708 8492
rect 19383 8452 19708 8480
rect 19383 8449 19395 8452
rect 19337 8443 19395 8449
rect 19702 8440 19708 8452
rect 19760 8480 19766 8492
rect 19886 8480 19892 8492
rect 19760 8452 19892 8480
rect 19760 8440 19766 8452
rect 19886 8440 19892 8452
rect 19944 8440 19950 8492
rect 20070 8480 20076 8492
rect 20031 8452 20076 8480
rect 20070 8440 20076 8452
rect 20128 8440 20134 8492
rect 20254 8480 20260 8492
rect 20215 8452 20260 8480
rect 20254 8440 20260 8452
rect 20312 8440 20318 8492
rect 21726 8480 21732 8492
rect 21687 8452 21732 8480
rect 21726 8440 21732 8452
rect 21784 8440 21790 8492
rect 5399 8384 6040 8412
rect 6641 8415 6699 8421
rect 5399 8381 5411 8384
rect 5353 8375 5411 8381
rect 6641 8381 6653 8415
rect 6687 8412 6699 8415
rect 7190 8412 7196 8424
rect 6687 8384 7196 8412
rect 6687 8381 6699 8384
rect 6641 8375 6699 8381
rect 7190 8372 7196 8384
rect 7248 8372 7254 8424
rect 8297 8415 8355 8421
rect 8297 8381 8309 8415
rect 8343 8412 8355 8415
rect 8478 8412 8484 8424
rect 8343 8384 8484 8412
rect 8343 8381 8355 8384
rect 8297 8375 8355 8381
rect 8478 8372 8484 8384
rect 8536 8412 8542 8424
rect 8846 8412 8852 8424
rect 8536 8384 8852 8412
rect 8536 8372 8542 8384
rect 8846 8372 8852 8384
rect 8904 8372 8910 8424
rect 16390 8372 16396 8424
rect 16448 8412 16454 8424
rect 16761 8415 16819 8421
rect 16761 8412 16773 8415
rect 16448 8384 16773 8412
rect 16448 8372 16454 8384
rect 16761 8381 16773 8384
rect 16807 8381 16819 8415
rect 16761 8375 16819 8381
rect 18782 8372 18788 8424
rect 18840 8412 18846 8424
rect 19426 8412 19432 8424
rect 18840 8384 19432 8412
rect 18840 8372 18846 8384
rect 19426 8372 19432 8384
rect 19484 8412 19490 8424
rect 19981 8415 20039 8421
rect 19981 8412 19993 8415
rect 19484 8384 19993 8412
rect 19484 8372 19490 8384
rect 19981 8381 19993 8384
rect 20027 8381 20039 8415
rect 19981 8375 20039 8381
rect 21358 8372 21364 8424
rect 21416 8412 21422 8424
rect 21545 8415 21603 8421
rect 21545 8412 21557 8415
rect 21416 8384 21557 8412
rect 21416 8372 21422 8384
rect 21545 8381 21557 8384
rect 21591 8381 21603 8415
rect 21545 8375 21603 8381
rect 21634 8372 21640 8424
rect 21692 8412 21698 8424
rect 25317 8415 25375 8421
rect 21692 8384 21737 8412
rect 21692 8372 21698 8384
rect 25317 8381 25329 8415
rect 25363 8412 25375 8415
rect 25774 8412 25780 8424
rect 25363 8384 25780 8412
rect 25363 8381 25375 8384
rect 25317 8375 25375 8381
rect 25774 8372 25780 8384
rect 25832 8372 25838 8424
rect 26418 8412 26424 8424
rect 26379 8384 26424 8412
rect 26418 8372 26424 8384
rect 26476 8412 26482 8424
rect 26973 8415 27031 8421
rect 26973 8412 26985 8415
rect 26476 8384 26985 8412
rect 26476 8372 26482 8384
rect 26973 8381 26985 8384
rect 27019 8381 27031 8415
rect 26973 8375 27031 8381
rect 27338 8372 27344 8424
rect 27396 8412 27402 8424
rect 27525 8415 27583 8421
rect 27525 8412 27537 8415
rect 27396 8384 27537 8412
rect 27396 8372 27402 8384
rect 27525 8381 27537 8384
rect 27571 8412 27583 8415
rect 28077 8415 28135 8421
rect 28077 8412 28089 8415
rect 27571 8384 28089 8412
rect 27571 8381 27583 8384
rect 27525 8375 27583 8381
rect 28077 8381 28089 8384
rect 28123 8381 28135 8415
rect 28077 8375 28135 8381
rect 2130 8344 2136 8356
rect 2091 8316 2136 8344
rect 2130 8304 2136 8316
rect 2188 8304 2194 8356
rect 4157 8347 4215 8353
rect 4157 8313 4169 8347
rect 4203 8313 4215 8347
rect 4157 8307 4215 8313
rect 1765 8279 1823 8285
rect 1765 8245 1777 8279
rect 1811 8276 1823 8279
rect 2314 8276 2320 8288
rect 1811 8248 2320 8276
rect 1811 8245 1823 8248
rect 1765 8239 1823 8245
rect 2314 8236 2320 8248
rect 2372 8236 2378 8288
rect 3694 8236 3700 8288
rect 3752 8276 3758 8288
rect 4172 8276 4200 8307
rect 4706 8304 4712 8356
rect 4764 8344 4770 8356
rect 4893 8347 4951 8353
rect 4893 8344 4905 8347
rect 4764 8316 4905 8344
rect 4764 8304 4770 8316
rect 4893 8313 4905 8316
rect 4939 8344 4951 8347
rect 6546 8344 6552 8356
rect 4939 8316 6552 8344
rect 4939 8313 4951 8316
rect 4893 8307 4951 8313
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 17497 8347 17555 8353
rect 17497 8313 17509 8347
rect 17543 8344 17555 8347
rect 18509 8347 18567 8353
rect 18509 8344 18521 8347
rect 17543 8316 18521 8344
rect 17543 8313 17555 8316
rect 17497 8307 17555 8313
rect 18509 8313 18521 8316
rect 18555 8344 18567 8347
rect 21085 8347 21143 8353
rect 18555 8316 19656 8344
rect 18555 8313 18567 8316
rect 18509 8307 18567 8313
rect 5258 8276 5264 8288
rect 3752 8248 4200 8276
rect 5219 8248 5264 8276
rect 3752 8236 3758 8248
rect 5258 8236 5264 8248
rect 5316 8236 5322 8288
rect 8386 8236 8392 8288
rect 8444 8276 8450 8288
rect 8757 8279 8815 8285
rect 8757 8276 8769 8279
rect 8444 8248 8769 8276
rect 8444 8236 8450 8248
rect 8757 8245 8769 8248
rect 8803 8245 8815 8279
rect 16390 8276 16396 8288
rect 16351 8248 16396 8276
rect 8757 8239 8815 8245
rect 16390 8236 16396 8248
rect 16448 8236 16454 8288
rect 17862 8236 17868 8288
rect 17920 8276 17926 8288
rect 18049 8279 18107 8285
rect 18049 8276 18061 8279
rect 17920 8248 18061 8276
rect 17920 8236 17926 8248
rect 18049 8245 18061 8248
rect 18095 8245 18107 8279
rect 18414 8276 18420 8288
rect 18375 8248 18420 8276
rect 18049 8239 18107 8245
rect 18414 8236 18420 8248
rect 18472 8236 18478 8288
rect 19628 8285 19656 8316
rect 21085 8313 21097 8347
rect 21131 8344 21143 8347
rect 21652 8344 21680 8372
rect 21131 8316 21680 8344
rect 21131 8313 21143 8316
rect 21085 8307 21143 8313
rect 19613 8279 19671 8285
rect 19613 8245 19625 8279
rect 19659 8245 19671 8279
rect 25498 8276 25504 8288
rect 25459 8248 25504 8276
rect 19613 8239 19671 8245
rect 25498 8236 25504 8248
rect 25556 8236 25562 8288
rect 1104 8186 28888 8208
rect 1104 8134 10982 8186
rect 11034 8134 11046 8186
rect 11098 8134 11110 8186
rect 11162 8134 11174 8186
rect 11226 8134 20982 8186
rect 21034 8134 21046 8186
rect 21098 8134 21110 8186
rect 21162 8134 21174 8186
rect 21226 8134 28888 8186
rect 1104 8112 28888 8134
rect 1670 8072 1676 8084
rect 1631 8044 1676 8072
rect 1670 8032 1676 8044
rect 1728 8032 1734 8084
rect 1762 8032 1768 8084
rect 1820 8072 1826 8084
rect 1949 8075 2007 8081
rect 1949 8072 1961 8075
rect 1820 8044 1961 8072
rect 1820 8032 1826 8044
rect 1949 8041 1961 8044
rect 1995 8041 2007 8075
rect 1949 8035 2007 8041
rect 2866 8032 2872 8084
rect 2924 8072 2930 8084
rect 3694 8072 3700 8084
rect 2924 8044 3700 8072
rect 2924 8032 2930 8044
rect 3694 8032 3700 8044
rect 3752 8072 3758 8084
rect 3789 8075 3847 8081
rect 3789 8072 3801 8075
rect 3752 8044 3801 8072
rect 3752 8032 3758 8044
rect 3789 8041 3801 8044
rect 3835 8041 3847 8075
rect 3789 8035 3847 8041
rect 3878 8032 3884 8084
rect 3936 8072 3942 8084
rect 4065 8075 4123 8081
rect 4065 8072 4077 8075
rect 3936 8044 4077 8072
rect 3936 8032 3942 8044
rect 4065 8041 4077 8044
rect 4111 8041 4123 8075
rect 4430 8072 4436 8084
rect 4391 8044 4436 8072
rect 4065 8035 4123 8041
rect 4430 8032 4436 8044
rect 4488 8032 4494 8084
rect 6365 8075 6423 8081
rect 6365 8041 6377 8075
rect 6411 8072 6423 8075
rect 6638 8072 6644 8084
rect 6411 8044 6644 8072
rect 6411 8041 6423 8044
rect 6365 8035 6423 8041
rect 6638 8032 6644 8044
rect 6696 8032 6702 8084
rect 6822 8072 6828 8084
rect 6783 8044 6828 8072
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 7374 8072 7380 8084
rect 7335 8044 7380 8072
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 16209 8075 16267 8081
rect 16209 8041 16221 8075
rect 16255 8072 16267 8075
rect 16298 8072 16304 8084
rect 16255 8044 16304 8072
rect 16255 8041 16267 8044
rect 16209 8035 16267 8041
rect 16298 8032 16304 8044
rect 16356 8032 16362 8084
rect 16577 8075 16635 8081
rect 16577 8041 16589 8075
rect 16623 8072 16635 8075
rect 17770 8072 17776 8084
rect 16623 8044 17776 8072
rect 16623 8041 16635 8044
rect 16577 8035 16635 8041
rect 17770 8032 17776 8044
rect 17828 8032 17834 8084
rect 18785 8075 18843 8081
rect 18785 8041 18797 8075
rect 18831 8072 18843 8075
rect 19150 8072 19156 8084
rect 18831 8044 19156 8072
rect 18831 8041 18843 8044
rect 18785 8035 18843 8041
rect 19150 8032 19156 8044
rect 19208 8032 19214 8084
rect 19334 8032 19340 8084
rect 19392 8072 19398 8084
rect 19705 8075 19763 8081
rect 19705 8072 19717 8075
rect 19392 8044 19717 8072
rect 19392 8032 19398 8044
rect 19705 8041 19717 8044
rect 19751 8072 19763 8075
rect 20346 8072 20352 8084
rect 19751 8044 20352 8072
rect 19751 8041 19763 8044
rect 19705 8035 19763 8041
rect 20346 8032 20352 8044
rect 20404 8032 20410 8084
rect 21269 8075 21327 8081
rect 21269 8041 21281 8075
rect 21315 8072 21327 8075
rect 21358 8072 21364 8084
rect 21315 8044 21364 8072
rect 21315 8041 21327 8044
rect 21269 8035 21327 8041
rect 21358 8032 21364 8044
rect 21416 8032 21422 8084
rect 21542 8072 21548 8084
rect 21503 8044 21548 8072
rect 21542 8032 21548 8044
rect 21600 8032 21606 8084
rect 21726 8032 21732 8084
rect 21784 8072 21790 8084
rect 21913 8075 21971 8081
rect 21913 8072 21925 8075
rect 21784 8044 21925 8072
rect 21784 8032 21790 8044
rect 21913 8041 21925 8044
rect 21959 8041 21971 8075
rect 21913 8035 21971 8041
rect 2406 7964 2412 8016
rect 2464 7964 2470 8016
rect 2682 7964 2688 8016
rect 2740 8004 2746 8016
rect 2740 7976 3096 8004
rect 2740 7964 2746 7976
rect 2314 7936 2320 7948
rect 2275 7908 2320 7936
rect 2314 7896 2320 7908
rect 2372 7896 2378 7948
rect 2424 7936 2452 7964
rect 2424 7908 2544 7936
rect 2406 7868 2412 7880
rect 2367 7840 2412 7868
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 2516 7877 2544 7908
rect 2501 7871 2559 7877
rect 2501 7837 2513 7871
rect 2547 7868 2559 7871
rect 2682 7868 2688 7880
rect 2547 7840 2688 7868
rect 2547 7837 2559 7840
rect 2501 7831 2559 7837
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 3068 7877 3096 7976
rect 3142 7964 3148 8016
rect 3200 8004 3206 8016
rect 3329 8007 3387 8013
rect 3329 8004 3341 8007
rect 3200 7976 3341 8004
rect 3200 7964 3206 7976
rect 3329 7973 3341 7976
rect 3375 7973 3387 8007
rect 4522 8004 4528 8016
rect 4435 7976 4528 8004
rect 3329 7967 3387 7973
rect 4522 7964 4528 7976
rect 4580 8004 4586 8016
rect 8938 8004 8944 8016
rect 4580 7976 8944 8004
rect 4580 7964 4586 7976
rect 8938 7964 8944 7976
rect 8996 7964 9002 8016
rect 19242 7964 19248 8016
rect 19300 8004 19306 8016
rect 19613 8007 19671 8013
rect 19613 8004 19625 8007
rect 19300 7976 19625 8004
rect 19300 7964 19306 7976
rect 19613 7973 19625 7976
rect 19659 7973 19671 8007
rect 20254 8004 20260 8016
rect 20215 7976 20260 8004
rect 19613 7967 19671 7973
rect 20254 7964 20260 7976
rect 20312 7964 20318 8016
rect 6730 7936 6736 7948
rect 6691 7908 6736 7936
rect 6730 7896 6736 7908
rect 6788 7896 6794 7948
rect 16574 7896 16580 7948
rect 16632 7936 16638 7948
rect 17034 7945 17040 7948
rect 16761 7939 16819 7945
rect 16761 7936 16773 7939
rect 16632 7908 16773 7936
rect 16632 7896 16638 7908
rect 16761 7905 16773 7908
rect 16807 7905 16819 7939
rect 17028 7936 17040 7945
rect 16995 7908 17040 7936
rect 16761 7899 16819 7905
rect 17028 7899 17040 7908
rect 17034 7896 17040 7899
rect 17092 7896 17098 7948
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3326 7868 3332 7880
rect 3099 7840 3332 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3326 7828 3332 7840
rect 3384 7828 3390 7880
rect 4706 7868 4712 7880
rect 4619 7840 4712 7868
rect 4706 7828 4712 7840
rect 4764 7868 4770 7880
rect 5258 7868 5264 7880
rect 4764 7840 5264 7868
rect 4764 7828 4770 7840
rect 5258 7828 5264 7840
rect 5316 7868 5322 7880
rect 6273 7871 6331 7877
rect 6273 7868 6285 7871
rect 5316 7840 6285 7868
rect 5316 7828 5322 7840
rect 6273 7837 6285 7840
rect 6319 7868 6331 7871
rect 6362 7868 6368 7880
rect 6319 7840 6368 7868
rect 6319 7837 6331 7840
rect 6273 7831 6331 7837
rect 6362 7828 6368 7840
rect 6420 7868 6426 7880
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 6420 7840 7021 7868
rect 6420 7828 6426 7840
rect 7009 7837 7021 7840
rect 7055 7868 7067 7871
rect 7466 7868 7472 7880
rect 7055 7840 7472 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 19058 7868 19064 7880
rect 19019 7840 19064 7868
rect 19058 7828 19064 7840
rect 19116 7828 19122 7880
rect 19794 7828 19800 7880
rect 19852 7868 19858 7880
rect 19889 7871 19947 7877
rect 19889 7868 19901 7871
rect 19852 7840 19901 7868
rect 19852 7828 19858 7840
rect 19889 7837 19901 7840
rect 19935 7868 19947 7871
rect 20272 7868 20300 7964
rect 26234 7896 26240 7948
rect 26292 7936 26298 7948
rect 26513 7939 26571 7945
rect 26513 7936 26525 7939
rect 26292 7908 26525 7936
rect 26292 7896 26298 7908
rect 26513 7905 26525 7908
rect 26559 7936 26571 7939
rect 26970 7936 26976 7948
rect 26559 7908 26976 7936
rect 26559 7905 26571 7908
rect 26513 7899 26571 7905
rect 26970 7896 26976 7908
rect 27028 7896 27034 7948
rect 19935 7840 20300 7868
rect 19935 7837 19947 7840
rect 19889 7831 19947 7837
rect 18414 7760 18420 7812
rect 18472 7800 18478 7812
rect 19245 7803 19303 7809
rect 19245 7800 19257 7803
rect 18472 7772 19257 7800
rect 18472 7760 18478 7772
rect 19245 7769 19257 7772
rect 19291 7769 19303 7803
rect 19245 7763 19303 7769
rect 7742 7732 7748 7744
rect 7703 7704 7748 7732
rect 7742 7692 7748 7704
rect 7800 7692 7806 7744
rect 8110 7692 8116 7744
rect 8168 7732 8174 7744
rect 8386 7732 8392 7744
rect 8168 7704 8392 7732
rect 8168 7692 8174 7704
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 18141 7735 18199 7741
rect 18141 7701 18153 7735
rect 18187 7732 18199 7735
rect 18690 7732 18696 7744
rect 18187 7704 18696 7732
rect 18187 7701 18199 7704
rect 18141 7695 18199 7701
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 26697 7735 26755 7741
rect 26697 7701 26709 7735
rect 26743 7732 26755 7735
rect 26786 7732 26792 7744
rect 26743 7704 26792 7732
rect 26743 7701 26755 7704
rect 26697 7695 26755 7701
rect 26786 7692 26792 7704
rect 26844 7692 26850 7744
rect 1104 7642 28888 7664
rect 1104 7590 5982 7642
rect 6034 7590 6046 7642
rect 6098 7590 6110 7642
rect 6162 7590 6174 7642
rect 6226 7590 15982 7642
rect 16034 7590 16046 7642
rect 16098 7590 16110 7642
rect 16162 7590 16174 7642
rect 16226 7590 25982 7642
rect 26034 7590 26046 7642
rect 26098 7590 26110 7642
rect 26162 7590 26174 7642
rect 26226 7590 28888 7642
rect 1104 7568 28888 7590
rect 2409 7531 2467 7537
rect 2409 7497 2421 7531
rect 2455 7528 2467 7531
rect 2682 7528 2688 7540
rect 2455 7500 2688 7528
rect 2455 7497 2467 7500
rect 2409 7491 2467 7497
rect 2682 7488 2688 7500
rect 2740 7488 2746 7540
rect 3510 7528 3516 7540
rect 3471 7500 3516 7528
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 3786 7528 3792 7540
rect 3747 7500 3792 7528
rect 3786 7488 3792 7500
rect 3844 7488 3850 7540
rect 4249 7531 4307 7537
rect 4249 7497 4261 7531
rect 4295 7528 4307 7531
rect 4430 7528 4436 7540
rect 4295 7500 4436 7528
rect 4295 7497 4307 7500
rect 4249 7491 4307 7497
rect 4430 7488 4436 7500
rect 4488 7488 4494 7540
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 5350 7528 5356 7540
rect 4580 7500 4625 7528
rect 5311 7500 5356 7528
rect 4580 7488 4586 7500
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 6270 7488 6276 7540
rect 6328 7528 6334 7540
rect 6457 7531 6515 7537
rect 6457 7528 6469 7531
rect 6328 7500 6469 7528
rect 6328 7488 6334 7500
rect 6457 7497 6469 7500
rect 6503 7528 6515 7531
rect 6549 7531 6607 7537
rect 6549 7528 6561 7531
rect 6503 7500 6561 7528
rect 6503 7497 6515 7500
rect 6457 7491 6515 7497
rect 6549 7497 6561 7500
rect 6595 7497 6607 7531
rect 6549 7491 6607 7497
rect 6730 7488 6736 7540
rect 6788 7528 6794 7540
rect 6917 7531 6975 7537
rect 6917 7528 6929 7531
rect 6788 7500 6929 7528
rect 6788 7488 6794 7500
rect 6917 7497 6929 7500
rect 6963 7528 6975 7531
rect 7929 7531 7987 7537
rect 7929 7528 7941 7531
rect 6963 7500 7941 7528
rect 6963 7497 6975 7500
rect 6917 7491 6975 7497
rect 7929 7497 7941 7500
rect 7975 7497 7987 7531
rect 7929 7491 7987 7497
rect 15933 7531 15991 7537
rect 15933 7497 15945 7531
rect 15979 7528 15991 7531
rect 16390 7528 16396 7540
rect 15979 7500 16396 7528
rect 15979 7497 15991 7500
rect 15933 7491 15991 7497
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 17405 7531 17463 7537
rect 17405 7528 17417 7531
rect 16632 7500 17417 7528
rect 16632 7488 16638 7500
rect 17405 7497 17417 7500
rect 17451 7497 17463 7531
rect 17405 7491 17463 7497
rect 17865 7531 17923 7537
rect 17865 7497 17877 7531
rect 17911 7528 17923 7531
rect 18414 7528 18420 7540
rect 17911 7500 18420 7528
rect 17911 7497 17923 7500
rect 17865 7491 17923 7497
rect 18414 7488 18420 7500
rect 18472 7488 18478 7540
rect 19242 7528 19248 7540
rect 19203 7500 19248 7528
rect 19242 7488 19248 7500
rect 19300 7488 19306 7540
rect 19337 7531 19395 7537
rect 19337 7497 19349 7531
rect 19383 7528 19395 7531
rect 19426 7528 19432 7540
rect 19383 7500 19432 7528
rect 19383 7497 19395 7500
rect 19337 7491 19395 7497
rect 19426 7488 19432 7500
rect 19484 7488 19490 7540
rect 20346 7528 20352 7540
rect 20307 7500 20352 7528
rect 20346 7488 20352 7500
rect 20404 7488 20410 7540
rect 26970 7528 26976 7540
rect 26931 7500 26976 7528
rect 26970 7488 26976 7500
rect 27028 7488 27034 7540
rect 4062 7420 4068 7472
rect 4120 7460 4126 7472
rect 4893 7463 4951 7469
rect 4893 7460 4905 7463
rect 4120 7432 4905 7460
rect 4120 7420 4126 7432
rect 4893 7429 4905 7432
rect 4939 7429 4951 7463
rect 4893 7423 4951 7429
rect 5905 7463 5963 7469
rect 5905 7429 5917 7463
rect 5951 7460 5963 7463
rect 6822 7460 6828 7472
rect 5951 7432 6828 7460
rect 5951 7429 5963 7432
rect 5905 7423 5963 7429
rect 6822 7420 6828 7432
rect 6880 7420 6886 7472
rect 17770 7420 17776 7472
rect 17828 7460 17834 7472
rect 18509 7463 18567 7469
rect 18509 7460 18521 7463
rect 17828 7432 18521 7460
rect 17828 7420 17834 7432
rect 18509 7429 18521 7432
rect 18555 7460 18567 7463
rect 19794 7460 19800 7472
rect 18555 7432 19800 7460
rect 18555 7429 18567 7432
rect 18509 7423 18567 7429
rect 19794 7420 19800 7432
rect 19852 7420 19858 7472
rect 26329 7463 26387 7469
rect 26329 7429 26341 7463
rect 26375 7460 26387 7463
rect 27430 7460 27436 7472
rect 26375 7432 27436 7460
rect 26375 7429 26387 7432
rect 26329 7423 26387 7429
rect 2038 7352 2044 7404
rect 2096 7352 2102 7404
rect 6273 7395 6331 7401
rect 6273 7361 6285 7395
rect 6319 7392 6331 7395
rect 7561 7395 7619 7401
rect 7561 7392 7573 7395
rect 6319 7364 7573 7392
rect 6319 7361 6331 7364
rect 6273 7355 6331 7361
rect 7561 7361 7573 7364
rect 7607 7392 7619 7395
rect 7742 7392 7748 7404
rect 7607 7364 7748 7392
rect 7607 7361 7619 7364
rect 7561 7355 7619 7361
rect 7742 7352 7748 7364
rect 7800 7392 7806 7404
rect 8202 7392 8208 7404
rect 7800 7364 8208 7392
rect 7800 7352 7806 7364
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 16301 7395 16359 7401
rect 16301 7361 16313 7395
rect 16347 7392 16359 7395
rect 17037 7395 17095 7401
rect 17037 7392 17049 7395
rect 16347 7364 17049 7392
rect 16347 7361 16359 7364
rect 16301 7355 16359 7361
rect 17037 7361 17049 7364
rect 17083 7392 17095 7395
rect 18690 7392 18696 7404
rect 17083 7364 18696 7392
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 18690 7352 18696 7364
rect 18748 7352 18754 7404
rect 19150 7352 19156 7404
rect 19208 7392 19214 7404
rect 19702 7392 19708 7404
rect 19208 7364 19708 7392
rect 19208 7352 19214 7364
rect 19702 7352 19708 7364
rect 19760 7392 19766 7404
rect 19889 7395 19947 7401
rect 19889 7392 19901 7395
rect 19760 7364 19901 7392
rect 19760 7352 19766 7364
rect 19889 7361 19901 7364
rect 19935 7361 19947 7395
rect 19889 7355 19947 7361
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7293 1455 7327
rect 2056 7324 2084 7352
rect 2501 7327 2559 7333
rect 2501 7324 2513 7327
rect 2056 7296 2513 7324
rect 1397 7287 1455 7293
rect 2501 7293 2513 7296
rect 2547 7324 2559 7327
rect 3053 7327 3111 7333
rect 3053 7324 3065 7327
rect 2547 7296 3065 7324
rect 2547 7293 2559 7296
rect 2501 7287 2559 7293
rect 3053 7293 3065 7296
rect 3099 7293 3111 7327
rect 3053 7287 3111 7293
rect 1412 7256 1440 7287
rect 3510 7284 3516 7336
rect 3568 7324 3574 7336
rect 3605 7327 3663 7333
rect 3605 7324 3617 7327
rect 3568 7296 3617 7324
rect 3568 7284 3574 7296
rect 3605 7293 3617 7296
rect 3651 7293 3663 7327
rect 3605 7287 3663 7293
rect 4709 7327 4767 7333
rect 4709 7293 4721 7327
rect 4755 7324 4767 7327
rect 5350 7324 5356 7336
rect 4755 7296 5356 7324
rect 4755 7293 4767 7296
rect 4709 7287 4767 7293
rect 5350 7284 5356 7296
rect 5408 7284 5414 7336
rect 6457 7327 6515 7333
rect 6457 7293 6469 7327
rect 6503 7324 6515 7327
rect 7377 7327 7435 7333
rect 7377 7324 7389 7327
rect 6503 7296 7389 7324
rect 6503 7293 6515 7296
rect 6457 7287 6515 7293
rect 7377 7293 7389 7296
rect 7423 7293 7435 7327
rect 7377 7287 7435 7293
rect 16390 7284 16396 7336
rect 16448 7324 16454 7336
rect 16761 7327 16819 7333
rect 16761 7324 16773 7327
rect 16448 7296 16773 7324
rect 16448 7284 16454 7296
rect 16761 7293 16773 7296
rect 16807 7293 16819 7327
rect 16761 7287 16819 7293
rect 16850 7284 16856 7336
rect 16908 7324 16914 7336
rect 17862 7324 17868 7336
rect 16908 7296 17868 7324
rect 16908 7284 16914 7296
rect 17862 7284 17868 7296
rect 17920 7284 17926 7336
rect 19426 7284 19432 7336
rect 19484 7324 19490 7336
rect 26436 7333 26464 7432
rect 27430 7420 27436 7432
rect 27488 7420 27494 7472
rect 19797 7327 19855 7333
rect 19797 7324 19809 7327
rect 19484 7296 19809 7324
rect 19484 7284 19490 7296
rect 19797 7293 19809 7296
rect 19843 7324 19855 7327
rect 26421 7327 26479 7333
rect 26421 7324 26433 7327
rect 19843 7296 26433 7324
rect 19843 7293 19855 7296
rect 19797 7287 19855 7293
rect 26421 7293 26433 7296
rect 26467 7293 26479 7327
rect 26421 7287 26479 7293
rect 27062 7284 27068 7336
rect 27120 7324 27126 7336
rect 27525 7327 27583 7333
rect 27525 7324 27537 7327
rect 27120 7296 27537 7324
rect 27120 7284 27126 7296
rect 27525 7293 27537 7296
rect 27571 7324 27583 7327
rect 28077 7327 28135 7333
rect 28077 7324 28089 7327
rect 27571 7296 28089 7324
rect 27571 7293 27583 7296
rect 27525 7287 27583 7293
rect 28077 7293 28089 7296
rect 28123 7293 28135 7327
rect 28077 7287 28135 7293
rect 2038 7256 2044 7268
rect 1412 7228 2044 7256
rect 2038 7216 2044 7228
rect 2096 7216 2102 7268
rect 18877 7259 18935 7265
rect 18877 7225 18889 7259
rect 18923 7256 18935 7259
rect 19610 7256 19616 7268
rect 18923 7228 19616 7256
rect 18923 7225 18935 7228
rect 18877 7219 18935 7225
rect 19610 7216 19616 7228
rect 19668 7256 19674 7268
rect 19705 7259 19763 7265
rect 19705 7256 19717 7259
rect 19668 7228 19717 7256
rect 19668 7216 19674 7228
rect 19705 7225 19717 7228
rect 19751 7225 19763 7259
rect 19705 7219 19763 7225
rect 1581 7191 1639 7197
rect 1581 7157 1593 7191
rect 1627 7188 1639 7191
rect 1670 7188 1676 7200
rect 1627 7160 1676 7188
rect 1627 7157 1639 7160
rect 1581 7151 1639 7157
rect 1670 7148 1676 7160
rect 1728 7148 1734 7200
rect 2682 7188 2688 7200
rect 2643 7160 2688 7188
rect 2682 7148 2688 7160
rect 2740 7148 2746 7200
rect 6914 7148 6920 7200
rect 6972 7188 6978 7200
rect 7285 7191 7343 7197
rect 7285 7188 7297 7191
rect 6972 7160 7297 7188
rect 6972 7148 6978 7160
rect 7285 7157 7297 7160
rect 7331 7188 7343 7191
rect 7834 7188 7840 7200
rect 7331 7160 7840 7188
rect 7331 7157 7343 7160
rect 7285 7151 7343 7157
rect 7834 7148 7840 7160
rect 7892 7148 7898 7200
rect 16390 7188 16396 7200
rect 16351 7160 16396 7188
rect 16390 7148 16396 7160
rect 16448 7148 16454 7200
rect 26326 7148 26332 7200
rect 26384 7188 26390 7200
rect 26605 7191 26663 7197
rect 26605 7188 26617 7191
rect 26384 7160 26617 7188
rect 26384 7148 26390 7160
rect 26605 7157 26617 7160
rect 26651 7157 26663 7191
rect 27706 7188 27712 7200
rect 27667 7160 27712 7188
rect 26605 7151 26663 7157
rect 27706 7148 27712 7160
rect 27764 7148 27770 7200
rect 1104 7098 28888 7120
rect 1104 7046 10982 7098
rect 11034 7046 11046 7098
rect 11098 7046 11110 7098
rect 11162 7046 11174 7098
rect 11226 7046 20982 7098
rect 21034 7046 21046 7098
rect 21098 7046 21110 7098
rect 21162 7046 21174 7098
rect 21226 7046 28888 7098
rect 1104 7024 28888 7046
rect 4341 6987 4399 6993
rect 4341 6953 4353 6987
rect 4387 6984 4399 6987
rect 4706 6984 4712 6996
rect 4387 6956 4712 6984
rect 4387 6953 4399 6956
rect 4341 6947 4399 6953
rect 4706 6944 4712 6956
rect 4764 6944 4770 6996
rect 6362 6984 6368 6996
rect 6323 6956 6368 6984
rect 6362 6944 6368 6956
rect 6420 6944 6426 6996
rect 16761 6987 16819 6993
rect 16761 6953 16773 6987
rect 16807 6984 16819 6987
rect 17034 6984 17040 6996
rect 16807 6956 17040 6984
rect 16807 6953 16819 6956
rect 16761 6947 16819 6953
rect 17034 6944 17040 6956
rect 17092 6944 17098 6996
rect 19426 6984 19432 6996
rect 19387 6956 19432 6984
rect 19426 6944 19432 6956
rect 19484 6944 19490 6996
rect 19702 6984 19708 6996
rect 19663 6956 19708 6984
rect 19702 6944 19708 6956
rect 19760 6944 19766 6996
rect 566 6876 572 6928
rect 624 6916 630 6928
rect 8662 6916 8668 6928
rect 624 6888 8668 6916
rect 624 6876 630 6888
rect 8662 6876 8668 6888
rect 8720 6876 8726 6928
rect 16850 6916 16856 6928
rect 16592 6888 16856 6916
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 2038 6848 2044 6860
rect 1443 6820 2044 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 2038 6808 2044 6820
rect 2096 6808 2102 6860
rect 2130 6808 2136 6860
rect 2188 6848 2194 6860
rect 2317 6851 2375 6857
rect 2317 6848 2329 6851
rect 2188 6820 2329 6848
rect 2188 6808 2194 6820
rect 2317 6817 2329 6820
rect 2363 6817 2375 6851
rect 2501 6851 2559 6857
rect 2501 6848 2513 6851
rect 2317 6811 2375 6817
rect 2424 6820 2513 6848
rect 1946 6780 1952 6792
rect 1907 6752 1952 6780
rect 1946 6740 1952 6752
rect 2004 6740 2010 6792
rect 2424 6724 2452 6820
rect 2501 6817 2513 6820
rect 2547 6817 2559 6851
rect 3050 6848 3056 6860
rect 3011 6820 3056 6848
rect 2501 6811 2559 6817
rect 3050 6808 3056 6820
rect 3108 6808 3114 6860
rect 3510 6848 3516 6860
rect 3471 6820 3516 6848
rect 3510 6808 3516 6820
rect 3568 6808 3574 6860
rect 15381 6851 15439 6857
rect 15381 6817 15393 6851
rect 15427 6848 15439 6851
rect 15470 6848 15476 6860
rect 15427 6820 15476 6848
rect 15427 6817 15439 6820
rect 15381 6811 15439 6817
rect 15470 6808 15476 6820
rect 15528 6848 15534 6860
rect 16390 6848 16396 6860
rect 15528 6820 16396 6848
rect 15528 6808 15534 6820
rect 16390 6808 16396 6820
rect 16448 6808 16454 6860
rect 16485 6851 16543 6857
rect 16485 6817 16497 6851
rect 16531 6848 16543 6851
rect 16592 6848 16620 6888
rect 16850 6876 16856 6888
rect 16908 6876 16914 6928
rect 26510 6848 26516 6860
rect 16531 6820 16620 6848
rect 26471 6820 26516 6848
rect 16531 6817 16543 6820
rect 16485 6811 16543 6817
rect 26510 6808 26516 6820
rect 26568 6808 26574 6860
rect 1394 6672 1400 6724
rect 1452 6712 1458 6724
rect 2406 6712 2412 6724
rect 1452 6684 2412 6712
rect 1452 6672 1458 6684
rect 2406 6672 2412 6684
rect 2464 6672 2470 6724
rect 2498 6672 2504 6724
rect 2556 6712 2562 6724
rect 2685 6715 2743 6721
rect 2685 6712 2697 6715
rect 2556 6684 2697 6712
rect 2556 6672 2562 6684
rect 2685 6681 2697 6684
rect 2731 6681 2743 6715
rect 2685 6675 2743 6681
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 6914 6644 6920 6656
rect 6875 6616 6920 6644
rect 6914 6604 6920 6616
rect 6972 6604 6978 6656
rect 15562 6644 15568 6656
rect 15523 6616 15568 6644
rect 15562 6604 15568 6616
rect 15620 6604 15626 6656
rect 26694 6644 26700 6656
rect 26655 6616 26700 6644
rect 26694 6604 26700 6616
rect 26752 6604 26758 6656
rect 1104 6554 28888 6576
rect 1104 6502 5982 6554
rect 6034 6502 6046 6554
rect 6098 6502 6110 6554
rect 6162 6502 6174 6554
rect 6226 6502 15982 6554
rect 16034 6502 16046 6554
rect 16098 6502 16110 6554
rect 16162 6502 16174 6554
rect 16226 6502 25982 6554
rect 26034 6502 26046 6554
rect 26098 6502 26110 6554
rect 26162 6502 26174 6554
rect 26226 6502 28888 6554
rect 1104 6480 28888 6502
rect 1486 6400 1492 6452
rect 1544 6440 1550 6452
rect 1581 6443 1639 6449
rect 1581 6440 1593 6443
rect 1544 6412 1593 6440
rect 1544 6400 1550 6412
rect 1581 6409 1593 6412
rect 1627 6409 1639 6443
rect 1581 6403 1639 6409
rect 2406 6400 2412 6452
rect 2464 6440 2470 6452
rect 3053 6443 3111 6449
rect 3053 6440 3065 6443
rect 2464 6412 3065 6440
rect 2464 6400 2470 6412
rect 3053 6409 3065 6412
rect 3099 6409 3111 6443
rect 15470 6440 15476 6452
rect 15431 6412 15476 6440
rect 3053 6403 3111 6409
rect 15470 6400 15476 6412
rect 15528 6400 15534 6452
rect 26510 6440 26516 6452
rect 26471 6412 26516 6440
rect 26510 6400 26516 6412
rect 26568 6400 26574 6452
rect 2038 6372 2044 6384
rect 1951 6344 2044 6372
rect 2038 6332 2044 6344
rect 2096 6372 2102 6384
rect 4522 6372 4528 6384
rect 2096 6344 4528 6372
rect 2096 6332 2102 6344
rect 4522 6332 4528 6344
rect 4580 6332 4586 6384
rect 2406 6304 2412 6316
rect 1412 6276 2412 6304
rect 1412 6245 1440 6276
rect 2406 6264 2412 6276
rect 2464 6264 2470 6316
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6205 1455 6239
rect 1397 6199 1455 6205
rect 2501 6239 2559 6245
rect 2501 6205 2513 6239
rect 2547 6236 2559 6239
rect 2590 6236 2596 6248
rect 2547 6208 2596 6236
rect 2547 6205 2559 6208
rect 2501 6199 2559 6205
rect 2590 6196 2596 6208
rect 2648 6196 2654 6248
rect 2682 6100 2688 6112
rect 2643 6072 2688 6100
rect 2682 6060 2688 6072
rect 2740 6060 2746 6112
rect 1104 6010 28888 6032
rect 1104 5958 10982 6010
rect 11034 5958 11046 6010
rect 11098 5958 11110 6010
rect 11162 5958 11174 6010
rect 11226 5958 20982 6010
rect 21034 5958 21046 6010
rect 21098 5958 21110 6010
rect 21162 5958 21174 6010
rect 21226 5958 28888 6010
rect 1104 5936 28888 5958
rect 2041 5899 2099 5905
rect 2041 5865 2053 5899
rect 2087 5896 2099 5899
rect 2314 5896 2320 5908
rect 2087 5868 2320 5896
rect 2087 5865 2099 5868
rect 2041 5859 2099 5865
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 2590 5896 2596 5908
rect 2551 5868 2596 5896
rect 2590 5856 2596 5868
rect 2648 5856 2654 5908
rect 1394 5760 1400 5772
rect 1355 5732 1400 5760
rect 1394 5720 1400 5732
rect 1452 5720 1458 5772
rect 1486 5516 1492 5568
rect 1544 5556 1550 5568
rect 1581 5559 1639 5565
rect 1581 5556 1593 5559
rect 1544 5528 1593 5556
rect 1544 5516 1550 5528
rect 1581 5525 1593 5528
rect 1627 5525 1639 5559
rect 1581 5519 1639 5525
rect 1104 5466 28888 5488
rect 1104 5414 5982 5466
rect 6034 5414 6046 5466
rect 6098 5414 6110 5466
rect 6162 5414 6174 5466
rect 6226 5414 15982 5466
rect 16034 5414 16046 5466
rect 16098 5414 16110 5466
rect 16162 5414 16174 5466
rect 16226 5414 25982 5466
rect 26034 5414 26046 5466
rect 26098 5414 26110 5466
rect 26162 5414 26174 5466
rect 26226 5414 28888 5466
rect 1104 5392 28888 5414
rect 1394 5312 1400 5364
rect 1452 5352 1458 5364
rect 1581 5355 1639 5361
rect 1581 5352 1593 5355
rect 1452 5324 1593 5352
rect 1452 5312 1458 5324
rect 1581 5321 1593 5324
rect 1627 5321 1639 5355
rect 1581 5315 1639 5321
rect 26418 5148 26424 5160
rect 26379 5120 26424 5148
rect 26418 5108 26424 5120
rect 26476 5148 26482 5160
rect 26973 5151 27031 5157
rect 26973 5148 26985 5151
rect 26476 5120 26985 5148
rect 26476 5108 26482 5120
rect 26973 5117 26985 5120
rect 27019 5117 27031 5151
rect 26973 5111 27031 5117
rect 26602 5012 26608 5024
rect 26563 4984 26608 5012
rect 26602 4972 26608 4984
rect 26660 4972 26666 5024
rect 1104 4922 28888 4944
rect 1104 4870 10982 4922
rect 11034 4870 11046 4922
rect 11098 4870 11110 4922
rect 11162 4870 11174 4922
rect 11226 4870 20982 4922
rect 21034 4870 21046 4922
rect 21098 4870 21110 4922
rect 21162 4870 21174 4922
rect 21226 4870 28888 4922
rect 1104 4848 28888 4870
rect 1104 4378 28888 4400
rect 1104 4326 5982 4378
rect 6034 4326 6046 4378
rect 6098 4326 6110 4378
rect 6162 4326 6174 4378
rect 6226 4326 15982 4378
rect 16034 4326 16046 4378
rect 16098 4326 16110 4378
rect 16162 4326 16174 4378
rect 16226 4326 25982 4378
rect 26034 4326 26046 4378
rect 26098 4326 26110 4378
rect 26162 4326 26174 4378
rect 26226 4326 28888 4378
rect 1104 4304 28888 4326
rect 1104 3834 28888 3856
rect 1104 3782 10982 3834
rect 11034 3782 11046 3834
rect 11098 3782 11110 3834
rect 11162 3782 11174 3834
rect 11226 3782 20982 3834
rect 21034 3782 21046 3834
rect 21098 3782 21110 3834
rect 21162 3782 21174 3834
rect 21226 3782 28888 3834
rect 1104 3760 28888 3782
rect 1104 3290 28888 3312
rect 1104 3238 5982 3290
rect 6034 3238 6046 3290
rect 6098 3238 6110 3290
rect 6162 3238 6174 3290
rect 6226 3238 15982 3290
rect 16034 3238 16046 3290
rect 16098 3238 16110 3290
rect 16162 3238 16174 3290
rect 16226 3238 25982 3290
rect 26034 3238 26046 3290
rect 26098 3238 26110 3290
rect 26162 3238 26174 3290
rect 26226 3238 28888 3290
rect 1104 3216 28888 3238
rect 2038 3176 2044 3188
rect 1999 3148 2044 3176
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 2038 2972 2044 2984
rect 1443 2944 2044 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 26418 2972 26424 2984
rect 26379 2944 26424 2972
rect 26418 2932 26424 2944
rect 26476 2972 26482 2984
rect 26973 2975 27031 2981
rect 26973 2972 26985 2975
rect 26476 2944 26985 2972
rect 26476 2932 26482 2944
rect 26973 2941 26985 2944
rect 27019 2941 27031 2975
rect 26973 2935 27031 2941
rect 1578 2836 1584 2848
rect 1539 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 26602 2836 26608 2848
rect 26563 2808 26608 2836
rect 26602 2796 26608 2808
rect 26660 2796 26666 2848
rect 1104 2746 28888 2768
rect 1104 2694 10982 2746
rect 11034 2694 11046 2746
rect 11098 2694 11110 2746
rect 11162 2694 11174 2746
rect 11226 2694 20982 2746
rect 21034 2694 21046 2746
rect 21098 2694 21110 2746
rect 21162 2694 21174 2746
rect 21226 2694 28888 2746
rect 1104 2672 28888 2694
rect 6365 2635 6423 2641
rect 6365 2601 6377 2635
rect 6411 2632 6423 2635
rect 6546 2632 6552 2644
rect 6411 2604 6552 2632
rect 6411 2601 6423 2604
rect 6365 2595 6423 2601
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 8294 2592 8300 2644
rect 8352 2632 8358 2644
rect 8573 2635 8631 2641
rect 8573 2632 8585 2635
rect 8352 2604 8585 2632
rect 8352 2592 8358 2604
rect 8573 2601 8585 2604
rect 8619 2601 8631 2635
rect 8573 2595 8631 2601
rect 7466 2505 7472 2508
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 7460 2496 7472 2505
rect 6779 2468 7472 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 7460 2459 7472 2468
rect 7466 2456 7472 2459
rect 7524 2456 7530 2508
rect 6546 2388 6552 2440
rect 6604 2428 6610 2440
rect 7193 2431 7251 2437
rect 7193 2428 7205 2431
rect 6604 2400 7205 2428
rect 6604 2388 6610 2400
rect 7193 2397 7205 2400
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 1104 2202 28888 2224
rect 1104 2150 5982 2202
rect 6034 2150 6046 2202
rect 6098 2150 6110 2202
rect 6162 2150 6174 2202
rect 6226 2150 15982 2202
rect 16034 2150 16046 2202
rect 16098 2150 16110 2202
rect 16162 2150 16174 2202
rect 16226 2150 25982 2202
rect 26034 2150 26046 2202
rect 26098 2150 26110 2202
rect 26162 2150 26174 2202
rect 26226 2150 28888 2202
rect 1104 2128 28888 2150
rect 24854 1980 24860 2032
rect 24912 2020 24918 2032
rect 26142 2020 26148 2032
rect 24912 1992 26148 2020
rect 24912 1980 24918 1992
rect 26142 1980 26148 1992
rect 26200 1980 26206 2032
<< via1 >>
rect 3516 22788 3568 22840
rect 10600 22788 10652 22840
rect 3424 22516 3476 22568
rect 7472 22516 7524 22568
rect 5982 21734 6034 21786
rect 6046 21734 6098 21786
rect 6110 21734 6162 21786
rect 6174 21734 6226 21786
rect 15982 21734 16034 21786
rect 16046 21734 16098 21786
rect 16110 21734 16162 21786
rect 16174 21734 16226 21786
rect 25982 21734 26034 21786
rect 26046 21734 26098 21786
rect 26110 21734 26162 21786
rect 26174 21734 26226 21786
rect 3792 21632 3844 21684
rect 4804 21632 4856 21684
rect 10982 21190 11034 21242
rect 11046 21190 11098 21242
rect 11110 21190 11162 21242
rect 11174 21190 11226 21242
rect 20982 21190 21034 21242
rect 21046 21190 21098 21242
rect 21110 21190 21162 21242
rect 21174 21190 21226 21242
rect 14004 21088 14056 21140
rect 19616 21088 19668 21140
rect 29000 21088 29052 21140
rect 12164 20995 12216 21004
rect 12164 20961 12173 20995
rect 12173 20961 12207 20995
rect 12207 20961 12216 20995
rect 12164 20952 12216 20961
rect 17132 20952 17184 21004
rect 17960 20952 18012 21004
rect 19616 20952 19668 21004
rect 24032 20952 24084 21004
rect 26884 20952 26936 21004
rect 4068 20816 4120 20868
rect 5632 20816 5684 20868
rect 18696 20816 18748 20868
rect 21732 20816 21784 20868
rect 25688 20816 25740 20868
rect 5080 20791 5132 20800
rect 5080 20757 5089 20791
rect 5089 20757 5123 20791
rect 5123 20757 5132 20791
rect 5080 20748 5132 20757
rect 9772 20748 9824 20800
rect 12808 20748 12860 20800
rect 18236 20791 18288 20800
rect 18236 20757 18245 20791
rect 18245 20757 18279 20791
rect 18279 20757 18288 20791
rect 18236 20748 18288 20757
rect 21272 20748 21324 20800
rect 25780 20748 25832 20800
rect 5982 20646 6034 20698
rect 6046 20646 6098 20698
rect 6110 20646 6162 20698
rect 6174 20646 6226 20698
rect 15982 20646 16034 20698
rect 16046 20646 16098 20698
rect 16110 20646 16162 20698
rect 16174 20646 16226 20698
rect 25982 20646 26034 20698
rect 26046 20646 26098 20698
rect 26110 20646 26162 20698
rect 26174 20646 26226 20698
rect 940 20544 992 20596
rect 2688 20544 2740 20596
rect 8208 20544 8260 20596
rect 10232 20544 10284 20596
rect 15844 20544 15896 20596
rect 17776 20544 17828 20596
rect 20352 20587 20404 20596
rect 20352 20553 20361 20587
rect 20361 20553 20395 20587
rect 20395 20553 20404 20587
rect 20352 20544 20404 20553
rect 25228 20544 25280 20596
rect 26884 20587 26936 20596
rect 26884 20553 26893 20587
rect 26893 20553 26927 20587
rect 26927 20553 26936 20587
rect 26884 20544 26936 20553
rect 12164 20476 12216 20528
rect 25412 20519 25464 20528
rect 25412 20485 25421 20519
rect 25421 20485 25455 20519
rect 25455 20485 25464 20519
rect 25412 20476 25464 20485
rect 5080 20408 5132 20460
rect 2044 20340 2096 20392
rect 4896 20383 4948 20392
rect 4896 20349 4905 20383
rect 4905 20349 4939 20383
rect 4939 20349 4948 20383
rect 13636 20408 13688 20460
rect 18696 20451 18748 20460
rect 18696 20417 18705 20451
rect 18705 20417 18739 20451
rect 18739 20417 18748 20451
rect 18696 20408 18748 20417
rect 4896 20340 4948 20349
rect 2320 20204 2372 20256
rect 4160 20204 4212 20256
rect 10784 20272 10836 20324
rect 12624 20340 12676 20392
rect 12808 20383 12860 20392
rect 12808 20349 12817 20383
rect 12817 20349 12851 20383
rect 12851 20349 12860 20383
rect 12808 20340 12860 20349
rect 13820 20340 13872 20392
rect 16672 20383 16724 20392
rect 16672 20349 16681 20383
rect 16681 20349 16715 20383
rect 16715 20349 16724 20383
rect 16672 20340 16724 20349
rect 17776 20383 17828 20392
rect 17776 20349 17785 20383
rect 17785 20349 17819 20383
rect 17819 20349 17828 20383
rect 17776 20340 17828 20349
rect 18328 20272 18380 20324
rect 4988 20247 5040 20256
rect 4988 20213 4997 20247
rect 4997 20213 5031 20247
rect 5031 20213 5040 20247
rect 4988 20204 5040 20213
rect 7380 20247 7432 20256
rect 7380 20213 7389 20247
rect 7389 20213 7423 20247
rect 7423 20213 7432 20247
rect 7380 20204 7432 20213
rect 9680 20247 9732 20256
rect 9680 20213 9689 20247
rect 9689 20213 9723 20247
rect 9723 20213 9732 20247
rect 9680 20204 9732 20213
rect 12624 20204 12676 20256
rect 17132 20204 17184 20256
rect 17500 20247 17552 20256
rect 17500 20213 17509 20247
rect 17509 20213 17543 20247
rect 17543 20213 17552 20247
rect 17500 20204 17552 20213
rect 18144 20247 18196 20256
rect 18144 20213 18153 20247
rect 18153 20213 18187 20247
rect 18187 20213 18196 20247
rect 18144 20204 18196 20213
rect 18420 20204 18472 20256
rect 19616 20247 19668 20256
rect 19616 20213 19625 20247
rect 19625 20213 19659 20247
rect 19659 20213 19668 20247
rect 19616 20204 19668 20213
rect 20536 20204 20588 20256
rect 21824 20204 21876 20256
rect 24768 20247 24820 20256
rect 24768 20213 24777 20247
rect 24777 20213 24811 20247
rect 24811 20213 24820 20247
rect 24768 20204 24820 20213
rect 25780 20247 25832 20256
rect 25780 20213 25789 20247
rect 25789 20213 25823 20247
rect 25823 20213 25832 20247
rect 25780 20204 25832 20213
rect 26700 20204 26752 20256
rect 10982 20102 11034 20154
rect 11046 20102 11098 20154
rect 11110 20102 11162 20154
rect 11174 20102 11226 20154
rect 20982 20102 21034 20154
rect 21046 20102 21098 20154
rect 21110 20102 21162 20154
rect 21174 20102 21226 20154
rect 4436 20043 4488 20052
rect 4436 20009 4445 20043
rect 4445 20009 4479 20043
rect 4479 20009 4488 20043
rect 4436 20000 4488 20009
rect 5080 20000 5132 20052
rect 5632 20043 5684 20052
rect 5632 20009 5641 20043
rect 5641 20009 5675 20043
rect 5675 20009 5684 20043
rect 5632 20000 5684 20009
rect 11796 20000 11848 20052
rect 16672 20043 16724 20052
rect 16672 20009 16681 20043
rect 16681 20009 16715 20043
rect 16715 20009 16724 20043
rect 16672 20000 16724 20009
rect 17592 20043 17644 20052
rect 17592 20009 17601 20043
rect 17601 20009 17635 20043
rect 17635 20009 17644 20043
rect 17592 20000 17644 20009
rect 17500 19932 17552 19984
rect 18696 19932 18748 19984
rect 4068 19864 4120 19916
rect 12164 19864 12216 19916
rect 19616 19864 19668 19916
rect 27252 19864 27304 19916
rect 5724 19839 5776 19848
rect 5724 19805 5733 19839
rect 5733 19805 5767 19839
rect 5767 19805 5776 19839
rect 5724 19796 5776 19805
rect 11428 19839 11480 19848
rect 11428 19805 11437 19839
rect 11437 19805 11471 19839
rect 11471 19805 11480 19839
rect 11428 19796 11480 19805
rect 17684 19839 17736 19848
rect 17684 19805 17693 19839
rect 17693 19805 17727 19839
rect 17727 19805 17736 19839
rect 17684 19796 17736 19805
rect 17776 19839 17828 19848
rect 17776 19805 17785 19839
rect 17785 19805 17819 19839
rect 17819 19805 17828 19839
rect 19248 19839 19300 19848
rect 17776 19796 17828 19805
rect 19248 19805 19257 19839
rect 19257 19805 19291 19839
rect 19291 19805 19300 19839
rect 19248 19796 19300 19805
rect 26976 19839 27028 19848
rect 10968 19728 11020 19780
rect 19156 19728 19208 19780
rect 26976 19805 26985 19839
rect 26985 19805 27019 19839
rect 27019 19805 27028 19839
rect 26976 19796 27028 19805
rect 27436 19796 27488 19848
rect 3884 19660 3936 19712
rect 5356 19660 5408 19712
rect 5540 19660 5592 19712
rect 10876 19703 10928 19712
rect 10876 19669 10885 19703
rect 10885 19669 10919 19703
rect 10919 19669 10928 19703
rect 10876 19660 10928 19669
rect 12992 19703 13044 19712
rect 12992 19669 13001 19703
rect 13001 19669 13035 19703
rect 13035 19669 13044 19703
rect 12992 19660 13044 19669
rect 15108 19703 15160 19712
rect 15108 19669 15117 19703
rect 15117 19669 15151 19703
rect 15151 19669 15160 19703
rect 15108 19660 15160 19669
rect 15568 19660 15620 19712
rect 18328 19660 18380 19712
rect 19616 19660 19668 19712
rect 25412 19703 25464 19712
rect 25412 19669 25421 19703
rect 25421 19669 25455 19703
rect 25455 19669 25464 19703
rect 25412 19660 25464 19669
rect 26516 19703 26568 19712
rect 26516 19669 26525 19703
rect 26525 19669 26559 19703
rect 26559 19669 26568 19703
rect 26516 19660 26568 19669
rect 5982 19558 6034 19610
rect 6046 19558 6098 19610
rect 6110 19558 6162 19610
rect 6174 19558 6226 19610
rect 15982 19558 16034 19610
rect 16046 19558 16098 19610
rect 16110 19558 16162 19610
rect 16174 19558 16226 19610
rect 25982 19558 26034 19610
rect 26046 19558 26098 19610
rect 26110 19558 26162 19610
rect 26174 19558 26226 19610
rect 5080 19456 5132 19508
rect 5632 19456 5684 19508
rect 6736 19456 6788 19508
rect 10784 19499 10836 19508
rect 10784 19465 10793 19499
rect 10793 19465 10827 19499
rect 10827 19465 10836 19499
rect 10784 19456 10836 19465
rect 13636 19456 13688 19508
rect 13912 19499 13964 19508
rect 13912 19465 13921 19499
rect 13921 19465 13955 19499
rect 13955 19465 13964 19499
rect 13912 19456 13964 19465
rect 17592 19456 17644 19508
rect 18696 19456 18748 19508
rect 3700 19320 3752 19372
rect 4988 19320 5040 19372
rect 5356 19320 5408 19372
rect 10876 19320 10928 19372
rect 11336 19363 11388 19372
rect 5448 19295 5500 19304
rect 5448 19261 5457 19295
rect 5457 19261 5491 19295
rect 5491 19261 5500 19295
rect 5448 19252 5500 19261
rect 8300 19252 8352 19304
rect 10140 19252 10192 19304
rect 10968 19252 11020 19304
rect 11336 19329 11345 19363
rect 11345 19329 11379 19363
rect 11379 19329 11388 19363
rect 11336 19320 11388 19329
rect 15568 19363 15620 19372
rect 15568 19329 15577 19363
rect 15577 19329 15611 19363
rect 15611 19329 15620 19363
rect 15568 19320 15620 19329
rect 11888 19252 11940 19304
rect 12532 19295 12584 19304
rect 12532 19261 12548 19295
rect 12548 19261 12582 19295
rect 12582 19261 12584 19295
rect 14832 19295 14884 19304
rect 12532 19252 12584 19261
rect 14832 19261 14841 19295
rect 14841 19261 14875 19295
rect 14875 19261 14884 19295
rect 14832 19252 14884 19261
rect 4068 19184 4120 19236
rect 5724 19184 5776 19236
rect 12256 19184 12308 19236
rect 12716 19184 12768 19236
rect 14924 19184 14976 19236
rect 3884 19159 3936 19168
rect 3884 19125 3893 19159
rect 3893 19125 3927 19159
rect 3927 19125 3936 19159
rect 3884 19116 3936 19125
rect 4436 19159 4488 19168
rect 4436 19125 4445 19159
rect 4445 19125 4479 19159
rect 4479 19125 4488 19159
rect 4436 19116 4488 19125
rect 4620 19116 4672 19168
rect 6828 19159 6880 19168
rect 6828 19125 6837 19159
rect 6837 19125 6871 19159
rect 6871 19125 6880 19159
rect 6828 19116 6880 19125
rect 9036 19159 9088 19168
rect 9036 19125 9045 19159
rect 9045 19125 9079 19159
rect 9079 19125 9088 19159
rect 9036 19116 9088 19125
rect 10416 19116 10468 19168
rect 11336 19116 11388 19168
rect 11796 19116 11848 19168
rect 12532 19116 12584 19168
rect 12992 19116 13044 19168
rect 15016 19159 15068 19168
rect 15016 19125 15025 19159
rect 15025 19125 15059 19159
rect 15059 19125 15068 19159
rect 15016 19116 15068 19125
rect 18604 19252 18656 19304
rect 19156 19252 19208 19304
rect 17684 19184 17736 19236
rect 19248 19184 19300 19236
rect 16396 19116 16448 19168
rect 17776 19116 17828 19168
rect 18880 19116 18932 19168
rect 19800 19227 19852 19236
rect 19800 19193 19834 19227
rect 19834 19193 19852 19227
rect 19800 19184 19852 19193
rect 19892 19116 19944 19168
rect 20720 19116 20772 19168
rect 24308 19116 24360 19168
rect 25412 19252 25464 19304
rect 25872 19252 25924 19304
rect 27436 19252 27488 19304
rect 25412 19116 25464 19168
rect 27252 19159 27304 19168
rect 27252 19125 27261 19159
rect 27261 19125 27295 19159
rect 27295 19125 27304 19159
rect 27252 19116 27304 19125
rect 27620 19159 27672 19168
rect 27620 19125 27629 19159
rect 27629 19125 27663 19159
rect 27663 19125 27672 19159
rect 27620 19116 27672 19125
rect 10982 19014 11034 19066
rect 11046 19014 11098 19066
rect 11110 19014 11162 19066
rect 11174 19014 11226 19066
rect 20982 19014 21034 19066
rect 21046 19014 21098 19066
rect 21110 19014 21162 19066
rect 21174 19014 21226 19066
rect 2412 18955 2464 18964
rect 2412 18921 2421 18955
rect 2421 18921 2455 18955
rect 2455 18921 2464 18955
rect 2412 18912 2464 18921
rect 4068 18912 4120 18964
rect 5632 18912 5684 18964
rect 6092 18955 6144 18964
rect 6092 18921 6101 18955
rect 6101 18921 6135 18955
rect 6135 18921 6144 18955
rect 6092 18912 6144 18921
rect 7196 18955 7248 18964
rect 7196 18921 7205 18955
rect 7205 18921 7239 18955
rect 7239 18921 7248 18955
rect 7196 18912 7248 18921
rect 7656 18955 7708 18964
rect 7656 18921 7665 18955
rect 7665 18921 7699 18955
rect 7699 18921 7708 18955
rect 7656 18912 7708 18921
rect 9772 18955 9824 18964
rect 9772 18921 9781 18955
rect 9781 18921 9815 18955
rect 9815 18921 9824 18955
rect 9772 18912 9824 18921
rect 10140 18955 10192 18964
rect 10140 18921 10149 18955
rect 10149 18921 10183 18955
rect 10183 18921 10192 18955
rect 10140 18912 10192 18921
rect 11336 18912 11388 18964
rect 12716 18955 12768 18964
rect 12716 18921 12725 18955
rect 12725 18921 12759 18955
rect 12759 18921 12768 18955
rect 12716 18912 12768 18921
rect 13912 18912 13964 18964
rect 18236 18912 18288 18964
rect 18696 18912 18748 18964
rect 4896 18844 4948 18896
rect 5540 18844 5592 18896
rect 11428 18844 11480 18896
rect 19248 18912 19300 18964
rect 20536 18912 20588 18964
rect 23388 18912 23440 18964
rect 24860 18955 24912 18964
rect 24860 18921 24869 18955
rect 24869 18921 24903 18955
rect 24903 18921 24912 18955
rect 24860 18912 24912 18921
rect 26516 18912 26568 18964
rect 2228 18819 2280 18828
rect 2228 18785 2237 18819
rect 2237 18785 2271 18819
rect 2271 18785 2280 18819
rect 2228 18776 2280 18785
rect 7564 18819 7616 18828
rect 7564 18785 7573 18819
rect 7573 18785 7607 18819
rect 7607 18785 7616 18819
rect 7564 18776 7616 18785
rect 10232 18819 10284 18828
rect 10232 18785 10241 18819
rect 10241 18785 10275 18819
rect 10275 18785 10284 18819
rect 10232 18776 10284 18785
rect 12532 18776 12584 18828
rect 16764 18819 16816 18828
rect 16764 18785 16798 18819
rect 16798 18785 16816 18819
rect 16764 18776 16816 18785
rect 19064 18776 19116 18828
rect 4712 18751 4764 18760
rect 4712 18717 4721 18751
rect 4721 18717 4755 18751
rect 4755 18717 4764 18751
rect 4712 18708 4764 18717
rect 6920 18708 6972 18760
rect 7840 18708 7892 18760
rect 10324 18751 10376 18760
rect 10324 18717 10333 18751
rect 10333 18717 10367 18751
rect 10367 18717 10376 18751
rect 10324 18708 10376 18717
rect 16488 18751 16540 18760
rect 16488 18717 16497 18751
rect 16497 18717 16531 18751
rect 16531 18717 16540 18751
rect 16488 18708 16540 18717
rect 19432 18751 19484 18760
rect 19432 18717 19441 18751
rect 19441 18717 19475 18751
rect 19475 18717 19484 18751
rect 19432 18708 19484 18717
rect 19800 18844 19852 18896
rect 20168 18844 20220 18896
rect 22468 18819 22520 18828
rect 20720 18708 20772 18760
rect 21456 18751 21508 18760
rect 21456 18717 21465 18751
rect 21465 18717 21499 18751
rect 21499 18717 21508 18751
rect 22468 18785 22477 18819
rect 22477 18785 22511 18819
rect 22511 18785 22520 18819
rect 22468 18776 22520 18785
rect 21456 18708 21508 18717
rect 22652 18708 22704 18760
rect 25504 18776 25556 18828
rect 26516 18776 26568 18828
rect 25412 18751 25464 18760
rect 25412 18717 25421 18751
rect 25421 18717 25455 18751
rect 25455 18717 25464 18751
rect 25412 18708 25464 18717
rect 25872 18708 25924 18760
rect 1860 18615 1912 18624
rect 1860 18581 1869 18615
rect 1869 18581 1903 18615
rect 1903 18581 1912 18615
rect 1860 18572 1912 18581
rect 3884 18572 3936 18624
rect 7104 18572 7156 18624
rect 8576 18615 8628 18624
rect 8576 18581 8585 18615
rect 8585 18581 8619 18615
rect 8619 18581 8628 18615
rect 8576 18572 8628 18581
rect 9036 18572 9088 18624
rect 10784 18615 10836 18624
rect 10784 18581 10793 18615
rect 10793 18581 10827 18615
rect 10827 18581 10836 18615
rect 10784 18572 10836 18581
rect 14924 18572 14976 18624
rect 17868 18615 17920 18624
rect 17868 18581 17877 18615
rect 17877 18581 17911 18615
rect 17911 18581 17920 18615
rect 17868 18572 17920 18581
rect 19984 18615 20036 18624
rect 19984 18581 19993 18615
rect 19993 18581 20027 18615
rect 20027 18581 20036 18615
rect 19984 18572 20036 18581
rect 22100 18572 22152 18624
rect 27344 18572 27396 18624
rect 5982 18470 6034 18522
rect 6046 18470 6098 18522
rect 6110 18470 6162 18522
rect 6174 18470 6226 18522
rect 15982 18470 16034 18522
rect 16046 18470 16098 18522
rect 16110 18470 16162 18522
rect 16174 18470 16226 18522
rect 25982 18470 26034 18522
rect 26046 18470 26098 18522
rect 26110 18470 26162 18522
rect 26174 18470 26226 18522
rect 3976 18368 4028 18420
rect 5448 18368 5500 18420
rect 7840 18411 7892 18420
rect 7840 18377 7849 18411
rect 7849 18377 7883 18411
rect 7883 18377 7892 18411
rect 7840 18368 7892 18377
rect 10232 18368 10284 18420
rect 11888 18368 11940 18420
rect 17684 18368 17736 18420
rect 19616 18411 19668 18420
rect 19616 18377 19625 18411
rect 19625 18377 19659 18411
rect 19659 18377 19668 18411
rect 19616 18368 19668 18377
rect 25504 18368 25556 18420
rect 7564 18300 7616 18352
rect 10324 18300 10376 18352
rect 10600 18343 10652 18352
rect 10600 18309 10609 18343
rect 10609 18309 10643 18343
rect 10643 18309 10652 18343
rect 10600 18300 10652 18309
rect 16764 18300 16816 18352
rect 19984 18300 20036 18352
rect 25872 18343 25924 18352
rect 3884 18275 3936 18284
rect 3884 18241 3893 18275
rect 3893 18241 3927 18275
rect 3927 18241 3936 18275
rect 3884 18232 3936 18241
rect 4160 18232 4212 18284
rect 4344 18232 4396 18284
rect 7288 18232 7340 18284
rect 9036 18275 9088 18284
rect 9036 18241 9045 18275
rect 9045 18241 9079 18275
rect 9079 18241 9088 18275
rect 9036 18232 9088 18241
rect 11428 18275 11480 18284
rect 11428 18241 11437 18275
rect 11437 18241 11471 18275
rect 11471 18241 11480 18275
rect 11428 18232 11480 18241
rect 12532 18232 12584 18284
rect 13084 18275 13136 18284
rect 3700 18207 3752 18216
rect 3700 18173 3709 18207
rect 3709 18173 3743 18207
rect 3743 18173 3752 18207
rect 3700 18164 3752 18173
rect 9588 18164 9640 18216
rect 10600 18164 10652 18216
rect 11152 18207 11204 18216
rect 11152 18173 11161 18207
rect 11161 18173 11195 18207
rect 11195 18173 11204 18207
rect 11152 18164 11204 18173
rect 5264 18139 5316 18148
rect 1676 18028 1728 18080
rect 2504 18028 2556 18080
rect 2688 18028 2740 18080
rect 3608 18028 3660 18080
rect 4252 18028 4304 18080
rect 5264 18105 5273 18139
rect 5273 18105 5307 18139
rect 5307 18105 5316 18139
rect 5264 18096 5316 18105
rect 7104 18096 7156 18148
rect 8944 18139 8996 18148
rect 4988 18028 5040 18080
rect 5448 18028 5500 18080
rect 7196 18071 7248 18080
rect 7196 18037 7205 18071
rect 7205 18037 7239 18071
rect 7239 18037 7248 18071
rect 7196 18028 7248 18037
rect 7932 18028 7984 18080
rect 8944 18105 8953 18139
rect 8953 18105 8987 18139
rect 8987 18105 8996 18139
rect 8944 18096 8996 18105
rect 10692 18096 10744 18148
rect 13084 18241 13093 18275
rect 13093 18241 13127 18275
rect 13127 18241 13136 18275
rect 13084 18232 13136 18241
rect 18144 18232 18196 18284
rect 18604 18275 18656 18284
rect 18604 18241 18613 18275
rect 18613 18241 18647 18275
rect 18647 18241 18656 18275
rect 25872 18309 25881 18343
rect 25881 18309 25915 18343
rect 25915 18309 25924 18343
rect 25872 18300 25924 18309
rect 18604 18232 18656 18241
rect 20168 18275 20220 18284
rect 20168 18241 20177 18275
rect 20177 18241 20211 18275
rect 20211 18241 20220 18275
rect 20168 18232 20220 18241
rect 21640 18232 21692 18284
rect 22100 18275 22152 18284
rect 22100 18241 22109 18275
rect 22109 18241 22143 18275
rect 22143 18241 22152 18275
rect 22100 18232 22152 18241
rect 13912 18096 13964 18148
rect 8484 18071 8536 18080
rect 8484 18037 8493 18071
rect 8493 18037 8527 18071
rect 8527 18037 8536 18071
rect 8484 18028 8536 18037
rect 8576 18028 8628 18080
rect 10784 18028 10836 18080
rect 12992 18028 13044 18080
rect 18236 18164 18288 18216
rect 18880 18164 18932 18216
rect 20260 18164 20312 18216
rect 22008 18164 22060 18216
rect 19064 18139 19116 18148
rect 19064 18105 19073 18139
rect 19073 18105 19107 18139
rect 19107 18105 19116 18139
rect 19064 18096 19116 18105
rect 20352 18096 20404 18148
rect 21272 18096 21324 18148
rect 22100 18096 22152 18148
rect 22468 18096 22520 18148
rect 24676 18096 24728 18148
rect 15292 18028 15344 18080
rect 15568 18071 15620 18080
rect 15568 18037 15577 18071
rect 15577 18037 15611 18071
rect 15611 18037 15620 18071
rect 15568 18028 15620 18037
rect 15844 18028 15896 18080
rect 16488 18071 16540 18080
rect 16488 18037 16497 18071
rect 16497 18037 16531 18071
rect 16531 18037 16540 18071
rect 16488 18028 16540 18037
rect 19432 18071 19484 18080
rect 19432 18037 19441 18071
rect 19441 18037 19475 18071
rect 19475 18037 19484 18071
rect 19432 18028 19484 18037
rect 20720 18028 20772 18080
rect 21548 18071 21600 18080
rect 21548 18037 21557 18071
rect 21557 18037 21591 18071
rect 21591 18037 21600 18071
rect 21548 18028 21600 18037
rect 21916 18028 21968 18080
rect 22652 18071 22704 18080
rect 22652 18037 22661 18071
rect 22661 18037 22695 18071
rect 22695 18037 22704 18071
rect 22652 18028 22704 18037
rect 24308 18071 24360 18080
rect 24308 18037 24317 18071
rect 24317 18037 24351 18071
rect 24351 18037 24360 18071
rect 24308 18028 24360 18037
rect 26240 18028 26292 18080
rect 27344 18071 27396 18080
rect 27344 18037 27353 18071
rect 27353 18037 27387 18071
rect 27387 18037 27396 18071
rect 27344 18028 27396 18037
rect 27528 18028 27580 18080
rect 10982 17926 11034 17978
rect 11046 17926 11098 17978
rect 11110 17926 11162 17978
rect 11174 17926 11226 17978
rect 20982 17926 21034 17978
rect 21046 17926 21098 17978
rect 21110 17926 21162 17978
rect 21174 17926 21226 17978
rect 2228 17824 2280 17876
rect 3700 17824 3752 17876
rect 4344 17867 4396 17876
rect 4344 17833 4353 17867
rect 4353 17833 4387 17867
rect 4387 17833 4396 17867
rect 4344 17824 4396 17833
rect 4712 17867 4764 17876
rect 4712 17833 4721 17867
rect 4721 17833 4755 17867
rect 4755 17833 4764 17867
rect 4712 17824 4764 17833
rect 5540 17824 5592 17876
rect 6828 17824 6880 17876
rect 7564 17824 7616 17876
rect 8208 17824 8260 17876
rect 8484 17824 8536 17876
rect 9404 17867 9456 17876
rect 9404 17833 9413 17867
rect 9413 17833 9447 17867
rect 9447 17833 9456 17867
rect 9404 17824 9456 17833
rect 11428 17824 11480 17876
rect 12164 17867 12216 17876
rect 4160 17756 4212 17808
rect 5356 17756 5408 17808
rect 7288 17756 7340 17808
rect 8392 17799 8444 17808
rect 8392 17765 8401 17799
rect 8401 17765 8435 17799
rect 8435 17765 8444 17799
rect 8392 17756 8444 17765
rect 10784 17756 10836 17808
rect 12164 17833 12173 17867
rect 12173 17833 12207 17867
rect 12207 17833 12216 17867
rect 12164 17824 12216 17833
rect 13728 17824 13780 17876
rect 13084 17756 13136 17808
rect 13820 17756 13872 17808
rect 20076 17824 20128 17876
rect 20260 17867 20312 17876
rect 20260 17833 20269 17867
rect 20269 17833 20303 17867
rect 20303 17833 20312 17867
rect 20260 17824 20312 17833
rect 22100 17824 22152 17876
rect 25412 17824 25464 17876
rect 26332 17824 26384 17876
rect 26516 17867 26568 17876
rect 26516 17833 26525 17867
rect 26525 17833 26559 17867
rect 26559 17833 26568 17867
rect 26516 17824 26568 17833
rect 19800 17756 19852 17808
rect 21456 17756 21508 17808
rect 22468 17756 22520 17808
rect 25596 17756 25648 17808
rect 2136 17731 2188 17740
rect 2136 17697 2145 17731
rect 2145 17697 2179 17731
rect 2179 17697 2188 17731
rect 2136 17688 2188 17697
rect 2688 17688 2740 17740
rect 4712 17688 4764 17740
rect 7656 17688 7708 17740
rect 8208 17688 8260 17740
rect 9588 17688 9640 17740
rect 9772 17688 9824 17740
rect 14004 17731 14056 17740
rect 14004 17697 14013 17731
rect 14013 17697 14047 17731
rect 14047 17697 14056 17731
rect 14004 17688 14056 17697
rect 16396 17688 16448 17740
rect 21272 17731 21324 17740
rect 21272 17697 21281 17731
rect 21281 17697 21315 17731
rect 21315 17697 21324 17731
rect 21272 17688 21324 17697
rect 25688 17688 25740 17740
rect 1860 17620 1912 17672
rect 3148 17620 3200 17672
rect 7472 17620 7524 17672
rect 8668 17663 8720 17672
rect 8668 17629 8677 17663
rect 8677 17629 8711 17663
rect 8711 17629 8720 17663
rect 8668 17620 8720 17629
rect 11520 17620 11572 17672
rect 12716 17663 12768 17672
rect 12716 17629 12725 17663
rect 12725 17629 12759 17663
rect 12759 17629 12768 17663
rect 12716 17620 12768 17629
rect 14188 17663 14240 17672
rect 14188 17629 14197 17663
rect 14197 17629 14231 17663
rect 14231 17629 14240 17663
rect 14188 17620 14240 17629
rect 15292 17620 15344 17672
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 17868 17620 17920 17672
rect 21364 17663 21416 17672
rect 21364 17629 21373 17663
rect 21373 17629 21407 17663
rect 21407 17629 21416 17663
rect 21364 17620 21416 17629
rect 21456 17663 21508 17672
rect 21456 17629 21465 17663
rect 21465 17629 21499 17663
rect 21499 17629 21508 17663
rect 21456 17620 21508 17629
rect 22376 17620 22428 17672
rect 24860 17620 24912 17672
rect 26148 17620 26200 17672
rect 27436 17620 27488 17672
rect 11244 17552 11296 17604
rect 19340 17552 19392 17604
rect 22100 17552 22152 17604
rect 2780 17527 2832 17536
rect 2780 17493 2789 17527
rect 2789 17493 2823 17527
rect 2823 17493 2832 17527
rect 2780 17484 2832 17493
rect 11520 17484 11572 17536
rect 12992 17527 13044 17536
rect 12992 17493 13001 17527
rect 13001 17493 13035 17527
rect 13035 17493 13044 17527
rect 12992 17484 13044 17493
rect 21916 17527 21968 17536
rect 21916 17493 21925 17527
rect 21925 17493 21959 17527
rect 21959 17493 21968 17527
rect 21916 17484 21968 17493
rect 24124 17484 24176 17536
rect 24676 17484 24728 17536
rect 25320 17527 25372 17536
rect 25320 17493 25329 17527
rect 25329 17493 25363 17527
rect 25363 17493 25372 17527
rect 25320 17484 25372 17493
rect 27620 17527 27672 17536
rect 27620 17493 27629 17527
rect 27629 17493 27663 17527
rect 27663 17493 27672 17527
rect 27620 17484 27672 17493
rect 5982 17382 6034 17434
rect 6046 17382 6098 17434
rect 6110 17382 6162 17434
rect 6174 17382 6226 17434
rect 15982 17382 16034 17434
rect 16046 17382 16098 17434
rect 16110 17382 16162 17434
rect 16174 17382 16226 17434
rect 25982 17382 26034 17434
rect 26046 17382 26098 17434
rect 26110 17382 26162 17434
rect 26174 17382 26226 17434
rect 3148 17323 3200 17332
rect 3148 17289 3157 17323
rect 3157 17289 3191 17323
rect 3191 17289 3200 17323
rect 3148 17280 3200 17289
rect 5356 17280 5408 17332
rect 6644 17323 6696 17332
rect 6644 17289 6653 17323
rect 6653 17289 6687 17323
rect 6687 17289 6696 17323
rect 6644 17280 6696 17289
rect 8668 17280 8720 17332
rect 9772 17280 9824 17332
rect 10784 17323 10836 17332
rect 10784 17289 10793 17323
rect 10793 17289 10827 17323
rect 10827 17289 10836 17323
rect 10784 17280 10836 17289
rect 11796 17323 11848 17332
rect 11796 17289 11805 17323
rect 11805 17289 11839 17323
rect 11839 17289 11848 17323
rect 11796 17280 11848 17289
rect 12992 17280 13044 17332
rect 14188 17280 14240 17332
rect 16396 17323 16448 17332
rect 16396 17289 16405 17323
rect 16405 17289 16439 17323
rect 16439 17289 16448 17323
rect 16396 17280 16448 17289
rect 18328 17323 18380 17332
rect 18328 17289 18337 17323
rect 18337 17289 18371 17323
rect 18371 17289 18380 17323
rect 18328 17280 18380 17289
rect 19800 17323 19852 17332
rect 19800 17289 19809 17323
rect 19809 17289 19843 17323
rect 19843 17289 19852 17323
rect 19800 17280 19852 17289
rect 21456 17280 21508 17332
rect 22468 17280 22520 17332
rect 25688 17323 25740 17332
rect 25688 17289 25697 17323
rect 25697 17289 25731 17323
rect 25731 17289 25740 17323
rect 25688 17280 25740 17289
rect 9588 17212 9640 17264
rect 11336 17187 11388 17196
rect 11336 17153 11345 17187
rect 11345 17153 11379 17187
rect 11379 17153 11388 17187
rect 11336 17144 11388 17153
rect 12716 17144 12768 17196
rect 1492 17076 1544 17128
rect 2412 17076 2464 17128
rect 2780 17076 2832 17128
rect 4344 17076 4396 17128
rect 8208 17076 8260 17128
rect 11152 17119 11204 17128
rect 11152 17085 11161 17119
rect 11161 17085 11195 17119
rect 11195 17085 11204 17119
rect 11152 17076 11204 17085
rect 11796 17076 11848 17128
rect 4712 17008 4764 17060
rect 7472 17008 7524 17060
rect 1860 16940 1912 16992
rect 2780 16940 2832 16992
rect 3700 16983 3752 16992
rect 3700 16949 3709 16983
rect 3709 16949 3743 16983
rect 3743 16949 3752 16983
rect 3700 16940 3752 16949
rect 9496 17008 9548 17060
rect 11244 17051 11296 17060
rect 11244 17017 11253 17051
rect 11253 17017 11287 17051
rect 11287 17017 11296 17051
rect 11244 17008 11296 17017
rect 12992 17008 13044 17060
rect 8208 16983 8260 16992
rect 8208 16949 8217 16983
rect 8217 16949 8251 16983
rect 8251 16949 8260 16983
rect 8208 16940 8260 16949
rect 12256 16983 12308 16992
rect 12256 16949 12265 16983
rect 12265 16949 12299 16983
rect 12299 16949 12308 16983
rect 12256 16940 12308 16949
rect 14924 17144 14976 17196
rect 19064 17144 19116 17196
rect 24676 17212 24728 17264
rect 27436 17280 27488 17332
rect 25596 17144 25648 17196
rect 13820 16940 13872 16992
rect 18604 17076 18656 17128
rect 20812 17076 20864 17128
rect 22376 17076 22428 17128
rect 24308 17076 24360 17128
rect 26240 17076 26292 17128
rect 15476 17008 15528 17060
rect 21916 17008 21968 17060
rect 24124 17008 24176 17060
rect 26332 17008 26384 17060
rect 15200 16940 15252 16992
rect 17500 16983 17552 16992
rect 17500 16949 17509 16983
rect 17509 16949 17543 16983
rect 17543 16949 17552 16983
rect 18696 16983 18748 16992
rect 17500 16940 17552 16949
rect 18696 16949 18705 16983
rect 18705 16949 18739 16983
rect 18739 16949 18748 16983
rect 18696 16940 18748 16949
rect 19892 16940 19944 16992
rect 20812 16940 20864 16992
rect 22468 16983 22520 16992
rect 22468 16949 22477 16983
rect 22477 16949 22511 16983
rect 22511 16949 22520 16983
rect 22468 16940 22520 16949
rect 27528 16983 27580 16992
rect 27528 16949 27537 16983
rect 27537 16949 27571 16983
rect 27571 16949 27580 16983
rect 27528 16940 27580 16949
rect 10982 16838 11034 16890
rect 11046 16838 11098 16890
rect 11110 16838 11162 16890
rect 11174 16838 11226 16890
rect 20982 16838 21034 16890
rect 21046 16838 21098 16890
rect 21110 16838 21162 16890
rect 21174 16838 21226 16890
rect 2136 16736 2188 16788
rect 2228 16736 2280 16788
rect 3700 16736 3752 16788
rect 4712 16736 4764 16788
rect 3148 16668 3200 16720
rect 3424 16668 3476 16720
rect 2044 16643 2096 16652
rect 2044 16609 2053 16643
rect 2053 16609 2087 16643
rect 2087 16609 2096 16643
rect 2044 16600 2096 16609
rect 8484 16736 8536 16788
rect 11336 16736 11388 16788
rect 13084 16736 13136 16788
rect 13820 16736 13872 16788
rect 17224 16736 17276 16788
rect 18420 16779 18472 16788
rect 18420 16745 18429 16779
rect 18429 16745 18463 16779
rect 18463 16745 18472 16779
rect 18420 16736 18472 16745
rect 21364 16736 21416 16788
rect 22468 16736 22520 16788
rect 24676 16779 24728 16788
rect 24676 16745 24685 16779
rect 24685 16745 24719 16779
rect 24719 16745 24728 16779
rect 24676 16736 24728 16745
rect 24860 16779 24912 16788
rect 24860 16745 24869 16779
rect 24869 16745 24903 16779
rect 24903 16745 24912 16779
rect 24860 16736 24912 16745
rect 25320 16779 25372 16788
rect 25320 16745 25329 16779
rect 25329 16745 25363 16779
rect 25363 16745 25372 16779
rect 25320 16736 25372 16745
rect 5632 16711 5684 16720
rect 5632 16677 5666 16711
rect 5666 16677 5684 16711
rect 5632 16668 5684 16677
rect 8300 16668 8352 16720
rect 10784 16668 10836 16720
rect 16580 16668 16632 16720
rect 21180 16668 21232 16720
rect 25228 16711 25280 16720
rect 25228 16677 25237 16711
rect 25237 16677 25271 16711
rect 25271 16677 25280 16711
rect 25228 16668 25280 16677
rect 5356 16643 5408 16652
rect 5356 16609 5365 16643
rect 5365 16609 5399 16643
rect 5399 16609 5408 16643
rect 5356 16600 5408 16609
rect 7564 16643 7616 16652
rect 7564 16609 7573 16643
rect 7573 16609 7607 16643
rect 7607 16609 7616 16643
rect 7564 16600 7616 16609
rect 8024 16600 8076 16652
rect 8760 16600 8812 16652
rect 9588 16600 9640 16652
rect 10416 16600 10468 16652
rect 11520 16600 11572 16652
rect 13820 16600 13872 16652
rect 15476 16600 15528 16652
rect 15660 16643 15712 16652
rect 15660 16609 15669 16643
rect 15669 16609 15703 16643
rect 15703 16609 15712 16643
rect 15660 16600 15712 16609
rect 16304 16600 16356 16652
rect 16672 16643 16724 16652
rect 16672 16609 16681 16643
rect 16681 16609 16715 16643
rect 16715 16609 16724 16643
rect 16672 16600 16724 16609
rect 18788 16643 18840 16652
rect 18788 16609 18797 16643
rect 18797 16609 18831 16643
rect 18831 16609 18840 16643
rect 18788 16600 18840 16609
rect 21640 16600 21692 16652
rect 23572 16643 23624 16652
rect 23572 16609 23581 16643
rect 23581 16609 23615 16643
rect 23615 16609 23624 16643
rect 23572 16600 23624 16609
rect 26884 16643 26936 16652
rect 26884 16609 26893 16643
rect 26893 16609 26927 16643
rect 26927 16609 26936 16643
rect 26884 16600 26936 16609
rect 26976 16643 27028 16652
rect 26976 16609 26985 16643
rect 26985 16609 27019 16643
rect 27019 16609 27028 16643
rect 26976 16600 27028 16609
rect 2136 16575 2188 16584
rect 2136 16541 2145 16575
rect 2145 16541 2179 16575
rect 2179 16541 2188 16575
rect 2136 16532 2188 16541
rect 2872 16532 2924 16584
rect 2412 16464 2464 16516
rect 9036 16532 9088 16584
rect 10232 16575 10284 16584
rect 10232 16541 10241 16575
rect 10241 16541 10275 16575
rect 10275 16541 10284 16575
rect 10232 16532 10284 16541
rect 11428 16575 11480 16584
rect 11428 16541 11437 16575
rect 11437 16541 11471 16575
rect 11471 16541 11480 16575
rect 11428 16532 11480 16541
rect 14464 16532 14516 16584
rect 15108 16532 15160 16584
rect 17408 16575 17460 16584
rect 17408 16541 17417 16575
rect 17417 16541 17451 16575
rect 17451 16541 17460 16575
rect 17408 16532 17460 16541
rect 17592 16532 17644 16584
rect 19064 16575 19116 16584
rect 19064 16541 19073 16575
rect 19073 16541 19107 16575
rect 19107 16541 19116 16575
rect 19064 16532 19116 16541
rect 20812 16532 20864 16584
rect 24676 16532 24728 16584
rect 25872 16532 25924 16584
rect 16856 16507 16908 16516
rect 16856 16473 16865 16507
rect 16865 16473 16899 16507
rect 16899 16473 16908 16507
rect 16856 16464 16908 16473
rect 24124 16507 24176 16516
rect 24124 16473 24133 16507
rect 24133 16473 24167 16507
rect 24167 16473 24176 16507
rect 24124 16464 24176 16473
rect 2688 16439 2740 16448
rect 2688 16405 2697 16439
rect 2697 16405 2731 16439
rect 2731 16405 2740 16439
rect 2688 16396 2740 16405
rect 3700 16439 3752 16448
rect 3700 16405 3709 16439
rect 3709 16405 3743 16439
rect 3743 16405 3752 16439
rect 3700 16396 3752 16405
rect 4528 16439 4580 16448
rect 4528 16405 4537 16439
rect 4537 16405 4571 16439
rect 4571 16405 4580 16439
rect 4528 16396 4580 16405
rect 6368 16396 6420 16448
rect 11060 16396 11112 16448
rect 17868 16396 17920 16448
rect 18144 16439 18196 16448
rect 18144 16405 18153 16439
rect 18153 16405 18187 16439
rect 18187 16405 18196 16439
rect 18144 16396 18196 16405
rect 22560 16396 22612 16448
rect 23480 16439 23532 16448
rect 23480 16405 23489 16439
rect 23489 16405 23523 16439
rect 23523 16405 23532 16439
rect 23480 16396 23532 16405
rect 26332 16396 26384 16448
rect 5982 16294 6034 16346
rect 6046 16294 6098 16346
rect 6110 16294 6162 16346
rect 6174 16294 6226 16346
rect 15982 16294 16034 16346
rect 16046 16294 16098 16346
rect 16110 16294 16162 16346
rect 16174 16294 16226 16346
rect 25982 16294 26034 16346
rect 26046 16294 26098 16346
rect 26110 16294 26162 16346
rect 26174 16294 26226 16346
rect 2872 16235 2924 16244
rect 2872 16201 2881 16235
rect 2881 16201 2915 16235
rect 2915 16201 2924 16235
rect 2872 16192 2924 16201
rect 4344 16192 4396 16244
rect 5356 16235 5408 16244
rect 5356 16201 5365 16235
rect 5365 16201 5399 16235
rect 5399 16201 5408 16235
rect 5356 16192 5408 16201
rect 5632 16192 5684 16244
rect 8208 16192 8260 16244
rect 9496 16192 9548 16244
rect 10784 16235 10836 16244
rect 10784 16201 10793 16235
rect 10793 16201 10827 16235
rect 10827 16201 10836 16235
rect 10784 16192 10836 16201
rect 11796 16235 11848 16244
rect 11796 16201 11805 16235
rect 11805 16201 11839 16235
rect 11839 16201 11848 16235
rect 11796 16192 11848 16201
rect 12440 16235 12492 16244
rect 12440 16201 12449 16235
rect 12449 16201 12483 16235
rect 12483 16201 12492 16235
rect 12440 16192 12492 16201
rect 13084 16192 13136 16244
rect 15476 16192 15528 16244
rect 17408 16192 17460 16244
rect 21272 16192 21324 16244
rect 24584 16235 24636 16244
rect 24584 16201 24593 16235
rect 24593 16201 24627 16235
rect 24627 16201 24636 16235
rect 24584 16192 24636 16201
rect 25228 16192 25280 16244
rect 25688 16192 25740 16244
rect 28080 16235 28132 16244
rect 28080 16201 28089 16235
rect 28089 16201 28123 16235
rect 28123 16201 28132 16235
rect 28080 16192 28132 16201
rect 2688 16056 2740 16108
rect 1492 15988 1544 16040
rect 3424 15988 3476 16040
rect 5448 15988 5500 16040
rect 8116 15988 8168 16040
rect 1584 15920 1636 15972
rect 4252 15920 4304 15972
rect 11060 16056 11112 16108
rect 11336 16099 11388 16108
rect 11336 16065 11345 16099
rect 11345 16065 11379 16099
rect 11379 16065 11388 16099
rect 11336 16056 11388 16065
rect 12348 16056 12400 16108
rect 16304 16124 16356 16176
rect 21640 16124 21692 16176
rect 21916 16124 21968 16176
rect 21548 16056 21600 16108
rect 24676 16124 24728 16176
rect 25964 16167 26016 16176
rect 25964 16133 25973 16167
rect 25973 16133 26007 16167
rect 26007 16133 26016 16167
rect 25964 16124 26016 16133
rect 10600 15988 10652 16040
rect 11612 15988 11664 16040
rect 14464 16031 14516 16040
rect 14464 15997 14498 16031
rect 14498 15997 14516 16031
rect 8392 15920 8444 15972
rect 1768 15895 1820 15904
rect 1768 15861 1777 15895
rect 1777 15861 1811 15895
rect 1811 15861 1820 15895
rect 1768 15852 1820 15861
rect 2504 15852 2556 15904
rect 6092 15895 6144 15904
rect 6092 15861 6101 15895
rect 6101 15861 6135 15895
rect 6135 15861 6144 15895
rect 6092 15852 6144 15861
rect 8760 15852 8812 15904
rect 10416 15852 10468 15904
rect 10784 15852 10836 15904
rect 11796 15920 11848 15972
rect 11612 15852 11664 15904
rect 12348 15920 12400 15972
rect 13084 15920 13136 15972
rect 14464 15988 14516 15997
rect 17868 15988 17920 16040
rect 18144 15988 18196 16040
rect 23480 15988 23532 16040
rect 24768 15988 24820 16040
rect 26148 16031 26200 16040
rect 26148 15997 26157 16031
rect 26157 15997 26191 16031
rect 26191 15997 26200 16031
rect 26148 15988 26200 15997
rect 26424 16031 26476 16040
rect 26424 15997 26458 16031
rect 26458 15997 26476 16031
rect 26424 15988 26476 15997
rect 27528 15988 27580 16040
rect 15292 15920 15344 15972
rect 16488 15920 16540 15972
rect 22192 15920 22244 15972
rect 23204 15920 23256 15972
rect 12900 15895 12952 15904
rect 12900 15861 12909 15895
rect 12909 15861 12943 15895
rect 12943 15861 12952 15895
rect 12900 15852 12952 15861
rect 16580 15895 16632 15904
rect 16580 15861 16589 15895
rect 16589 15861 16623 15895
rect 16623 15861 16632 15895
rect 16580 15852 16632 15861
rect 17592 15852 17644 15904
rect 18512 15852 18564 15904
rect 19984 15895 20036 15904
rect 19984 15861 19993 15895
rect 19993 15861 20027 15895
rect 20027 15861 20036 15895
rect 19984 15852 20036 15861
rect 20812 15852 20864 15904
rect 21916 15852 21968 15904
rect 22560 15852 22612 15904
rect 27344 15852 27396 15904
rect 10982 15750 11034 15802
rect 11046 15750 11098 15802
rect 11110 15750 11162 15802
rect 11174 15750 11226 15802
rect 20982 15750 21034 15802
rect 21046 15750 21098 15802
rect 21110 15750 21162 15802
rect 21174 15750 21226 15802
rect 2780 15648 2832 15700
rect 4528 15691 4580 15700
rect 4528 15657 4537 15691
rect 4537 15657 4571 15691
rect 4571 15657 4580 15691
rect 4528 15648 4580 15657
rect 8116 15648 8168 15700
rect 8300 15648 8352 15700
rect 8576 15691 8628 15700
rect 8576 15657 8585 15691
rect 8585 15657 8619 15691
rect 8619 15657 8628 15691
rect 8576 15648 8628 15657
rect 9680 15691 9732 15700
rect 9680 15657 9689 15691
rect 9689 15657 9723 15691
rect 9723 15657 9732 15691
rect 9680 15648 9732 15657
rect 8392 15580 8444 15632
rect 10232 15648 10284 15700
rect 14464 15691 14516 15700
rect 14464 15657 14473 15691
rect 14473 15657 14507 15691
rect 14507 15657 14516 15691
rect 14464 15648 14516 15657
rect 17224 15691 17276 15700
rect 17224 15657 17233 15691
rect 17233 15657 17267 15691
rect 17267 15657 17276 15691
rect 17224 15648 17276 15657
rect 19064 15648 19116 15700
rect 21364 15648 21416 15700
rect 21640 15648 21692 15700
rect 23204 15691 23256 15700
rect 23204 15657 23213 15691
rect 23213 15657 23247 15691
rect 23247 15657 23256 15691
rect 23204 15648 23256 15657
rect 24768 15691 24820 15700
rect 24768 15657 24777 15691
rect 24777 15657 24811 15691
rect 24811 15657 24820 15691
rect 24768 15648 24820 15657
rect 25872 15691 25924 15700
rect 25872 15657 25881 15691
rect 25881 15657 25915 15691
rect 25915 15657 25924 15691
rect 25872 15648 25924 15657
rect 27528 15691 27580 15700
rect 27528 15657 27537 15691
rect 27537 15657 27571 15691
rect 27571 15657 27580 15691
rect 27528 15648 27580 15657
rect 11336 15580 11388 15632
rect 12164 15580 12216 15632
rect 15568 15623 15620 15632
rect 15568 15589 15602 15623
rect 15602 15589 15620 15623
rect 15568 15580 15620 15589
rect 1492 15555 1544 15564
rect 1492 15521 1501 15555
rect 1501 15521 1535 15555
rect 1535 15521 1544 15555
rect 1492 15512 1544 15521
rect 2596 15512 2648 15564
rect 4436 15555 4488 15564
rect 4436 15521 4445 15555
rect 4445 15521 4479 15555
rect 4479 15521 4488 15555
rect 4436 15512 4488 15521
rect 6368 15512 6420 15564
rect 9680 15512 9732 15564
rect 17408 15512 17460 15564
rect 18512 15555 18564 15564
rect 18512 15521 18535 15555
rect 18535 15521 18564 15555
rect 18512 15512 18564 15521
rect 20628 15512 20680 15564
rect 23572 15555 23624 15564
rect 23572 15521 23581 15555
rect 23581 15521 23615 15555
rect 23615 15521 23624 15555
rect 23572 15512 23624 15521
rect 24676 15555 24728 15564
rect 24676 15521 24685 15555
rect 24685 15521 24719 15555
rect 24719 15521 24728 15555
rect 24676 15512 24728 15521
rect 25596 15512 25648 15564
rect 27436 15512 27488 15564
rect 3700 15444 3752 15496
rect 4620 15487 4672 15496
rect 4620 15453 4629 15487
rect 4629 15453 4663 15487
rect 4663 15453 4672 15487
rect 4620 15444 4672 15453
rect 5448 15444 5500 15496
rect 9772 15444 9824 15496
rect 10324 15487 10376 15496
rect 10324 15453 10333 15487
rect 10333 15453 10367 15487
rect 10367 15453 10376 15487
rect 10324 15444 10376 15453
rect 11428 15444 11480 15496
rect 11796 15487 11848 15496
rect 11796 15453 11805 15487
rect 11805 15453 11839 15487
rect 11839 15453 11848 15487
rect 11796 15444 11848 15453
rect 15292 15487 15344 15496
rect 15292 15453 15301 15487
rect 15301 15453 15335 15487
rect 15335 15453 15344 15487
rect 15292 15444 15344 15453
rect 3884 15351 3936 15360
rect 3884 15317 3893 15351
rect 3893 15317 3927 15351
rect 3927 15317 3936 15351
rect 3884 15308 3936 15317
rect 5632 15351 5684 15360
rect 5632 15317 5641 15351
rect 5641 15317 5675 15351
rect 5675 15317 5684 15351
rect 5632 15308 5684 15317
rect 10784 15351 10836 15360
rect 10784 15317 10793 15351
rect 10793 15317 10827 15351
rect 10827 15317 10836 15351
rect 10784 15308 10836 15317
rect 14096 15308 14148 15360
rect 16488 15308 16540 15360
rect 17868 15308 17920 15360
rect 18236 15308 18288 15360
rect 20536 15308 20588 15360
rect 20720 15351 20772 15360
rect 20720 15317 20729 15351
rect 20729 15317 20763 15351
rect 20763 15317 20772 15351
rect 21916 15444 21968 15496
rect 23664 15487 23716 15496
rect 23664 15453 23673 15487
rect 23673 15453 23707 15487
rect 23707 15453 23716 15487
rect 23664 15444 23716 15453
rect 25228 15487 25280 15496
rect 23480 15376 23532 15428
rect 25228 15453 25237 15487
rect 25237 15453 25271 15487
rect 25271 15453 25280 15487
rect 25228 15444 25280 15453
rect 25320 15376 25372 15428
rect 25872 15444 25924 15496
rect 26148 15487 26200 15496
rect 24308 15351 24360 15360
rect 20720 15308 20772 15317
rect 24308 15317 24317 15351
rect 24317 15317 24351 15351
rect 24351 15317 24360 15351
rect 26148 15453 26157 15487
rect 26157 15453 26191 15487
rect 26191 15453 26200 15487
rect 26148 15444 26200 15453
rect 26608 15444 26660 15496
rect 27528 15444 27580 15496
rect 26516 15351 26568 15360
rect 24308 15308 24360 15317
rect 26516 15317 26525 15351
rect 26525 15317 26559 15351
rect 26559 15317 26568 15351
rect 26516 15308 26568 15317
rect 5982 15206 6034 15258
rect 6046 15206 6098 15258
rect 6110 15206 6162 15258
rect 6174 15206 6226 15258
rect 15982 15206 16034 15258
rect 16046 15206 16098 15258
rect 16110 15206 16162 15258
rect 16174 15206 16226 15258
rect 25982 15206 26034 15258
rect 26046 15206 26098 15258
rect 26110 15206 26162 15258
rect 26174 15206 26226 15258
rect 2044 15104 2096 15156
rect 5448 15104 5500 15156
rect 7564 15104 7616 15156
rect 9772 15104 9824 15156
rect 11520 15147 11572 15156
rect 11520 15113 11529 15147
rect 11529 15113 11563 15147
rect 11563 15113 11572 15147
rect 11520 15104 11572 15113
rect 12164 15147 12216 15156
rect 12164 15113 12173 15147
rect 12173 15113 12207 15147
rect 12207 15113 12216 15147
rect 12164 15104 12216 15113
rect 14096 15104 14148 15156
rect 20628 15104 20680 15156
rect 22192 15104 22244 15156
rect 3516 15079 3568 15088
rect 3516 15045 3525 15079
rect 3525 15045 3559 15079
rect 3559 15045 3568 15079
rect 3516 15036 3568 15045
rect 7656 15079 7708 15088
rect 7656 15045 7665 15079
rect 7665 15045 7699 15079
rect 7699 15045 7708 15079
rect 7656 15036 7708 15045
rect 8300 15036 8352 15088
rect 9220 15079 9272 15088
rect 9220 15045 9229 15079
rect 9229 15045 9263 15079
rect 9263 15045 9272 15079
rect 9220 15036 9272 15045
rect 2596 15011 2648 15020
rect 2596 14977 2605 15011
rect 2605 14977 2639 15011
rect 2639 14977 2648 15011
rect 2596 14968 2648 14977
rect 3884 14968 3936 15020
rect 6368 14968 6420 15020
rect 7288 15011 7340 15020
rect 7288 14977 7297 15011
rect 7297 14977 7331 15011
rect 7331 14977 7340 15011
rect 7288 14968 7340 14977
rect 1952 14900 2004 14952
rect 2688 14900 2740 14952
rect 4252 14900 4304 14952
rect 7196 14900 7248 14952
rect 8392 15011 8444 15020
rect 8392 14977 8401 15011
rect 8401 14977 8435 15011
rect 8435 14977 8444 15011
rect 8392 14968 8444 14977
rect 11796 14968 11848 15020
rect 13084 14968 13136 15020
rect 13544 15011 13596 15020
rect 13544 14977 13553 15011
rect 13553 14977 13587 15011
rect 13587 14977 13596 15011
rect 13544 14968 13596 14977
rect 14280 15011 14332 15020
rect 14280 14977 14289 15011
rect 14289 14977 14323 15011
rect 14323 14977 14332 15011
rect 15568 15036 15620 15088
rect 15844 15079 15896 15088
rect 15844 15045 15853 15079
rect 15853 15045 15887 15079
rect 15887 15045 15896 15079
rect 15844 15036 15896 15045
rect 17592 15036 17644 15088
rect 14280 14968 14332 14977
rect 15108 15011 15160 15020
rect 15108 14977 15117 15011
rect 15117 14977 15151 15011
rect 15151 14977 15160 15011
rect 15108 14968 15160 14977
rect 16488 14968 16540 15020
rect 19156 15011 19208 15020
rect 19156 14977 19165 15011
rect 19165 14977 19199 15011
rect 19199 14977 19208 15011
rect 19156 14968 19208 14977
rect 21640 14968 21692 15020
rect 22836 14968 22888 15020
rect 23204 15011 23256 15020
rect 23204 14977 23213 15011
rect 23213 14977 23247 15011
rect 23247 14977 23256 15011
rect 23204 14968 23256 14977
rect 13268 14943 13320 14952
rect 13268 14909 13277 14943
rect 13277 14909 13311 14943
rect 13311 14909 13320 14943
rect 13268 14900 13320 14909
rect 14832 14943 14884 14952
rect 14832 14909 14841 14943
rect 14841 14909 14875 14943
rect 14875 14909 14884 14943
rect 14832 14900 14884 14909
rect 15292 14900 15344 14952
rect 17868 14900 17920 14952
rect 22008 14943 22060 14952
rect 22008 14909 22017 14943
rect 22017 14909 22051 14943
rect 22051 14909 22060 14943
rect 22008 14900 22060 14909
rect 5908 14832 5960 14884
rect 9496 14832 9548 14884
rect 14004 14832 14056 14884
rect 2964 14807 3016 14816
rect 2964 14773 2973 14807
rect 2973 14773 3007 14807
rect 3007 14773 3016 14807
rect 2964 14764 3016 14773
rect 3792 14764 3844 14816
rect 3976 14807 4028 14816
rect 3976 14773 3985 14807
rect 3985 14773 4019 14807
rect 4019 14773 4028 14807
rect 3976 14764 4028 14773
rect 4804 14764 4856 14816
rect 5172 14807 5224 14816
rect 5172 14773 5181 14807
rect 5181 14773 5215 14807
rect 5215 14773 5224 14807
rect 5172 14764 5224 14773
rect 5448 14764 5500 14816
rect 6368 14764 6420 14816
rect 6644 14764 6696 14816
rect 7840 14764 7892 14816
rect 11336 14764 11388 14816
rect 12900 14764 12952 14816
rect 16672 14832 16724 14884
rect 18604 14832 18656 14884
rect 23572 14832 23624 14884
rect 16488 14807 16540 14816
rect 16488 14773 16497 14807
rect 16497 14773 16531 14807
rect 16531 14773 16540 14807
rect 16488 14764 16540 14773
rect 17408 14807 17460 14816
rect 17408 14773 17417 14807
rect 17417 14773 17451 14807
rect 17451 14773 17460 14807
rect 17408 14764 17460 14773
rect 17868 14807 17920 14816
rect 17868 14773 17877 14807
rect 17877 14773 17911 14807
rect 17911 14773 17920 14807
rect 17868 14764 17920 14773
rect 18512 14807 18564 14816
rect 18512 14773 18521 14807
rect 18521 14773 18555 14807
rect 18555 14773 18564 14807
rect 18512 14764 18564 14773
rect 18972 14807 19024 14816
rect 18972 14773 18981 14807
rect 18981 14773 19015 14807
rect 19015 14773 19024 14807
rect 18972 14764 19024 14773
rect 19892 14807 19944 14816
rect 19892 14773 19901 14807
rect 19901 14773 19935 14807
rect 19935 14773 19944 14807
rect 20444 14807 20496 14816
rect 19892 14764 19944 14773
rect 20444 14773 20453 14807
rect 20453 14773 20487 14807
rect 20487 14773 20496 14807
rect 20444 14764 20496 14773
rect 20536 14807 20588 14816
rect 20536 14773 20545 14807
rect 20545 14773 20579 14807
rect 20579 14773 20588 14807
rect 20536 14764 20588 14773
rect 21272 14764 21324 14816
rect 21732 14764 21784 14816
rect 22928 14807 22980 14816
rect 22928 14773 22937 14807
rect 22937 14773 22971 14807
rect 22971 14773 22980 14807
rect 22928 14764 22980 14773
rect 27344 15011 27396 15020
rect 27344 14977 27353 15011
rect 27353 14977 27387 15011
rect 27387 14977 27396 15011
rect 27344 14968 27396 14977
rect 24308 14943 24360 14952
rect 24308 14909 24317 14943
rect 24317 14909 24351 14943
rect 24351 14909 24360 14943
rect 24308 14900 24360 14909
rect 26516 14900 26568 14952
rect 24400 14832 24452 14884
rect 27620 14832 27672 14884
rect 25136 14764 25188 14816
rect 25688 14807 25740 14816
rect 25688 14773 25697 14807
rect 25697 14773 25731 14807
rect 25731 14773 25740 14807
rect 25688 14764 25740 14773
rect 26608 14807 26660 14816
rect 26608 14773 26617 14807
rect 26617 14773 26651 14807
rect 26651 14773 26660 14807
rect 26608 14764 26660 14773
rect 26792 14807 26844 14816
rect 26792 14773 26801 14807
rect 26801 14773 26835 14807
rect 26835 14773 26844 14807
rect 26792 14764 26844 14773
rect 27344 14764 27396 14816
rect 10982 14662 11034 14714
rect 11046 14662 11098 14714
rect 11110 14662 11162 14714
rect 11174 14662 11226 14714
rect 20982 14662 21034 14714
rect 21046 14662 21098 14714
rect 21110 14662 21162 14714
rect 21174 14662 21226 14714
rect 2136 14560 2188 14612
rect 2044 14424 2096 14476
rect 2780 14560 2832 14612
rect 2964 14603 3016 14612
rect 2964 14569 2973 14603
rect 2973 14569 3007 14603
rect 3007 14569 3016 14603
rect 2964 14560 3016 14569
rect 3976 14560 4028 14612
rect 4620 14603 4672 14612
rect 4620 14569 4629 14603
rect 4629 14569 4663 14603
rect 4663 14569 4672 14603
rect 4620 14560 4672 14569
rect 4804 14560 4856 14612
rect 5908 14560 5960 14612
rect 7564 14560 7616 14612
rect 8484 14603 8536 14612
rect 8484 14569 8493 14603
rect 8493 14569 8527 14603
rect 8527 14569 8536 14603
rect 8484 14560 8536 14569
rect 12164 14560 12216 14612
rect 13268 14560 13320 14612
rect 13728 14560 13780 14612
rect 14096 14603 14148 14612
rect 14096 14569 14105 14603
rect 14105 14569 14139 14603
rect 14139 14569 14148 14603
rect 14096 14560 14148 14569
rect 16488 14560 16540 14612
rect 17132 14603 17184 14612
rect 17132 14569 17141 14603
rect 17141 14569 17175 14603
rect 17175 14569 17184 14603
rect 17132 14560 17184 14569
rect 18236 14603 18288 14612
rect 18236 14569 18245 14603
rect 18245 14569 18279 14603
rect 18279 14569 18288 14603
rect 18236 14560 18288 14569
rect 18512 14560 18564 14612
rect 20260 14560 20312 14612
rect 20628 14560 20680 14612
rect 21916 14560 21968 14612
rect 22836 14603 22888 14612
rect 22836 14569 22845 14603
rect 22845 14569 22879 14603
rect 22879 14569 22888 14603
rect 22836 14560 22888 14569
rect 23480 14603 23532 14612
rect 23480 14569 23489 14603
rect 23489 14569 23523 14603
rect 23523 14569 23532 14603
rect 23480 14560 23532 14569
rect 23756 14603 23808 14612
rect 23756 14569 23765 14603
rect 23765 14569 23799 14603
rect 23799 14569 23808 14603
rect 23756 14560 23808 14569
rect 26516 14560 26568 14612
rect 27252 14560 27304 14612
rect 5632 14492 5684 14544
rect 16396 14535 16448 14544
rect 16396 14501 16405 14535
rect 16405 14501 16439 14535
rect 16439 14501 16448 14535
rect 16396 14492 16448 14501
rect 19156 14492 19208 14544
rect 26424 14492 26476 14544
rect 4712 14424 4764 14476
rect 5540 14424 5592 14476
rect 9220 14424 9272 14476
rect 2412 14399 2464 14408
rect 2412 14365 2421 14399
rect 2421 14365 2455 14399
rect 2455 14365 2464 14399
rect 2412 14356 2464 14365
rect 3884 14356 3936 14408
rect 8300 14356 8352 14408
rect 9404 14356 9456 14408
rect 10324 14424 10376 14476
rect 11336 14467 11388 14476
rect 11336 14433 11370 14467
rect 11370 14433 11388 14467
rect 11336 14424 11388 14433
rect 14004 14467 14056 14476
rect 14004 14433 14013 14467
rect 14013 14433 14047 14467
rect 14047 14433 14056 14467
rect 14004 14424 14056 14433
rect 15660 14467 15712 14476
rect 15660 14433 15669 14467
rect 15669 14433 15703 14467
rect 15703 14433 15712 14467
rect 15660 14424 15712 14433
rect 16304 14424 16356 14476
rect 16488 14424 16540 14476
rect 19340 14424 19392 14476
rect 19708 14467 19760 14476
rect 19708 14433 19717 14467
rect 19717 14433 19751 14467
rect 19751 14433 19760 14467
rect 19708 14424 19760 14433
rect 22192 14424 22244 14476
rect 23480 14424 23532 14476
rect 26884 14467 26936 14476
rect 26884 14433 26893 14467
rect 26893 14433 26927 14467
rect 26927 14433 26936 14467
rect 26884 14424 26936 14433
rect 1676 14331 1728 14340
rect 1676 14297 1685 14331
rect 1685 14297 1719 14331
rect 1719 14297 1728 14331
rect 1676 14288 1728 14297
rect 2688 14288 2740 14340
rect 6736 14288 6788 14340
rect 7472 14288 7524 14340
rect 1492 14220 1544 14272
rect 2596 14220 2648 14272
rect 2964 14220 3016 14272
rect 4252 14263 4304 14272
rect 4252 14229 4261 14263
rect 4261 14229 4295 14263
rect 4295 14229 4304 14263
rect 4252 14220 4304 14229
rect 6828 14263 6880 14272
rect 6828 14229 6837 14263
rect 6837 14229 6871 14263
rect 6871 14229 6880 14263
rect 6828 14220 6880 14229
rect 7840 14263 7892 14272
rect 7840 14229 7849 14263
rect 7849 14229 7883 14263
rect 7883 14229 7892 14263
rect 7840 14220 7892 14229
rect 9128 14263 9180 14272
rect 9128 14229 9137 14263
rect 9137 14229 9171 14263
rect 9171 14229 9180 14263
rect 9128 14220 9180 14229
rect 9496 14263 9548 14272
rect 9496 14229 9505 14263
rect 9505 14229 9539 14263
rect 9539 14229 9548 14263
rect 9496 14220 9548 14229
rect 10324 14263 10376 14272
rect 10324 14229 10333 14263
rect 10333 14229 10367 14263
rect 10367 14229 10376 14263
rect 10324 14220 10376 14229
rect 10876 14263 10928 14272
rect 10876 14229 10885 14263
rect 10885 14229 10919 14263
rect 10919 14229 10928 14263
rect 10876 14220 10928 14229
rect 13820 14356 13872 14408
rect 15844 14399 15896 14408
rect 15844 14365 15853 14399
rect 15853 14365 15887 14399
rect 15887 14365 15896 14399
rect 15844 14356 15896 14365
rect 16764 14356 16816 14408
rect 17776 14399 17828 14408
rect 17776 14365 17785 14399
rect 17785 14365 17819 14399
rect 17819 14365 17828 14399
rect 17776 14356 17828 14365
rect 20076 14356 20128 14408
rect 20812 14356 20864 14408
rect 13544 14288 13596 14340
rect 23848 14356 23900 14408
rect 26976 14399 27028 14408
rect 11428 14220 11480 14272
rect 16672 14263 16724 14272
rect 16672 14229 16681 14263
rect 16681 14229 16715 14263
rect 16715 14229 16724 14263
rect 16672 14220 16724 14229
rect 18512 14263 18564 14272
rect 18512 14229 18521 14263
rect 18521 14229 18555 14263
rect 18555 14229 18564 14263
rect 18512 14220 18564 14229
rect 18972 14220 19024 14272
rect 19248 14263 19300 14272
rect 19248 14229 19257 14263
rect 19257 14229 19291 14263
rect 19291 14229 19300 14263
rect 19248 14220 19300 14229
rect 21088 14263 21140 14272
rect 21088 14229 21097 14263
rect 21097 14229 21131 14263
rect 21131 14229 21140 14263
rect 21088 14220 21140 14229
rect 26976 14365 26985 14399
rect 26985 14365 27019 14399
rect 27019 14365 27028 14399
rect 26976 14356 27028 14365
rect 27712 14288 27764 14340
rect 24308 14220 24360 14272
rect 25872 14220 25924 14272
rect 26332 14220 26384 14272
rect 26884 14220 26936 14272
rect 27160 14220 27212 14272
rect 5982 14118 6034 14170
rect 6046 14118 6098 14170
rect 6110 14118 6162 14170
rect 6174 14118 6226 14170
rect 15982 14118 16034 14170
rect 16046 14118 16098 14170
rect 16110 14118 16162 14170
rect 16174 14118 16226 14170
rect 25982 14118 26034 14170
rect 26046 14118 26098 14170
rect 26110 14118 26162 14170
rect 26174 14118 26226 14170
rect 2044 14059 2096 14068
rect 2044 14025 2053 14059
rect 2053 14025 2087 14059
rect 2087 14025 2096 14059
rect 2044 14016 2096 14025
rect 2412 14059 2464 14068
rect 2412 14025 2421 14059
rect 2421 14025 2455 14059
rect 2455 14025 2464 14059
rect 2412 14016 2464 14025
rect 4712 14016 4764 14068
rect 5264 14016 5316 14068
rect 5540 14016 5592 14068
rect 6552 14059 6604 14068
rect 6552 14025 6561 14059
rect 6561 14025 6595 14059
rect 6595 14025 6604 14059
rect 6552 14016 6604 14025
rect 8300 14059 8352 14068
rect 8300 14025 8309 14059
rect 8309 14025 8343 14059
rect 8343 14025 8352 14059
rect 8300 14016 8352 14025
rect 9588 14016 9640 14068
rect 10324 14016 10376 14068
rect 14740 14059 14792 14068
rect 14740 14025 14749 14059
rect 14749 14025 14783 14059
rect 14783 14025 14792 14059
rect 14740 14016 14792 14025
rect 16488 14059 16540 14068
rect 16488 14025 16497 14059
rect 16497 14025 16531 14059
rect 16531 14025 16540 14059
rect 16488 14016 16540 14025
rect 20076 14059 20128 14068
rect 20076 14025 20085 14059
rect 20085 14025 20119 14059
rect 20119 14025 20128 14059
rect 20076 14016 20128 14025
rect 21364 14016 21416 14068
rect 22008 14016 22060 14068
rect 23480 14059 23532 14068
rect 23480 14025 23489 14059
rect 23489 14025 23523 14059
rect 23523 14025 23532 14059
rect 23480 14016 23532 14025
rect 24216 14059 24268 14068
rect 24216 14025 24225 14059
rect 24225 14025 24259 14059
rect 24259 14025 24268 14059
rect 24216 14016 24268 14025
rect 25320 14059 25372 14068
rect 25320 14025 25329 14059
rect 25329 14025 25363 14059
rect 25363 14025 25372 14059
rect 25320 14016 25372 14025
rect 27712 14059 27764 14068
rect 27712 14025 27721 14059
rect 27721 14025 27755 14059
rect 27755 14025 27764 14059
rect 27712 14016 27764 14025
rect 1860 13948 1912 14000
rect 2596 13923 2648 13932
rect 2596 13889 2605 13923
rect 2605 13889 2639 13923
rect 2639 13889 2648 13923
rect 2596 13880 2648 13889
rect 1676 13812 1728 13864
rect 2872 13787 2924 13796
rect 2872 13753 2906 13787
rect 2906 13753 2924 13787
rect 2872 13744 2924 13753
rect 6276 13948 6328 14000
rect 10600 13991 10652 14000
rect 10600 13957 10609 13991
rect 10609 13957 10643 13991
rect 10643 13957 10652 13991
rect 10600 13948 10652 13957
rect 13820 13991 13872 14000
rect 13820 13957 13829 13991
rect 13829 13957 13863 13991
rect 13863 13957 13872 13991
rect 13820 13948 13872 13957
rect 16672 13948 16724 14000
rect 19432 13991 19484 14000
rect 19432 13957 19441 13991
rect 19441 13957 19475 13991
rect 19475 13957 19484 13991
rect 19432 13948 19484 13957
rect 26976 13948 27028 14000
rect 6368 13880 6420 13932
rect 9496 13880 9548 13932
rect 10416 13880 10468 13932
rect 5540 13855 5592 13864
rect 5540 13821 5549 13855
rect 5549 13821 5583 13855
rect 5583 13821 5592 13855
rect 5540 13812 5592 13821
rect 6552 13812 6604 13864
rect 5724 13744 5776 13796
rect 6736 13744 6788 13796
rect 3884 13676 3936 13728
rect 4528 13676 4580 13728
rect 5908 13676 5960 13728
rect 7012 13676 7064 13728
rect 7104 13676 7156 13728
rect 8208 13812 8260 13864
rect 9128 13812 9180 13864
rect 8576 13676 8628 13728
rect 10324 13812 10376 13864
rect 10876 13880 10928 13932
rect 11428 13880 11480 13932
rect 15844 13880 15896 13932
rect 11888 13855 11940 13864
rect 11888 13821 11897 13855
rect 11897 13821 11931 13855
rect 11931 13821 11940 13855
rect 11888 13812 11940 13821
rect 13084 13812 13136 13864
rect 14740 13812 14792 13864
rect 15752 13812 15804 13864
rect 16028 13855 16080 13864
rect 16028 13821 16037 13855
rect 16037 13821 16071 13855
rect 16071 13821 16080 13855
rect 16028 13812 16080 13821
rect 16304 13812 16356 13864
rect 16396 13812 16448 13864
rect 16764 13855 16816 13864
rect 16764 13821 16773 13855
rect 16773 13821 16807 13855
rect 16807 13821 16816 13855
rect 16764 13812 16816 13821
rect 17776 13812 17828 13864
rect 21088 13855 21140 13864
rect 11520 13744 11572 13796
rect 12716 13787 12768 13796
rect 12716 13753 12750 13787
rect 12750 13753 12768 13787
rect 12716 13744 12768 13753
rect 14188 13744 14240 13796
rect 17408 13744 17460 13796
rect 10232 13719 10284 13728
rect 10232 13685 10241 13719
rect 10241 13685 10275 13719
rect 10275 13685 10284 13719
rect 10232 13676 10284 13685
rect 10876 13676 10928 13728
rect 14924 13676 14976 13728
rect 15568 13676 15620 13728
rect 16580 13676 16632 13728
rect 17132 13676 17184 13728
rect 17868 13744 17920 13796
rect 18236 13744 18288 13796
rect 20812 13676 20864 13728
rect 21088 13821 21097 13855
rect 21097 13821 21131 13855
rect 21131 13821 21140 13855
rect 21088 13812 21140 13821
rect 23480 13880 23532 13932
rect 25688 13880 25740 13932
rect 24676 13855 24728 13864
rect 24676 13821 24685 13855
rect 24685 13821 24719 13855
rect 24719 13821 24728 13855
rect 24676 13812 24728 13821
rect 22100 13744 22152 13796
rect 22192 13676 22244 13728
rect 23848 13676 23900 13728
rect 25872 13812 25924 13864
rect 24584 13719 24636 13728
rect 24584 13685 24593 13719
rect 24593 13685 24627 13719
rect 24627 13685 24636 13719
rect 24584 13676 24636 13685
rect 27160 13719 27212 13728
rect 27160 13685 27169 13719
rect 27169 13685 27203 13719
rect 27203 13685 27212 13719
rect 27160 13676 27212 13685
rect 10982 13574 11034 13626
rect 11046 13574 11098 13626
rect 11110 13574 11162 13626
rect 11174 13574 11226 13626
rect 20982 13574 21034 13626
rect 21046 13574 21098 13626
rect 21110 13574 21162 13626
rect 21174 13574 21226 13626
rect 2504 13472 2556 13524
rect 4528 13515 4580 13524
rect 4528 13481 4537 13515
rect 4537 13481 4571 13515
rect 4571 13481 4580 13515
rect 4528 13472 4580 13481
rect 6368 13472 6420 13524
rect 3884 13447 3936 13456
rect 3884 13413 3893 13447
rect 3893 13413 3927 13447
rect 3927 13413 3936 13447
rect 3884 13404 3936 13413
rect 6920 13472 6972 13524
rect 9772 13472 9824 13524
rect 10048 13515 10100 13524
rect 10048 13481 10057 13515
rect 10057 13481 10091 13515
rect 10091 13481 10100 13515
rect 10048 13472 10100 13481
rect 10232 13472 10284 13524
rect 11336 13472 11388 13524
rect 11520 13515 11572 13524
rect 11520 13481 11529 13515
rect 11529 13481 11563 13515
rect 11563 13481 11572 13515
rect 11520 13472 11572 13481
rect 11796 13472 11848 13524
rect 13728 13472 13780 13524
rect 14096 13515 14148 13524
rect 14096 13481 14105 13515
rect 14105 13481 14139 13515
rect 14139 13481 14148 13515
rect 14096 13472 14148 13481
rect 16672 13472 16724 13524
rect 18236 13472 18288 13524
rect 19248 13472 19300 13524
rect 20260 13515 20312 13524
rect 20260 13481 20269 13515
rect 20269 13481 20303 13515
rect 20303 13481 20312 13515
rect 20260 13472 20312 13481
rect 20720 13472 20772 13524
rect 22744 13515 22796 13524
rect 22744 13481 22753 13515
rect 22753 13481 22787 13515
rect 22787 13481 22796 13515
rect 22744 13472 22796 13481
rect 23204 13472 23256 13524
rect 23480 13472 23532 13524
rect 24492 13472 24544 13524
rect 25872 13515 25924 13524
rect 25872 13481 25881 13515
rect 25881 13481 25915 13515
rect 25915 13481 25924 13515
rect 25872 13472 25924 13481
rect 27620 13515 27672 13524
rect 27620 13481 27629 13515
rect 27629 13481 27663 13515
rect 27663 13481 27672 13515
rect 27620 13472 27672 13481
rect 1492 13379 1544 13388
rect 1492 13345 1501 13379
rect 1501 13345 1535 13379
rect 1535 13345 1544 13379
rect 1492 13336 1544 13345
rect 2320 13336 2372 13388
rect 4620 13336 4672 13388
rect 6828 13404 6880 13456
rect 7380 13447 7432 13456
rect 7380 13413 7414 13447
rect 7414 13413 7432 13447
rect 7380 13404 7432 13413
rect 14924 13447 14976 13456
rect 14924 13413 14933 13447
rect 14933 13413 14967 13447
rect 14967 13413 14976 13447
rect 14924 13404 14976 13413
rect 19616 13447 19668 13456
rect 19616 13413 19625 13447
rect 19625 13413 19659 13447
rect 19659 13413 19668 13447
rect 19616 13404 19668 13413
rect 20904 13404 20956 13456
rect 21364 13404 21416 13456
rect 24584 13404 24636 13456
rect 2872 13243 2924 13252
rect 2872 13209 2881 13243
rect 2881 13209 2915 13243
rect 2915 13209 2924 13243
rect 2872 13200 2924 13209
rect 4804 13268 4856 13320
rect 5816 13336 5868 13388
rect 6368 13336 6420 13388
rect 7012 13336 7064 13388
rect 5540 13268 5592 13320
rect 6828 13268 6880 13320
rect 11336 13336 11388 13388
rect 11428 13336 11480 13388
rect 11796 13336 11848 13388
rect 5172 13200 5224 13252
rect 10416 13268 10468 13320
rect 11980 13311 12032 13320
rect 11980 13277 11989 13311
rect 11989 13277 12023 13311
rect 12023 13277 12032 13311
rect 11980 13268 12032 13277
rect 13912 13336 13964 13388
rect 15660 13336 15712 13388
rect 17500 13336 17552 13388
rect 14188 13311 14240 13320
rect 14188 13277 14197 13311
rect 14197 13277 14231 13311
rect 14231 13277 14240 13311
rect 14188 13268 14240 13277
rect 19708 13311 19760 13320
rect 12716 13200 12768 13252
rect 5816 13175 5868 13184
rect 5816 13141 5825 13175
rect 5825 13141 5859 13175
rect 5859 13141 5868 13175
rect 5816 13132 5868 13141
rect 7104 13132 7156 13184
rect 8024 13132 8076 13184
rect 8852 13132 8904 13184
rect 10968 13132 11020 13184
rect 12624 13175 12676 13184
rect 12624 13141 12633 13175
rect 12633 13141 12667 13175
rect 12667 13141 12676 13175
rect 12624 13132 12676 13141
rect 13636 13175 13688 13184
rect 13636 13141 13645 13175
rect 13645 13141 13679 13175
rect 13679 13141 13688 13175
rect 13636 13132 13688 13141
rect 15108 13132 15160 13184
rect 15384 13132 15436 13184
rect 15844 13132 15896 13184
rect 16304 13175 16356 13184
rect 16304 13141 16313 13175
rect 16313 13141 16347 13175
rect 16347 13141 16356 13175
rect 16304 13132 16356 13141
rect 19708 13277 19717 13311
rect 19717 13277 19751 13311
rect 19751 13277 19760 13311
rect 19708 13268 19760 13277
rect 19800 13311 19852 13320
rect 19800 13277 19809 13311
rect 19809 13277 19843 13311
rect 19843 13277 19852 13311
rect 19800 13268 19852 13277
rect 23756 13379 23808 13388
rect 23756 13345 23765 13379
rect 23765 13345 23799 13379
rect 23799 13345 23808 13379
rect 23756 13336 23808 13345
rect 24676 13379 24728 13388
rect 24676 13345 24685 13379
rect 24685 13345 24719 13379
rect 24719 13345 24728 13379
rect 24676 13336 24728 13345
rect 25688 13336 25740 13388
rect 27528 13336 27580 13388
rect 21640 13311 21692 13320
rect 21640 13277 21649 13311
rect 21649 13277 21683 13311
rect 21683 13277 21692 13311
rect 21640 13268 21692 13277
rect 21732 13268 21784 13320
rect 23204 13311 23256 13320
rect 23204 13277 23213 13311
rect 23213 13277 23247 13311
rect 23247 13277 23256 13311
rect 23204 13268 23256 13277
rect 25320 13268 25372 13320
rect 25872 13268 25924 13320
rect 26976 13311 27028 13320
rect 26976 13277 26985 13311
rect 26985 13277 27019 13311
rect 27019 13277 27028 13311
rect 26976 13268 27028 13277
rect 27160 13311 27212 13320
rect 27160 13277 27169 13311
rect 27169 13277 27203 13311
rect 27203 13277 27212 13311
rect 27160 13268 27212 13277
rect 23388 13200 23440 13252
rect 25596 13200 25648 13252
rect 26424 13200 26476 13252
rect 17132 13132 17184 13184
rect 17776 13132 17828 13184
rect 18328 13132 18380 13184
rect 22192 13175 22244 13184
rect 22192 13141 22201 13175
rect 22201 13141 22235 13175
rect 22235 13141 22244 13175
rect 22192 13132 22244 13141
rect 24308 13175 24360 13184
rect 24308 13141 24317 13175
rect 24317 13141 24351 13175
rect 24351 13141 24360 13175
rect 24308 13132 24360 13141
rect 25320 13175 25372 13184
rect 25320 13141 25329 13175
rect 25329 13141 25363 13175
rect 25363 13141 25372 13175
rect 25320 13132 25372 13141
rect 26332 13132 26384 13184
rect 5982 13030 6034 13082
rect 6046 13030 6098 13082
rect 6110 13030 6162 13082
rect 6174 13030 6226 13082
rect 15982 13030 16034 13082
rect 16046 13030 16098 13082
rect 16110 13030 16162 13082
rect 16174 13030 16226 13082
rect 25982 13030 26034 13082
rect 26046 13030 26098 13082
rect 26110 13030 26162 13082
rect 26174 13030 26226 13082
rect 572 12928 624 12980
rect 4620 12928 4672 12980
rect 4804 12971 4856 12980
rect 4804 12937 4813 12971
rect 4813 12937 4847 12971
rect 4847 12937 4856 12971
rect 4804 12928 4856 12937
rect 5540 12928 5592 12980
rect 7012 12928 7064 12980
rect 3056 12860 3108 12912
rect 4988 12860 5040 12912
rect 6184 12860 6236 12912
rect 6920 12860 6972 12912
rect 1492 12792 1544 12844
rect 4068 12792 4120 12844
rect 4528 12792 4580 12844
rect 5632 12792 5684 12844
rect 6552 12792 6604 12844
rect 11520 12928 11572 12980
rect 11980 12928 12032 12980
rect 14096 12928 14148 12980
rect 15844 12928 15896 12980
rect 17500 12971 17552 12980
rect 10876 12860 10928 12912
rect 11704 12860 11756 12912
rect 12164 12903 12216 12912
rect 12164 12869 12173 12903
rect 12173 12869 12207 12903
rect 12207 12869 12216 12903
rect 12164 12860 12216 12869
rect 14740 12903 14792 12912
rect 14740 12869 14749 12903
rect 14749 12869 14783 12903
rect 14783 12869 14792 12903
rect 14740 12860 14792 12869
rect 15108 12860 15160 12912
rect 10968 12792 11020 12844
rect 11980 12792 12032 12844
rect 2228 12724 2280 12776
rect 5172 12724 5224 12776
rect 7564 12767 7616 12776
rect 7564 12733 7573 12767
rect 7573 12733 7607 12767
rect 7607 12733 7616 12767
rect 7564 12724 7616 12733
rect 8852 12724 8904 12776
rect 12348 12792 12400 12844
rect 12624 12792 12676 12844
rect 16488 12860 16540 12912
rect 15384 12792 15436 12844
rect 16672 12792 16724 12844
rect 13912 12724 13964 12776
rect 15108 12724 15160 12776
rect 16580 12724 16632 12776
rect 17500 12937 17509 12971
rect 17509 12937 17543 12971
rect 17543 12937 17552 12971
rect 17500 12928 17552 12937
rect 19708 12928 19760 12980
rect 21916 12928 21968 12980
rect 22100 12928 22152 12980
rect 23020 12971 23072 12980
rect 23020 12937 23029 12971
rect 23029 12937 23063 12971
rect 23063 12937 23072 12971
rect 23020 12928 23072 12937
rect 23204 12928 23256 12980
rect 24492 12928 24544 12980
rect 25688 12971 25740 12980
rect 25688 12937 25697 12971
rect 25697 12937 25731 12971
rect 25731 12937 25740 12971
rect 25688 12928 25740 12937
rect 27160 12928 27212 12980
rect 17040 12835 17092 12844
rect 17040 12801 17049 12835
rect 17049 12801 17083 12835
rect 17083 12801 17092 12835
rect 20076 12860 20128 12912
rect 23756 12860 23808 12912
rect 17040 12792 17092 12801
rect 23204 12792 23256 12844
rect 24768 12860 24820 12912
rect 25872 12860 25924 12912
rect 17132 12724 17184 12776
rect 18328 12767 18380 12776
rect 18328 12733 18362 12767
rect 18362 12733 18380 12767
rect 5724 12656 5776 12708
rect 7472 12699 7524 12708
rect 7472 12665 7481 12699
rect 7481 12665 7515 12699
rect 7515 12665 7524 12699
rect 7472 12656 7524 12665
rect 16120 12656 16172 12708
rect 18328 12724 18380 12733
rect 20720 12767 20772 12776
rect 20720 12733 20729 12767
rect 20729 12733 20763 12767
rect 20763 12733 20772 12767
rect 20720 12724 20772 12733
rect 23112 12724 23164 12776
rect 23296 12724 23348 12776
rect 24400 12835 24452 12844
rect 24400 12801 24409 12835
rect 24409 12801 24443 12835
rect 24443 12801 24452 12835
rect 24400 12792 24452 12801
rect 27252 12792 27304 12844
rect 26148 12767 26200 12776
rect 26148 12733 26157 12767
rect 26157 12733 26191 12767
rect 26191 12733 26200 12767
rect 26148 12724 26200 12733
rect 26424 12767 26476 12776
rect 26424 12733 26458 12767
rect 26458 12733 26476 12767
rect 26424 12724 26476 12733
rect 27528 12724 27580 12776
rect 19248 12656 19300 12708
rect 19892 12656 19944 12708
rect 23480 12656 23532 12708
rect 24676 12656 24728 12708
rect 26976 12656 27028 12708
rect 27252 12656 27304 12708
rect 2320 12588 2372 12640
rect 2504 12588 2556 12640
rect 3424 12588 3476 12640
rect 5172 12631 5224 12640
rect 5172 12597 5181 12631
rect 5181 12597 5215 12631
rect 5215 12597 5224 12631
rect 5172 12588 5224 12597
rect 7288 12588 7340 12640
rect 10784 12631 10836 12640
rect 10784 12597 10793 12631
rect 10793 12597 10827 12631
rect 10827 12597 10836 12631
rect 10784 12588 10836 12597
rect 12440 12631 12492 12640
rect 12440 12597 12449 12631
rect 12449 12597 12483 12631
rect 12483 12597 12492 12631
rect 12440 12588 12492 12597
rect 12716 12588 12768 12640
rect 12992 12588 13044 12640
rect 17132 12588 17184 12640
rect 19340 12588 19392 12640
rect 23756 12631 23808 12640
rect 23756 12597 23765 12631
rect 23765 12597 23799 12631
rect 23799 12597 23808 12631
rect 23756 12588 23808 12597
rect 27160 12588 27212 12640
rect 10982 12486 11034 12538
rect 11046 12486 11098 12538
rect 11110 12486 11162 12538
rect 11174 12486 11226 12538
rect 20982 12486 21034 12538
rect 21046 12486 21098 12538
rect 21110 12486 21162 12538
rect 21174 12486 21226 12538
rect 2228 12427 2280 12436
rect 2228 12393 2237 12427
rect 2237 12393 2271 12427
rect 2271 12393 2280 12427
rect 2228 12384 2280 12393
rect 3700 12384 3752 12436
rect 5816 12384 5868 12436
rect 7012 12427 7064 12436
rect 7012 12393 7021 12427
rect 7021 12393 7055 12427
rect 7055 12393 7064 12427
rect 7012 12384 7064 12393
rect 7104 12427 7156 12436
rect 7104 12393 7113 12427
rect 7113 12393 7147 12427
rect 7147 12393 7156 12427
rect 7104 12384 7156 12393
rect 8208 12384 8260 12436
rect 8852 12427 8904 12436
rect 8852 12393 8861 12427
rect 8861 12393 8895 12427
rect 8895 12393 8904 12427
rect 8852 12384 8904 12393
rect 10416 12384 10468 12436
rect 10784 12384 10836 12436
rect 11796 12384 11848 12436
rect 12716 12384 12768 12436
rect 14004 12427 14056 12436
rect 14004 12393 14013 12427
rect 14013 12393 14047 12427
rect 14047 12393 14056 12427
rect 14004 12384 14056 12393
rect 15108 12384 15160 12436
rect 5172 12316 5224 12368
rect 5724 12316 5776 12368
rect 10876 12359 10928 12368
rect 10876 12325 10910 12359
rect 10910 12325 10928 12359
rect 10876 12316 10928 12325
rect 11428 12316 11480 12368
rect 12348 12316 12400 12368
rect 14188 12316 14240 12368
rect 15844 12384 15896 12436
rect 17040 12427 17092 12436
rect 17040 12393 17049 12427
rect 17049 12393 17083 12427
rect 17083 12393 17092 12427
rect 17040 12384 17092 12393
rect 18328 12384 18380 12436
rect 19616 12384 19668 12436
rect 19800 12384 19852 12436
rect 21732 12384 21784 12436
rect 22744 12384 22796 12436
rect 23112 12384 23164 12436
rect 26516 12384 26568 12436
rect 26976 12427 27028 12436
rect 26976 12393 26985 12427
rect 26985 12393 27019 12427
rect 27019 12393 27028 12427
rect 26976 12384 27028 12393
rect 16120 12316 16172 12368
rect 16304 12316 16356 12368
rect 1676 12180 1728 12232
rect 2412 12087 2464 12096
rect 2412 12053 2421 12087
rect 2421 12053 2455 12087
rect 2455 12053 2464 12087
rect 2412 12044 2464 12053
rect 2872 12291 2924 12300
rect 2872 12257 2881 12291
rect 2881 12257 2915 12291
rect 2915 12257 2924 12291
rect 2872 12248 2924 12257
rect 4160 12248 4212 12300
rect 6368 12248 6420 12300
rect 6644 12248 6696 12300
rect 7564 12291 7616 12300
rect 7564 12257 7573 12291
rect 7573 12257 7607 12291
rect 7607 12257 7616 12291
rect 15936 12291 15988 12300
rect 7564 12248 7616 12257
rect 15936 12257 15945 12291
rect 15945 12257 15979 12291
rect 15979 12257 15988 12291
rect 15936 12248 15988 12257
rect 16488 12248 16540 12300
rect 17132 12291 17184 12300
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 17776 12248 17828 12300
rect 21548 12316 21600 12368
rect 3516 12180 3568 12232
rect 5908 12223 5960 12232
rect 5908 12189 5917 12223
rect 5917 12189 5951 12223
rect 5951 12189 5960 12223
rect 5908 12180 5960 12189
rect 5080 12112 5132 12164
rect 7656 12223 7708 12232
rect 7656 12189 7665 12223
rect 7665 12189 7699 12223
rect 7699 12189 7708 12223
rect 10600 12223 10652 12232
rect 7656 12180 7708 12189
rect 10600 12189 10609 12223
rect 10609 12189 10643 12223
rect 10643 12189 10652 12223
rect 10600 12180 10652 12189
rect 16672 12180 16724 12232
rect 16948 12180 17000 12232
rect 22192 12248 22244 12300
rect 23848 12316 23900 12368
rect 26148 12359 26200 12368
rect 26148 12325 26157 12359
rect 26157 12325 26191 12359
rect 26191 12325 26200 12359
rect 26148 12316 26200 12325
rect 23480 12248 23532 12300
rect 24400 12248 24452 12300
rect 25320 12291 25372 12300
rect 25320 12257 25329 12291
rect 25329 12257 25363 12291
rect 25363 12257 25372 12291
rect 25320 12248 25372 12257
rect 25596 12248 25648 12300
rect 26516 12248 26568 12300
rect 23388 12223 23440 12232
rect 23388 12189 23397 12223
rect 23397 12189 23431 12223
rect 23431 12189 23440 12223
rect 23388 12180 23440 12189
rect 27160 12223 27212 12232
rect 27160 12189 27169 12223
rect 27169 12189 27203 12223
rect 27203 12189 27212 12223
rect 27160 12180 27212 12189
rect 6552 12112 6604 12164
rect 21640 12112 21692 12164
rect 3884 12087 3936 12096
rect 3884 12053 3893 12087
rect 3893 12053 3927 12087
rect 3927 12053 3936 12087
rect 3884 12044 3936 12053
rect 4252 12087 4304 12096
rect 4252 12053 4261 12087
rect 4261 12053 4295 12087
rect 4295 12053 4304 12087
rect 4252 12044 4304 12053
rect 4620 12087 4672 12096
rect 4620 12053 4629 12087
rect 4629 12053 4663 12087
rect 4663 12053 4672 12087
rect 4620 12044 4672 12053
rect 5540 12044 5592 12096
rect 8116 12087 8168 12096
rect 8116 12053 8125 12087
rect 8125 12053 8159 12087
rect 8159 12053 8168 12087
rect 8116 12044 8168 12053
rect 10232 12087 10284 12096
rect 10232 12053 10241 12087
rect 10241 12053 10275 12087
rect 10275 12053 10284 12087
rect 10232 12044 10284 12053
rect 20168 12044 20220 12096
rect 24952 12044 25004 12096
rect 25872 12044 25924 12096
rect 5982 11942 6034 11994
rect 6046 11942 6098 11994
rect 6110 11942 6162 11994
rect 6174 11942 6226 11994
rect 15982 11942 16034 11994
rect 16046 11942 16098 11994
rect 16110 11942 16162 11994
rect 16174 11942 16226 11994
rect 25982 11942 26034 11994
rect 26046 11942 26098 11994
rect 26110 11942 26162 11994
rect 26174 11942 26226 11994
rect 2504 11840 2556 11892
rect 4160 11883 4212 11892
rect 4160 11849 4169 11883
rect 4169 11849 4203 11883
rect 4203 11849 4212 11883
rect 4160 11840 4212 11849
rect 5080 11883 5132 11892
rect 5080 11849 5089 11883
rect 5089 11849 5123 11883
rect 5123 11849 5132 11883
rect 5080 11840 5132 11849
rect 6368 11840 6420 11892
rect 6644 11883 6696 11892
rect 6644 11849 6653 11883
rect 6653 11849 6687 11883
rect 6687 11849 6696 11883
rect 6644 11840 6696 11849
rect 7564 11840 7616 11892
rect 9220 11840 9272 11892
rect 9404 11883 9456 11892
rect 9404 11849 9413 11883
rect 9413 11849 9447 11883
rect 9447 11849 9456 11883
rect 9404 11840 9456 11849
rect 10048 11883 10100 11892
rect 10048 11849 10057 11883
rect 10057 11849 10091 11883
rect 10091 11849 10100 11883
rect 10048 11840 10100 11849
rect 10600 11840 10652 11892
rect 11888 11840 11940 11892
rect 15384 11840 15436 11892
rect 15844 11840 15896 11892
rect 16396 11883 16448 11892
rect 16396 11849 16405 11883
rect 16405 11849 16439 11883
rect 16439 11849 16448 11883
rect 16396 11840 16448 11849
rect 17132 11840 17184 11892
rect 17776 11883 17828 11892
rect 17776 11849 17785 11883
rect 17785 11849 17819 11883
rect 17819 11849 17828 11883
rect 17776 11840 17828 11849
rect 19892 11840 19944 11892
rect 21548 11840 21600 11892
rect 9956 11815 10008 11824
rect 9956 11781 9965 11815
rect 9965 11781 9999 11815
rect 9999 11781 10008 11815
rect 11428 11815 11480 11824
rect 9956 11772 10008 11781
rect 7380 11747 7432 11756
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7380 11704 7432 11713
rect 7564 11704 7616 11756
rect 8116 11704 8168 11756
rect 8852 11704 8904 11756
rect 2228 11636 2280 11688
rect 7104 11636 7156 11688
rect 7288 11679 7340 11688
rect 7288 11645 7297 11679
rect 7297 11645 7331 11679
rect 7331 11645 7340 11679
rect 11428 11781 11437 11815
rect 11437 11781 11471 11815
rect 11471 11781 11480 11815
rect 11428 11772 11480 11781
rect 20996 11772 21048 11824
rect 22744 11772 22796 11824
rect 10600 11747 10652 11756
rect 10600 11713 10609 11747
rect 10609 11713 10643 11747
rect 10643 11713 10652 11747
rect 10600 11704 10652 11713
rect 10784 11704 10836 11756
rect 17040 11747 17092 11756
rect 17040 11713 17049 11747
rect 17049 11713 17083 11747
rect 17083 11713 17092 11747
rect 17040 11704 17092 11713
rect 19800 11704 19852 11756
rect 21364 11704 21416 11756
rect 7288 11636 7340 11645
rect 19340 11636 19392 11688
rect 4804 11568 4856 11620
rect 5264 11568 5316 11620
rect 5724 11568 5776 11620
rect 2228 11500 2280 11552
rect 3424 11500 3476 11552
rect 5172 11543 5224 11552
rect 5172 11509 5181 11543
rect 5181 11509 5215 11543
rect 5215 11509 5224 11543
rect 5172 11500 5224 11509
rect 5540 11543 5592 11552
rect 5540 11509 5549 11543
rect 5549 11509 5583 11543
rect 5583 11509 5592 11543
rect 5540 11500 5592 11509
rect 9220 11568 9272 11620
rect 11796 11611 11848 11620
rect 11796 11577 11805 11611
rect 11805 11577 11839 11611
rect 11839 11577 11848 11611
rect 11796 11568 11848 11577
rect 16488 11568 16540 11620
rect 19248 11568 19300 11620
rect 8852 11543 8904 11552
rect 8852 11509 8861 11543
rect 8861 11509 8895 11543
rect 8895 11509 8904 11543
rect 8852 11500 8904 11509
rect 10508 11543 10560 11552
rect 10508 11509 10517 11543
rect 10517 11509 10551 11543
rect 10551 11509 10560 11543
rect 10508 11500 10560 11509
rect 15752 11500 15804 11552
rect 16856 11543 16908 11552
rect 16856 11509 16865 11543
rect 16865 11509 16899 11543
rect 16899 11509 16908 11543
rect 18420 11543 18472 11552
rect 16856 11500 16908 11509
rect 18420 11509 18429 11543
rect 18429 11509 18463 11543
rect 18463 11509 18472 11543
rect 18420 11500 18472 11509
rect 18880 11543 18932 11552
rect 18880 11509 18889 11543
rect 18889 11509 18923 11543
rect 18923 11509 18932 11543
rect 18880 11500 18932 11509
rect 19708 11500 19760 11552
rect 20168 11568 20220 11620
rect 23204 11840 23256 11892
rect 24032 11883 24084 11892
rect 24032 11849 24041 11883
rect 24041 11849 24075 11883
rect 24075 11849 24084 11883
rect 24032 11840 24084 11849
rect 26516 11840 26568 11892
rect 26976 11883 27028 11892
rect 24676 11772 24728 11824
rect 26976 11849 26985 11883
rect 26985 11849 27019 11883
rect 27019 11849 27028 11883
rect 26976 11840 27028 11849
rect 27160 11840 27212 11892
rect 27068 11772 27120 11824
rect 24952 11704 25004 11756
rect 23388 11611 23440 11620
rect 23388 11577 23397 11611
rect 23397 11577 23431 11611
rect 23431 11577 23440 11611
rect 23388 11568 23440 11577
rect 24768 11636 24820 11688
rect 25872 11636 25924 11688
rect 26976 11636 27028 11688
rect 26516 11568 26568 11620
rect 22652 11543 22704 11552
rect 22652 11509 22661 11543
rect 22661 11509 22695 11543
rect 22695 11509 22704 11543
rect 22652 11500 22704 11509
rect 23848 11543 23900 11552
rect 23848 11509 23857 11543
rect 23857 11509 23891 11543
rect 23891 11509 23900 11543
rect 23848 11500 23900 11509
rect 24952 11500 25004 11552
rect 27344 11543 27396 11552
rect 27344 11509 27353 11543
rect 27353 11509 27387 11543
rect 27387 11509 27396 11543
rect 27344 11500 27396 11509
rect 10982 11398 11034 11450
rect 11046 11398 11098 11450
rect 11110 11398 11162 11450
rect 11174 11398 11226 11450
rect 20982 11398 21034 11450
rect 21046 11398 21098 11450
rect 21110 11398 21162 11450
rect 21174 11398 21226 11450
rect 2872 11296 2924 11348
rect 3516 11339 3568 11348
rect 3516 11305 3525 11339
rect 3525 11305 3559 11339
rect 3559 11305 3568 11339
rect 3516 11296 3568 11305
rect 7656 11296 7708 11348
rect 8392 11339 8444 11348
rect 8392 11305 8401 11339
rect 8401 11305 8435 11339
rect 8435 11305 8444 11339
rect 8392 11296 8444 11305
rect 9312 11339 9364 11348
rect 9312 11305 9321 11339
rect 9321 11305 9355 11339
rect 9355 11305 9364 11339
rect 9312 11296 9364 11305
rect 1400 11228 1452 11280
rect 2596 11228 2648 11280
rect 2780 11271 2832 11280
rect 2780 11237 2789 11271
rect 2789 11237 2823 11271
rect 2823 11237 2832 11271
rect 2780 11228 2832 11237
rect 3332 11228 3384 11280
rect 5448 11228 5500 11280
rect 6276 11228 6328 11280
rect 7564 11228 7616 11280
rect 10508 11296 10560 11348
rect 11336 11296 11388 11348
rect 12348 11296 12400 11348
rect 16856 11296 16908 11348
rect 16948 11296 17000 11348
rect 18880 11296 18932 11348
rect 22192 11296 22244 11348
rect 23480 11339 23532 11348
rect 23480 11305 23489 11339
rect 23489 11305 23523 11339
rect 23523 11305 23532 11339
rect 23480 11296 23532 11305
rect 12532 11228 12584 11280
rect 16304 11228 16356 11280
rect 4068 11203 4120 11212
rect 4068 11169 4077 11203
rect 4077 11169 4111 11203
rect 4111 11169 4120 11203
rect 4068 11160 4120 11169
rect 5724 11203 5776 11212
rect 5724 11169 5758 11203
rect 5758 11169 5776 11203
rect 5724 11160 5776 11169
rect 8300 11203 8352 11212
rect 8300 11169 8309 11203
rect 8309 11169 8343 11203
rect 8343 11169 8352 11203
rect 8300 11160 8352 11169
rect 10416 11160 10468 11212
rect 15476 11160 15528 11212
rect 17684 11160 17736 11212
rect 20812 11228 20864 11280
rect 22008 11228 22060 11280
rect 23756 11296 23808 11348
rect 24676 11339 24728 11348
rect 24676 11305 24685 11339
rect 24685 11305 24719 11339
rect 24719 11305 24728 11339
rect 24676 11296 24728 11305
rect 24952 11339 25004 11348
rect 24952 11305 24961 11339
rect 24961 11305 24995 11339
rect 24995 11305 25004 11339
rect 24952 11296 25004 11305
rect 26332 11339 26384 11348
rect 26332 11305 26341 11339
rect 26341 11305 26375 11339
rect 26375 11305 26384 11339
rect 26332 11296 26384 11305
rect 26516 11339 26568 11348
rect 26516 11305 26525 11339
rect 26525 11305 26559 11339
rect 26559 11305 26568 11339
rect 26516 11296 26568 11305
rect 2872 11135 2924 11144
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 2228 10999 2280 11008
rect 2228 10965 2237 10999
rect 2237 10965 2271 10999
rect 2271 10965 2280 10999
rect 2228 10956 2280 10965
rect 2320 10956 2372 11008
rect 4068 11024 4120 11076
rect 10692 11135 10744 11144
rect 7932 11067 7984 11076
rect 7932 11033 7941 11067
rect 7941 11033 7975 11067
rect 7975 11033 7984 11067
rect 7932 11024 7984 11033
rect 8300 11024 8352 11076
rect 10692 11101 10701 11135
rect 10701 11101 10735 11135
rect 10735 11101 10744 11135
rect 10692 11092 10744 11101
rect 10876 11135 10928 11144
rect 10876 11101 10885 11135
rect 10885 11101 10919 11135
rect 10919 11101 10928 11135
rect 10876 11092 10928 11101
rect 10600 11024 10652 11076
rect 11796 11024 11848 11076
rect 16948 11092 17000 11144
rect 17960 11092 18012 11144
rect 19800 11135 19852 11144
rect 19800 11101 19809 11135
rect 19809 11101 19843 11135
rect 19843 11101 19852 11135
rect 19800 11092 19852 11101
rect 23296 11160 23348 11212
rect 24308 11160 24360 11212
rect 25136 11160 25188 11212
rect 20812 11092 20864 11144
rect 21916 11092 21968 11144
rect 22100 11092 22152 11144
rect 24216 11135 24268 11144
rect 24216 11101 24225 11135
rect 24225 11101 24259 11135
rect 24259 11101 24268 11135
rect 24216 11092 24268 11101
rect 24860 11092 24912 11144
rect 27160 11092 27212 11144
rect 20628 11024 20680 11076
rect 21824 11024 21876 11076
rect 22284 11024 22336 11076
rect 25320 11024 25372 11076
rect 25412 11024 25464 11076
rect 4436 10956 4488 11008
rect 4804 10956 4856 11008
rect 4988 10999 5040 11008
rect 4988 10965 4997 10999
rect 4997 10965 5031 10999
rect 5031 10965 5040 10999
rect 4988 10956 5040 10965
rect 15752 10956 15804 11008
rect 18236 10956 18288 11008
rect 5982 10854 6034 10906
rect 6046 10854 6098 10906
rect 6110 10854 6162 10906
rect 6174 10854 6226 10906
rect 15982 10854 16034 10906
rect 16046 10854 16098 10906
rect 16110 10854 16162 10906
rect 16174 10854 16226 10906
rect 25982 10854 26034 10906
rect 26046 10854 26098 10906
rect 26110 10854 26162 10906
rect 26174 10854 26226 10906
rect 2688 10795 2740 10804
rect 2688 10761 2697 10795
rect 2697 10761 2731 10795
rect 2731 10761 2740 10795
rect 2688 10752 2740 10761
rect 3332 10752 3384 10804
rect 4160 10795 4212 10804
rect 4160 10761 4169 10795
rect 4169 10761 4203 10795
rect 4203 10761 4212 10795
rect 4160 10752 4212 10761
rect 5356 10752 5408 10804
rect 6828 10795 6880 10804
rect 6828 10761 6837 10795
rect 6837 10761 6871 10795
rect 6871 10761 6880 10795
rect 6828 10752 6880 10761
rect 10508 10752 10560 10804
rect 10876 10752 10928 10804
rect 11796 10795 11848 10804
rect 11796 10761 11805 10795
rect 11805 10761 11839 10795
rect 11839 10761 11848 10795
rect 11796 10752 11848 10761
rect 12348 10752 12400 10804
rect 12532 10752 12584 10804
rect 15384 10795 15436 10804
rect 15384 10761 15393 10795
rect 15393 10761 15427 10795
rect 15427 10761 15436 10795
rect 15384 10752 15436 10761
rect 15568 10752 15620 10804
rect 16304 10752 16356 10804
rect 17960 10752 18012 10804
rect 19800 10752 19852 10804
rect 21916 10752 21968 10804
rect 22008 10752 22060 10804
rect 22192 10752 22244 10804
rect 23388 10795 23440 10804
rect 23388 10761 23397 10795
rect 23397 10761 23431 10795
rect 23431 10761 23440 10795
rect 23388 10752 23440 10761
rect 24860 10752 24912 10804
rect 25136 10752 25188 10804
rect 26424 10795 26476 10804
rect 26424 10761 26433 10795
rect 26433 10761 26467 10795
rect 26467 10761 26476 10795
rect 26424 10752 26476 10761
rect 2872 10684 2924 10736
rect 3516 10616 3568 10668
rect 5724 10616 5776 10668
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 2228 10548 2280 10600
rect 3148 10548 3200 10600
rect 4252 10591 4304 10600
rect 4252 10557 4261 10591
rect 4261 10557 4295 10591
rect 4295 10557 4304 10591
rect 4252 10548 4304 10557
rect 4528 10591 4580 10600
rect 4528 10557 4562 10591
rect 4562 10557 4580 10591
rect 4528 10548 4580 10557
rect 4988 10548 5040 10600
rect 10692 10616 10744 10668
rect 15844 10684 15896 10736
rect 18144 10684 18196 10736
rect 16948 10659 17000 10668
rect 16948 10625 16957 10659
rect 16957 10625 16991 10659
rect 16991 10625 17000 10659
rect 16948 10616 17000 10625
rect 18328 10616 18380 10668
rect 26884 10659 26936 10668
rect 8392 10591 8444 10600
rect 8392 10557 8401 10591
rect 8401 10557 8435 10591
rect 8435 10557 8444 10591
rect 8392 10548 8444 10557
rect 10600 10591 10652 10600
rect 10600 10557 10609 10591
rect 10609 10557 10643 10591
rect 10643 10557 10652 10591
rect 10600 10548 10652 10557
rect 17592 10548 17644 10600
rect 18696 10548 18748 10600
rect 19708 10548 19760 10600
rect 20076 10591 20128 10600
rect 20076 10557 20110 10591
rect 20110 10557 20128 10591
rect 20076 10548 20128 10557
rect 23388 10548 23440 10600
rect 26884 10625 26893 10659
rect 26893 10625 26927 10659
rect 26927 10625 26936 10659
rect 26884 10616 26936 10625
rect 27160 10616 27212 10668
rect 27528 10616 27580 10668
rect 23940 10591 23992 10600
rect 23940 10557 23974 10591
rect 23974 10557 23992 10591
rect 2320 10480 2372 10532
rect 5080 10480 5132 10532
rect 1860 10412 1912 10464
rect 3148 10455 3200 10464
rect 3148 10421 3157 10455
rect 3157 10421 3191 10455
rect 3191 10421 3200 10455
rect 3148 10412 3200 10421
rect 4252 10412 4304 10464
rect 4804 10412 4856 10464
rect 5724 10480 5776 10532
rect 7196 10523 7248 10532
rect 7196 10489 7205 10523
rect 7205 10489 7239 10523
rect 7239 10489 7248 10523
rect 7196 10480 7248 10489
rect 10416 10480 10468 10532
rect 16672 10480 16724 10532
rect 18144 10480 18196 10532
rect 19156 10480 19208 10532
rect 23940 10548 23992 10557
rect 24216 10548 24268 10600
rect 26792 10591 26844 10600
rect 26792 10557 26801 10591
rect 26801 10557 26835 10591
rect 26835 10557 26844 10591
rect 26792 10548 26844 10557
rect 6184 10455 6236 10464
rect 6184 10421 6193 10455
rect 6193 10421 6227 10455
rect 6227 10421 6236 10455
rect 6184 10412 6236 10421
rect 8300 10455 8352 10464
rect 8300 10421 8309 10455
rect 8309 10421 8343 10455
rect 8343 10421 8352 10455
rect 8300 10412 8352 10421
rect 8668 10412 8720 10464
rect 10324 10412 10376 10464
rect 19708 10455 19760 10464
rect 19708 10421 19717 10455
rect 19717 10421 19751 10455
rect 19751 10421 19760 10455
rect 19708 10412 19760 10421
rect 24860 10480 24912 10532
rect 10982 10310 11034 10362
rect 11046 10310 11098 10362
rect 11110 10310 11162 10362
rect 11174 10310 11226 10362
rect 20982 10310 21034 10362
rect 21046 10310 21098 10362
rect 21110 10310 21162 10362
rect 21174 10310 21226 10362
rect 1952 10251 2004 10260
rect 1952 10217 1961 10251
rect 1961 10217 1995 10251
rect 1995 10217 2004 10251
rect 1952 10208 2004 10217
rect 2320 10251 2372 10260
rect 2320 10217 2329 10251
rect 2329 10217 2363 10251
rect 2363 10217 2372 10251
rect 2320 10208 2372 10217
rect 2412 10208 2464 10260
rect 3516 10251 3568 10260
rect 2872 10140 2924 10192
rect 3516 10217 3525 10251
rect 3525 10217 3559 10251
rect 3559 10217 3568 10251
rect 3516 10208 3568 10217
rect 4068 10208 4120 10260
rect 4436 10251 4488 10260
rect 4436 10217 4445 10251
rect 4445 10217 4479 10251
rect 4479 10217 4488 10251
rect 4436 10208 4488 10217
rect 5080 10251 5132 10260
rect 5080 10217 5089 10251
rect 5089 10217 5123 10251
rect 5123 10217 5132 10251
rect 5080 10208 5132 10217
rect 5632 10251 5684 10260
rect 4528 10140 4580 10192
rect 3056 10072 3108 10124
rect 3976 10072 4028 10124
rect 5632 10217 5641 10251
rect 5641 10217 5675 10251
rect 5675 10217 5684 10251
rect 5632 10208 5684 10217
rect 5724 10208 5776 10260
rect 6000 10251 6052 10260
rect 6000 10217 6009 10251
rect 6009 10217 6043 10251
rect 6043 10217 6052 10251
rect 6000 10208 6052 10217
rect 6552 10208 6604 10260
rect 7196 10208 7248 10260
rect 8484 10208 8536 10260
rect 9220 10208 9272 10260
rect 10600 10251 10652 10260
rect 10600 10217 10609 10251
rect 10609 10217 10643 10251
rect 10643 10217 10652 10251
rect 10600 10208 10652 10217
rect 15476 10208 15528 10260
rect 16672 10208 16724 10260
rect 17132 10251 17184 10260
rect 17132 10217 17141 10251
rect 17141 10217 17175 10251
rect 17175 10217 17184 10251
rect 17132 10208 17184 10217
rect 18328 10208 18380 10260
rect 19248 10251 19300 10260
rect 19248 10217 19257 10251
rect 19257 10217 19291 10251
rect 19291 10217 19300 10251
rect 19248 10208 19300 10217
rect 20076 10208 20128 10260
rect 20628 10208 20680 10260
rect 22008 10208 22060 10260
rect 23756 10208 23808 10260
rect 24400 10251 24452 10260
rect 24400 10217 24409 10251
rect 24409 10217 24443 10251
rect 24443 10217 24452 10251
rect 24400 10208 24452 10217
rect 25320 10208 25372 10260
rect 26700 10208 26752 10260
rect 26976 10251 27028 10260
rect 26976 10217 26985 10251
rect 26985 10217 27019 10251
rect 27019 10217 27028 10251
rect 26976 10208 27028 10217
rect 6092 10183 6144 10192
rect 6092 10149 6101 10183
rect 6101 10149 6135 10183
rect 6135 10149 6144 10183
rect 6092 10140 6144 10149
rect 6184 10140 6236 10192
rect 2136 9936 2188 9988
rect 3148 9936 3200 9988
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 18696 10140 18748 10192
rect 19064 10140 19116 10192
rect 20352 10140 20404 10192
rect 21180 10140 21232 10192
rect 23296 10140 23348 10192
rect 6920 10072 6972 10124
rect 17408 10072 17460 10124
rect 19156 10115 19208 10124
rect 19156 10081 19165 10115
rect 19165 10081 19199 10115
rect 19199 10081 19208 10115
rect 19156 10072 19208 10081
rect 19340 10072 19392 10124
rect 19524 10072 19576 10124
rect 23940 10072 23992 10124
rect 24124 10072 24176 10124
rect 25320 10115 25372 10124
rect 25320 10081 25329 10115
rect 25329 10081 25363 10115
rect 25363 10081 25372 10115
rect 25320 10072 25372 10081
rect 26792 10072 26844 10124
rect 6460 10004 6512 10056
rect 6644 10004 6696 10056
rect 3976 9936 4028 9988
rect 7196 9979 7248 9988
rect 7196 9945 7205 9979
rect 7205 9945 7239 9979
rect 7239 9945 7248 9979
rect 7196 9936 7248 9945
rect 8116 10004 8168 10056
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 17316 10047 17368 10056
rect 17316 10013 17325 10047
rect 17325 10013 17359 10047
rect 17359 10013 17368 10047
rect 17316 10004 17368 10013
rect 18236 10004 18288 10056
rect 18972 10004 19024 10056
rect 20168 10004 20220 10056
rect 21824 10004 21876 10056
rect 23112 10004 23164 10056
rect 27160 10047 27212 10056
rect 27160 10013 27169 10047
rect 27169 10013 27203 10047
rect 27203 10013 27212 10047
rect 27160 10004 27212 10013
rect 3884 9911 3936 9920
rect 3884 9877 3893 9911
rect 3893 9877 3927 9911
rect 3927 9877 3936 9911
rect 3884 9868 3936 9877
rect 16672 9911 16724 9920
rect 16672 9877 16681 9911
rect 16681 9877 16715 9911
rect 16715 9877 16724 9911
rect 16672 9868 16724 9877
rect 25596 9868 25648 9920
rect 5982 9766 6034 9818
rect 6046 9766 6098 9818
rect 6110 9766 6162 9818
rect 6174 9766 6226 9818
rect 15982 9766 16034 9818
rect 16046 9766 16098 9818
rect 16110 9766 16162 9818
rect 16174 9766 16226 9818
rect 25982 9766 26034 9818
rect 26046 9766 26098 9818
rect 26110 9766 26162 9818
rect 26174 9766 26226 9818
rect 2412 9664 2464 9716
rect 1952 9528 2004 9580
rect 2228 9571 2280 9580
rect 2228 9537 2237 9571
rect 2237 9537 2271 9571
rect 2271 9537 2280 9571
rect 2228 9528 2280 9537
rect 2964 9528 3016 9580
rect 3516 9664 3568 9716
rect 4528 9707 4580 9716
rect 4528 9673 4537 9707
rect 4537 9673 4571 9707
rect 4571 9673 4580 9707
rect 4528 9664 4580 9673
rect 5724 9664 5776 9716
rect 6368 9664 6420 9716
rect 6092 9596 6144 9648
rect 8116 9596 8168 9648
rect 15752 9596 15804 9648
rect 17132 9664 17184 9716
rect 19156 9664 19208 9716
rect 19064 9596 19116 9648
rect 21180 9664 21232 9716
rect 22008 9664 22060 9716
rect 24124 9707 24176 9716
rect 24124 9673 24133 9707
rect 24133 9673 24167 9707
rect 24167 9673 24176 9707
rect 24124 9664 24176 9673
rect 25320 9664 25372 9716
rect 26976 9664 27028 9716
rect 25504 9639 25556 9648
rect 4804 9460 4856 9512
rect 5816 9528 5868 9580
rect 15936 9571 15988 9580
rect 15936 9537 15945 9571
rect 15945 9537 15979 9571
rect 15979 9537 15988 9571
rect 16856 9571 16908 9580
rect 15936 9528 15988 9537
rect 16856 9537 16865 9571
rect 16865 9537 16899 9571
rect 16899 9537 16908 9571
rect 16856 9528 16908 9537
rect 17316 9528 17368 9580
rect 17776 9528 17828 9580
rect 25504 9605 25513 9639
rect 25513 9605 25547 9639
rect 25547 9605 25556 9639
rect 25504 9596 25556 9605
rect 1492 9392 1544 9444
rect 1676 9392 1728 9444
rect 1952 9435 2004 9444
rect 1952 9401 1961 9435
rect 1961 9401 1995 9435
rect 1995 9401 2004 9435
rect 1952 9392 2004 9401
rect 3424 9435 3476 9444
rect 3424 9401 3458 9435
rect 3458 9401 3476 9435
rect 3424 9392 3476 9401
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 5816 9367 5868 9376
rect 5816 9333 5825 9367
rect 5825 9333 5859 9367
rect 5859 9333 5868 9367
rect 5816 9324 5868 9333
rect 6460 9324 6512 9376
rect 18512 9503 18564 9512
rect 18512 9469 18521 9503
rect 18521 9469 18555 9503
rect 18555 9469 18564 9503
rect 18512 9460 18564 9469
rect 7104 9392 7156 9444
rect 15476 9392 15528 9444
rect 19892 9460 19944 9512
rect 24216 9503 24268 9512
rect 24216 9469 24225 9503
rect 24225 9469 24259 9503
rect 24259 9469 24268 9503
rect 24216 9460 24268 9469
rect 25228 9460 25280 9512
rect 27252 9596 27304 9648
rect 27528 9503 27580 9512
rect 19708 9392 19760 9444
rect 27528 9469 27537 9503
rect 27537 9469 27571 9503
rect 27571 9469 27580 9503
rect 27528 9460 27580 9469
rect 26792 9392 26844 9444
rect 7472 9324 7524 9376
rect 16396 9367 16448 9376
rect 16396 9333 16405 9367
rect 16405 9333 16439 9367
rect 16439 9333 16448 9367
rect 16396 9324 16448 9333
rect 17408 9367 17460 9376
rect 17408 9333 17417 9367
rect 17417 9333 17451 9367
rect 17451 9333 17460 9367
rect 17408 9324 17460 9333
rect 17776 9367 17828 9376
rect 17776 9333 17785 9367
rect 17785 9333 17819 9367
rect 17819 9333 17828 9367
rect 17776 9324 17828 9333
rect 19248 9367 19300 9376
rect 19248 9333 19257 9367
rect 19257 9333 19291 9367
rect 19291 9333 19300 9367
rect 19248 9324 19300 9333
rect 20260 9324 20312 9376
rect 22100 9367 22152 9376
rect 22100 9333 22109 9367
rect 22109 9333 22143 9367
rect 22143 9333 22152 9367
rect 24400 9367 24452 9376
rect 22100 9324 22152 9333
rect 24400 9333 24409 9367
rect 24409 9333 24443 9367
rect 24443 9333 24452 9367
rect 24400 9324 24452 9333
rect 26884 9324 26936 9376
rect 27804 9324 27856 9376
rect 10982 9222 11034 9274
rect 11046 9222 11098 9274
rect 11110 9222 11162 9274
rect 11174 9222 11226 9274
rect 20982 9222 21034 9274
rect 21046 9222 21098 9274
rect 21110 9222 21162 9274
rect 21174 9222 21226 9274
rect 1952 9120 2004 9172
rect 3424 9120 3476 9172
rect 4712 9120 4764 9172
rect 6092 9163 6144 9172
rect 6092 9129 6101 9163
rect 6101 9129 6135 9163
rect 6135 9129 6144 9163
rect 6092 9120 6144 9129
rect 7012 9120 7064 9172
rect 7380 9120 7432 9172
rect 7748 9120 7800 9172
rect 15476 9163 15528 9172
rect 15476 9129 15485 9163
rect 15485 9129 15519 9163
rect 15519 9129 15528 9163
rect 15476 9120 15528 9129
rect 18972 9120 19024 9172
rect 20720 9120 20772 9172
rect 21548 9120 21600 9172
rect 27160 9163 27212 9172
rect 27160 9129 27169 9163
rect 27169 9129 27203 9163
rect 27203 9129 27212 9163
rect 27160 9120 27212 9129
rect 1492 9052 1544 9104
rect 2780 9052 2832 9104
rect 4160 9052 4212 9104
rect 21456 9052 21508 9104
rect 5264 8984 5316 9036
rect 17776 8984 17828 9036
rect 19524 8984 19576 9036
rect 25320 9027 25372 9036
rect 25320 8993 25329 9027
rect 25329 8993 25363 9027
rect 25363 8993 25372 9027
rect 25320 8984 25372 8993
rect 26516 9027 26568 9036
rect 26516 8993 26525 9027
rect 26525 8993 26559 9027
rect 26559 8993 26568 9027
rect 26516 8984 26568 8993
rect 2228 8916 2280 8968
rect 2964 8916 3016 8968
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 7104 8916 7156 8968
rect 16488 8959 16540 8968
rect 6828 8848 6880 8900
rect 16488 8925 16497 8959
rect 16497 8925 16531 8959
rect 16531 8925 16540 8959
rect 16488 8916 16540 8925
rect 19708 8959 19760 8968
rect 19708 8925 19717 8959
rect 19717 8925 19751 8959
rect 19751 8925 19760 8959
rect 19708 8916 19760 8925
rect 19892 8959 19944 8968
rect 19892 8925 19901 8959
rect 19901 8925 19935 8959
rect 19935 8925 19944 8959
rect 19892 8916 19944 8925
rect 20812 8848 20864 8900
rect 21824 8916 21876 8968
rect 22100 8916 22152 8968
rect 21732 8848 21784 8900
rect 2136 8780 2188 8832
rect 8208 8780 8260 8832
rect 17868 8823 17920 8832
rect 17868 8789 17877 8823
rect 17877 8789 17911 8823
rect 17911 8789 17920 8823
rect 17868 8780 17920 8789
rect 18788 8823 18840 8832
rect 18788 8789 18797 8823
rect 18797 8789 18831 8823
rect 18831 8789 18840 8823
rect 18788 8780 18840 8789
rect 19340 8780 19392 8832
rect 20076 8780 20128 8832
rect 25504 8823 25556 8832
rect 25504 8789 25513 8823
rect 25513 8789 25547 8823
rect 25547 8789 25556 8823
rect 25504 8780 25556 8789
rect 25872 8780 25924 8832
rect 5982 8678 6034 8730
rect 6046 8678 6098 8730
rect 6110 8678 6162 8730
rect 6174 8678 6226 8730
rect 15982 8678 16034 8730
rect 16046 8678 16098 8730
rect 16110 8678 16162 8730
rect 16174 8678 16226 8730
rect 25982 8678 26034 8730
rect 26046 8678 26098 8730
rect 26110 8678 26162 8730
rect 26174 8678 26226 8730
rect 1492 8576 1544 8628
rect 4068 8576 4120 8628
rect 2780 8551 2832 8560
rect 2780 8517 2789 8551
rect 2789 8517 2823 8551
rect 2823 8517 2832 8551
rect 5540 8551 5592 8560
rect 2780 8508 2832 8517
rect 5540 8517 5549 8551
rect 5549 8517 5583 8551
rect 5583 8517 5592 8551
rect 5540 8508 5592 8517
rect 1584 8440 1636 8492
rect 1952 8440 2004 8492
rect 2688 8440 2740 8492
rect 3516 8440 3568 8492
rect 4252 8483 4304 8492
rect 4252 8449 4261 8483
rect 4261 8449 4295 8483
rect 4295 8449 4304 8483
rect 4252 8440 4304 8449
rect 5264 8440 5316 8492
rect 1676 8372 1728 8424
rect 2964 8372 3016 8424
rect 6552 8576 6604 8628
rect 6736 8576 6788 8628
rect 7748 8576 7800 8628
rect 16488 8576 16540 8628
rect 21456 8576 21508 8628
rect 22100 8576 22152 8628
rect 25320 8576 25372 8628
rect 25780 8576 25832 8628
rect 26516 8576 26568 8628
rect 27712 8619 27764 8628
rect 27712 8585 27721 8619
rect 27721 8585 27755 8619
rect 27755 8585 27764 8619
rect 27712 8576 27764 8585
rect 21640 8508 21692 8560
rect 26240 8508 26292 8560
rect 26608 8551 26660 8560
rect 26608 8517 26617 8551
rect 26617 8517 26651 8551
rect 26651 8517 26660 8551
rect 26608 8508 26660 8517
rect 7472 8483 7524 8492
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 8208 8440 8260 8492
rect 16672 8440 16724 8492
rect 17040 8483 17092 8492
rect 17040 8449 17049 8483
rect 17049 8449 17083 8483
rect 17083 8449 17092 8483
rect 17040 8440 17092 8449
rect 17868 8440 17920 8492
rect 19708 8440 19760 8492
rect 19892 8440 19944 8492
rect 20076 8483 20128 8492
rect 20076 8449 20085 8483
rect 20085 8449 20119 8483
rect 20119 8449 20128 8483
rect 20076 8440 20128 8449
rect 20260 8483 20312 8492
rect 20260 8449 20269 8483
rect 20269 8449 20303 8483
rect 20303 8449 20312 8483
rect 20260 8440 20312 8449
rect 21732 8483 21784 8492
rect 21732 8449 21741 8483
rect 21741 8449 21775 8483
rect 21775 8449 21784 8483
rect 21732 8440 21784 8449
rect 7196 8415 7248 8424
rect 7196 8381 7205 8415
rect 7205 8381 7239 8415
rect 7239 8381 7248 8415
rect 7196 8372 7248 8381
rect 8484 8372 8536 8424
rect 8852 8415 8904 8424
rect 8852 8381 8861 8415
rect 8861 8381 8895 8415
rect 8895 8381 8904 8415
rect 8852 8372 8904 8381
rect 16396 8372 16448 8424
rect 18788 8372 18840 8424
rect 19432 8372 19484 8424
rect 21364 8372 21416 8424
rect 21640 8415 21692 8424
rect 21640 8381 21649 8415
rect 21649 8381 21683 8415
rect 21683 8381 21692 8415
rect 21640 8372 21692 8381
rect 25780 8372 25832 8424
rect 26424 8415 26476 8424
rect 26424 8381 26433 8415
rect 26433 8381 26467 8415
rect 26467 8381 26476 8415
rect 26424 8372 26476 8381
rect 27344 8372 27396 8424
rect 2136 8347 2188 8356
rect 2136 8313 2145 8347
rect 2145 8313 2179 8347
rect 2179 8313 2188 8347
rect 2136 8304 2188 8313
rect 2320 8236 2372 8288
rect 3700 8236 3752 8288
rect 4712 8304 4764 8356
rect 6552 8304 6604 8356
rect 5264 8279 5316 8288
rect 5264 8245 5273 8279
rect 5273 8245 5307 8279
rect 5307 8245 5316 8279
rect 5264 8236 5316 8245
rect 8392 8236 8444 8288
rect 16396 8279 16448 8288
rect 16396 8245 16405 8279
rect 16405 8245 16439 8279
rect 16439 8245 16448 8279
rect 16396 8236 16448 8245
rect 17868 8236 17920 8288
rect 18420 8279 18472 8288
rect 18420 8245 18429 8279
rect 18429 8245 18463 8279
rect 18463 8245 18472 8279
rect 18420 8236 18472 8245
rect 25504 8279 25556 8288
rect 25504 8245 25513 8279
rect 25513 8245 25547 8279
rect 25547 8245 25556 8279
rect 25504 8236 25556 8245
rect 10982 8134 11034 8186
rect 11046 8134 11098 8186
rect 11110 8134 11162 8186
rect 11174 8134 11226 8186
rect 20982 8134 21034 8186
rect 21046 8134 21098 8186
rect 21110 8134 21162 8186
rect 21174 8134 21226 8186
rect 1676 8075 1728 8084
rect 1676 8041 1685 8075
rect 1685 8041 1719 8075
rect 1719 8041 1728 8075
rect 1676 8032 1728 8041
rect 1768 8032 1820 8084
rect 2872 8032 2924 8084
rect 3700 8032 3752 8084
rect 3884 8032 3936 8084
rect 4436 8075 4488 8084
rect 4436 8041 4445 8075
rect 4445 8041 4479 8075
rect 4479 8041 4488 8075
rect 4436 8032 4488 8041
rect 6644 8032 6696 8084
rect 6828 8075 6880 8084
rect 6828 8041 6837 8075
rect 6837 8041 6871 8075
rect 6871 8041 6880 8075
rect 6828 8032 6880 8041
rect 7380 8075 7432 8084
rect 7380 8041 7389 8075
rect 7389 8041 7423 8075
rect 7423 8041 7432 8075
rect 7380 8032 7432 8041
rect 16304 8032 16356 8084
rect 17776 8032 17828 8084
rect 19156 8032 19208 8084
rect 19340 8032 19392 8084
rect 20352 8032 20404 8084
rect 21364 8032 21416 8084
rect 21548 8075 21600 8084
rect 21548 8041 21557 8075
rect 21557 8041 21591 8075
rect 21591 8041 21600 8075
rect 21548 8032 21600 8041
rect 21732 8032 21784 8084
rect 2412 7964 2464 8016
rect 2688 7964 2740 8016
rect 2320 7939 2372 7948
rect 2320 7905 2329 7939
rect 2329 7905 2363 7939
rect 2363 7905 2372 7939
rect 2320 7896 2372 7905
rect 2412 7871 2464 7880
rect 2412 7837 2421 7871
rect 2421 7837 2455 7871
rect 2455 7837 2464 7871
rect 2412 7828 2464 7837
rect 2688 7828 2740 7880
rect 3148 7964 3200 8016
rect 4528 8007 4580 8016
rect 4528 7973 4537 8007
rect 4537 7973 4571 8007
rect 4571 7973 4580 8007
rect 4528 7964 4580 7973
rect 8944 7964 8996 8016
rect 19248 7964 19300 8016
rect 20260 8007 20312 8016
rect 20260 7973 20269 8007
rect 20269 7973 20303 8007
rect 20303 7973 20312 8007
rect 20260 7964 20312 7973
rect 6736 7939 6788 7948
rect 6736 7905 6745 7939
rect 6745 7905 6779 7939
rect 6779 7905 6788 7939
rect 6736 7896 6788 7905
rect 16580 7896 16632 7948
rect 17040 7939 17092 7948
rect 17040 7905 17074 7939
rect 17074 7905 17092 7939
rect 17040 7896 17092 7905
rect 3332 7828 3384 7880
rect 4712 7871 4764 7880
rect 4712 7837 4721 7871
rect 4721 7837 4755 7871
rect 4755 7837 4764 7871
rect 4712 7828 4764 7837
rect 5264 7828 5316 7880
rect 6368 7828 6420 7880
rect 7472 7828 7524 7880
rect 19064 7871 19116 7880
rect 19064 7837 19073 7871
rect 19073 7837 19107 7871
rect 19107 7837 19116 7871
rect 19064 7828 19116 7837
rect 19800 7828 19852 7880
rect 26240 7896 26292 7948
rect 26976 7896 27028 7948
rect 18420 7760 18472 7812
rect 7748 7735 7800 7744
rect 7748 7701 7757 7735
rect 7757 7701 7791 7735
rect 7791 7701 7800 7735
rect 7748 7692 7800 7701
rect 8116 7692 8168 7744
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 8392 7692 8444 7701
rect 18696 7692 18748 7744
rect 26792 7692 26844 7744
rect 5982 7590 6034 7642
rect 6046 7590 6098 7642
rect 6110 7590 6162 7642
rect 6174 7590 6226 7642
rect 15982 7590 16034 7642
rect 16046 7590 16098 7642
rect 16110 7590 16162 7642
rect 16174 7590 16226 7642
rect 25982 7590 26034 7642
rect 26046 7590 26098 7642
rect 26110 7590 26162 7642
rect 26174 7590 26226 7642
rect 2688 7488 2740 7540
rect 3516 7531 3568 7540
rect 3516 7497 3525 7531
rect 3525 7497 3559 7531
rect 3559 7497 3568 7531
rect 3516 7488 3568 7497
rect 3792 7531 3844 7540
rect 3792 7497 3801 7531
rect 3801 7497 3835 7531
rect 3835 7497 3844 7531
rect 3792 7488 3844 7497
rect 4436 7488 4488 7540
rect 4528 7531 4580 7540
rect 4528 7497 4537 7531
rect 4537 7497 4571 7531
rect 4571 7497 4580 7531
rect 5356 7531 5408 7540
rect 4528 7488 4580 7497
rect 5356 7497 5365 7531
rect 5365 7497 5399 7531
rect 5399 7497 5408 7531
rect 5356 7488 5408 7497
rect 6276 7488 6328 7540
rect 6736 7488 6788 7540
rect 16396 7488 16448 7540
rect 16580 7488 16632 7540
rect 18420 7488 18472 7540
rect 19248 7531 19300 7540
rect 19248 7497 19257 7531
rect 19257 7497 19291 7531
rect 19291 7497 19300 7531
rect 19248 7488 19300 7497
rect 19432 7488 19484 7540
rect 20352 7531 20404 7540
rect 20352 7497 20361 7531
rect 20361 7497 20395 7531
rect 20395 7497 20404 7531
rect 20352 7488 20404 7497
rect 26976 7531 27028 7540
rect 26976 7497 26985 7531
rect 26985 7497 27019 7531
rect 27019 7497 27028 7531
rect 26976 7488 27028 7497
rect 4068 7420 4120 7472
rect 6828 7420 6880 7472
rect 17776 7420 17828 7472
rect 19800 7420 19852 7472
rect 2044 7352 2096 7404
rect 7748 7352 7800 7404
rect 8208 7352 8260 7404
rect 18696 7352 18748 7404
rect 19156 7352 19208 7404
rect 19708 7352 19760 7404
rect 3516 7284 3568 7336
rect 5356 7284 5408 7336
rect 16396 7284 16448 7336
rect 16856 7327 16908 7336
rect 16856 7293 16865 7327
rect 16865 7293 16899 7327
rect 16899 7293 16908 7327
rect 16856 7284 16908 7293
rect 17868 7284 17920 7336
rect 19432 7284 19484 7336
rect 27436 7420 27488 7472
rect 27068 7284 27120 7336
rect 2044 7259 2096 7268
rect 2044 7225 2053 7259
rect 2053 7225 2087 7259
rect 2087 7225 2096 7259
rect 2044 7216 2096 7225
rect 19616 7216 19668 7268
rect 1676 7148 1728 7200
rect 2688 7191 2740 7200
rect 2688 7157 2697 7191
rect 2697 7157 2731 7191
rect 2731 7157 2740 7191
rect 2688 7148 2740 7157
rect 6920 7148 6972 7200
rect 7840 7148 7892 7200
rect 16396 7191 16448 7200
rect 16396 7157 16405 7191
rect 16405 7157 16439 7191
rect 16439 7157 16448 7191
rect 16396 7148 16448 7157
rect 26332 7148 26384 7200
rect 27712 7191 27764 7200
rect 27712 7157 27721 7191
rect 27721 7157 27755 7191
rect 27755 7157 27764 7191
rect 27712 7148 27764 7157
rect 10982 7046 11034 7098
rect 11046 7046 11098 7098
rect 11110 7046 11162 7098
rect 11174 7046 11226 7098
rect 20982 7046 21034 7098
rect 21046 7046 21098 7098
rect 21110 7046 21162 7098
rect 21174 7046 21226 7098
rect 4712 6944 4764 6996
rect 6368 6987 6420 6996
rect 6368 6953 6377 6987
rect 6377 6953 6411 6987
rect 6411 6953 6420 6987
rect 6368 6944 6420 6953
rect 17040 6944 17092 6996
rect 19432 6987 19484 6996
rect 19432 6953 19441 6987
rect 19441 6953 19475 6987
rect 19475 6953 19484 6987
rect 19432 6944 19484 6953
rect 19708 6987 19760 6996
rect 19708 6953 19717 6987
rect 19717 6953 19751 6987
rect 19751 6953 19760 6987
rect 19708 6944 19760 6953
rect 572 6876 624 6928
rect 8668 6876 8720 6928
rect 2044 6808 2096 6860
rect 2136 6808 2188 6860
rect 1952 6783 2004 6792
rect 1952 6749 1961 6783
rect 1961 6749 1995 6783
rect 1995 6749 2004 6783
rect 1952 6740 2004 6749
rect 3056 6851 3108 6860
rect 3056 6817 3065 6851
rect 3065 6817 3099 6851
rect 3099 6817 3108 6851
rect 3056 6808 3108 6817
rect 3516 6851 3568 6860
rect 3516 6817 3525 6851
rect 3525 6817 3559 6851
rect 3559 6817 3568 6851
rect 3516 6808 3568 6817
rect 15476 6808 15528 6860
rect 16396 6808 16448 6860
rect 16856 6876 16908 6928
rect 26516 6851 26568 6860
rect 26516 6817 26525 6851
rect 26525 6817 26559 6851
rect 26559 6817 26568 6851
rect 26516 6808 26568 6817
rect 1400 6672 1452 6724
rect 2412 6672 2464 6724
rect 2504 6672 2556 6724
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 6920 6647 6972 6656
rect 6920 6613 6929 6647
rect 6929 6613 6963 6647
rect 6963 6613 6972 6647
rect 6920 6604 6972 6613
rect 15568 6647 15620 6656
rect 15568 6613 15577 6647
rect 15577 6613 15611 6647
rect 15611 6613 15620 6647
rect 15568 6604 15620 6613
rect 26700 6647 26752 6656
rect 26700 6613 26709 6647
rect 26709 6613 26743 6647
rect 26743 6613 26752 6647
rect 26700 6604 26752 6613
rect 5982 6502 6034 6554
rect 6046 6502 6098 6554
rect 6110 6502 6162 6554
rect 6174 6502 6226 6554
rect 15982 6502 16034 6554
rect 16046 6502 16098 6554
rect 16110 6502 16162 6554
rect 16174 6502 16226 6554
rect 25982 6502 26034 6554
rect 26046 6502 26098 6554
rect 26110 6502 26162 6554
rect 26174 6502 26226 6554
rect 1492 6400 1544 6452
rect 2412 6400 2464 6452
rect 15476 6443 15528 6452
rect 15476 6409 15485 6443
rect 15485 6409 15519 6443
rect 15519 6409 15528 6443
rect 15476 6400 15528 6409
rect 26516 6443 26568 6452
rect 26516 6409 26525 6443
rect 26525 6409 26559 6443
rect 26559 6409 26568 6443
rect 26516 6400 26568 6409
rect 2044 6375 2096 6384
rect 2044 6341 2053 6375
rect 2053 6341 2087 6375
rect 2087 6341 2096 6375
rect 2044 6332 2096 6341
rect 4528 6332 4580 6384
rect 2412 6307 2464 6316
rect 2412 6273 2421 6307
rect 2421 6273 2455 6307
rect 2455 6273 2464 6307
rect 2412 6264 2464 6273
rect 2596 6196 2648 6248
rect 2688 6103 2740 6112
rect 2688 6069 2697 6103
rect 2697 6069 2731 6103
rect 2731 6069 2740 6103
rect 2688 6060 2740 6069
rect 10982 5958 11034 6010
rect 11046 5958 11098 6010
rect 11110 5958 11162 6010
rect 11174 5958 11226 6010
rect 20982 5958 21034 6010
rect 21046 5958 21098 6010
rect 21110 5958 21162 6010
rect 21174 5958 21226 6010
rect 2320 5856 2372 5908
rect 2596 5899 2648 5908
rect 2596 5865 2605 5899
rect 2605 5865 2639 5899
rect 2639 5865 2648 5899
rect 2596 5856 2648 5865
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 1492 5516 1544 5568
rect 5982 5414 6034 5466
rect 6046 5414 6098 5466
rect 6110 5414 6162 5466
rect 6174 5414 6226 5466
rect 15982 5414 16034 5466
rect 16046 5414 16098 5466
rect 16110 5414 16162 5466
rect 16174 5414 16226 5466
rect 25982 5414 26034 5466
rect 26046 5414 26098 5466
rect 26110 5414 26162 5466
rect 26174 5414 26226 5466
rect 1400 5312 1452 5364
rect 26424 5151 26476 5160
rect 26424 5117 26433 5151
rect 26433 5117 26467 5151
rect 26467 5117 26476 5151
rect 26424 5108 26476 5117
rect 26608 5015 26660 5024
rect 26608 4981 26617 5015
rect 26617 4981 26651 5015
rect 26651 4981 26660 5015
rect 26608 4972 26660 4981
rect 10982 4870 11034 4922
rect 11046 4870 11098 4922
rect 11110 4870 11162 4922
rect 11174 4870 11226 4922
rect 20982 4870 21034 4922
rect 21046 4870 21098 4922
rect 21110 4870 21162 4922
rect 21174 4870 21226 4922
rect 5982 4326 6034 4378
rect 6046 4326 6098 4378
rect 6110 4326 6162 4378
rect 6174 4326 6226 4378
rect 15982 4326 16034 4378
rect 16046 4326 16098 4378
rect 16110 4326 16162 4378
rect 16174 4326 16226 4378
rect 25982 4326 26034 4378
rect 26046 4326 26098 4378
rect 26110 4326 26162 4378
rect 26174 4326 26226 4378
rect 10982 3782 11034 3834
rect 11046 3782 11098 3834
rect 11110 3782 11162 3834
rect 11174 3782 11226 3834
rect 20982 3782 21034 3834
rect 21046 3782 21098 3834
rect 21110 3782 21162 3834
rect 21174 3782 21226 3834
rect 5982 3238 6034 3290
rect 6046 3238 6098 3290
rect 6110 3238 6162 3290
rect 6174 3238 6226 3290
rect 15982 3238 16034 3290
rect 16046 3238 16098 3290
rect 16110 3238 16162 3290
rect 16174 3238 16226 3290
rect 25982 3238 26034 3290
rect 26046 3238 26098 3290
rect 26110 3238 26162 3290
rect 26174 3238 26226 3290
rect 2044 3179 2096 3188
rect 2044 3145 2053 3179
rect 2053 3145 2087 3179
rect 2087 3145 2096 3179
rect 2044 3136 2096 3145
rect 2044 2932 2096 2984
rect 26424 2975 26476 2984
rect 26424 2941 26433 2975
rect 26433 2941 26467 2975
rect 26467 2941 26476 2975
rect 26424 2932 26476 2941
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 26608 2839 26660 2848
rect 26608 2805 26617 2839
rect 26617 2805 26651 2839
rect 26651 2805 26660 2839
rect 26608 2796 26660 2805
rect 10982 2694 11034 2746
rect 11046 2694 11098 2746
rect 11110 2694 11162 2746
rect 11174 2694 11226 2746
rect 20982 2694 21034 2746
rect 21046 2694 21098 2746
rect 21110 2694 21162 2746
rect 21174 2694 21226 2746
rect 6552 2592 6604 2644
rect 8300 2592 8352 2644
rect 7472 2499 7524 2508
rect 7472 2465 7506 2499
rect 7506 2465 7524 2499
rect 7472 2456 7524 2465
rect 6552 2388 6604 2440
rect 5982 2150 6034 2202
rect 6046 2150 6098 2202
rect 6110 2150 6162 2202
rect 6174 2150 6226 2202
rect 15982 2150 16034 2202
rect 16046 2150 16098 2202
rect 16110 2150 16162 2202
rect 16174 2150 16226 2202
rect 25982 2150 26034 2202
rect 26046 2150 26098 2202
rect 26110 2150 26162 2202
rect 26174 2150 26226 2202
rect 24860 1980 24912 2032
rect 26148 1980 26200 2032
<< metal2 >>
rect 938 23520 994 24000
rect 2778 23520 2834 24000
rect 3514 23624 3570 23633
rect 3514 23559 3570 23568
rect 952 20602 980 23520
rect 2792 20618 2820 23520
rect 3422 23080 3478 23089
rect 3422 23015 3478 23024
rect 3436 22574 3464 23015
rect 3528 22846 3556 23559
rect 4618 23520 4674 24000
rect 6550 23520 6606 24000
rect 8390 23520 8446 24000
rect 10230 23520 10286 24000
rect 12162 23520 12218 24000
rect 14002 23520 14058 24000
rect 15934 23520 15990 24000
rect 17774 23520 17830 24000
rect 19614 23520 19670 24000
rect 21546 23520 21602 24000
rect 23386 23520 23442 24000
rect 25042 23624 25098 23633
rect 25042 23559 25098 23568
rect 3516 22840 3568 22846
rect 3516 22782 3568 22788
rect 3424 22568 3476 22574
rect 3424 22510 3476 22516
rect 3238 22400 3294 22409
rect 3238 22335 3294 22344
rect 2700 20602 2820 20618
rect 940 20596 992 20602
rect 940 20538 992 20544
rect 2688 20596 2820 20602
rect 2740 20590 2820 20596
rect 2962 20632 3018 20641
rect 2962 20567 3018 20576
rect 2688 20538 2740 20544
rect 2044 20392 2096 20398
rect 1964 20340 2044 20346
rect 1964 20334 2096 20340
rect 1964 20318 2084 20334
rect 1860 18624 1912 18630
rect 1860 18566 1912 18572
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1492 17128 1544 17134
rect 1492 17070 1544 17076
rect 1504 16046 1532 17070
rect 1492 16040 1544 16046
rect 1492 15982 1544 15988
rect 1504 15570 1532 15982
rect 1584 15972 1636 15978
rect 1584 15914 1636 15920
rect 1492 15564 1544 15570
rect 1492 15506 1544 15512
rect 1504 14278 1532 15506
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1504 13394 1532 14214
rect 1596 13433 1624 15914
rect 1688 14521 1716 18022
rect 1872 17678 1900 18566
rect 1860 17672 1912 17678
rect 1860 17614 1912 17620
rect 1872 16998 1900 17614
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1964 16810 1992 20318
rect 2320 20256 2372 20262
rect 2320 20198 2372 20204
rect 2228 18828 2280 18834
rect 2228 18770 2280 18776
rect 2240 17882 2268 18770
rect 2228 17876 2280 17882
rect 2228 17818 2280 17824
rect 2136 17740 2188 17746
rect 2136 17682 2188 17688
rect 1872 16782 1992 16810
rect 2148 16794 2176 17682
rect 2136 16788 2188 16794
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1780 15745 1808 15846
rect 1766 15736 1822 15745
rect 1766 15671 1822 15680
rect 1674 14512 1730 14521
rect 1674 14447 1730 14456
rect 1676 14340 1728 14346
rect 1676 14282 1728 14288
rect 1688 13870 1716 14282
rect 1872 14090 1900 16782
rect 2136 16730 2188 16736
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 2056 15473 2084 16594
rect 2136 16584 2188 16590
rect 2240 16572 2268 16730
rect 2188 16544 2268 16572
rect 2136 16526 2188 16532
rect 2042 15464 2098 15473
rect 2042 15399 2098 15408
rect 2056 15162 2084 15399
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 1952 14952 2004 14958
rect 1952 14894 2004 14900
rect 1780 14062 1900 14090
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1582 13424 1638 13433
rect 1492 13388 1544 13394
rect 1582 13359 1638 13368
rect 1492 13330 1544 13336
rect 572 12980 624 12986
rect 572 12922 624 12928
rect 584 12889 612 12922
rect 570 12880 626 12889
rect 1504 12850 1532 13330
rect 570 12815 626 12824
rect 1492 12844 1544 12850
rect 1492 12786 1544 12792
rect 1676 12232 1728 12238
rect 1490 12200 1546 12209
rect 1676 12174 1728 12180
rect 1490 12135 1546 12144
rect 1400 11280 1452 11286
rect 1400 11222 1452 11228
rect 1412 10606 1440 11222
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1504 9704 1532 12135
rect 1412 9676 1532 9704
rect 572 6928 624 6934
rect 572 6870 624 6876
rect 584 3369 612 6870
rect 1412 6730 1440 9676
rect 1688 9450 1716 12174
rect 1492 9444 1544 9450
rect 1492 9386 1544 9392
rect 1676 9444 1728 9450
rect 1676 9386 1728 9392
rect 1504 9110 1532 9386
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1492 9104 1544 9110
rect 1492 9046 1544 9052
rect 1504 8634 1532 9046
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 1596 8498 1624 9318
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1688 8090 1716 8366
rect 1780 8090 1808 14062
rect 1860 14000 1912 14006
rect 1860 13942 1912 13948
rect 1964 13954 1992 14894
rect 2148 14618 2176 16526
rect 2332 16402 2360 20198
rect 2410 19544 2466 19553
rect 2410 19479 2466 19488
rect 2424 18970 2452 19479
rect 2412 18964 2464 18970
rect 2412 18906 2464 18912
rect 2504 18080 2556 18086
rect 2504 18022 2556 18028
rect 2688 18080 2740 18086
rect 2688 18022 2740 18028
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 2424 16522 2452 17070
rect 2412 16516 2464 16522
rect 2412 16458 2464 16464
rect 2240 16374 2360 16402
rect 2136 14612 2188 14618
rect 2136 14554 2188 14560
rect 2240 14498 2268 16374
rect 2516 15910 2544 18022
rect 2700 17746 2728 18022
rect 2688 17740 2740 17746
rect 2688 17682 2740 17688
rect 2780 17536 2832 17542
rect 2780 17478 2832 17484
rect 2792 17134 2820 17478
rect 2780 17128 2832 17134
rect 2780 17070 2832 17076
rect 2780 16992 2832 16998
rect 2780 16934 2832 16940
rect 2688 16448 2740 16454
rect 2688 16390 2740 16396
rect 2700 16114 2728 16390
rect 2688 16108 2740 16114
rect 2688 16050 2740 16056
rect 2504 15904 2556 15910
rect 2504 15846 2556 15852
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 2148 14470 2268 14498
rect 2056 14074 2084 14418
rect 2044 14068 2096 14074
rect 2044 14010 2096 14016
rect 1872 10690 1900 13942
rect 1964 13926 2084 13954
rect 2056 12209 2084 13926
rect 2042 12200 2098 12209
rect 2042 12135 2098 12144
rect 1872 10662 2084 10690
rect 1950 10568 2006 10577
rect 1950 10503 2006 10512
rect 1860 10464 1912 10470
rect 1860 10406 1912 10412
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1490 7440 1546 7449
rect 1490 7375 1546 7384
rect 1400 6724 1452 6730
rect 1400 6666 1452 6672
rect 1504 6458 1532 7375
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1492 6452 1544 6458
rect 1492 6394 1544 6400
rect 1596 6361 1624 6598
rect 1582 6352 1638 6361
rect 1582 6287 1638 6296
rect 1398 5808 1454 5817
rect 1398 5743 1400 5752
rect 1452 5743 1454 5752
rect 1400 5714 1452 5720
rect 1412 5370 1440 5714
rect 1688 5681 1716 7142
rect 1674 5672 1730 5681
rect 1674 5607 1730 5616
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 570 3360 626 3369
rect 570 3295 626 3304
rect 1504 1465 1532 5510
rect 1872 4457 1900 10406
rect 1964 10266 1992 10503
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 1964 9602 1992 10202
rect 2056 9704 2084 10662
rect 2148 9994 2176 14470
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2424 14074 2452 14350
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2516 13530 2544 15846
rect 2700 15586 2728 16050
rect 2792 15706 2820 16934
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2884 16250 2912 16526
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2608 15570 2728 15586
rect 2596 15564 2728 15570
rect 2648 15558 2728 15564
rect 2596 15506 2648 15512
rect 2608 15026 2636 15506
rect 2884 15450 2912 16186
rect 2700 15422 2912 15450
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2700 14958 2728 15422
rect 2688 14952 2740 14958
rect 2976 14906 3004 20567
rect 3054 17776 3110 17785
rect 3054 17711 3110 17720
rect 2688 14894 2740 14900
rect 2792 14878 3004 14906
rect 2792 14618 2820 14878
rect 2964 14816 3016 14822
rect 2964 14758 3016 14764
rect 2976 14618 3004 14758
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 2686 14376 2742 14385
rect 2686 14311 2688 14320
rect 2740 14311 2742 14320
rect 2688 14282 2740 14288
rect 2596 14272 2648 14278
rect 2596 14214 2648 14220
rect 2608 13938 2636 14214
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2240 12442 2268 12718
rect 2332 12646 2360 13330
rect 2792 13025 2820 14554
rect 2976 14278 3004 14554
rect 2964 14272 3016 14278
rect 2964 14214 3016 14220
rect 2872 13796 2924 13802
rect 2872 13738 2924 13744
rect 2884 13258 2912 13738
rect 2872 13252 2924 13258
rect 2872 13194 2924 13200
rect 3068 13138 3096 17711
rect 3148 17672 3200 17678
rect 3148 17614 3200 17620
rect 3160 17338 3188 17614
rect 3148 17332 3200 17338
rect 3148 17274 3200 17280
rect 3160 16726 3188 17274
rect 3148 16720 3200 16726
rect 3148 16662 3200 16668
rect 3146 16008 3202 16017
rect 3146 15943 3202 15952
rect 2884 13110 3096 13138
rect 2778 13016 2834 13025
rect 2778 12951 2834 12960
rect 2320 12640 2372 12646
rect 2320 12582 2372 12588
rect 2504 12640 2556 12646
rect 2884 12594 2912 13110
rect 3056 12912 3108 12918
rect 2962 12880 3018 12889
rect 3056 12854 3108 12860
rect 2962 12815 3018 12824
rect 2504 12582 2556 12588
rect 2228 12436 2280 12442
rect 2228 12378 2280 12384
rect 2240 11694 2268 12378
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2228 11688 2280 11694
rect 2424 11665 2452 12038
rect 2516 11898 2544 12582
rect 2608 12566 2912 12594
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2228 11630 2280 11636
rect 2410 11656 2466 11665
rect 2410 11591 2466 11600
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2240 11014 2268 11494
rect 2228 11008 2280 11014
rect 2228 10950 2280 10956
rect 2320 11008 2372 11014
rect 2320 10950 2372 10956
rect 2240 10606 2268 10950
rect 2228 10600 2280 10606
rect 2228 10542 2280 10548
rect 2332 10538 2360 10950
rect 2320 10532 2372 10538
rect 2320 10474 2372 10480
rect 2332 10266 2360 10474
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2136 9988 2188 9994
rect 2136 9930 2188 9936
rect 2424 9722 2452 10202
rect 2412 9716 2464 9722
rect 2056 9676 2360 9704
rect 1964 9586 2084 9602
rect 1952 9580 2084 9586
rect 2004 9574 2084 9580
rect 1952 9522 2004 9528
rect 1950 9480 2006 9489
rect 1950 9415 1952 9424
rect 2004 9415 2006 9424
rect 1952 9386 2004 9392
rect 1964 9178 1992 9386
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1964 6798 1992 8434
rect 2056 7410 2084 9574
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2240 8974 2268 9522
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2136 8832 2188 8838
rect 2136 8774 2188 8780
rect 2148 8362 2176 8774
rect 2332 8650 2360 9676
rect 2412 9658 2464 9664
rect 2516 8786 2544 11834
rect 2608 11286 2636 12566
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 2884 11354 2912 12242
rect 2976 11801 3004 12815
rect 2962 11792 3018 11801
rect 2962 11727 3018 11736
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2596 11280 2648 11286
rect 2780 11280 2832 11286
rect 2596 11222 2648 11228
rect 2686 11248 2742 11257
rect 2780 11222 2832 11228
rect 2686 11183 2742 11192
rect 2700 10810 2728 11183
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2792 9738 2820 11222
rect 2872 11144 2924 11150
rect 3068 11132 3096 12854
rect 2924 11104 3096 11132
rect 2872 11086 2924 11092
rect 2884 10742 2912 11086
rect 2872 10736 2924 10742
rect 2872 10678 2924 10684
rect 3160 10606 3188 15943
rect 3252 10713 3280 22335
rect 3790 21856 3846 21865
rect 3790 21791 3846 21800
rect 3804 21690 3832 21791
rect 3792 21684 3844 21690
rect 3792 21626 3844 21632
rect 4066 21312 4122 21321
rect 4066 21247 4122 21256
rect 4080 20874 4108 21247
rect 4068 20868 4120 20874
rect 4068 20810 4120 20816
rect 4160 20256 4212 20262
rect 3988 20216 4160 20244
rect 3884 19712 3936 19718
rect 3884 19654 3936 19660
rect 3700 19372 3752 19378
rect 3700 19314 3752 19320
rect 3712 19281 3740 19314
rect 3698 19272 3754 19281
rect 3698 19207 3754 19216
rect 3896 19174 3924 19654
rect 3884 19168 3936 19174
rect 3882 19136 3884 19145
rect 3936 19136 3938 19145
rect 3882 19071 3938 19080
rect 3790 18864 3846 18873
rect 3790 18799 3846 18808
rect 3514 18320 3570 18329
rect 3514 18255 3570 18264
rect 3698 18320 3754 18329
rect 3698 18255 3754 18264
rect 3330 17912 3386 17921
rect 3330 17847 3386 17856
rect 3344 11286 3372 17847
rect 3424 16720 3476 16726
rect 3528 16697 3556 18255
rect 3712 18222 3740 18255
rect 3700 18216 3752 18222
rect 3700 18158 3752 18164
rect 3608 18080 3660 18086
rect 3608 18022 3660 18028
rect 3424 16662 3476 16668
rect 3514 16688 3570 16697
rect 3436 16046 3464 16662
rect 3514 16623 3570 16632
rect 3424 16040 3476 16046
rect 3424 15982 3476 15988
rect 3516 15088 3568 15094
rect 3514 15056 3516 15065
rect 3568 15056 3570 15065
rect 3514 14991 3570 15000
rect 3620 15008 3648 18022
rect 3712 17882 3740 18158
rect 3700 17876 3752 17882
rect 3700 17818 3752 17824
rect 3700 16992 3752 16998
rect 3700 16934 3752 16940
rect 3712 16794 3740 16934
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 3700 16448 3752 16454
rect 3700 16390 3752 16396
rect 3712 15502 3740 16390
rect 3804 16017 3832 18799
rect 3884 18624 3936 18630
rect 3884 18566 3936 18572
rect 3896 18290 3924 18566
rect 3988 18426 4016 20216
rect 4160 20198 4212 20204
rect 4434 20088 4490 20097
rect 4434 20023 4436 20032
rect 4488 20023 4490 20032
rect 4436 19994 4488 20000
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 4080 19242 4108 19858
rect 4632 19553 4660 23520
rect 5956 21788 6252 21808
rect 6012 21786 6036 21788
rect 6092 21786 6116 21788
rect 6172 21786 6196 21788
rect 6034 21734 6036 21786
rect 6098 21734 6110 21786
rect 6172 21734 6174 21786
rect 6012 21732 6036 21734
rect 6092 21732 6116 21734
rect 6172 21732 6196 21734
rect 5956 21712 6252 21732
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 4618 19544 4674 19553
rect 4618 19479 4674 19488
rect 4068 19236 4120 19242
rect 4068 19178 4120 19184
rect 4080 18970 4108 19178
rect 4436 19168 4488 19174
rect 4436 19110 4488 19116
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 3884 18284 3936 18290
rect 3884 18226 3936 18232
rect 4160 18284 4212 18290
rect 4160 18226 4212 18232
rect 4344 18284 4396 18290
rect 4344 18226 4396 18232
rect 4172 17814 4200 18226
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 4264 17921 4292 18022
rect 4250 17912 4306 17921
rect 4356 17882 4384 18226
rect 4250 17847 4306 17856
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4160 17808 4212 17814
rect 4160 17750 4212 17756
rect 4356 17134 4384 17818
rect 4448 17785 4476 19110
rect 4434 17776 4490 17785
rect 4434 17711 4490 17720
rect 4344 17128 4396 17134
rect 4344 17070 4396 17076
rect 4158 16824 4214 16833
rect 4158 16759 4214 16768
rect 3790 16008 3846 16017
rect 3846 15966 3924 15994
rect 3790 15943 3846 15952
rect 3790 15872 3846 15881
rect 3790 15807 3846 15816
rect 3700 15496 3752 15502
rect 3700 15438 3752 15444
rect 3620 14980 3740 15008
rect 3606 14512 3662 14521
rect 3606 14447 3662 14456
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 3436 12458 3464 12582
rect 3427 12430 3464 12458
rect 3427 12322 3455 12430
rect 3427 12294 3464 12322
rect 3436 11558 3464 12294
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3332 11280 3384 11286
rect 3332 11222 3384 11228
rect 3344 10810 3372 11222
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3238 10704 3294 10713
rect 3238 10639 3294 10648
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 3160 10305 3188 10406
rect 3146 10296 3202 10305
rect 3146 10231 3202 10240
rect 2872 10192 2924 10198
rect 2872 10134 2924 10140
rect 2240 8622 2360 8650
rect 2424 8758 2544 8786
rect 2608 9710 2820 9738
rect 2136 8356 2188 8362
rect 2136 8298 2188 8304
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 2042 7304 2098 7313
rect 2042 7239 2044 7248
rect 2096 7239 2098 7248
rect 2044 7210 2096 7216
rect 2148 6866 2176 8298
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 2056 6390 2084 6802
rect 2044 6384 2096 6390
rect 2044 6326 2096 6332
rect 2240 5137 2268 8622
rect 2320 8288 2372 8294
rect 2320 8230 2372 8236
rect 2332 7954 2360 8230
rect 2424 8022 2452 8758
rect 2502 8664 2558 8673
rect 2502 8599 2558 8608
rect 2412 8016 2464 8022
rect 2412 7958 2464 7964
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2332 5914 2360 7890
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2424 7041 2452 7822
rect 2410 7032 2466 7041
rect 2410 6967 2466 6976
rect 2516 6730 2544 8599
rect 2412 6724 2464 6730
rect 2412 6666 2464 6672
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 2424 6458 2452 6666
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2410 6352 2466 6361
rect 2410 6287 2412 6296
rect 2464 6287 2466 6296
rect 2412 6258 2464 6264
rect 2608 6254 2636 9710
rect 2780 9104 2832 9110
rect 2780 9046 2832 9052
rect 2792 8566 2820 9046
rect 2780 8560 2832 8566
rect 2780 8502 2832 8508
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2700 8022 2728 8434
rect 2778 8392 2834 8401
rect 2778 8327 2834 8336
rect 2688 8016 2740 8022
rect 2688 7958 2740 7964
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2700 7546 2728 7822
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 2700 6905 2728 7142
rect 2686 6896 2742 6905
rect 2686 6831 2742 6840
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2608 5914 2636 6190
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2596 5908 2648 5914
rect 2596 5850 2648 5856
rect 2226 5128 2282 5137
rect 2226 5063 2282 5072
rect 1858 4448 1914 4457
rect 1858 4383 1914 4392
rect 2042 4040 2098 4049
rect 2042 3975 2098 3984
rect 2056 3194 2084 3975
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2056 2990 2084 3130
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1596 2689 1624 2790
rect 1582 2680 1638 2689
rect 1582 2615 1638 2624
rect 1490 1456 1546 1465
rect 1490 1391 1546 1400
rect 2700 921 2728 6054
rect 2792 2145 2820 8327
rect 2884 8090 2912 10134
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2976 8974 3004 9522
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2976 8430 3004 8910
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 3068 6866 3096 10066
rect 3146 10024 3202 10033
rect 3146 9959 3148 9968
rect 3200 9959 3202 9968
rect 3148 9930 3200 9936
rect 3160 8022 3188 9930
rect 3252 9489 3280 10639
rect 3436 9625 3464 11494
rect 3528 11354 3556 12174
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3528 10674 3556 11290
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3528 10266 3556 10610
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3528 9722 3556 10202
rect 3516 9716 3568 9722
rect 3516 9658 3568 9664
rect 3422 9616 3478 9625
rect 3344 9574 3422 9602
rect 3238 9480 3294 9489
rect 3238 9415 3294 9424
rect 3148 8016 3200 8022
rect 3148 7958 3200 7964
rect 3344 7886 3372 9574
rect 3422 9551 3478 9560
rect 3424 9444 3476 9450
rect 3424 9386 3476 9392
rect 3436 9178 3464 9386
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3528 7546 3556 8434
rect 3620 8129 3648 14447
rect 3712 13977 3740 14980
rect 3804 14822 3832 15807
rect 3896 15609 3924 15966
rect 3882 15600 3938 15609
rect 3882 15535 3938 15544
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 4066 15328 4122 15337
rect 3896 15026 3924 15302
rect 4066 15263 4122 15272
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3698 13968 3754 13977
rect 3698 13903 3754 13912
rect 3712 12442 3740 13903
rect 3804 13297 3832 14758
rect 3896 14414 3924 14962
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3988 14618 4016 14758
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 3896 13734 3924 14350
rect 3884 13728 3936 13734
rect 4080 13705 4108 15263
rect 3884 13670 3936 13676
rect 4066 13696 4122 13705
rect 3896 13462 3924 13670
rect 4066 13631 4122 13640
rect 3884 13456 3936 13462
rect 3884 13398 3936 13404
rect 3790 13288 3846 13297
rect 3790 13223 3846 13232
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 4080 12345 4108 12786
rect 4066 12336 4122 12345
rect 4172 12306 4200 16759
rect 4356 16250 4384 17070
rect 4528 16448 4580 16454
rect 4528 16390 4580 16396
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 4252 15972 4304 15978
rect 4252 15914 4304 15920
rect 4264 14958 4292 15914
rect 4540 15745 4568 16390
rect 4632 15881 4660 19110
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4816 18714 4844 21626
rect 5632 20868 5684 20874
rect 5632 20810 5684 20816
rect 5080 20800 5132 20806
rect 5080 20742 5132 20748
rect 5092 20466 5120 20742
rect 5080 20460 5132 20466
rect 5080 20402 5132 20408
rect 4896 20392 4948 20398
rect 4896 20334 4948 20340
rect 4908 18902 4936 20334
rect 4988 20256 5040 20262
rect 4988 20198 5040 20204
rect 5000 19378 5028 20198
rect 5092 20058 5120 20402
rect 5644 20058 5672 20810
rect 5956 20700 6252 20720
rect 6012 20698 6036 20700
rect 6092 20698 6116 20700
rect 6172 20698 6196 20700
rect 6034 20646 6036 20698
rect 6098 20646 6110 20698
rect 6172 20646 6174 20698
rect 6012 20644 6036 20646
rect 6092 20644 6116 20646
rect 6172 20644 6196 20646
rect 5956 20624 6252 20644
rect 6564 20097 6592 23520
rect 8404 23474 8432 23520
rect 8312 23446 8432 23474
rect 7472 22568 7524 22574
rect 7472 22510 7524 22516
rect 7380 20256 7432 20262
rect 7378 20224 7380 20233
rect 7432 20224 7434 20233
rect 7378 20159 7434 20168
rect 6550 20088 6606 20097
rect 5080 20052 5132 20058
rect 5080 19994 5132 20000
rect 5632 20052 5684 20058
rect 6550 20023 6606 20032
rect 5632 19994 5684 20000
rect 5356 19712 5408 19718
rect 5356 19654 5408 19660
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5080 19508 5132 19514
rect 5080 19450 5132 19456
rect 4988 19372 5040 19378
rect 4988 19314 5040 19320
rect 5092 19009 5120 19450
rect 5368 19378 5396 19654
rect 5356 19372 5408 19378
rect 5356 19314 5408 19320
rect 5078 19000 5134 19009
rect 5078 18935 5134 18944
rect 4896 18896 4948 18902
rect 4896 18838 4948 18844
rect 4724 17882 4752 18702
rect 4816 18686 4936 18714
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 4724 17746 4752 17818
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 4724 17066 4752 17682
rect 4712 17060 4764 17066
rect 4712 17002 4764 17008
rect 4724 16794 4752 17002
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4618 15872 4674 15881
rect 4618 15807 4674 15816
rect 4526 15736 4582 15745
rect 4526 15671 4528 15680
rect 4580 15671 4582 15680
rect 4528 15642 4580 15648
rect 4632 15586 4660 15807
rect 4436 15564 4488 15570
rect 4436 15506 4488 15512
rect 4540 15558 4660 15586
rect 4448 15065 4476 15506
rect 4434 15056 4490 15065
rect 4434 14991 4490 15000
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4066 12271 4122 12280
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3896 11801 3924 12038
rect 4172 11898 4200 12242
rect 4264 12186 4292 14214
rect 4540 14113 4568 15558
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4632 14618 4660 15438
rect 4710 14920 4766 14929
rect 4710 14855 4766 14864
rect 4620 14612 4672 14618
rect 4620 14554 4672 14560
rect 4724 14482 4752 14855
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4816 14618 4844 14758
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4526 14104 4582 14113
rect 4724 14074 4752 14418
rect 4526 14039 4582 14048
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4540 13530 4568 13670
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4540 12850 4568 13466
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4632 12986 4660 13330
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4816 12986 4844 13262
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4264 12158 4384 12186
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 3882 11792 3938 11801
rect 3882 11727 3938 11736
rect 4068 11212 4120 11218
rect 4120 11172 4200 11200
rect 4068 11154 4120 11160
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 4080 10441 4108 11018
rect 4172 10810 4200 11172
rect 4264 11121 4292 12038
rect 4250 11112 4306 11121
rect 4250 11047 4306 11056
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4066 10432 4122 10441
rect 4066 10367 4122 10376
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 3976 10124 4028 10130
rect 3976 10066 4028 10072
rect 3988 9994 4016 10066
rect 3976 9988 4028 9994
rect 3976 9930 4028 9936
rect 3884 9920 3936 9926
rect 3790 9888 3846 9897
rect 3884 9862 3936 9868
rect 3790 9823 3846 9832
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3606 8120 3662 8129
rect 3712 8090 3740 8230
rect 3606 8055 3662 8064
rect 3700 8084 3752 8090
rect 3700 8026 3752 8032
rect 3804 7546 3832 9823
rect 3896 8090 3924 9862
rect 4080 8634 4108 10202
rect 4172 9110 4200 10746
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4264 10470 4292 10542
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4250 9480 4306 9489
rect 4250 9415 4306 9424
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4264 8498 4292 9415
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3528 7342 3556 7482
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3514 7032 3570 7041
rect 3514 6967 3570 6976
rect 3528 6866 3556 6967
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 3516 6860 3568 6866
rect 3516 6802 3568 6808
rect 3698 3496 3754 3505
rect 3698 3431 3754 3440
rect 2778 2136 2834 2145
rect 2778 2071 2834 2080
rect 2686 912 2742 921
rect 2686 847 2742 856
rect 3712 480 3740 3431
rect 3698 0 3754 480
rect 4080 377 4108 7414
rect 4356 3913 4384 12158
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4436 11008 4488 11014
rect 4436 10950 4488 10956
rect 4448 10266 4476 10950
rect 4528 10600 4580 10606
rect 4528 10542 4580 10548
rect 4436 10260 4488 10266
rect 4436 10202 4488 10208
rect 4540 10198 4568 10542
rect 4632 10305 4660 12038
rect 4804 11620 4856 11626
rect 4804 11562 4856 11568
rect 4816 11014 4844 11562
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4816 10470 4844 10950
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4618 10296 4674 10305
rect 4618 10231 4674 10240
rect 4528 10192 4580 10198
rect 4528 10134 4580 10140
rect 4540 9722 4568 10134
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4724 9178 4752 9998
rect 4816 9518 4844 10406
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4434 9072 4490 9081
rect 4434 9007 4490 9016
rect 4448 8090 4476 9007
rect 4712 8968 4764 8974
rect 4816 8956 4844 9454
rect 4908 9081 4936 18686
rect 5264 18148 5316 18154
rect 5264 18090 5316 18096
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 5000 12918 5028 18022
rect 5276 17649 5304 18090
rect 5368 17814 5396 19314
rect 5448 19304 5500 19310
rect 5552 19292 5580 19654
rect 5644 19514 5672 19994
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 5632 19508 5684 19514
rect 5632 19450 5684 19456
rect 5500 19264 5580 19292
rect 5448 19246 5500 19252
rect 5460 18426 5488 19246
rect 5736 19242 5764 19790
rect 5956 19612 6252 19632
rect 6012 19610 6036 19612
rect 6092 19610 6116 19612
rect 6172 19610 6196 19612
rect 6034 19558 6036 19610
rect 6098 19558 6110 19610
rect 6172 19558 6174 19610
rect 6012 19556 6036 19558
rect 6092 19556 6116 19558
rect 6172 19556 6196 19558
rect 5956 19536 6252 19556
rect 6736 19508 6788 19514
rect 6736 19450 6788 19456
rect 6090 19272 6146 19281
rect 5724 19236 5776 19242
rect 6090 19207 6146 19216
rect 5724 19178 5776 19184
rect 5632 18964 5684 18970
rect 5632 18906 5684 18912
rect 5540 18896 5592 18902
rect 5540 18838 5592 18844
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 5448 18080 5500 18086
rect 5448 18022 5500 18028
rect 5356 17808 5408 17814
rect 5356 17750 5408 17756
rect 5078 17640 5134 17649
rect 5078 17575 5134 17584
rect 5262 17640 5318 17649
rect 5262 17575 5318 17584
rect 5092 16017 5120 17575
rect 5368 17338 5396 17750
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5368 16250 5396 16594
rect 5460 16425 5488 18022
rect 5552 17882 5580 18838
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5644 16726 5672 18906
rect 5632 16720 5684 16726
rect 5632 16662 5684 16668
rect 5446 16416 5502 16425
rect 5446 16351 5502 16360
rect 5644 16250 5672 16662
rect 5356 16244 5408 16250
rect 5632 16244 5684 16250
rect 5408 16204 5488 16232
rect 5356 16186 5408 16192
rect 5460 16046 5488 16204
rect 5632 16186 5684 16192
rect 5736 16153 5764 19178
rect 6104 18970 6132 19207
rect 6092 18964 6144 18970
rect 6092 18906 6144 18912
rect 5956 18524 6252 18544
rect 6012 18522 6036 18524
rect 6092 18522 6116 18524
rect 6172 18522 6196 18524
rect 6034 18470 6036 18522
rect 6098 18470 6110 18522
rect 6172 18470 6174 18522
rect 6012 18468 6036 18470
rect 6092 18468 6116 18470
rect 6172 18468 6196 18470
rect 5956 18448 6252 18468
rect 5956 17436 6252 17456
rect 6012 17434 6036 17436
rect 6092 17434 6116 17436
rect 6172 17434 6196 17436
rect 6034 17382 6036 17434
rect 6098 17382 6110 17434
rect 6172 17382 6174 17434
rect 6012 17380 6036 17382
rect 6092 17380 6116 17382
rect 6172 17380 6196 17382
rect 5956 17360 6252 17380
rect 6642 17368 6698 17377
rect 6642 17303 6644 17312
rect 6696 17303 6698 17312
rect 6644 17274 6696 17280
rect 5814 17096 5870 17105
rect 5814 17031 5870 17040
rect 5722 16144 5778 16153
rect 5722 16079 5778 16088
rect 5448 16040 5500 16046
rect 5078 16008 5134 16017
rect 5448 15982 5500 15988
rect 5078 15943 5134 15952
rect 5354 15736 5410 15745
rect 5354 15671 5410 15680
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5184 13258 5212 14758
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 5172 13252 5224 13258
rect 5172 13194 5224 13200
rect 4988 12912 5040 12918
rect 4988 12854 5040 12860
rect 5184 12782 5212 13194
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5184 12374 5212 12582
rect 5172 12368 5224 12374
rect 5172 12310 5224 12316
rect 5080 12164 5132 12170
rect 5080 12106 5132 12112
rect 5092 11898 5120 12106
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 5276 11626 5304 14010
rect 5264 11620 5316 11626
rect 5264 11562 5316 11568
rect 5172 11552 5224 11558
rect 5170 11520 5172 11529
rect 5224 11520 5226 11529
rect 5170 11455 5226 11464
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 5000 10606 5028 10950
rect 5368 10810 5396 15671
rect 5460 15502 5488 15982
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5460 15162 5488 15438
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5460 15008 5488 15098
rect 5460 14980 5580 15008
rect 5448 14816 5500 14822
rect 5446 14784 5448 14793
rect 5500 14784 5502 14793
rect 5446 14719 5502 14728
rect 5460 11286 5488 14719
rect 5552 14482 5580 14980
rect 5644 14550 5672 15302
rect 5632 14544 5684 14550
rect 5632 14486 5684 14492
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5552 14074 5580 14418
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5552 13326 5580 13806
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5538 13016 5594 13025
rect 5538 12951 5540 12960
rect 5592 12951 5594 12960
rect 5540 12922 5592 12928
rect 5644 12850 5672 14486
rect 5724 13796 5776 13802
rect 5724 13738 5776 13744
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5736 12714 5764 13738
rect 5828 13394 5856 17031
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 5956 16348 6252 16368
rect 6012 16346 6036 16348
rect 6092 16346 6116 16348
rect 6172 16346 6196 16348
rect 6034 16294 6036 16346
rect 6098 16294 6110 16346
rect 6172 16294 6174 16346
rect 6012 16292 6036 16294
rect 6092 16292 6116 16294
rect 6172 16292 6196 16294
rect 5956 16272 6252 16292
rect 6092 15904 6144 15910
rect 6092 15846 6144 15852
rect 6104 15473 6132 15846
rect 6380 15570 6408 16390
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 6090 15464 6146 15473
rect 6090 15399 6146 15408
rect 5956 15260 6252 15280
rect 6012 15258 6036 15260
rect 6092 15258 6116 15260
rect 6172 15258 6196 15260
rect 6034 15206 6036 15258
rect 6098 15206 6110 15258
rect 6172 15206 6174 15258
rect 6012 15204 6036 15206
rect 6092 15204 6116 15206
rect 6172 15204 6196 15206
rect 5956 15184 6252 15204
rect 6380 15026 6408 15506
rect 6368 15020 6420 15026
rect 6368 14962 6420 14968
rect 5908 14884 5960 14890
rect 5908 14826 5960 14832
rect 5920 14618 5948 14826
rect 6380 14822 6408 14962
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 5956 14172 6252 14192
rect 6012 14170 6036 14172
rect 6092 14170 6116 14172
rect 6172 14170 6196 14172
rect 6034 14118 6036 14170
rect 6098 14118 6110 14170
rect 6172 14118 6174 14170
rect 6012 14116 6036 14118
rect 6092 14116 6116 14118
rect 6172 14116 6196 14118
rect 5956 14096 6252 14116
rect 6276 14000 6328 14006
rect 6276 13942 6328 13948
rect 5908 13728 5960 13734
rect 5908 13670 5960 13676
rect 5920 13433 5948 13670
rect 5906 13424 5962 13433
rect 5816 13388 5868 13394
rect 5906 13359 5962 13368
rect 5816 13330 5868 13336
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5828 12889 5856 13126
rect 5956 13084 6252 13104
rect 6012 13082 6036 13084
rect 6092 13082 6116 13084
rect 6172 13082 6196 13084
rect 6034 13030 6036 13082
rect 6098 13030 6110 13082
rect 6172 13030 6174 13082
rect 6012 13028 6036 13030
rect 6092 13028 6116 13030
rect 6172 13028 6196 13030
rect 5956 13008 6252 13028
rect 6184 12912 6236 12918
rect 5814 12880 5870 12889
rect 5814 12815 5870 12824
rect 6182 12880 6184 12889
rect 6236 12880 6238 12889
rect 6182 12815 6238 12824
rect 5724 12708 5776 12714
rect 5724 12650 5776 12656
rect 5816 12436 5868 12442
rect 5816 12378 5868 12384
rect 5724 12368 5776 12374
rect 5724 12310 5776 12316
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5552 11558 5580 12038
rect 5736 11626 5764 12310
rect 5724 11620 5776 11626
rect 5724 11562 5776 11568
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5552 11393 5580 11494
rect 5538 11384 5594 11393
rect 5538 11319 5594 11328
rect 5448 11280 5500 11286
rect 5448 11222 5500 11228
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5736 10674 5764 11154
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 4988 10600 5040 10606
rect 4988 10542 5040 10548
rect 5736 10538 5764 10610
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 5724 10532 5776 10538
rect 5724 10474 5776 10480
rect 5092 10266 5120 10474
rect 5630 10296 5686 10305
rect 5080 10260 5132 10266
rect 5630 10231 5632 10240
rect 5080 10202 5132 10208
rect 5684 10231 5686 10240
rect 5724 10260 5776 10266
rect 5632 10202 5684 10208
rect 5724 10202 5776 10208
rect 5736 9722 5764 10202
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5828 9586 5856 12378
rect 5908 12232 5960 12238
rect 5906 12200 5908 12209
rect 6288 12209 6316 13942
rect 6380 13938 6408 14758
rect 6550 14648 6606 14657
rect 6550 14583 6606 14592
rect 6564 14074 6592 14583
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6380 13530 6408 13874
rect 6564 13870 6592 14010
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6458 13696 6514 13705
rect 6458 13631 6514 13640
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6380 12306 6408 13330
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 5960 12200 5962 12209
rect 5906 12135 5962 12144
rect 6274 12200 6330 12209
rect 6274 12135 6330 12144
rect 5956 11996 6252 12016
rect 6012 11994 6036 11996
rect 6092 11994 6116 11996
rect 6172 11994 6196 11996
rect 6034 11942 6036 11994
rect 6098 11942 6110 11994
rect 6172 11942 6174 11994
rect 6012 11940 6036 11942
rect 6092 11940 6116 11942
rect 6172 11940 6196 11942
rect 5956 11920 6252 11940
rect 6380 11937 6408 12242
rect 6366 11928 6422 11937
rect 6366 11863 6368 11872
rect 6420 11863 6422 11872
rect 6368 11834 6420 11840
rect 6380 11803 6408 11834
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 5956 10908 6252 10928
rect 6012 10906 6036 10908
rect 6092 10906 6116 10908
rect 6172 10906 6196 10908
rect 6034 10854 6036 10906
rect 6098 10854 6110 10906
rect 6172 10854 6174 10906
rect 6012 10852 6036 10854
rect 6092 10852 6116 10854
rect 6172 10852 6196 10854
rect 5956 10832 6252 10852
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 5998 10296 6054 10305
rect 5998 10231 6000 10240
rect 6052 10231 6054 10240
rect 6000 10202 6052 10208
rect 6196 10198 6224 10406
rect 6092 10192 6144 10198
rect 6090 10160 6092 10169
rect 6184 10192 6236 10198
rect 6144 10160 6146 10169
rect 6184 10134 6236 10140
rect 6090 10095 6146 10104
rect 5956 9820 6252 9840
rect 6012 9818 6036 9820
rect 6092 9818 6116 9820
rect 6172 9818 6196 9820
rect 6034 9766 6036 9818
rect 6098 9766 6110 9818
rect 6172 9766 6174 9818
rect 6012 9764 6036 9766
rect 6092 9764 6116 9766
rect 6172 9764 6196 9766
rect 5956 9744 6252 9764
rect 6092 9648 6144 9654
rect 6092 9590 6144 9596
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5816 9376 5868 9382
rect 5814 9344 5816 9353
rect 5868 9344 5870 9353
rect 5814 9279 5870 9288
rect 6104 9178 6132 9590
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 4894 9072 4950 9081
rect 4894 9007 4950 9016
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 4764 8928 4844 8956
rect 4712 8910 4764 8916
rect 4724 8362 4752 8910
rect 5276 8498 5304 8978
rect 5956 8732 6252 8752
rect 6012 8730 6036 8732
rect 6092 8730 6116 8732
rect 6172 8730 6196 8732
rect 6034 8678 6036 8730
rect 6098 8678 6110 8730
rect 6172 8678 6174 8730
rect 6012 8676 6036 8678
rect 6092 8676 6116 8678
rect 6172 8676 6196 8678
rect 5956 8656 6252 8676
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 5276 8294 5304 8434
rect 5552 8401 5580 8502
rect 5538 8392 5594 8401
rect 5538 8327 5594 8336
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4448 7546 4476 8026
rect 4528 8016 4580 8022
rect 4528 7958 4580 7964
rect 4540 7546 4568 7958
rect 5276 7886 5304 8230
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5354 7848 5410 7857
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4540 6390 4568 7482
rect 4724 7002 4752 7822
rect 5354 7783 5410 7792
rect 5368 7546 5396 7783
rect 5956 7644 6252 7664
rect 6012 7642 6036 7644
rect 6092 7642 6116 7644
rect 6172 7642 6196 7644
rect 6034 7590 6036 7642
rect 6098 7590 6110 7642
rect 6172 7590 6174 7642
rect 6012 7588 6036 7590
rect 6092 7588 6116 7590
rect 6172 7588 6196 7590
rect 5956 7568 6252 7588
rect 6288 7546 6316 11222
rect 6366 10160 6422 10169
rect 6472 10146 6500 13631
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6564 12170 6592 12786
rect 6656 12306 6684 14758
rect 6748 14521 6776 19450
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 7194 19136 7250 19145
rect 6840 18329 6868 19110
rect 7194 19071 7250 19080
rect 7208 18970 7236 19071
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 7010 18728 7066 18737
rect 6826 18320 6882 18329
rect 6826 18255 6882 18264
rect 6932 18170 6960 18702
rect 7010 18663 7066 18672
rect 6840 18142 6960 18170
rect 6840 17882 6868 18142
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6734 14512 6790 14521
rect 6734 14447 6790 14456
rect 6736 14340 6788 14346
rect 6736 14282 6788 14288
rect 6748 13802 6776 14282
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 6840 13462 6868 14214
rect 7024 13852 7052 18663
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 7116 18154 7144 18566
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 7104 18148 7156 18154
rect 7104 18090 7156 18096
rect 7116 16289 7144 18090
rect 7196 18080 7248 18086
rect 7196 18022 7248 18028
rect 7102 16280 7158 16289
rect 7102 16215 7158 16224
rect 7208 15609 7236 18022
rect 7300 17814 7328 18226
rect 7288 17808 7340 17814
rect 7484 17785 7512 22510
rect 8208 20596 8260 20602
rect 8312 20584 8340 23446
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 8260 20556 8340 20584
rect 8208 20538 8260 20544
rect 9680 20256 9732 20262
rect 9310 20224 9366 20233
rect 9680 20198 9732 20204
rect 9310 20159 9366 20168
rect 8300 19304 8352 19310
rect 8220 19264 8300 19292
rect 7654 19000 7710 19009
rect 7654 18935 7656 18944
rect 7708 18935 7710 18944
rect 7656 18906 7708 18912
rect 7564 18828 7616 18834
rect 7564 18770 7616 18776
rect 7576 18358 7604 18770
rect 7564 18352 7616 18358
rect 7564 18294 7616 18300
rect 7576 17882 7604 18294
rect 7564 17876 7616 17882
rect 7564 17818 7616 17824
rect 7288 17750 7340 17756
rect 7470 17776 7526 17785
rect 7668 17746 7696 18906
rect 7840 18760 7892 18766
rect 7840 18702 7892 18708
rect 7852 18426 7880 18702
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 7932 18080 7984 18086
rect 7932 18022 7984 18028
rect 7470 17711 7526 17720
rect 7656 17740 7708 17746
rect 7656 17682 7708 17688
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7484 17066 7512 17614
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7194 15600 7250 15609
rect 7194 15535 7250 15544
rect 7286 15056 7342 15065
rect 7286 14991 7288 15000
rect 7340 14991 7342 15000
rect 7288 14962 7340 14968
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 6932 13824 7052 13852
rect 6932 13530 6960 13824
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6828 13456 6880 13462
rect 6828 13398 6880 13404
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6840 12730 6868 13262
rect 6932 12918 6960 13466
rect 7024 13394 7052 13670
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 7024 12986 7052 13330
rect 7116 13190 7144 13670
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 6918 12744 6974 12753
rect 6840 12702 6918 12730
rect 6918 12679 6974 12688
rect 6644 12300 6696 12306
rect 6644 12242 6696 12248
rect 6552 12164 6604 12170
rect 6552 12106 6604 12112
rect 6656 11898 6684 12242
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6826 11792 6882 11801
rect 6826 11727 6882 11736
rect 6840 10810 6868 11727
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6552 10260 6604 10266
rect 6932 10248 6960 12679
rect 7024 12442 7052 12922
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7116 11694 7144 12378
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7208 10690 7236 14894
rect 7484 14346 7512 17002
rect 7944 16833 7972 18022
rect 8220 17882 8248 19264
rect 8300 19246 8352 19252
rect 9034 19272 9090 19281
rect 9034 19207 9090 19216
rect 9048 19174 9076 19207
rect 9036 19168 9088 19174
rect 9036 19110 9088 19116
rect 8576 18624 8628 18630
rect 9036 18624 9088 18630
rect 8576 18566 8628 18572
rect 8942 18592 8998 18601
rect 8588 18086 8616 18566
rect 9036 18566 9088 18572
rect 8942 18527 8998 18536
rect 8956 18154 8984 18527
rect 9048 18290 9076 18566
rect 9036 18284 9088 18290
rect 9036 18226 9088 18232
rect 8944 18148 8996 18154
rect 8944 18090 8996 18096
rect 8484 18080 8536 18086
rect 8484 18022 8536 18028
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8942 18048 8998 18057
rect 8496 17882 8524 18022
rect 8208 17876 8260 17882
rect 8208 17818 8260 17824
rect 8484 17876 8536 17882
rect 8484 17818 8536 17824
rect 8392 17808 8444 17814
rect 8298 17776 8354 17785
rect 8208 17740 8260 17746
rect 8392 17750 8444 17756
rect 8298 17711 8354 17720
rect 8208 17682 8260 17688
rect 8220 17134 8248 17682
rect 8208 17128 8260 17134
rect 8022 17096 8078 17105
rect 8208 17070 8260 17076
rect 8022 17031 8078 17040
rect 7930 16824 7986 16833
rect 7930 16759 7986 16768
rect 7654 16688 7710 16697
rect 7564 16652 7616 16658
rect 8036 16658 8064 17031
rect 8220 16998 8248 17070
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 8220 16810 8248 16934
rect 8128 16782 8248 16810
rect 7654 16623 7710 16632
rect 8024 16652 8076 16658
rect 7564 16594 7616 16600
rect 7576 15162 7604 16594
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7576 14618 7604 15098
rect 7668 15094 7696 16623
rect 8024 16594 8076 16600
rect 8128 16046 8156 16782
rect 8312 16726 8340 17711
rect 8404 17377 8432 17750
rect 8390 17368 8446 17377
rect 8390 17303 8446 17312
rect 8484 16788 8536 16794
rect 8484 16730 8536 16736
rect 8300 16720 8352 16726
rect 8220 16668 8300 16674
rect 8220 16662 8352 16668
rect 8220 16646 8340 16662
rect 8220 16250 8248 16646
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8116 16040 8168 16046
rect 8116 15982 8168 15988
rect 8128 15706 8156 15982
rect 8392 15972 8444 15978
rect 8392 15914 8444 15920
rect 8116 15700 8168 15706
rect 8116 15642 8168 15648
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8312 15094 8340 15642
rect 8404 15638 8432 15914
rect 8392 15632 8444 15638
rect 8392 15574 8444 15580
rect 7656 15088 7708 15094
rect 7656 15030 7708 15036
rect 8300 15088 8352 15094
rect 8300 15030 8352 15036
rect 8404 15026 8432 15574
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 7840 14816 7892 14822
rect 7840 14758 7892 14764
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7562 14376 7618 14385
rect 7472 14340 7524 14346
rect 7562 14311 7618 14320
rect 7472 14282 7524 14288
rect 7576 14113 7604 14311
rect 7852 14278 7880 14758
rect 8496 14618 8524 16730
rect 8588 15706 8616 18022
rect 8942 17983 8998 17992
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8680 17338 8708 17614
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8760 16652 8812 16658
rect 8760 16594 8812 16600
rect 8772 15910 8800 16594
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7562 14104 7618 14113
rect 7562 14039 7618 14048
rect 7380 13456 7432 13462
rect 7380 13398 7432 13404
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7300 11801 7328 12582
rect 7286 11792 7342 11801
rect 7392 11762 7420 13398
rect 7576 12782 7604 14039
rect 7852 13433 7880 14214
rect 8312 14074 8340 14350
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 7654 13424 7710 13433
rect 7654 13359 7710 13368
rect 7838 13424 7894 13433
rect 7838 13359 7894 13368
rect 7668 13002 7696 13359
rect 7746 13016 7802 13025
rect 7668 12974 7746 13002
rect 7746 12951 7802 12960
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 7484 12481 7512 12650
rect 7470 12472 7526 12481
rect 7470 12407 7526 12416
rect 7562 12336 7618 12345
rect 7562 12271 7564 12280
rect 7616 12271 7618 12280
rect 7564 12242 7616 12248
rect 7576 12073 7604 12242
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7562 12064 7618 12073
rect 7562 11999 7618 12008
rect 7576 11898 7604 11999
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7286 11727 7342 11736
rect 7380 11756 7432 11762
rect 7300 11694 7328 11727
rect 7380 11698 7432 11704
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7576 11286 7604 11698
rect 7668 11354 7696 12174
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7564 11280 7616 11286
rect 7564 11222 7616 11228
rect 7208 10662 7328 10690
rect 7196 10532 7248 10538
rect 7196 10474 7248 10480
rect 7208 10266 7236 10474
rect 7196 10260 7248 10266
rect 6932 10220 7052 10248
rect 6552 10202 6604 10208
rect 6422 10118 6500 10146
rect 6366 10095 6422 10104
rect 6380 9722 6408 10095
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6472 9382 6500 9998
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6472 8514 6500 9318
rect 6564 8634 6592 10202
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6644 10056 6696 10062
rect 6932 10010 6960 10066
rect 6644 9998 6696 10004
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6472 8486 6592 8514
rect 6564 8362 6592 8486
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 5368 7342 5396 7482
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 6380 7002 6408 7822
rect 4712 6996 4764 7002
rect 4712 6938 4764 6944
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 5956 6556 6252 6576
rect 6012 6554 6036 6556
rect 6092 6554 6116 6556
rect 6172 6554 6196 6556
rect 6034 6502 6036 6554
rect 6098 6502 6110 6554
rect 6172 6502 6174 6554
rect 6012 6500 6036 6502
rect 6092 6500 6116 6502
rect 6172 6500 6196 6502
rect 5956 6480 6252 6500
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 5956 5468 6252 5488
rect 6012 5466 6036 5468
rect 6092 5466 6116 5468
rect 6172 5466 6196 5468
rect 6034 5414 6036 5466
rect 6098 5414 6110 5466
rect 6172 5414 6174 5466
rect 6012 5412 6036 5414
rect 6092 5412 6116 5414
rect 6172 5412 6196 5414
rect 5956 5392 6252 5412
rect 5956 4380 6252 4400
rect 6012 4378 6036 4380
rect 6092 4378 6116 4380
rect 6172 4378 6196 4380
rect 6034 4326 6036 4378
rect 6098 4326 6110 4378
rect 6172 4326 6174 4378
rect 6012 4324 6036 4326
rect 6092 4324 6116 4326
rect 6172 4324 6196 4326
rect 5956 4304 6252 4324
rect 4342 3904 4398 3913
rect 4342 3839 4398 3848
rect 5956 3292 6252 3312
rect 6012 3290 6036 3292
rect 6092 3290 6116 3292
rect 6172 3290 6196 3292
rect 6034 3238 6036 3290
rect 6098 3238 6110 3290
rect 6172 3238 6174 3290
rect 6012 3236 6036 3238
rect 6092 3236 6116 3238
rect 6172 3236 6196 3238
rect 5956 3216 6252 3236
rect 6564 2650 6592 8298
rect 6656 8090 6684 9998
rect 6748 9982 6960 10010
rect 6748 8634 6776 9982
rect 7024 9178 7052 10220
rect 7196 10202 7248 10208
rect 7194 10024 7250 10033
rect 7194 9959 7196 9968
rect 7248 9959 7250 9968
rect 7196 9930 7248 9936
rect 7300 9874 7328 10662
rect 7208 9846 7328 9874
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 7116 8974 7144 9386
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6840 8090 6868 8842
rect 7208 8430 7236 9846
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7196 8424 7248 8430
rect 7194 8392 7196 8401
rect 7248 8392 7250 8401
rect 7194 8327 7250 8336
rect 7392 8090 7420 9114
rect 7484 8498 7512 9318
rect 7760 9178 7788 12951
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7760 8634 7788 9114
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6748 7546 6776 7890
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6840 7478 6868 8026
rect 7392 7857 7420 8026
rect 7484 7886 7512 8434
rect 7472 7880 7524 7886
rect 7378 7848 7434 7857
rect 7472 7822 7524 7828
rect 7378 7783 7434 7792
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 7760 7410 7788 7686
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7852 7206 7880 13359
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 6932 6662 6960 7142
rect 7944 7041 7972 11018
rect 8036 8106 8064 13126
rect 8220 12442 8248 13806
rect 8576 13728 8628 13734
rect 8576 13670 8628 13676
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8128 11762 8156 12038
rect 8116 11756 8168 11762
rect 8116 11698 8168 11704
rect 8390 11656 8446 11665
rect 8390 11591 8446 11600
rect 8404 11354 8432 11591
rect 8392 11348 8444 11354
rect 8444 11308 8524 11336
rect 8392 11290 8444 11296
rect 8298 11248 8354 11257
rect 8298 11183 8300 11192
rect 8352 11183 8354 11192
rect 8300 11154 8352 11160
rect 8300 11076 8352 11082
rect 8300 11018 8352 11024
rect 8312 10470 8340 11018
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8128 9654 8156 9998
rect 8116 9648 8168 9654
rect 8312 9625 8340 10406
rect 8404 10305 8432 10542
rect 8390 10296 8446 10305
rect 8496 10266 8524 11308
rect 8390 10231 8446 10240
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8588 9636 8616 13670
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8116 9590 8168 9596
rect 8298 9616 8354 9625
rect 8298 9551 8354 9560
rect 8496 9608 8616 9636
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8220 8498 8248 8774
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8036 8078 8156 8106
rect 8128 7750 8156 8078
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 7930 7032 7986 7041
rect 7930 6967 7986 6976
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6932 5817 6960 6598
rect 6918 5808 6974 5817
rect 6918 5743 6974 5752
rect 8128 4049 8156 7686
rect 8220 7410 8248 8434
rect 8496 8430 8524 9608
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8404 7857 8432 8230
rect 8390 7848 8446 7857
rect 8390 7783 8446 7792
rect 8404 7750 8432 7783
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8220 7290 8248 7346
rect 8220 7262 8340 7290
rect 8114 4040 8170 4049
rect 8114 3975 8170 3984
rect 8312 2650 8340 7262
rect 8680 6934 8708 10406
rect 8772 9761 8800 15846
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8864 12782 8892 13126
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8864 12442 8892 12718
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8864 11762 8892 12378
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8852 11552 8904 11558
rect 8850 11520 8852 11529
rect 8904 11520 8906 11529
rect 8850 11455 8906 11464
rect 8956 10577 8984 17983
rect 9048 16590 9076 18226
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 9220 15088 9272 15094
rect 9220 15030 9272 15036
rect 9232 14482 9260 15030
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9140 13870 9168 14214
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9220 11892 9272 11898
rect 9324 11880 9352 20159
rect 9586 19544 9642 19553
rect 9586 19479 9642 19488
rect 9600 19417 9628 19479
rect 9586 19408 9642 19417
rect 9586 19343 9642 19352
rect 9588 18216 9640 18222
rect 9586 18184 9588 18193
rect 9640 18184 9642 18193
rect 9586 18119 9642 18128
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9416 17241 9444 17818
rect 9588 17740 9640 17746
rect 9588 17682 9640 17688
rect 9600 17270 9628 17682
rect 9588 17264 9640 17270
rect 9402 17232 9458 17241
rect 9588 17206 9640 17212
rect 9402 17167 9458 17176
rect 9496 17060 9548 17066
rect 9496 17002 9548 17008
rect 9508 16697 9536 17002
rect 9494 16688 9550 16697
rect 9494 16623 9550 16632
rect 9588 16652 9640 16658
rect 9508 16250 9536 16623
rect 9588 16594 9640 16600
rect 9496 16244 9548 16250
rect 9416 16204 9496 16232
rect 9416 14414 9444 16204
rect 9496 16186 9548 16192
rect 9600 15450 9628 16594
rect 9692 15706 9720 20198
rect 9784 18970 9812 20742
rect 10244 20602 10272 23520
rect 12176 23474 12204 23520
rect 12084 23446 12204 23474
rect 10600 22840 10652 22846
rect 10600 22782 10652 22788
rect 10232 20596 10284 20602
rect 10232 20538 10284 20544
rect 10140 19304 10192 19310
rect 10140 19246 10192 19252
rect 10152 18970 10180 19246
rect 10416 19168 10468 19174
rect 10336 19128 10416 19156
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 10232 18828 10284 18834
rect 10232 18770 10284 18776
rect 10244 18426 10272 18770
rect 10336 18766 10364 19128
rect 10416 19110 10468 19116
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 10336 18358 10364 18702
rect 10612 18358 10640 22782
rect 10956 21244 11252 21264
rect 11012 21242 11036 21244
rect 11092 21242 11116 21244
rect 11172 21242 11196 21244
rect 11034 21190 11036 21242
rect 11098 21190 11110 21242
rect 11172 21190 11174 21242
rect 11012 21188 11036 21190
rect 11092 21188 11116 21190
rect 11172 21188 11196 21190
rect 10956 21168 11252 21188
rect 10784 20324 10836 20330
rect 10784 20266 10836 20272
rect 10796 19514 10824 20266
rect 10956 20156 11252 20176
rect 11012 20154 11036 20156
rect 11092 20154 11116 20156
rect 11172 20154 11196 20156
rect 11034 20102 11036 20154
rect 11098 20102 11110 20154
rect 11172 20102 11174 20154
rect 11012 20100 11036 20102
rect 11092 20100 11116 20102
rect 11172 20100 11196 20102
rect 10956 20080 11252 20100
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 10968 19780 11020 19786
rect 10968 19722 11020 19728
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10784 19508 10836 19514
rect 10784 19450 10836 19456
rect 10888 19378 10916 19654
rect 10876 19372 10928 19378
rect 10876 19314 10928 19320
rect 10980 19310 11008 19722
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 11348 19174 11376 19314
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 10956 19068 11252 19088
rect 11012 19066 11036 19068
rect 11092 19066 11116 19068
rect 11172 19066 11196 19068
rect 11034 19014 11036 19066
rect 11098 19014 11110 19066
rect 11172 19014 11174 19066
rect 11012 19012 11036 19014
rect 11092 19012 11116 19014
rect 11172 19012 11196 19014
rect 10956 18992 11252 19012
rect 11348 18970 11376 19110
rect 11336 18964 11388 18970
rect 11336 18906 11388 18912
rect 11440 18902 11468 19790
rect 11808 19174 11836 19994
rect 11888 19304 11940 19310
rect 12084 19281 12112 23446
rect 14016 21146 14044 23520
rect 15948 23474 15976 23520
rect 15856 23446 15976 23474
rect 14004 21140 14056 21146
rect 14004 21082 14056 21088
rect 12164 21004 12216 21010
rect 12164 20946 12216 20952
rect 12176 20534 12204 20946
rect 12808 20800 12860 20806
rect 12808 20742 12860 20748
rect 12164 20528 12216 20534
rect 12164 20470 12216 20476
rect 12820 20398 12848 20742
rect 15856 20602 15884 23446
rect 15956 21788 16252 21808
rect 16012 21786 16036 21788
rect 16092 21786 16116 21788
rect 16172 21786 16196 21788
rect 16034 21734 16036 21786
rect 16098 21734 16110 21786
rect 16172 21734 16174 21786
rect 16012 21732 16036 21734
rect 16092 21732 16116 21734
rect 16172 21732 16196 21734
rect 15956 21712 16252 21732
rect 17132 21004 17184 21010
rect 17132 20946 17184 20952
rect 15956 20700 16252 20720
rect 16012 20698 16036 20700
rect 16092 20698 16116 20700
rect 16172 20698 16196 20700
rect 16034 20646 16036 20698
rect 16098 20646 16110 20698
rect 16172 20646 16174 20698
rect 16012 20644 16036 20646
rect 16092 20644 16116 20646
rect 16172 20644 16196 20646
rect 15956 20624 16252 20644
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 13636 20460 13688 20466
rect 13636 20402 13688 20408
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 12636 20262 12664 20334
rect 12624 20256 12676 20262
rect 12624 20198 12676 20204
rect 12164 19916 12216 19922
rect 12164 19858 12216 19864
rect 11888 19246 11940 19252
rect 12070 19272 12126 19281
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11428 18896 11480 18902
rect 10782 18864 10838 18873
rect 11428 18838 11480 18844
rect 11702 18864 11758 18873
rect 10782 18799 10838 18808
rect 10796 18630 10824 18799
rect 10784 18624 10836 18630
rect 10784 18566 10836 18572
rect 10324 18352 10376 18358
rect 10324 18294 10376 18300
rect 10600 18352 10652 18358
rect 10600 18294 10652 18300
rect 10612 18222 10640 18294
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 10692 18148 10744 18154
rect 10692 18090 10744 18096
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 9784 17338 9812 17682
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 9954 16008 10010 16017
rect 9954 15943 10010 15952
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9692 15450 9720 15506
rect 9600 15422 9720 15450
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9496 14884 9548 14890
rect 9496 14826 9548 14832
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9508 14278 9536 14826
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9508 13938 9536 14214
rect 9600 14074 9628 15422
rect 9784 15162 9812 15438
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9784 13530 9812 15098
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9402 12200 9458 12209
rect 9402 12135 9458 12144
rect 9416 11898 9444 12135
rect 9272 11852 9352 11880
rect 9404 11892 9456 11898
rect 9220 11834 9272 11840
rect 9404 11834 9456 11840
rect 9968 11830 9996 15943
rect 10244 15706 10272 16526
rect 10428 15910 10456 16594
rect 10506 16280 10562 16289
rect 10506 16215 10562 16224
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10336 14482 10364 15438
rect 10428 14793 10456 15846
rect 10414 14784 10470 14793
rect 10414 14719 10470 14728
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10324 14272 10376 14278
rect 10428 14249 10456 14719
rect 10324 14214 10376 14220
rect 10414 14240 10470 14249
rect 10336 14074 10364 14214
rect 10414 14175 10470 14184
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10336 13870 10364 14010
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10324 13864 10376 13870
rect 10428 13841 10456 13874
rect 10324 13806 10376 13812
rect 10414 13832 10470 13841
rect 10414 13767 10470 13776
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 10244 13530 10272 13670
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10060 11898 10088 13466
rect 10428 13326 10456 13767
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10428 12442 10456 13262
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 9956 11824 10008 11830
rect 10244 11801 10272 12038
rect 9956 11766 10008 11772
rect 10230 11792 10286 11801
rect 10230 11727 10286 11736
rect 10520 11642 10548 16215
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 10612 15745 10640 15982
rect 10704 15881 10732 18090
rect 10796 18086 10824 18566
rect 11150 18320 11206 18329
rect 11440 18290 11468 18838
rect 11702 18799 11758 18808
rect 11716 18601 11744 18799
rect 11808 18737 11836 19110
rect 11794 18728 11850 18737
rect 11794 18663 11850 18672
rect 11702 18592 11758 18601
rect 11702 18527 11758 18536
rect 11808 18465 11836 18663
rect 11794 18456 11850 18465
rect 11900 18426 11928 19246
rect 12070 19207 12126 19216
rect 11794 18391 11850 18400
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11150 18255 11206 18264
rect 11428 18284 11480 18290
rect 11164 18222 11192 18255
rect 11428 18226 11480 18232
rect 11152 18216 11204 18222
rect 11152 18158 11204 18164
rect 10784 18080 10836 18086
rect 10782 18048 10784 18057
rect 10836 18048 10838 18057
rect 10782 17983 10838 17992
rect 10956 17980 11252 18000
rect 11012 17978 11036 17980
rect 11092 17978 11116 17980
rect 11172 17978 11196 17980
rect 11034 17926 11036 17978
rect 11098 17926 11110 17978
rect 11172 17926 11174 17978
rect 11012 17924 11036 17926
rect 11092 17924 11116 17926
rect 11172 17924 11196 17926
rect 10956 17904 11252 17924
rect 11440 17882 11468 18226
rect 12176 17882 12204 19858
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12256 19236 12308 19242
rect 12256 19178 12308 19184
rect 12268 18816 12296 19178
rect 12544 19174 12572 19246
rect 12716 19236 12768 19242
rect 12716 19178 12768 19184
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12544 18834 12572 19110
rect 12728 18970 12756 19178
rect 13004 19174 13032 19654
rect 13648 19514 13676 20402
rect 13820 20392 13872 20398
rect 13740 20340 13820 20346
rect 13740 20334 13872 20340
rect 16672 20392 16724 20398
rect 16672 20334 16724 20340
rect 13740 20318 13860 20334
rect 13636 19508 13688 19514
rect 13636 19450 13688 19456
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 12716 18964 12768 18970
rect 12716 18906 12768 18912
rect 12532 18828 12584 18834
rect 12268 18788 12480 18816
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 12164 17876 12216 17882
rect 12164 17818 12216 17824
rect 10784 17808 10836 17814
rect 10784 17750 10836 17756
rect 10796 17338 10824 17750
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11794 17640 11850 17649
rect 11244 17604 11296 17610
rect 11244 17546 11296 17552
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 11150 17232 11206 17241
rect 11150 17167 11206 17176
rect 11164 17134 11192 17167
rect 11152 17128 11204 17134
rect 11256 17105 11284 17546
rect 11532 17542 11560 17614
rect 11794 17575 11850 17584
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11152 17070 11204 17076
rect 11242 17096 11298 17105
rect 11242 17031 11244 17040
rect 11296 17031 11298 17040
rect 11244 17002 11296 17008
rect 10956 16892 11252 16912
rect 11012 16890 11036 16892
rect 11092 16890 11116 16892
rect 11172 16890 11196 16892
rect 11034 16838 11036 16890
rect 11098 16838 11110 16890
rect 11172 16838 11174 16890
rect 11012 16836 11036 16838
rect 11092 16836 11116 16838
rect 11172 16836 11196 16838
rect 10956 16816 11252 16836
rect 11348 16794 11376 17138
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 10784 16720 10836 16726
rect 11348 16697 11376 16730
rect 10784 16662 10836 16668
rect 11334 16688 11390 16697
rect 10796 16250 10824 16662
rect 11532 16658 11560 17478
rect 11808 17338 11836 17575
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11808 17134 11836 17274
rect 11796 17128 11848 17134
rect 11610 17096 11666 17105
rect 11796 17070 11848 17076
rect 11610 17031 11666 17040
rect 11334 16623 11390 16632
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 11428 16584 11480 16590
rect 11428 16526 11480 16532
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 11072 16114 11100 16390
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 10784 15904 10836 15910
rect 10690 15872 10746 15881
rect 10784 15846 10836 15852
rect 10690 15807 10746 15816
rect 10598 15736 10654 15745
rect 10598 15671 10654 15680
rect 10600 14000 10652 14006
rect 10598 13968 10600 13977
rect 10652 13968 10654 13977
rect 10598 13903 10654 13912
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10612 11898 10640 12174
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 10428 11614 10548 11642
rect 8942 10568 8998 10577
rect 8942 10503 8998 10512
rect 9232 10266 9260 11562
rect 9310 11384 9366 11393
rect 9310 11319 9312 11328
rect 9364 11319 9366 11328
rect 9312 11290 9364 11296
rect 10428 11218 10456 11614
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10520 11354 10548 11494
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10428 10538 10456 11154
rect 10520 10810 10548 11290
rect 10612 11082 10640 11698
rect 10704 11150 10732 15807
rect 10796 15366 10824 15846
rect 10956 15804 11252 15824
rect 11012 15802 11036 15804
rect 11092 15802 11116 15804
rect 11172 15802 11196 15804
rect 11034 15750 11036 15802
rect 11098 15750 11110 15802
rect 11172 15750 11174 15802
rect 11012 15748 11036 15750
rect 11092 15748 11116 15750
rect 11172 15748 11196 15750
rect 10956 15728 11252 15748
rect 11348 15638 11376 16050
rect 11336 15632 11388 15638
rect 11336 15574 11388 15580
rect 11440 15502 11468 16526
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 10796 12753 10824 15302
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 10956 14716 11252 14736
rect 11012 14714 11036 14716
rect 11092 14714 11116 14716
rect 11172 14714 11196 14716
rect 11034 14662 11036 14714
rect 11098 14662 11110 14714
rect 11172 14662 11174 14714
rect 11012 14660 11036 14662
rect 11092 14660 11116 14662
rect 11172 14660 11196 14662
rect 10956 14640 11252 14660
rect 11348 14482 11376 14758
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10888 13938 10916 14214
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10888 13172 10916 13670
rect 10956 13628 11252 13648
rect 11012 13626 11036 13628
rect 11092 13626 11116 13628
rect 11172 13626 11196 13628
rect 11034 13574 11036 13626
rect 11098 13574 11110 13626
rect 11172 13574 11174 13626
rect 11012 13572 11036 13574
rect 11092 13572 11116 13574
rect 11172 13572 11196 13574
rect 10956 13552 11252 13572
rect 11348 13530 11376 14418
rect 11440 14278 11468 15438
rect 11532 15162 11560 16594
rect 11624 16046 11652 17031
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 11794 16280 11850 16289
rect 11794 16215 11796 16224
rect 11848 16215 11850 16224
rect 11796 16186 11848 16192
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11702 16008 11758 16017
rect 11808 15978 11836 16186
rect 11702 15943 11758 15952
rect 11796 15972 11848 15978
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11520 15156 11572 15162
rect 11520 15098 11572 15104
rect 11428 14272 11480 14278
rect 11428 14214 11480 14220
rect 11428 13932 11480 13938
rect 11428 13874 11480 13880
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11440 13394 11468 13874
rect 11520 13796 11572 13802
rect 11520 13738 11572 13744
rect 11532 13530 11560 13738
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 11428 13388 11480 13394
rect 11428 13330 11480 13336
rect 10968 13184 11020 13190
rect 10888 13144 10968 13172
rect 10968 13126 11020 13132
rect 10876 12912 10928 12918
rect 10876 12854 10928 12860
rect 10782 12744 10838 12753
rect 10782 12679 10838 12688
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10796 12442 10824 12582
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 10796 11762 10824 12378
rect 10888 12374 10916 12854
rect 10980 12850 11008 13126
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 10956 12540 11252 12560
rect 11012 12538 11036 12540
rect 11092 12538 11116 12540
rect 11172 12538 11196 12540
rect 11034 12486 11036 12538
rect 11098 12486 11110 12538
rect 11172 12486 11174 12538
rect 11012 12484 11036 12486
rect 11092 12484 11116 12486
rect 11172 12484 11196 12486
rect 10956 12464 11252 12484
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10888 11150 10916 12310
rect 10956 11452 11252 11472
rect 11012 11450 11036 11452
rect 11092 11450 11116 11452
rect 11172 11450 11196 11452
rect 11034 11398 11036 11450
rect 11098 11398 11110 11450
rect 11172 11398 11174 11450
rect 11012 11396 11036 11398
rect 11092 11396 11116 11398
rect 11172 11396 11196 11398
rect 10956 11376 11252 11396
rect 11348 11354 11376 13330
rect 11624 13025 11652 15846
rect 11716 15473 11744 15943
rect 11796 15914 11848 15920
rect 12164 15632 12216 15638
rect 12164 15574 12216 15580
rect 11796 15496 11848 15502
rect 11702 15464 11758 15473
rect 11796 15438 11848 15444
rect 11702 15399 11758 15408
rect 11808 15026 11836 15438
rect 12176 15162 12204 15574
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 12176 14618 12204 15098
rect 12164 14612 12216 14618
rect 12164 14554 12216 14560
rect 11794 14512 11850 14521
rect 11794 14447 11850 14456
rect 11808 13530 11836 14447
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11796 13524 11848 13530
rect 11716 13484 11796 13512
rect 11610 13016 11666 13025
rect 11520 12980 11572 12986
rect 11610 12951 11666 12960
rect 11520 12922 11572 12928
rect 11428 12368 11480 12374
rect 11428 12310 11480 12316
rect 11440 11830 11468 12310
rect 11428 11824 11480 11830
rect 11428 11766 11480 11772
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 10598 10840 10654 10849
rect 10508 10804 10560 10810
rect 10598 10775 10654 10784
rect 10508 10746 10560 10752
rect 10612 10606 10640 10775
rect 10704 10674 10732 11086
rect 10888 10810 10916 11086
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10600 10600 10652 10606
rect 10600 10542 10652 10548
rect 10416 10532 10468 10538
rect 10416 10474 10468 10480
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 10336 10062 10364 10406
rect 10612 10266 10640 10542
rect 10956 10364 11252 10384
rect 11012 10362 11036 10364
rect 11092 10362 11116 10364
rect 11172 10362 11196 10364
rect 11034 10310 11036 10362
rect 11098 10310 11110 10362
rect 11172 10310 11174 10362
rect 11012 10308 11036 10310
rect 11092 10308 11116 10310
rect 11172 10308 11196 10310
rect 10956 10288 11252 10308
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10324 10056 10376 10062
rect 10322 10024 10324 10033
rect 10376 10024 10378 10033
rect 10322 9959 10378 9968
rect 8758 9752 8814 9761
rect 8758 9687 8814 9696
rect 8772 9636 8800 9687
rect 8772 9608 8892 9636
rect 8864 8616 8892 9608
rect 10956 9276 11252 9296
rect 11012 9274 11036 9276
rect 11092 9274 11116 9276
rect 11172 9274 11196 9276
rect 11034 9222 11036 9274
rect 11098 9222 11110 9274
rect 11172 9222 11174 9274
rect 11012 9220 11036 9222
rect 11092 9220 11116 9222
rect 11172 9220 11196 9222
rect 10956 9200 11252 9220
rect 8864 8588 8984 8616
rect 8850 8528 8906 8537
rect 8850 8463 8906 8472
rect 8864 8430 8892 8463
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8956 8022 8984 8588
rect 10956 8188 11252 8208
rect 11012 8186 11036 8188
rect 11092 8186 11116 8188
rect 11172 8186 11196 8188
rect 11034 8134 11036 8186
rect 11098 8134 11110 8186
rect 11172 8134 11174 8186
rect 11012 8132 11036 8134
rect 11092 8132 11116 8134
rect 11172 8132 11196 8134
rect 10956 8112 11252 8132
rect 8944 8016 8996 8022
rect 8944 7958 8996 7964
rect 11532 7313 11560 12922
rect 11716 12918 11744 13484
rect 11796 13466 11848 13472
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 11808 12442 11836 13330
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11900 11898 11928 13806
rect 11980 13320 12032 13326
rect 11978 13288 11980 13297
rect 12032 13288 12034 13297
rect 11978 13223 12034 13232
rect 11992 12986 12020 13223
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 12164 12912 12216 12918
rect 12162 12880 12164 12889
rect 12268 12900 12296 16934
rect 12452 16250 12480 18788
rect 12532 18770 12584 18776
rect 12544 18290 12572 18770
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 12992 18080 13044 18086
rect 12992 18022 13044 18028
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12728 17202 12756 17614
rect 13004 17542 13032 18022
rect 13096 17814 13124 18226
rect 13740 17882 13768 20318
rect 16684 20058 16712 20334
rect 17144 20262 17172 20946
rect 17788 20602 17816 23520
rect 19628 21146 19656 23520
rect 20956 21244 21252 21264
rect 21012 21242 21036 21244
rect 21092 21242 21116 21244
rect 21172 21242 21196 21244
rect 21034 21190 21036 21242
rect 21098 21190 21110 21242
rect 21172 21190 21174 21242
rect 21012 21188 21036 21190
rect 21092 21188 21116 21190
rect 21172 21188 21196 21190
rect 20956 21168 21252 21188
rect 19616 21140 19668 21146
rect 19616 21082 19668 21088
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 19616 21004 19668 21010
rect 19616 20946 19668 20952
rect 17776 20596 17828 20602
rect 17776 20538 17828 20544
rect 17972 20482 18000 20946
rect 18696 20868 18748 20874
rect 18696 20810 18748 20816
rect 18236 20800 18288 20806
rect 18236 20742 18288 20748
rect 17788 20454 18000 20482
rect 17788 20398 17816 20454
rect 17776 20392 17828 20398
rect 17774 20360 17776 20369
rect 17828 20360 17830 20369
rect 17774 20295 17830 20304
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 15382 19816 15438 19825
rect 15382 19751 15438 19760
rect 15108 19712 15160 19718
rect 14278 19680 14334 19689
rect 15108 19654 15160 19660
rect 14278 19615 14334 19624
rect 13912 19508 13964 19514
rect 13912 19450 13964 19456
rect 13924 18970 13952 19450
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13924 18154 13952 18906
rect 13912 18148 13964 18154
rect 13912 18090 13964 18096
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13084 17808 13136 17814
rect 13084 17750 13136 17756
rect 13820 17808 13872 17814
rect 13820 17750 13872 17756
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 13004 17338 13032 17478
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12992 17060 13044 17066
rect 12992 17002 13044 17008
rect 13004 16697 13032 17002
rect 13096 16794 13124 17750
rect 13266 17232 13322 17241
rect 13266 17167 13322 17176
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 12990 16688 13046 16697
rect 12990 16623 13046 16632
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12348 16108 12400 16114
rect 12348 16050 12400 16056
rect 12360 16017 12388 16050
rect 12346 16008 12402 16017
rect 12346 15943 12348 15952
rect 12400 15943 12402 15952
rect 12348 15914 12400 15920
rect 12900 15904 12952 15910
rect 12898 15872 12900 15881
rect 12952 15872 12954 15881
rect 12898 15807 12954 15816
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12716 13796 12768 13802
rect 12716 13738 12768 13744
rect 12728 13258 12756 13738
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12216 12880 12296 12900
rect 12218 12872 12296 12880
rect 11980 12844 12032 12850
rect 12636 12850 12664 13126
rect 12162 12815 12218 12824
rect 12348 12844 12400 12850
rect 11980 12786 12032 12792
rect 12348 12786 12400 12792
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11794 11656 11850 11665
rect 11794 11591 11796 11600
rect 11848 11591 11850 11600
rect 11796 11562 11848 11568
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11808 10810 11836 11018
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11992 10169 12020 12786
rect 12360 12374 12388 12786
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12348 12368 12400 12374
rect 12348 12310 12400 12316
rect 12348 11348 12400 11354
rect 12452 11336 12480 12582
rect 12728 12442 12756 12582
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12912 11937 12940 14758
rect 13004 12646 13032 16623
rect 13096 16250 13124 16730
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 13084 15972 13136 15978
rect 13084 15914 13136 15920
rect 13096 15026 13124 15914
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 13096 13870 13124 14962
rect 13280 14958 13308 17167
rect 13832 16998 13860 17750
rect 14004 17740 14056 17746
rect 14004 17682 14056 17688
rect 13820 16992 13872 16998
rect 13740 16940 13820 16946
rect 13740 16934 13872 16940
rect 13740 16918 13860 16934
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 13280 14618 13308 14894
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13280 14113 13308 14554
rect 13556 14346 13584 14962
rect 13740 14618 13768 16918
rect 14016 16833 14044 17682
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14200 17338 14228 17614
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 13818 16824 13874 16833
rect 13818 16759 13820 16768
rect 13872 16759 13874 16768
rect 14002 16824 14058 16833
rect 14002 16759 14058 16768
rect 13820 16730 13872 16736
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13832 14414 13860 16594
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 14108 15162 14136 15302
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 14004 14884 14056 14890
rect 14004 14826 14056 14832
rect 14016 14482 14044 14826
rect 14108 14618 14136 15098
rect 14292 15026 14320 19615
rect 14832 19304 14884 19310
rect 14832 19246 14884 19252
rect 14844 18873 14872 19246
rect 14924 19236 14976 19242
rect 14924 19178 14976 19184
rect 14830 18864 14886 18873
rect 14830 18799 14886 18808
rect 14936 18630 14964 19178
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 14924 18624 14976 18630
rect 14924 18566 14976 18572
rect 14936 17202 14964 18566
rect 15028 18057 15056 19110
rect 15014 18048 15070 18057
rect 15014 17983 15070 17992
rect 14924 17196 14976 17202
rect 14924 17138 14976 17144
rect 15120 16590 15148 19654
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15304 17678 15332 18022
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15200 16992 15252 16998
rect 15304 16980 15332 17614
rect 15252 16952 15332 16980
rect 15200 16934 15252 16940
rect 14464 16584 14516 16590
rect 14464 16526 14516 16532
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 14476 16046 14504 16526
rect 14464 16040 14516 16046
rect 14464 15982 14516 15988
rect 14476 15706 14504 15982
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 15120 15026 15148 16526
rect 15304 15978 15332 16952
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 15304 15502 15332 15914
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 15304 14958 15332 15438
rect 14832 14952 14884 14958
rect 15292 14952 15344 14958
rect 14832 14894 14884 14900
rect 15198 14920 15254 14929
rect 14844 14657 14872 14894
rect 15292 14894 15344 14900
rect 15198 14855 15254 14864
rect 14830 14648 14886 14657
rect 14096 14612 14148 14618
rect 14830 14583 14886 14592
rect 14096 14554 14148 14560
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 13820 14408 13872 14414
rect 13740 14356 13820 14362
rect 13740 14350 13872 14356
rect 13544 14340 13596 14346
rect 13544 14282 13596 14288
rect 13740 14334 13860 14350
rect 13266 14104 13322 14113
rect 13266 14039 13322 14048
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 13740 13530 13768 14334
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13832 13841 13860 13942
rect 13818 13832 13874 13841
rect 13818 13767 13874 13776
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13648 12889 13676 13126
rect 13634 12880 13690 12889
rect 13634 12815 13690 12824
rect 13924 12782 13952 13330
rect 13912 12776 13964 12782
rect 13910 12744 13912 12753
rect 13964 12744 13966 12753
rect 13910 12679 13966 12688
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 14016 12442 14044 14418
rect 14738 14240 14794 14249
rect 14738 14175 14794 14184
rect 14752 14074 14780 14175
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14752 13870 14780 14010
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14188 13796 14240 13802
rect 14188 13738 14240 13744
rect 14094 13560 14150 13569
rect 14094 13495 14096 13504
rect 14148 13495 14150 13504
rect 14096 13466 14148 13472
rect 14108 13025 14136 13466
rect 14200 13326 14228 13738
rect 14924 13728 14976 13734
rect 14924 13670 14976 13676
rect 14936 13462 14964 13670
rect 14924 13456 14976 13462
rect 14922 13424 14924 13433
rect 14976 13424 14978 13433
rect 14922 13359 14978 13368
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14094 13016 14150 13025
rect 14094 12951 14096 12960
rect 14148 12951 14150 12960
rect 14096 12922 14148 12928
rect 14108 12891 14136 12922
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 14200 12374 14228 13262
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15120 12918 15148 13126
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 15108 12912 15160 12918
rect 15108 12854 15160 12860
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 14752 12073 14780 12854
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15120 12442 15148 12718
rect 15212 12617 15240 14855
rect 15396 13190 15424 19751
rect 15568 19712 15620 19718
rect 15568 19654 15620 19660
rect 15580 19378 15608 19654
rect 15956 19612 16252 19632
rect 16012 19610 16036 19612
rect 16092 19610 16116 19612
rect 16172 19610 16196 19612
rect 16034 19558 16036 19610
rect 16098 19558 16110 19610
rect 16172 19558 16174 19610
rect 16012 19556 16036 19558
rect 16092 19556 16116 19558
rect 16172 19556 16196 19558
rect 15956 19536 16252 19556
rect 15568 19372 15620 19378
rect 15568 19314 15620 19320
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 16408 18601 16436 19110
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16394 18592 16450 18601
rect 15956 18524 16252 18544
rect 16394 18527 16450 18536
rect 16012 18522 16036 18524
rect 16092 18522 16116 18524
rect 16172 18522 16196 18524
rect 16034 18470 16036 18522
rect 16098 18470 16110 18522
rect 16172 18470 16174 18522
rect 16012 18468 16036 18470
rect 16092 18468 16116 18470
rect 16172 18468 16196 18470
rect 15956 18448 16252 18468
rect 16500 18086 16528 18702
rect 16776 18358 16804 18770
rect 16764 18352 16816 18358
rect 16764 18294 16816 18300
rect 15568 18080 15620 18086
rect 15568 18022 15620 18028
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16670 18048 16726 18057
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15488 16658 15516 17002
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15488 16250 15516 16594
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15580 15638 15608 18022
rect 15658 17776 15714 17785
rect 15658 17711 15714 17720
rect 15672 16658 15700 17711
rect 15856 17678 15884 18022
rect 16670 17983 16726 17992
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15956 17436 16252 17456
rect 16012 17434 16036 17436
rect 16092 17434 16116 17436
rect 16172 17434 16196 17436
rect 16034 17382 16036 17434
rect 16098 17382 16110 17434
rect 16172 17382 16174 17434
rect 16012 17380 16036 17382
rect 16092 17380 16116 17382
rect 16172 17380 16196 17382
rect 15956 17360 16252 17380
rect 16408 17338 16436 17682
rect 16578 17504 16634 17513
rect 16578 17439 16634 17448
rect 16396 17332 16448 17338
rect 16396 17274 16448 17280
rect 16592 16726 16620 17439
rect 16580 16720 16632 16726
rect 16580 16662 16632 16668
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16316 16561 16344 16594
rect 16302 16552 16358 16561
rect 16302 16487 16358 16496
rect 15956 16348 16252 16368
rect 16012 16346 16036 16348
rect 16092 16346 16116 16348
rect 16172 16346 16196 16348
rect 16034 16294 16036 16346
rect 16098 16294 16110 16346
rect 16172 16294 16174 16346
rect 16012 16292 16036 16294
rect 16092 16292 16116 16294
rect 16172 16292 16196 16294
rect 15956 16272 16252 16292
rect 16316 16182 16344 16487
rect 16304 16176 16356 16182
rect 16304 16118 16356 16124
rect 16488 15972 16540 15978
rect 16488 15914 16540 15920
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 15580 15094 15608 15574
rect 16500 15366 16528 15914
rect 16592 15910 16620 16662
rect 16684 16658 16712 17983
rect 16854 16824 16910 16833
rect 16854 16759 16910 16768
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16868 16522 16896 16759
rect 16856 16516 16908 16522
rect 16856 16458 16908 16464
rect 16580 15904 16632 15910
rect 16580 15846 16632 15852
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 15956 15260 16252 15280
rect 16012 15258 16036 15260
rect 16092 15258 16116 15260
rect 16172 15258 16196 15260
rect 16034 15206 16036 15258
rect 16098 15206 16110 15258
rect 16172 15206 16174 15258
rect 16012 15204 16036 15206
rect 16092 15204 16116 15206
rect 16172 15204 16196 15206
rect 15956 15184 16252 15204
rect 15568 15088 15620 15094
rect 15568 15030 15620 15036
rect 15844 15088 15896 15094
rect 15844 15030 15896 15036
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15568 13728 15620 13734
rect 15566 13696 15568 13705
rect 15620 13696 15622 13705
rect 15566 13631 15622 13640
rect 15384 13184 15436 13190
rect 15290 13152 15346 13161
rect 15384 13126 15436 13132
rect 15290 13087 15346 13096
rect 15198 12608 15254 12617
rect 15198 12543 15254 12552
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15304 12209 15332 13087
rect 15474 12880 15530 12889
rect 15384 12844 15436 12850
rect 15474 12815 15530 12824
rect 15384 12786 15436 12792
rect 15290 12200 15346 12209
rect 15290 12135 15346 12144
rect 14738 12064 14794 12073
rect 14738 11999 14794 12008
rect 12898 11928 12954 11937
rect 15396 11898 15424 12786
rect 12898 11863 12954 11872
rect 15384 11892 15436 11898
rect 12400 11308 12480 11336
rect 12348 11290 12400 11296
rect 12360 10810 12388 11290
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12544 10810 12572 11222
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 11978 10160 12034 10169
rect 11978 10095 12034 10104
rect 11518 7304 11574 7313
rect 11518 7239 11574 7248
rect 10956 7100 11252 7120
rect 11012 7098 11036 7100
rect 11092 7098 11116 7100
rect 11172 7098 11196 7100
rect 11034 7046 11036 7098
rect 11098 7046 11110 7098
rect 11172 7046 11174 7098
rect 11012 7044 11036 7046
rect 11092 7044 11116 7046
rect 11172 7044 11196 7046
rect 10956 7024 11252 7044
rect 8668 6928 8720 6934
rect 8668 6870 8720 6876
rect 10956 6012 11252 6032
rect 11012 6010 11036 6012
rect 11092 6010 11116 6012
rect 11172 6010 11196 6012
rect 11034 5958 11036 6010
rect 11098 5958 11110 6010
rect 11172 5958 11174 6010
rect 11012 5956 11036 5958
rect 11092 5956 11116 5958
rect 11172 5956 11196 5958
rect 10956 5936 11252 5956
rect 12912 5273 12940 11863
rect 15384 11834 15436 11840
rect 14278 11792 14334 11801
rect 14278 11727 14334 11736
rect 14292 10849 14320 11727
rect 14278 10840 14334 10849
rect 15396 10810 15424 11834
rect 15488 11218 15516 12815
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 14278 10775 14334 10784
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15488 10266 15516 11154
rect 15580 10810 15608 13631
rect 15672 13394 15700 14418
rect 15856 14414 15884 15030
rect 16500 15026 16528 15302
rect 16488 15020 16540 15026
rect 16408 14980 16488 15008
rect 16408 14550 16436 14980
rect 16488 14962 16540 14968
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16500 14618 16528 14758
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15856 13938 15884 14350
rect 15956 14172 16252 14192
rect 16012 14170 16036 14172
rect 16092 14170 16116 14172
rect 16172 14170 16196 14172
rect 16034 14118 16036 14170
rect 16098 14118 16110 14170
rect 16172 14118 16174 14170
rect 16012 14116 16036 14118
rect 16092 14116 16116 14118
rect 16172 14116 16196 14118
rect 15956 14096 16252 14116
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 16316 13870 16344 14418
rect 16500 14074 16528 14418
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 16028 13864 16080 13870
rect 16028 13806 16080 13812
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15672 12753 15700 13330
rect 15764 12866 15792 13806
rect 16040 13569 16068 13806
rect 16026 13560 16082 13569
rect 16026 13495 16082 13504
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 15856 12986 15884 13126
rect 15956 13084 16252 13104
rect 16012 13082 16036 13084
rect 16092 13082 16116 13084
rect 16172 13082 16196 13084
rect 16034 13030 16036 13082
rect 16098 13030 16110 13082
rect 16172 13030 16174 13082
rect 16012 13028 16036 13030
rect 16092 13028 16116 13030
rect 16172 13028 16196 13030
rect 15956 13008 16252 13028
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 16210 12880 16266 12889
rect 15764 12838 16210 12866
rect 16210 12815 16266 12824
rect 15658 12744 15714 12753
rect 15658 12679 15714 12688
rect 16120 12708 16172 12714
rect 16120 12650 16172 12656
rect 15842 12608 15898 12617
rect 15842 12543 15898 12552
rect 15856 12442 15884 12543
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15856 11898 15884 12378
rect 16132 12374 16160 12650
rect 16120 12368 16172 12374
rect 15934 12336 15990 12345
rect 16120 12310 16172 12316
rect 15934 12271 15936 12280
rect 15988 12271 15990 12280
rect 15936 12242 15988 12248
rect 16224 12186 16252 12815
rect 16316 12374 16344 13126
rect 16304 12368 16356 12374
rect 16304 12310 16356 12316
rect 16224 12158 16344 12186
rect 15956 11996 16252 12016
rect 16012 11994 16036 11996
rect 16092 11994 16116 11996
rect 16172 11994 16196 11996
rect 16034 11942 16036 11994
rect 16098 11942 16110 11994
rect 16172 11942 16174 11994
rect 16012 11940 16036 11942
rect 16092 11940 16116 11942
rect 16172 11940 16196 11942
rect 15956 11920 16252 11940
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15764 11014 15792 11494
rect 16316 11286 16344 12158
rect 16408 11898 16436 13806
rect 16500 12918 16528 14010
rect 16592 13852 16620 15846
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16684 14278 16712 14826
rect 17144 14618 17172 20198
rect 17512 19990 17540 20198
rect 17592 20052 17644 20058
rect 17592 19994 17644 20000
rect 17500 19984 17552 19990
rect 17500 19926 17552 19932
rect 17604 19514 17632 19994
rect 17972 19961 18000 20454
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 17958 19952 18014 19961
rect 17958 19887 18014 19896
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 17696 19242 17724 19790
rect 17684 19236 17736 19242
rect 17684 19178 17736 19184
rect 17696 18426 17724 19178
rect 17788 19174 17816 19790
rect 17776 19168 17828 19174
rect 17828 19116 17908 19122
rect 17776 19110 17908 19116
rect 17788 19094 17908 19110
rect 17880 18630 17908 19094
rect 17868 18624 17920 18630
rect 17868 18566 17920 18572
rect 17684 18420 17736 18426
rect 17684 18362 17736 18368
rect 17880 18034 17908 18566
rect 18156 18290 18184 20198
rect 18248 18970 18276 20742
rect 18708 20466 18736 20810
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18328 20324 18380 20330
rect 18328 20266 18380 20272
rect 18340 19718 18368 20266
rect 18420 20256 18472 20262
rect 18420 20198 18472 20204
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 18236 18964 18288 18970
rect 18236 18906 18288 18912
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 18248 18222 18276 18906
rect 18236 18216 18288 18222
rect 18236 18158 18288 18164
rect 17880 18006 18184 18034
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 17236 15706 17264 16730
rect 17512 16697 17540 16934
rect 17498 16688 17554 16697
rect 17498 16623 17554 16632
rect 17408 16584 17460 16590
rect 17408 16526 17460 16532
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17420 16250 17448 16526
rect 17408 16244 17460 16250
rect 17408 16186 17460 16192
rect 17604 15910 17632 16526
rect 17880 16454 17908 17614
rect 18156 16454 18184 18006
rect 18340 17338 18368 19654
rect 18328 17332 18380 17338
rect 18328 17274 18380 17280
rect 18432 16794 18460 20198
rect 18708 19990 18736 20402
rect 19628 20262 19656 20946
rect 21272 20800 21324 20806
rect 21272 20742 21324 20748
rect 20350 20632 20406 20641
rect 20350 20567 20352 20576
rect 20404 20567 20406 20576
rect 20352 20538 20404 20544
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 18696 19984 18748 19990
rect 18696 19926 18748 19932
rect 18708 19514 18736 19926
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19248 19848 19300 19854
rect 19248 19790 19300 19796
rect 19156 19780 19208 19786
rect 19156 19722 19208 19728
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 18604 19304 18656 19310
rect 18604 19246 18656 19252
rect 18616 18290 18644 19246
rect 18708 18970 18736 19450
rect 19168 19310 19196 19722
rect 19156 19304 19208 19310
rect 19154 19272 19156 19281
rect 19208 19272 19210 19281
rect 19260 19242 19288 19790
rect 19628 19718 19656 19858
rect 19616 19712 19668 19718
rect 19616 19654 19668 19660
rect 19154 19207 19210 19216
rect 19248 19236 19300 19242
rect 19168 19181 19196 19207
rect 19248 19178 19300 19184
rect 18880 19168 18932 19174
rect 18880 19110 18932 19116
rect 18696 18964 18748 18970
rect 18696 18906 18748 18912
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18892 18222 18920 19110
rect 19260 18970 19288 19178
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19430 18864 19486 18873
rect 19064 18828 19116 18834
rect 19430 18799 19486 18808
rect 19064 18770 19116 18776
rect 18880 18216 18932 18222
rect 19076 18193 19104 18770
rect 19444 18766 19472 18799
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 18880 18158 18932 18164
rect 19062 18184 19118 18193
rect 19062 18119 19064 18128
rect 19116 18119 19118 18128
rect 19064 18090 19116 18096
rect 19444 18086 19472 18702
rect 19628 18426 19656 19654
rect 19800 19236 19852 19242
rect 19800 19178 19852 19184
rect 19812 18902 19840 19178
rect 19892 19168 19944 19174
rect 19892 19110 19944 19116
rect 19800 18896 19852 18902
rect 19800 18838 19852 18844
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 19432 18080 19484 18086
rect 19430 18048 19432 18057
rect 19484 18048 19486 18057
rect 19430 17983 19486 17992
rect 19800 17808 19852 17814
rect 19154 17776 19210 17785
rect 19800 17750 19852 17756
rect 19154 17711 19210 17720
rect 19064 17196 19116 17202
rect 19064 17138 19116 17144
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 17868 16448 17920 16454
rect 17868 16390 17920 16396
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 17880 16046 17908 16390
rect 18156 16046 18184 16390
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17224 15700 17276 15706
rect 17224 15642 17276 15648
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 17420 14822 17448 15506
rect 17604 15094 17632 15846
rect 17880 15366 17908 15982
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18524 15570 18552 15846
rect 18512 15564 18564 15570
rect 18512 15506 18564 15512
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 18236 15360 18288 15366
rect 18236 15302 18288 15308
rect 17592 15088 17644 15094
rect 17592 15030 17644 15036
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16684 14006 16712 14214
rect 16672 14000 16724 14006
rect 16672 13942 16724 13948
rect 16776 13870 16804 14350
rect 16764 13864 16816 13870
rect 16592 13824 16712 13852
rect 16580 13728 16632 13734
rect 16684 13716 16712 13824
rect 16764 13806 16816 13812
rect 17420 13802 17448 14758
rect 17498 13832 17554 13841
rect 17408 13796 17460 13802
rect 17498 13767 17554 13776
rect 17408 13738 17460 13744
rect 17132 13728 17184 13734
rect 16684 13688 16804 13716
rect 16580 13670 16632 13676
rect 16488 12912 16540 12918
rect 16488 12854 16540 12860
rect 16592 12782 16620 13670
rect 16672 13524 16724 13530
rect 16672 13466 16724 13472
rect 16684 12850 16712 13466
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16580 12776 16632 12782
rect 16486 12744 16542 12753
rect 16580 12718 16632 12724
rect 16486 12679 16542 12688
rect 16500 12424 16528 12679
rect 16500 12396 16620 12424
rect 16592 12345 16620 12396
rect 16578 12336 16634 12345
rect 16488 12300 16540 12306
rect 16578 12271 16634 12280
rect 16488 12242 16540 12248
rect 16396 11892 16448 11898
rect 16396 11834 16448 11840
rect 16500 11626 16528 12242
rect 16684 12238 16712 12786
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16670 12064 16726 12073
rect 16670 11999 16726 12008
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 16304 11280 16356 11286
rect 16304 11222 16356 11228
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15764 10826 15792 10950
rect 15956 10908 16252 10928
rect 16012 10906 16036 10908
rect 16092 10906 16116 10908
rect 16172 10906 16196 10908
rect 16034 10854 16036 10906
rect 16098 10854 16110 10906
rect 16172 10854 16174 10906
rect 16012 10852 16036 10854
rect 16092 10852 16116 10854
rect 16172 10852 16196 10854
rect 15956 10832 16252 10852
rect 15568 10804 15620 10810
rect 15764 10798 15884 10826
rect 16316 10810 16344 11222
rect 16500 10962 16528 11562
rect 16500 10934 16620 10962
rect 15568 10746 15620 10752
rect 15856 10742 15884 10798
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 15844 10736 15896 10742
rect 15844 10678 15896 10684
rect 15476 10260 15528 10266
rect 15476 10202 15528 10208
rect 15956 9820 16252 9840
rect 16012 9818 16036 9820
rect 16092 9818 16116 9820
rect 16172 9818 16196 9820
rect 16034 9766 16036 9818
rect 16098 9766 16110 9818
rect 16172 9766 16174 9818
rect 16012 9764 16036 9766
rect 16092 9764 16116 9766
rect 16172 9764 16196 9766
rect 15750 9752 15806 9761
rect 15956 9744 16252 9764
rect 15750 9687 15806 9696
rect 15764 9654 15792 9687
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15948 9489 15976 9522
rect 15934 9480 15990 9489
rect 15476 9444 15528 9450
rect 15934 9415 15990 9424
rect 15476 9386 15528 9392
rect 15488 9178 15516 9386
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 16486 9344 16542 9353
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15956 8732 16252 8752
rect 16012 8730 16036 8732
rect 16092 8730 16116 8732
rect 16172 8730 16196 8732
rect 16034 8678 16036 8730
rect 16098 8678 16110 8730
rect 16172 8678 16174 8730
rect 16012 8676 16036 8678
rect 16092 8676 16116 8678
rect 16172 8676 16196 8678
rect 15956 8656 16252 8676
rect 16408 8430 16436 9318
rect 16486 9279 16542 9288
rect 16500 8974 16528 9279
rect 16592 9217 16620 10934
rect 16684 10538 16712 11999
rect 16672 10532 16724 10538
rect 16672 10474 16724 10480
rect 16684 10266 16712 10474
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16578 9208 16634 9217
rect 16578 9143 16634 9152
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16500 8634 16528 8910
rect 16488 8628 16540 8634
rect 16540 8588 16620 8616
rect 16488 8570 16540 8576
rect 16396 8424 16448 8430
rect 16316 8372 16396 8378
rect 16316 8366 16448 8372
rect 16316 8350 16436 8366
rect 16316 8090 16344 8350
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 15956 7644 16252 7664
rect 16012 7642 16036 7644
rect 16092 7642 16116 7644
rect 16172 7642 16196 7644
rect 16034 7590 16036 7642
rect 16098 7590 16110 7642
rect 16172 7590 16174 7642
rect 16012 7588 16036 7590
rect 16092 7588 16116 7590
rect 16172 7588 16196 7590
rect 15956 7568 16252 7588
rect 16408 7546 16436 8230
rect 16592 7954 16620 8588
rect 16684 8498 16712 9862
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16592 7546 16620 7890
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16408 7342 16436 7482
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16408 6866 16436 7142
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 15488 6458 15516 6802
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 12898 5264 12954 5273
rect 12898 5199 12954 5208
rect 10956 4924 11252 4944
rect 11012 4922 11036 4924
rect 11092 4922 11116 4924
rect 11172 4922 11196 4924
rect 11034 4870 11036 4922
rect 11098 4870 11110 4922
rect 11172 4870 11174 4922
rect 11012 4868 11036 4870
rect 11092 4868 11116 4870
rect 11172 4868 11196 4870
rect 10956 4848 11252 4868
rect 10956 3836 11252 3856
rect 11012 3834 11036 3836
rect 11092 3834 11116 3836
rect 11172 3834 11196 3836
rect 11034 3782 11036 3834
rect 11098 3782 11110 3834
rect 11172 3782 11174 3834
rect 11012 3780 11036 3782
rect 11092 3780 11116 3782
rect 11172 3780 11196 3782
rect 10956 3760 11252 3780
rect 15580 3505 15608 6598
rect 15956 6556 16252 6576
rect 16012 6554 16036 6556
rect 16092 6554 16116 6556
rect 16172 6554 16196 6556
rect 16034 6502 16036 6554
rect 16098 6502 16110 6554
rect 16172 6502 16174 6554
rect 16012 6500 16036 6502
rect 16092 6500 16116 6502
rect 16172 6500 16196 6502
rect 15956 6480 16252 6500
rect 16776 6361 16804 13688
rect 17132 13670 17184 13676
rect 17144 13190 17172 13670
rect 17512 13394 17540 13767
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 17052 12442 17080 12786
rect 17144 12782 17172 13126
rect 17512 12986 17540 13330
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 17144 12646 17172 12718
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16868 11354 16896 11494
rect 16960 11354 16988 12174
rect 17052 11762 17080 12378
rect 17144 12306 17172 12582
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17144 11898 17172 12242
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16960 11150 16988 11290
rect 17604 11200 17632 15030
rect 17880 14958 17908 15302
rect 18142 15056 18198 15065
rect 18142 14991 18198 15000
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17880 14822 17908 14894
rect 17868 14816 17920 14822
rect 17868 14758 17920 14764
rect 17776 14408 17828 14414
rect 17776 14350 17828 14356
rect 17788 13870 17816 14350
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17788 13190 17816 13806
rect 17880 13802 17908 14758
rect 17868 13796 17920 13802
rect 17868 13738 17920 13744
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 17788 12306 17816 13126
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 17788 11898 17816 12242
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17684 11212 17736 11218
rect 17604 11172 17684 11200
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16960 10674 16988 11086
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 17604 10606 17632 11172
rect 17684 11154 17736 11160
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 17972 10810 18000 11086
rect 17960 10804 18012 10810
rect 17960 10746 18012 10752
rect 18156 10742 18184 14991
rect 18248 14618 18276 15302
rect 18616 15065 18644 17070
rect 18696 16992 18748 16998
rect 18696 16934 18748 16940
rect 18708 15201 18736 16934
rect 18788 16652 18840 16658
rect 18788 16594 18840 16600
rect 18800 15881 18828 16594
rect 19076 16590 19104 17138
rect 19168 17105 19196 17711
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19352 17377 19380 17546
rect 19338 17368 19394 17377
rect 19812 17338 19840 17750
rect 19338 17303 19394 17312
rect 19800 17332 19852 17338
rect 19800 17274 19852 17280
rect 19154 17096 19210 17105
rect 19154 17031 19210 17040
rect 19904 16998 19932 19110
rect 20548 18970 20576 20198
rect 20956 20156 21252 20176
rect 21012 20154 21036 20156
rect 21092 20154 21116 20156
rect 21172 20154 21196 20156
rect 21034 20102 21036 20154
rect 21098 20102 21110 20154
rect 21172 20102 21174 20154
rect 21012 20100 21036 20102
rect 21092 20100 21116 20102
rect 21172 20100 21196 20102
rect 20956 20080 21252 20100
rect 20718 19272 20774 19281
rect 20718 19207 20774 19216
rect 20732 19174 20760 19207
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20956 19068 21252 19088
rect 21012 19066 21036 19068
rect 21092 19066 21116 19068
rect 21172 19066 21196 19068
rect 21034 19014 21036 19066
rect 21098 19014 21110 19066
rect 21172 19014 21174 19066
rect 21012 19012 21036 19014
rect 21092 19012 21116 19014
rect 21172 19012 21196 19014
rect 20956 18992 21252 19012
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 20168 18896 20220 18902
rect 20168 18838 20220 18844
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19996 18358 20024 18566
rect 19984 18352 20036 18358
rect 19982 18320 19984 18329
rect 20036 18320 20038 18329
rect 20180 18290 20208 18838
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 19982 18255 20038 18264
rect 20168 18284 20220 18290
rect 19996 18229 20024 18255
rect 20168 18226 20220 18232
rect 20076 17876 20128 17882
rect 20180 17864 20208 18226
rect 20260 18216 20312 18222
rect 20260 18158 20312 18164
rect 20272 17882 20300 18158
rect 20352 18148 20404 18154
rect 20352 18090 20404 18096
rect 20128 17836 20208 17864
rect 20260 17876 20312 17882
rect 20076 17818 20128 17824
rect 20260 17818 20312 17824
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19064 16584 19116 16590
rect 19064 16526 19116 16532
rect 18786 15872 18842 15881
rect 18786 15807 18842 15816
rect 18970 15872 19026 15881
rect 18970 15807 19026 15816
rect 18694 15192 18750 15201
rect 18694 15127 18750 15136
rect 18602 15056 18658 15065
rect 18602 14991 18658 15000
rect 18604 14884 18656 14890
rect 18604 14826 18656 14832
rect 18512 14816 18564 14822
rect 18512 14758 18564 14764
rect 18524 14618 18552 14758
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18248 13802 18276 14554
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18236 13796 18288 13802
rect 18236 13738 18288 13744
rect 18248 13530 18276 13738
rect 18524 13705 18552 14214
rect 18510 13696 18566 13705
rect 18510 13631 18566 13640
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 18340 12782 18368 13126
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 18340 12442 18368 12718
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 18144 10736 18196 10742
rect 18144 10678 18196 10684
rect 17592 10600 17644 10606
rect 17130 10568 17186 10577
rect 17592 10542 17644 10548
rect 18156 10538 18184 10678
rect 17130 10503 17186 10512
rect 18144 10532 18196 10538
rect 17144 10266 17172 10503
rect 18144 10474 18196 10480
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 17144 9722 17172 10202
rect 17222 10160 17278 10169
rect 17222 10095 17278 10104
rect 17406 10160 17462 10169
rect 17406 10095 17408 10104
rect 17236 9761 17264 10095
rect 17460 10095 17462 10104
rect 17408 10066 17460 10072
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17222 9752 17278 9761
rect 17132 9716 17184 9722
rect 17222 9687 17278 9696
rect 17132 9658 17184 9664
rect 16854 9616 16910 9625
rect 17328 9586 17356 9998
rect 16854 9551 16856 9560
rect 16908 9551 16910 9560
rect 17316 9580 17368 9586
rect 16856 9522 16908 9528
rect 17316 9522 17368 9528
rect 17420 9382 17448 10066
rect 18248 10062 18276 10950
rect 18340 10674 18368 12378
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18432 11393 18460 11494
rect 18418 11384 18474 11393
rect 18418 11319 18474 11328
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18340 10266 18368 10610
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17788 9382 17816 9522
rect 18512 9512 18564 9518
rect 18512 9454 18564 9460
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17776 9376 17828 9382
rect 18524 9353 18552 9454
rect 17776 9318 17828 9324
rect 18510 9344 18566 9353
rect 17420 9081 17448 9318
rect 17406 9072 17462 9081
rect 17788 9042 17816 9318
rect 18510 9279 18566 9288
rect 17406 9007 17462 9016
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 17052 7954 17080 8434
rect 17788 8090 17816 8978
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17880 8498 17908 8774
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 18616 8401 18644 14826
rect 18708 10606 18736 15127
rect 18984 14906 19012 15807
rect 19076 15706 19104 16526
rect 19338 16144 19394 16153
rect 19338 16079 19394 16088
rect 19064 15700 19116 15706
rect 19064 15642 19116 15648
rect 19352 15609 19380 16079
rect 19984 15904 20036 15910
rect 19982 15872 19984 15881
rect 20036 15872 20038 15881
rect 19982 15807 20038 15816
rect 19338 15600 19394 15609
rect 19394 15558 19564 15586
rect 19338 15535 19394 15544
rect 19156 15020 19208 15026
rect 19156 14962 19208 14968
rect 19168 14929 19196 14962
rect 19154 14920 19210 14929
rect 18984 14878 19104 14906
rect 18972 14816 19024 14822
rect 18972 14758 19024 14764
rect 18984 14278 19012 14758
rect 18972 14272 19024 14278
rect 18972 14214 19024 14220
rect 18880 11552 18932 11558
rect 18880 11494 18932 11500
rect 18892 11354 18920 11494
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 18708 10198 18736 10542
rect 19076 10198 19104 14878
rect 19154 14855 19210 14864
rect 19168 14550 19196 14855
rect 19156 14544 19208 14550
rect 19156 14486 19208 14492
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19260 13977 19288 14214
rect 19246 13968 19302 13977
rect 19246 13903 19302 13912
rect 19352 13818 19380 14418
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 19444 13841 19472 13942
rect 19260 13790 19380 13818
rect 19430 13832 19486 13841
rect 19260 13530 19288 13790
rect 19430 13767 19486 13776
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19248 12708 19300 12714
rect 19248 12650 19300 12656
rect 19260 12424 19288 12650
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19352 12424 19380 12582
rect 19260 12396 19380 12424
rect 19352 11694 19380 12396
rect 19340 11688 19392 11694
rect 19340 11630 19392 11636
rect 19248 11620 19300 11626
rect 19248 11562 19300 11568
rect 19156 10532 19208 10538
rect 19156 10474 19208 10480
rect 18696 10192 18748 10198
rect 18696 10134 18748 10140
rect 19064 10192 19116 10198
rect 19064 10134 19116 10140
rect 18972 10056 19024 10062
rect 18972 9998 19024 10004
rect 18984 9178 19012 9998
rect 19076 9654 19104 10134
rect 19168 10130 19196 10474
rect 19260 10266 19288 11562
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 19536 10130 19564 15558
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19904 14657 19932 14758
rect 19890 14648 19946 14657
rect 19890 14583 19946 14592
rect 20260 14612 20312 14618
rect 20260 14554 20312 14560
rect 19706 14512 19762 14521
rect 19706 14447 19708 14456
rect 19760 14447 19762 14456
rect 19708 14418 19760 14424
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 20088 14113 20116 14350
rect 20074 14104 20130 14113
rect 20074 14039 20076 14048
rect 20128 14039 20130 14048
rect 20076 14010 20128 14016
rect 19614 13696 19670 13705
rect 19614 13631 19670 13640
rect 19628 13462 19656 13631
rect 20272 13530 20300 14554
rect 20364 14249 20392 18090
rect 20732 18086 20760 18702
rect 21284 18154 21312 20742
rect 21560 20641 21588 23520
rect 21732 20868 21784 20874
rect 21732 20810 21784 20816
rect 21546 20632 21602 20641
rect 21546 20567 21602 20576
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 21272 18148 21324 18154
rect 21272 18090 21324 18096
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20548 14822 20576 15302
rect 20640 15162 20668 15506
rect 20732 15473 20760 18022
rect 20956 17980 21252 18000
rect 21012 17978 21036 17980
rect 21092 17978 21116 17980
rect 21172 17978 21196 17980
rect 21034 17926 21036 17978
rect 21098 17926 21110 17978
rect 21172 17926 21174 17978
rect 21012 17924 21036 17926
rect 21092 17924 21116 17926
rect 21172 17924 21196 17926
rect 20956 17904 21252 17924
rect 21468 17814 21496 18702
rect 21640 18284 21692 18290
rect 21640 18226 21692 18232
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 21456 17808 21508 17814
rect 21456 17750 21508 17756
rect 21272 17740 21324 17746
rect 21272 17682 21324 17688
rect 20812 17128 20864 17134
rect 20812 17070 20864 17076
rect 20824 16998 20852 17070
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20824 16590 20852 16934
rect 20956 16892 21252 16912
rect 21012 16890 21036 16892
rect 21092 16890 21116 16892
rect 21172 16890 21196 16892
rect 21034 16838 21036 16890
rect 21098 16838 21110 16890
rect 21172 16838 21174 16890
rect 21012 16836 21036 16838
rect 21092 16836 21116 16838
rect 21172 16836 21196 16838
rect 20956 16816 21252 16836
rect 21180 16720 21232 16726
rect 21284 16674 21312 17682
rect 21364 17672 21416 17678
rect 21364 17614 21416 17620
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21376 16794 21404 17614
rect 21468 17338 21496 17614
rect 21456 17332 21508 17338
rect 21456 17274 21508 17280
rect 21364 16788 21416 16794
rect 21364 16730 21416 16736
rect 21232 16668 21312 16674
rect 21180 16662 21312 16668
rect 21192 16646 21312 16662
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20824 15910 20852 16526
rect 21284 16250 21312 16646
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20718 15464 20774 15473
rect 20718 15399 20774 15408
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20350 14240 20406 14249
rect 20350 14175 20406 14184
rect 20260 13524 20312 13530
rect 20260 13466 20312 13472
rect 19616 13456 19668 13462
rect 19616 13398 19668 13404
rect 19628 13025 19656 13398
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19800 13320 19852 13326
rect 19800 13262 19852 13268
rect 19614 13016 19670 13025
rect 19720 12986 19748 13262
rect 19614 12951 19670 12960
rect 19708 12980 19760 12986
rect 19628 12442 19656 12951
rect 19708 12922 19760 12928
rect 19720 12889 19748 12922
rect 19706 12880 19762 12889
rect 19706 12815 19762 12824
rect 19812 12442 19840 13262
rect 20076 12912 20128 12918
rect 20076 12854 20128 12860
rect 19892 12708 19944 12714
rect 19892 12650 19944 12656
rect 19616 12436 19668 12442
rect 19616 12378 19668 12384
rect 19800 12436 19852 12442
rect 19800 12378 19852 12384
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 19168 9722 19196 10066
rect 19156 9716 19208 9722
rect 19156 9658 19208 9664
rect 19064 9648 19116 9654
rect 19064 9590 19116 9596
rect 18972 9172 19024 9178
rect 18972 9114 19024 9120
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18800 8430 18828 8774
rect 18788 8424 18840 8430
rect 18602 8392 18658 8401
rect 18788 8366 18840 8372
rect 18602 8327 18658 8336
rect 17868 8288 17920 8294
rect 17868 8230 17920 8236
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 17776 8084 17828 8090
rect 17776 8026 17828 8032
rect 17040 7948 17092 7954
rect 17040 7890 17092 7896
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16868 6934 16896 7278
rect 17052 7002 17080 7890
rect 17788 7478 17816 8026
rect 17776 7472 17828 7478
rect 17776 7414 17828 7420
rect 17880 7342 17908 8230
rect 18432 7818 18460 8230
rect 19168 8090 19196 9658
rect 19248 9376 19300 9382
rect 19352 9364 19380 10066
rect 19300 9336 19380 9364
rect 19248 9318 19300 9324
rect 19260 8673 19288 9318
rect 19524 9036 19576 9042
rect 19524 8978 19576 8984
rect 19340 8832 19392 8838
rect 19536 8809 19564 8978
rect 19340 8774 19392 8780
rect 19522 8800 19578 8809
rect 19246 8664 19302 8673
rect 19246 8599 19302 8608
rect 19246 8392 19302 8401
rect 19246 8327 19302 8336
rect 19156 8084 19208 8090
rect 19156 8026 19208 8032
rect 19064 7880 19116 7886
rect 19062 7848 19064 7857
rect 19116 7848 19118 7857
rect 18420 7812 18472 7818
rect 19062 7783 19118 7792
rect 18420 7754 18472 7760
rect 18432 7546 18460 7754
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18708 7410 18736 7686
rect 19168 7410 19196 8026
rect 19260 8022 19288 8327
rect 19352 8090 19380 8774
rect 19522 8735 19578 8744
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19248 8016 19300 8022
rect 19248 7958 19300 7964
rect 19260 7546 19288 7958
rect 19444 7546 19472 8366
rect 19536 7857 19564 8735
rect 19522 7848 19578 7857
rect 19522 7783 19578 7792
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 17040 6996 17092 7002
rect 17040 6938 17092 6944
rect 16856 6928 16908 6934
rect 16856 6870 16908 6876
rect 16762 6352 16818 6361
rect 16762 6287 16818 6296
rect 15956 5468 16252 5488
rect 16012 5466 16036 5468
rect 16092 5466 16116 5468
rect 16172 5466 16196 5468
rect 16034 5414 16036 5466
rect 16098 5414 16110 5466
rect 16172 5414 16174 5466
rect 16012 5412 16036 5414
rect 16092 5412 16116 5414
rect 16172 5412 16196 5414
rect 15956 5392 16252 5412
rect 15956 4380 16252 4400
rect 16012 4378 16036 4380
rect 16092 4378 16116 4380
rect 16172 4378 16196 4380
rect 16034 4326 16036 4378
rect 16098 4326 16110 4378
rect 16172 4326 16174 4378
rect 16012 4324 16036 4326
rect 16092 4324 16116 4326
rect 16172 4324 16196 4326
rect 15956 4304 16252 4324
rect 15566 3496 15622 3505
rect 15566 3431 15622 3440
rect 15956 3292 16252 3312
rect 16012 3290 16036 3292
rect 16092 3290 16116 3292
rect 16172 3290 16196 3292
rect 16034 3238 16036 3290
rect 16098 3238 16110 3290
rect 16172 3238 16174 3290
rect 16012 3236 16036 3238
rect 16092 3236 16116 3238
rect 16172 3236 16196 3238
rect 15956 3216 16252 3236
rect 10956 2748 11252 2768
rect 11012 2746 11036 2748
rect 11092 2746 11116 2748
rect 11172 2746 11196 2748
rect 11034 2694 11036 2746
rect 11098 2694 11110 2746
rect 11172 2694 11174 2746
rect 11012 2692 11036 2694
rect 11092 2692 11116 2694
rect 11172 2692 11196 2694
rect 10956 2672 11252 2692
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 6564 2446 6592 2586
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 6552 2440 6604 2446
rect 7484 2417 7512 2450
rect 6552 2382 6604 2388
rect 7470 2408 7526 2417
rect 7470 2343 7526 2352
rect 11150 2408 11206 2417
rect 11150 2343 11206 2352
rect 5956 2204 6252 2224
rect 6012 2202 6036 2204
rect 6092 2202 6116 2204
rect 6172 2202 6196 2204
rect 6034 2150 6036 2202
rect 6098 2150 6110 2202
rect 6172 2150 6174 2202
rect 6012 2148 6036 2150
rect 6092 2148 6116 2150
rect 6172 2148 6196 2150
rect 5956 2128 6252 2148
rect 11164 480 11192 2343
rect 15956 2204 16252 2224
rect 16012 2202 16036 2204
rect 16092 2202 16116 2204
rect 16172 2202 16196 2204
rect 16034 2150 16036 2202
rect 16098 2150 16110 2202
rect 16172 2150 16174 2202
rect 16012 2148 16036 2150
rect 16092 2148 16116 2150
rect 16172 2148 16196 2150
rect 15956 2128 16252 2148
rect 18708 480 18736 7346
rect 19260 7313 19288 7482
rect 19432 7336 19484 7342
rect 19246 7304 19302 7313
rect 19432 7278 19484 7284
rect 19246 7239 19302 7248
rect 19444 7002 19472 7278
rect 19628 7274 19656 12378
rect 19904 11898 19932 12650
rect 20088 12084 20116 12854
rect 20168 12096 20220 12102
rect 20088 12056 20168 12084
rect 20168 12038 20220 12044
rect 19892 11892 19944 11898
rect 19892 11834 19944 11840
rect 19800 11756 19852 11762
rect 19904 11744 19932 11834
rect 19852 11716 19932 11744
rect 19800 11698 19852 11704
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19720 10606 19748 11494
rect 19812 11150 19840 11698
rect 20180 11626 20208 12038
rect 20168 11620 20220 11626
rect 20168 11562 20220 11568
rect 19800 11144 19852 11150
rect 19800 11086 19852 11092
rect 19812 10810 19840 11086
rect 20074 10976 20130 10985
rect 20074 10911 20130 10920
rect 19800 10804 19852 10810
rect 19800 10746 19852 10752
rect 20088 10606 20116 10911
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 19720 10470 19748 10542
rect 19708 10464 19760 10470
rect 19708 10406 19760 10412
rect 19720 9450 19748 10406
rect 20088 10266 20116 10542
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 20180 10062 20208 11562
rect 20364 10198 20392 14175
rect 20456 10849 20484 14758
rect 20548 13433 20576 14758
rect 20640 14618 20668 15098
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20626 13560 20682 13569
rect 20732 13530 20760 15302
rect 20824 14414 20852 15846
rect 20956 15804 21252 15824
rect 21012 15802 21036 15804
rect 21092 15802 21116 15804
rect 21172 15802 21196 15804
rect 21034 15750 21036 15802
rect 21098 15750 21110 15802
rect 21172 15750 21174 15802
rect 21012 15748 21036 15750
rect 21092 15748 21116 15750
rect 21172 15748 21196 15750
rect 20956 15728 21252 15748
rect 21376 15706 21404 16730
rect 21454 16280 21510 16289
rect 21454 16215 21510 16224
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 21362 15464 21418 15473
rect 21362 15399 21418 15408
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 20956 14716 21252 14736
rect 21012 14714 21036 14716
rect 21092 14714 21116 14716
rect 21172 14714 21196 14716
rect 21034 14662 21036 14714
rect 21098 14662 21110 14714
rect 21172 14662 21174 14714
rect 21012 14660 21036 14662
rect 21092 14660 21116 14662
rect 21172 14660 21196 14662
rect 20956 14640 21252 14660
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 21088 14272 21140 14278
rect 21088 14214 21140 14220
rect 21100 13870 21128 14214
rect 21088 13864 21140 13870
rect 21088 13806 21140 13812
rect 20812 13728 20864 13734
rect 20812 13670 20864 13676
rect 20626 13495 20682 13504
rect 20720 13524 20772 13530
rect 20534 13424 20590 13433
rect 20640 13410 20668 13495
rect 20720 13466 20772 13472
rect 20640 13382 20760 13410
rect 20534 13359 20590 13368
rect 20732 13161 20760 13382
rect 20718 13152 20774 13161
rect 20718 13087 20774 13096
rect 20824 13002 20852 13670
rect 20956 13628 21252 13648
rect 21012 13626 21036 13628
rect 21092 13626 21116 13628
rect 21172 13626 21196 13628
rect 21034 13574 21036 13626
rect 21098 13574 21110 13626
rect 21172 13574 21174 13626
rect 21012 13572 21036 13574
rect 21092 13572 21116 13574
rect 21172 13572 21196 13574
rect 20956 13552 21252 13572
rect 20904 13456 20956 13462
rect 20904 13398 20956 13404
rect 20732 12974 20852 13002
rect 20732 12782 20760 12974
rect 20916 12866 20944 13398
rect 20824 12838 20944 12866
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 20824 11506 20852 12838
rect 21284 12696 21312 14758
rect 21376 14074 21404 15399
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 21468 13682 21496 16215
rect 21560 16114 21588 18022
rect 21652 16658 21680 18226
rect 21640 16652 21692 16658
rect 21640 16594 21692 16600
rect 21652 16182 21680 16594
rect 21640 16176 21692 16182
rect 21640 16118 21692 16124
rect 21548 16108 21600 16114
rect 21548 16050 21600 16056
rect 21652 15706 21680 16118
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 21652 15026 21680 15642
rect 21640 15020 21692 15026
rect 21640 14962 21692 14968
rect 21652 14634 21680 14962
rect 21744 14822 21772 20810
rect 21824 20256 21876 20262
rect 21824 20198 21876 20204
rect 21732 14816 21784 14822
rect 21732 14758 21784 14764
rect 21652 14606 21772 14634
rect 21376 13654 21496 13682
rect 21376 13462 21404 13654
rect 21454 13560 21510 13569
rect 21454 13495 21510 13504
rect 21364 13456 21416 13462
rect 21364 13398 21416 13404
rect 21468 12753 21496 13495
rect 21744 13326 21772 14606
rect 21640 13320 21692 13326
rect 21640 13262 21692 13268
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21546 13152 21602 13161
rect 21546 13087 21602 13096
rect 21454 12744 21510 12753
rect 21284 12668 21373 12696
rect 21454 12679 21510 12688
rect 21345 12594 21373 12668
rect 21284 12566 21373 12594
rect 20956 12540 21252 12560
rect 21012 12538 21036 12540
rect 21092 12538 21116 12540
rect 21172 12538 21196 12540
rect 21034 12486 21036 12538
rect 21098 12486 21110 12538
rect 21172 12486 21174 12538
rect 21012 12484 21036 12486
rect 21092 12484 21116 12486
rect 21172 12484 21196 12486
rect 20956 12464 21252 12484
rect 20994 12336 21050 12345
rect 20994 12271 21050 12280
rect 21008 11830 21036 12271
rect 20996 11824 21048 11830
rect 20996 11766 21048 11772
rect 20732 11478 20852 11506
rect 20628 11076 20680 11082
rect 20628 11018 20680 11024
rect 20442 10840 20498 10849
rect 20442 10775 20498 10784
rect 20640 10266 20668 11018
rect 20628 10260 20680 10266
rect 20628 10202 20680 10208
rect 20352 10192 20404 10198
rect 20352 10134 20404 10140
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 19892 9512 19944 9518
rect 19892 9454 19944 9460
rect 19708 9444 19760 9450
rect 19708 9386 19760 9392
rect 19904 8974 19932 9454
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19720 8537 19748 8910
rect 20076 8832 20128 8838
rect 20076 8774 20128 8780
rect 19706 8528 19762 8537
rect 20088 8498 20116 8774
rect 20272 8498 20300 9318
rect 20732 9178 20760 11478
rect 20956 11452 21252 11472
rect 21012 11450 21036 11452
rect 21092 11450 21116 11452
rect 21172 11450 21196 11452
rect 21034 11398 21036 11450
rect 21098 11398 21110 11450
rect 21172 11398 21174 11450
rect 21012 11396 21036 11398
rect 21092 11396 21116 11398
rect 21172 11396 21196 11398
rect 20810 11384 20866 11393
rect 20956 11376 21252 11396
rect 20810 11319 20866 11328
rect 20824 11286 20852 11319
rect 20812 11280 20864 11286
rect 20812 11222 20864 11228
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20824 8906 20852 11086
rect 20956 10364 21252 10384
rect 21012 10362 21036 10364
rect 21092 10362 21116 10364
rect 21172 10362 21196 10364
rect 21034 10310 21036 10362
rect 21098 10310 21110 10362
rect 21172 10310 21174 10362
rect 21012 10308 21036 10310
rect 21092 10308 21116 10310
rect 21172 10308 21196 10310
rect 20956 10288 21252 10308
rect 21180 10192 21232 10198
rect 21180 10134 21232 10140
rect 21192 9722 21220 10134
rect 21180 9716 21232 9722
rect 21180 9658 21232 9664
rect 21284 9625 21312 12566
rect 21560 12481 21588 13087
rect 21546 12472 21602 12481
rect 21546 12407 21602 12416
rect 21560 12374 21588 12407
rect 21548 12368 21600 12374
rect 21548 12310 21600 12316
rect 21560 11898 21588 12310
rect 21652 12170 21680 13262
rect 21744 12442 21772 13262
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21640 12164 21692 12170
rect 21640 12106 21692 12112
rect 21548 11892 21600 11898
rect 21600 11852 21680 11880
rect 21548 11834 21600 11840
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21270 9616 21326 9625
rect 21270 9551 21326 9560
rect 20956 9276 21252 9296
rect 21012 9274 21036 9276
rect 21092 9274 21116 9276
rect 21172 9274 21196 9276
rect 21034 9222 21036 9274
rect 21098 9222 21110 9274
rect 21172 9222 21174 9274
rect 21012 9220 21036 9222
rect 21092 9220 21116 9222
rect 21172 9220 21196 9222
rect 20956 9200 21252 9220
rect 20812 8900 20864 8906
rect 20812 8842 20864 8848
rect 19706 8463 19708 8472
rect 19760 8463 19762 8472
rect 19892 8492 19944 8498
rect 19708 8434 19760 8440
rect 19892 8434 19944 8440
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 20260 8492 20312 8498
rect 20260 8434 20312 8440
rect 19720 8403 19748 8434
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 19812 7478 19840 7822
rect 19800 7472 19852 7478
rect 19800 7414 19852 7420
rect 19708 7404 19760 7410
rect 19708 7346 19760 7352
rect 19616 7268 19668 7274
rect 19616 7210 19668 7216
rect 19720 7002 19748 7346
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19708 6996 19760 7002
rect 19708 6938 19760 6944
rect 19904 4049 19932 8434
rect 20272 8022 20300 8434
rect 21376 8430 21404 11698
rect 21454 9616 21510 9625
rect 21454 9551 21510 9560
rect 21468 9110 21496 9551
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 21456 9104 21508 9110
rect 21456 9046 21508 9052
rect 21468 8634 21496 9046
rect 21456 8628 21508 8634
rect 21456 8570 21508 8576
rect 21364 8424 21416 8430
rect 21364 8366 21416 8372
rect 20956 8188 21252 8208
rect 21012 8186 21036 8188
rect 21092 8186 21116 8188
rect 21172 8186 21196 8188
rect 21034 8134 21036 8186
rect 21098 8134 21110 8186
rect 21172 8134 21174 8186
rect 21012 8132 21036 8134
rect 21092 8132 21116 8134
rect 21172 8132 21196 8134
rect 20956 8112 21252 8132
rect 21376 8090 21404 8366
rect 21560 8090 21588 9114
rect 21652 8566 21680 11852
rect 21836 11082 21864 20198
rect 21914 19272 21970 19281
rect 21914 19207 21970 19216
rect 21928 18086 21956 19207
rect 23400 18970 23428 23520
rect 24032 21004 24084 21010
rect 24032 20946 24084 20952
rect 23388 18964 23440 18970
rect 23388 18906 23440 18912
rect 22468 18828 22520 18834
rect 22468 18770 22520 18776
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 22112 18290 22140 18566
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22008 18216 22060 18222
rect 22008 18158 22060 18164
rect 21916 18080 21968 18086
rect 21916 18022 21968 18028
rect 21928 17542 21956 18022
rect 21916 17536 21968 17542
rect 21914 17504 21916 17513
rect 21968 17504 21970 17513
rect 21914 17439 21970 17448
rect 21916 17060 21968 17066
rect 21916 17002 21968 17008
rect 21928 16182 21956 17002
rect 22020 16810 22048 18158
rect 22480 18154 22508 18770
rect 22652 18760 22704 18766
rect 22652 18702 22704 18708
rect 23846 18728 23902 18737
rect 22100 18148 22152 18154
rect 22100 18090 22152 18096
rect 22468 18148 22520 18154
rect 22468 18090 22520 18096
rect 22112 17882 22140 18090
rect 22664 18086 22692 18702
rect 23846 18663 23902 18672
rect 23110 18184 23166 18193
rect 23110 18119 23166 18128
rect 22652 18080 22704 18086
rect 22652 18022 22704 18028
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 22468 17808 22520 17814
rect 22468 17750 22520 17756
rect 22376 17672 22428 17678
rect 22376 17614 22428 17620
rect 22100 17604 22152 17610
rect 22100 17546 22152 17552
rect 22112 17105 22140 17546
rect 22388 17134 22416 17614
rect 22480 17338 22508 17750
rect 22664 17649 22692 18022
rect 22650 17640 22706 17649
rect 22650 17575 22706 17584
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 22376 17128 22428 17134
rect 22098 17096 22154 17105
rect 22376 17070 22428 17076
rect 22098 17031 22154 17040
rect 22480 16998 22508 17274
rect 22468 16992 22520 16998
rect 22468 16934 22520 16940
rect 22020 16782 22232 16810
rect 22480 16794 22508 16934
rect 22006 16688 22062 16697
rect 22006 16623 22062 16632
rect 21916 16176 21968 16182
rect 21916 16118 21968 16124
rect 21928 15910 21956 16118
rect 21916 15904 21968 15910
rect 21916 15846 21968 15852
rect 21928 15502 21956 15846
rect 21916 15496 21968 15502
rect 21916 15438 21968 15444
rect 21928 14618 21956 15438
rect 22020 14958 22048 16623
rect 22204 16130 22232 16782
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22560 16448 22612 16454
rect 22560 16390 22612 16396
rect 22204 16102 22508 16130
rect 22192 15972 22244 15978
rect 22192 15914 22244 15920
rect 22204 15162 22232 15914
rect 22192 15156 22244 15162
rect 22192 15098 22244 15104
rect 22008 14952 22060 14958
rect 22008 14894 22060 14900
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 22192 14476 22244 14482
rect 22192 14418 22244 14424
rect 22008 14068 22060 14074
rect 22008 14010 22060 14016
rect 21916 12980 21968 12986
rect 21916 12922 21968 12928
rect 21928 11150 21956 12922
rect 22020 12209 22048 14010
rect 22100 13796 22152 13802
rect 22100 13738 22152 13744
rect 22112 12986 22140 13738
rect 22204 13734 22232 14418
rect 22192 13728 22244 13734
rect 22192 13670 22244 13676
rect 22204 13190 22232 13670
rect 22192 13184 22244 13190
rect 22192 13126 22244 13132
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 22204 12306 22232 13126
rect 22192 12300 22244 12306
rect 22192 12242 22244 12248
rect 22006 12200 22062 12209
rect 22006 12135 22062 12144
rect 22204 11506 22232 12242
rect 22204 11478 22324 11506
rect 22192 11348 22244 11354
rect 22192 11290 22244 11296
rect 22008 11280 22060 11286
rect 22008 11222 22060 11228
rect 21916 11144 21968 11150
rect 21916 11086 21968 11092
rect 21824 11076 21876 11082
rect 21824 11018 21876 11024
rect 21928 10810 21956 11086
rect 22020 10810 22048 11222
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 21916 10804 21968 10810
rect 21916 10746 21968 10752
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 22008 10260 22060 10266
rect 22112 10248 22140 11086
rect 22204 10810 22232 11290
rect 22296 11082 22324 11478
rect 22284 11076 22336 11082
rect 22284 11018 22336 11024
rect 22192 10804 22244 10810
rect 22192 10746 22244 10752
rect 22060 10220 22140 10248
rect 22008 10202 22060 10208
rect 21824 10056 21876 10062
rect 21824 9998 21876 10004
rect 21836 8974 21864 9998
rect 22020 9722 22048 10202
rect 22480 10169 22508 16102
rect 22572 15910 22600 16390
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22664 13297 22692 17575
rect 22926 15192 22982 15201
rect 22926 15127 22982 15136
rect 22836 15020 22888 15026
rect 22836 14962 22888 14968
rect 22848 14618 22876 14962
rect 22940 14822 22968 15127
rect 22928 14816 22980 14822
rect 22928 14758 22980 14764
rect 22836 14612 22888 14618
rect 22836 14554 22888 14560
rect 22940 13841 22968 14758
rect 22926 13832 22982 13841
rect 22926 13767 22982 13776
rect 22744 13524 22796 13530
rect 22744 13466 22796 13472
rect 22756 13433 22784 13466
rect 22742 13424 22798 13433
rect 22742 13359 22798 13368
rect 22650 13288 22706 13297
rect 22650 13223 22706 13232
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 22744 12436 22796 12442
rect 22744 12378 22796 12384
rect 22756 12345 22784 12378
rect 22742 12336 22798 12345
rect 22742 12271 22798 12280
rect 22756 11830 22784 12271
rect 23032 12073 23060 12922
rect 23124 12866 23152 18119
rect 23570 16688 23626 16697
rect 23570 16623 23572 16632
rect 23624 16623 23626 16632
rect 23572 16594 23624 16600
rect 23480 16448 23532 16454
rect 23480 16390 23532 16396
rect 23492 16046 23520 16390
rect 23480 16040 23532 16046
rect 23386 16008 23442 16017
rect 23204 15972 23256 15978
rect 23480 15982 23532 15988
rect 23386 15943 23442 15952
rect 23204 15914 23256 15920
rect 23216 15706 23244 15914
rect 23204 15700 23256 15706
rect 23204 15642 23256 15648
rect 23202 15056 23258 15065
rect 23202 14991 23204 15000
rect 23256 14991 23258 15000
rect 23204 14962 23256 14968
rect 23202 13560 23258 13569
rect 23202 13495 23204 13504
rect 23256 13495 23258 13504
rect 23204 13466 23256 13472
rect 23216 13410 23244 13466
rect 23216 13382 23336 13410
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 23216 12986 23244 13262
rect 23204 12980 23256 12986
rect 23204 12922 23256 12928
rect 23124 12850 23244 12866
rect 23124 12844 23256 12850
rect 23124 12838 23204 12844
rect 23204 12786 23256 12792
rect 23112 12776 23164 12782
rect 23112 12718 23164 12724
rect 23124 12442 23152 12718
rect 23112 12436 23164 12442
rect 23112 12378 23164 12384
rect 23018 12064 23074 12073
rect 23018 11999 23074 12008
rect 23216 11898 23244 12786
rect 23308 12782 23336 13382
rect 23400 13258 23428 15943
rect 23572 15564 23624 15570
rect 23572 15506 23624 15512
rect 23480 15428 23532 15434
rect 23480 15370 23532 15376
rect 23492 14618 23520 15370
rect 23584 14890 23612 15506
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23676 15065 23704 15438
rect 23662 15056 23718 15065
rect 23662 14991 23718 15000
rect 23754 14920 23810 14929
rect 23572 14884 23624 14890
rect 23754 14855 23810 14864
rect 23572 14826 23624 14832
rect 23768 14618 23796 14855
rect 23480 14612 23532 14618
rect 23480 14554 23532 14560
rect 23756 14612 23808 14618
rect 23756 14554 23808 14560
rect 23860 14498 23888 18663
rect 23938 16552 23994 16561
rect 23938 16487 23994 16496
rect 23480 14476 23532 14482
rect 23480 14418 23532 14424
rect 23768 14470 23888 14498
rect 23492 14113 23520 14418
rect 23478 14104 23534 14113
rect 23478 14039 23480 14048
rect 23532 14039 23534 14048
rect 23480 14010 23532 14016
rect 23492 13938 23520 14010
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23492 13530 23520 13874
rect 23480 13524 23532 13530
rect 23480 13466 23532 13472
rect 23768 13394 23796 14470
rect 23848 14408 23900 14414
rect 23848 14350 23900 14356
rect 23860 13734 23888 14350
rect 23848 13728 23900 13734
rect 23848 13670 23900 13676
rect 23756 13388 23808 13394
rect 23756 13330 23808 13336
rect 23388 13252 23440 13258
rect 23388 13194 23440 13200
rect 23768 12918 23796 13330
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 23296 12776 23348 12782
rect 23296 12718 23348 12724
rect 23480 12708 23532 12714
rect 23480 12650 23532 12656
rect 23492 12424 23520 12650
rect 23756 12640 23808 12646
rect 23756 12582 23808 12588
rect 23308 12396 23520 12424
rect 23204 11892 23256 11898
rect 23204 11834 23256 11840
rect 22744 11824 22796 11830
rect 22744 11766 22796 11772
rect 22650 11656 22706 11665
rect 22650 11591 22706 11600
rect 22664 11558 22692 11591
rect 22652 11552 22704 11558
rect 22652 11494 22704 11500
rect 23308 11370 23336 12396
rect 23480 12300 23532 12306
rect 23480 12242 23532 12248
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 23400 11626 23428 12174
rect 23388 11620 23440 11626
rect 23388 11562 23440 11568
rect 23124 11342 23336 11370
rect 22466 10160 22522 10169
rect 22466 10095 22522 10104
rect 23124 10062 23152 11342
rect 23296 11212 23348 11218
rect 23296 11154 23348 11160
rect 23202 10840 23258 10849
rect 23202 10775 23258 10784
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 22008 9716 22060 9722
rect 22008 9658 22060 9664
rect 22100 9376 22152 9382
rect 22100 9318 22152 9324
rect 22112 8974 22140 9318
rect 23216 9217 23244 10775
rect 23308 10198 23336 11154
rect 23400 10810 23428 11562
rect 23492 11354 23520 12242
rect 23768 11354 23796 12582
rect 23860 12374 23888 13670
rect 23848 12368 23900 12374
rect 23848 12310 23900 12316
rect 23848 11552 23900 11558
rect 23848 11494 23900 11500
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23756 11348 23808 11354
rect 23756 11290 23808 11296
rect 23388 10804 23440 10810
rect 23388 10746 23440 10752
rect 23400 10606 23428 10746
rect 23388 10600 23440 10606
rect 23388 10542 23440 10548
rect 23768 10266 23796 11290
rect 23860 10985 23888 11494
rect 23846 10976 23902 10985
rect 23846 10911 23902 10920
rect 23952 10849 23980 16487
rect 24044 11898 24072 20946
rect 24768 20256 24820 20262
rect 24820 20216 24900 20244
rect 24768 20198 24820 20204
rect 24308 19168 24360 19174
rect 24308 19110 24360 19116
rect 24320 18086 24348 19110
rect 24872 18970 24900 20216
rect 24860 18964 24912 18970
rect 24860 18906 24912 18912
rect 25056 18329 25084 23559
rect 25226 23520 25282 24000
rect 27158 23520 27214 24000
rect 28998 23520 29054 24000
rect 25240 20602 25268 23520
rect 25594 23080 25650 23089
rect 25594 23015 25650 23024
rect 25608 20618 25636 23015
rect 25870 22400 25926 22409
rect 25870 22335 25926 22344
rect 25686 21584 25742 21593
rect 25686 21519 25742 21528
rect 25700 20874 25728 21519
rect 25778 21312 25834 21321
rect 25778 21247 25834 21256
rect 25688 20868 25740 20874
rect 25688 20810 25740 20816
rect 25792 20806 25820 21247
rect 25780 20800 25832 20806
rect 25780 20742 25832 20748
rect 25228 20596 25280 20602
rect 25228 20538 25280 20544
rect 25332 20590 25636 20618
rect 25226 19952 25282 19961
rect 25226 19887 25282 19896
rect 24490 18320 24546 18329
rect 24490 18255 24546 18264
rect 25042 18320 25098 18329
rect 25042 18255 25098 18264
rect 24308 18080 24360 18086
rect 24308 18022 24360 18028
rect 24214 17912 24270 17921
rect 24214 17847 24270 17856
rect 24124 17536 24176 17542
rect 24124 17478 24176 17484
rect 24136 17066 24164 17478
rect 24124 17060 24176 17066
rect 24124 17002 24176 17008
rect 24136 16522 24164 17002
rect 24124 16516 24176 16522
rect 24124 16458 24176 16464
rect 24228 16402 24256 17847
rect 24320 17134 24348 18022
rect 24308 17128 24360 17134
rect 24308 17070 24360 17076
rect 24136 16374 24256 16402
rect 24032 11892 24084 11898
rect 24032 11834 24084 11840
rect 23938 10840 23994 10849
rect 23938 10775 23994 10784
rect 24136 10713 24164 16374
rect 24308 15360 24360 15366
rect 24308 15302 24360 15308
rect 24320 14958 24348 15302
rect 24308 14952 24360 14958
rect 24308 14894 24360 14900
rect 24398 14920 24454 14929
rect 24214 14376 24270 14385
rect 24214 14311 24270 14320
rect 24228 14074 24256 14311
rect 24320 14278 24348 14894
rect 24398 14855 24400 14864
rect 24452 14855 24454 14864
rect 24400 14826 24452 14832
rect 24308 14272 24360 14278
rect 24308 14214 24360 14220
rect 24216 14068 24268 14074
rect 24216 14010 24268 14016
rect 24504 13530 24532 18255
rect 24676 18148 24728 18154
rect 24676 18090 24728 18096
rect 24688 17542 24716 18090
rect 24860 17672 24912 17678
rect 24860 17614 24912 17620
rect 24676 17536 24728 17542
rect 24676 17478 24728 17484
rect 24688 17270 24716 17478
rect 24676 17264 24728 17270
rect 24582 17232 24638 17241
rect 24676 17206 24728 17212
rect 24582 17167 24638 17176
rect 24596 16250 24624 17167
rect 24688 16794 24716 17206
rect 24872 16794 24900 17614
rect 24676 16788 24728 16794
rect 24676 16730 24728 16736
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 24688 16590 24716 16730
rect 25240 16726 25268 19887
rect 25332 18601 25360 20590
rect 25412 20528 25464 20534
rect 25410 20496 25412 20505
rect 25464 20496 25466 20505
rect 25410 20431 25466 20440
rect 25884 20346 25912 22335
rect 25956 21788 26252 21808
rect 26012 21786 26036 21788
rect 26092 21786 26116 21788
rect 26172 21786 26196 21788
rect 26034 21734 26036 21786
rect 26098 21734 26110 21786
rect 26172 21734 26174 21786
rect 26012 21732 26036 21734
rect 26092 21732 26116 21734
rect 26172 21732 26196 21734
rect 25956 21712 26252 21732
rect 26884 21004 26936 21010
rect 26884 20946 26936 20952
rect 25956 20700 26252 20720
rect 26012 20698 26036 20700
rect 26092 20698 26116 20700
rect 26172 20698 26196 20700
rect 26034 20646 26036 20698
rect 26098 20646 26110 20698
rect 26172 20646 26174 20698
rect 26012 20644 26036 20646
rect 26092 20644 26116 20646
rect 26172 20644 26196 20646
rect 25956 20624 26252 20644
rect 26896 20602 26924 20946
rect 26884 20596 26936 20602
rect 26884 20538 26936 20544
rect 27172 20505 27200 23520
rect 29012 21146 29040 23520
rect 29000 21140 29052 21146
rect 29000 21082 29052 21088
rect 27158 20496 27214 20505
rect 27158 20431 27214 20440
rect 25608 20318 25912 20346
rect 25412 19712 25464 19718
rect 25412 19654 25464 19660
rect 25424 19310 25452 19654
rect 25412 19304 25464 19310
rect 25412 19246 25464 19252
rect 25412 19168 25464 19174
rect 25412 19110 25464 19116
rect 25424 18766 25452 19110
rect 25504 18828 25556 18834
rect 25504 18770 25556 18776
rect 25412 18760 25464 18766
rect 25412 18702 25464 18708
rect 25318 18592 25374 18601
rect 25318 18527 25374 18536
rect 25332 17762 25360 18527
rect 25424 17882 25452 18702
rect 25516 18426 25544 18770
rect 25504 18420 25556 18426
rect 25504 18362 25556 18368
rect 25502 18320 25558 18329
rect 25502 18255 25558 18264
rect 25412 17876 25464 17882
rect 25412 17818 25464 17824
rect 25332 17734 25452 17762
rect 25320 17536 25372 17542
rect 25320 17478 25372 17484
rect 25332 16794 25360 17478
rect 25320 16788 25372 16794
rect 25320 16730 25372 16736
rect 25228 16720 25280 16726
rect 25228 16662 25280 16668
rect 24676 16584 24728 16590
rect 24676 16526 24728 16532
rect 24584 16244 24636 16250
rect 24584 16186 24636 16192
rect 24688 16182 24716 16526
rect 25240 16250 25268 16662
rect 25228 16244 25280 16250
rect 25228 16186 25280 16192
rect 24676 16176 24728 16182
rect 24676 16118 24728 16124
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24780 15706 24808 15982
rect 24950 15736 25006 15745
rect 24768 15700 24820 15706
rect 24950 15671 25006 15680
rect 24768 15642 24820 15648
rect 24674 15600 24730 15609
rect 24674 15535 24676 15544
rect 24728 15535 24730 15544
rect 24676 15506 24728 15512
rect 24858 15464 24914 15473
rect 24858 15399 24914 15408
rect 24766 15056 24822 15065
rect 24766 14991 24822 15000
rect 24676 13864 24728 13870
rect 24674 13832 24676 13841
rect 24728 13832 24730 13841
rect 24674 13767 24730 13776
rect 24584 13728 24636 13734
rect 24584 13670 24636 13676
rect 24492 13524 24544 13530
rect 24492 13466 24544 13472
rect 24308 13184 24360 13190
rect 24308 13126 24360 13132
rect 24320 11218 24348 13126
rect 24504 12986 24532 13466
rect 24596 13462 24624 13670
rect 24584 13456 24636 13462
rect 24584 13398 24636 13404
rect 24492 12980 24544 12986
rect 24492 12922 24544 12928
rect 24400 12844 24452 12850
rect 24400 12786 24452 12792
rect 24412 12306 24440 12786
rect 24596 12617 24624 13398
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24688 12714 24716 13330
rect 24780 12918 24808 14991
rect 24768 12912 24820 12918
rect 24768 12854 24820 12860
rect 24676 12708 24728 12714
rect 24676 12650 24728 12656
rect 24582 12608 24638 12617
rect 24582 12543 24638 12552
rect 24400 12300 24452 12306
rect 24400 12242 24452 12248
rect 24582 12200 24638 12209
rect 24582 12135 24638 12144
rect 24308 11212 24360 11218
rect 24308 11154 24360 11160
rect 24216 11144 24268 11150
rect 24216 11086 24268 11092
rect 24122 10704 24178 10713
rect 24122 10639 24178 10648
rect 23940 10600 23992 10606
rect 23940 10542 23992 10548
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 23296 10192 23348 10198
rect 23296 10134 23348 10140
rect 23952 10130 23980 10542
rect 24136 10130 24164 10639
rect 24228 10606 24256 11086
rect 24216 10600 24268 10606
rect 24216 10542 24268 10548
rect 24398 10432 24454 10441
rect 24398 10367 24454 10376
rect 24412 10266 24440 10367
rect 24400 10260 24452 10266
rect 24400 10202 24452 10208
rect 23940 10124 23992 10130
rect 23940 10066 23992 10072
rect 24124 10124 24176 10130
rect 24124 10066 24176 10072
rect 24136 9722 24164 10066
rect 24124 9716 24176 9722
rect 24124 9658 24176 9664
rect 24596 9625 24624 12135
rect 24676 11824 24728 11830
rect 24872 11801 24900 15399
rect 24964 13569 24992 15671
rect 25424 15609 25452 17734
rect 25410 15600 25466 15609
rect 25410 15535 25466 15544
rect 25228 15496 25280 15502
rect 25148 15456 25228 15484
rect 25148 14822 25176 15456
rect 25228 15438 25280 15444
rect 25320 15428 25372 15434
rect 25320 15370 25372 15376
rect 25136 14816 25188 14822
rect 25136 14758 25188 14764
rect 25042 14648 25098 14657
rect 25042 14583 25098 14592
rect 24950 13560 25006 13569
rect 24950 13495 25006 13504
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 24676 11766 24728 11772
rect 24858 11792 24914 11801
rect 24688 11354 24716 11766
rect 24964 11762 24992 12038
rect 24858 11727 24914 11736
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24768 11688 24820 11694
rect 24964 11642 24992 11698
rect 24768 11630 24820 11636
rect 24676 11348 24728 11354
rect 24676 11290 24728 11296
rect 24780 10792 24808 11630
rect 24872 11614 24992 11642
rect 24872 11150 24900 11614
rect 24952 11552 25004 11558
rect 24952 11494 25004 11500
rect 24964 11354 24992 11494
rect 24952 11348 25004 11354
rect 24952 11290 25004 11296
rect 24860 11144 24912 11150
rect 24860 11086 24912 11092
rect 24950 10976 25006 10985
rect 24950 10911 25006 10920
rect 24860 10804 24912 10810
rect 24780 10764 24860 10792
rect 24860 10746 24912 10752
rect 24964 10577 24992 10911
rect 24950 10568 25006 10577
rect 24860 10532 24912 10538
rect 24950 10503 25006 10512
rect 24860 10474 24912 10480
rect 24582 9616 24638 9625
rect 24582 9551 24638 9560
rect 24216 9512 24268 9518
rect 24214 9480 24216 9489
rect 24268 9480 24270 9489
rect 24214 9415 24270 9424
rect 24400 9376 24452 9382
rect 24398 9344 24400 9353
rect 24452 9344 24454 9353
rect 24398 9279 24454 9288
rect 23202 9208 23258 9217
rect 23202 9143 23258 9152
rect 21824 8968 21876 8974
rect 21824 8910 21876 8916
rect 22100 8968 22152 8974
rect 22100 8910 22152 8916
rect 21732 8900 21784 8906
rect 21732 8842 21784 8848
rect 21640 8560 21692 8566
rect 21640 8502 21692 8508
rect 21652 8430 21680 8502
rect 21744 8498 21772 8842
rect 22112 8634 22140 8910
rect 22100 8628 22152 8634
rect 22100 8570 22152 8576
rect 21732 8492 21784 8498
rect 21732 8434 21784 8440
rect 21640 8424 21692 8430
rect 21640 8366 21692 8372
rect 21744 8090 21772 8434
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 21364 8084 21416 8090
rect 21364 8026 21416 8032
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21732 8084 21784 8090
rect 21732 8026 21784 8032
rect 20260 8016 20312 8022
rect 20260 7958 20312 7964
rect 20364 7546 20392 8026
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20956 7100 21252 7120
rect 21012 7098 21036 7100
rect 21092 7098 21116 7100
rect 21172 7098 21196 7100
rect 21034 7046 21036 7098
rect 21098 7046 21110 7098
rect 21172 7046 21174 7098
rect 21012 7044 21036 7046
rect 21092 7044 21116 7046
rect 21172 7044 21196 7046
rect 20956 7024 21252 7044
rect 20956 6012 21252 6032
rect 21012 6010 21036 6012
rect 21092 6010 21116 6012
rect 21172 6010 21196 6012
rect 21034 5958 21036 6010
rect 21098 5958 21110 6010
rect 21172 5958 21174 6010
rect 21012 5956 21036 5958
rect 21092 5956 21116 5958
rect 21172 5956 21196 5958
rect 20956 5936 21252 5956
rect 20956 4924 21252 4944
rect 21012 4922 21036 4924
rect 21092 4922 21116 4924
rect 21172 4922 21196 4924
rect 21034 4870 21036 4922
rect 21098 4870 21110 4922
rect 21172 4870 21174 4922
rect 21012 4868 21036 4870
rect 21092 4868 21116 4870
rect 21172 4868 21196 4870
rect 20956 4848 21252 4868
rect 19890 4040 19946 4049
rect 19890 3975 19946 3984
rect 20956 3836 21252 3856
rect 21012 3834 21036 3836
rect 21092 3834 21116 3836
rect 21172 3834 21196 3836
rect 21034 3782 21036 3834
rect 21098 3782 21110 3834
rect 21172 3782 21174 3834
rect 21012 3780 21036 3782
rect 21092 3780 21116 3782
rect 21172 3780 21196 3782
rect 20956 3760 21252 3780
rect 20956 2748 21252 2768
rect 21012 2746 21036 2748
rect 21092 2746 21116 2748
rect 21172 2746 21196 2748
rect 21034 2694 21036 2746
rect 21098 2694 21110 2746
rect 21172 2694 21174 2746
rect 21012 2692 21036 2694
rect 21092 2692 21116 2694
rect 21172 2692 21196 2694
rect 20956 2672 21252 2692
rect 24872 2038 24900 10474
rect 25056 8809 25084 14583
rect 25148 11218 25176 14758
rect 25332 14074 25360 15370
rect 25320 14068 25372 14074
rect 25320 14010 25372 14016
rect 25516 13954 25544 18255
rect 25608 17814 25636 20318
rect 25780 20256 25832 20262
rect 25780 20198 25832 20204
rect 26700 20256 26752 20262
rect 26700 20198 26752 20204
rect 25596 17808 25648 17814
rect 25594 17776 25596 17785
rect 25648 17776 25650 17785
rect 25594 17711 25650 17720
rect 25688 17740 25740 17746
rect 25608 17202 25636 17711
rect 25688 17682 25740 17688
rect 25700 17338 25728 17682
rect 25688 17332 25740 17338
rect 25688 17274 25740 17280
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25688 16244 25740 16250
rect 25688 16186 25740 16192
rect 25700 15858 25728 16186
rect 25792 16017 25820 20198
rect 26516 19712 26568 19718
rect 26516 19654 26568 19660
rect 25956 19612 26252 19632
rect 26012 19610 26036 19612
rect 26092 19610 26116 19612
rect 26172 19610 26196 19612
rect 26034 19558 26036 19610
rect 26098 19558 26110 19610
rect 26172 19558 26174 19610
rect 26012 19556 26036 19558
rect 26092 19556 26116 19558
rect 26172 19556 26196 19558
rect 25956 19536 26252 19556
rect 25872 19304 25924 19310
rect 25872 19246 25924 19252
rect 25884 18766 25912 19246
rect 26528 18970 26556 19654
rect 26516 18964 26568 18970
rect 26516 18906 26568 18912
rect 26516 18828 26568 18834
rect 26516 18770 26568 18776
rect 25872 18760 25924 18766
rect 25872 18702 25924 18708
rect 25884 18358 25912 18702
rect 25956 18524 26252 18544
rect 26012 18522 26036 18524
rect 26092 18522 26116 18524
rect 26172 18522 26196 18524
rect 26034 18470 26036 18522
rect 26098 18470 26110 18522
rect 26172 18470 26174 18522
rect 26012 18468 26036 18470
rect 26092 18468 26116 18470
rect 26172 18468 26196 18470
rect 25956 18448 26252 18468
rect 25872 18352 25924 18358
rect 25872 18294 25924 18300
rect 26240 18080 26292 18086
rect 26160 18040 26240 18068
rect 26160 17678 26188 18040
rect 26240 18022 26292 18028
rect 26528 17882 26556 18770
rect 26332 17876 26384 17882
rect 26332 17818 26384 17824
rect 26516 17876 26568 17882
rect 26516 17818 26568 17824
rect 26148 17672 26200 17678
rect 26148 17614 26200 17620
rect 25956 17436 26252 17456
rect 26012 17434 26036 17436
rect 26092 17434 26116 17436
rect 26172 17434 26196 17436
rect 26034 17382 26036 17434
rect 26098 17382 26110 17434
rect 26172 17382 26174 17434
rect 26012 17380 26036 17382
rect 26092 17380 26116 17382
rect 26172 17380 26196 17382
rect 25956 17360 26252 17380
rect 26240 17128 26292 17134
rect 26240 17070 26292 17076
rect 25872 16584 25924 16590
rect 25872 16526 25924 16532
rect 25778 16008 25834 16017
rect 25778 15943 25834 15952
rect 25700 15830 25820 15858
rect 25596 15564 25648 15570
rect 25596 15506 25648 15512
rect 25240 13926 25544 13954
rect 25136 11212 25188 11218
rect 25136 11154 25188 11160
rect 25148 10810 25176 11154
rect 25240 10985 25268 13926
rect 25608 13569 25636 15506
rect 25688 14816 25740 14822
rect 25688 14758 25740 14764
rect 25700 13938 25728 14758
rect 25688 13932 25740 13938
rect 25688 13874 25740 13880
rect 25686 13696 25742 13705
rect 25686 13631 25742 13640
rect 25594 13560 25650 13569
rect 25594 13495 25650 13504
rect 25700 13394 25728 13631
rect 25688 13388 25740 13394
rect 25688 13330 25740 13336
rect 25320 13320 25372 13326
rect 25320 13262 25372 13268
rect 25332 13190 25360 13262
rect 25596 13252 25648 13258
rect 25596 13194 25648 13200
rect 25320 13184 25372 13190
rect 25320 13126 25372 13132
rect 25332 12306 25360 13126
rect 25608 12306 25636 13194
rect 25700 12986 25728 13330
rect 25688 12980 25740 12986
rect 25688 12922 25740 12928
rect 25320 12300 25372 12306
rect 25320 12242 25372 12248
rect 25596 12300 25648 12306
rect 25596 12242 25648 12248
rect 25332 11082 25360 12242
rect 25502 11112 25558 11121
rect 25320 11076 25372 11082
rect 25320 11018 25372 11024
rect 25412 11076 25464 11082
rect 25502 11047 25558 11056
rect 25412 11018 25464 11024
rect 25226 10976 25282 10985
rect 25226 10911 25282 10920
rect 25226 10840 25282 10849
rect 25136 10804 25188 10810
rect 25226 10775 25282 10784
rect 25136 10746 25188 10752
rect 25240 9518 25268 10775
rect 25332 10266 25360 11018
rect 25320 10260 25372 10266
rect 25320 10202 25372 10208
rect 25320 10124 25372 10130
rect 25320 10066 25372 10072
rect 25332 10033 25360 10066
rect 25318 10024 25374 10033
rect 25318 9959 25374 9968
rect 25332 9722 25360 9959
rect 25320 9716 25372 9722
rect 25320 9658 25372 9664
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 25318 9072 25374 9081
rect 25318 9007 25320 9016
rect 25372 9007 25374 9016
rect 25320 8978 25372 8984
rect 25042 8800 25098 8809
rect 25042 8735 25098 8744
rect 25332 8634 25360 8978
rect 25320 8628 25372 8634
rect 25320 8570 25372 8576
rect 25424 2417 25452 11018
rect 25516 9654 25544 11047
rect 25686 10704 25742 10713
rect 25686 10639 25742 10648
rect 25596 9920 25648 9926
rect 25596 9862 25648 9868
rect 25504 9648 25556 9654
rect 25504 9590 25556 9596
rect 25504 8832 25556 8838
rect 25504 8774 25556 8780
rect 25516 8537 25544 8774
rect 25502 8528 25558 8537
rect 25502 8463 25558 8472
rect 25504 8288 25556 8294
rect 25504 8230 25556 8236
rect 25516 8129 25544 8230
rect 25502 8120 25558 8129
rect 25502 8055 25558 8064
rect 25608 3505 25636 9862
rect 25700 3913 25728 10639
rect 25792 8634 25820 15830
rect 25884 15706 25912 16526
rect 26252 16436 26280 17070
rect 26344 17066 26372 17818
rect 26332 17060 26384 17066
rect 26332 17002 26384 17008
rect 26332 16448 26384 16454
rect 26252 16408 26332 16436
rect 26332 16390 26384 16396
rect 25956 16348 26252 16368
rect 26012 16346 26036 16348
rect 26092 16346 26116 16348
rect 26172 16346 26196 16348
rect 26034 16294 26036 16346
rect 26098 16294 26110 16346
rect 26172 16294 26174 16346
rect 26012 16292 26036 16294
rect 26092 16292 26116 16294
rect 26172 16292 26196 16294
rect 25956 16272 26252 16292
rect 26344 16232 26372 16390
rect 26252 16204 26372 16232
rect 25964 16176 26016 16182
rect 25962 16144 25964 16153
rect 26016 16144 26018 16153
rect 25962 16079 26018 16088
rect 26148 16040 26200 16046
rect 26252 16028 26280 16204
rect 26200 16000 26280 16028
rect 26424 16040 26476 16046
rect 26330 16008 26386 16017
rect 26148 15982 26200 15988
rect 25872 15700 25924 15706
rect 25872 15642 25924 15648
rect 25884 15502 25912 15642
rect 26160 15502 26188 15982
rect 26424 15982 26476 15988
rect 26330 15943 26386 15952
rect 25872 15496 25924 15502
rect 25872 15438 25924 15444
rect 26148 15496 26200 15502
rect 26148 15438 26200 15444
rect 25956 15260 26252 15280
rect 26012 15258 26036 15260
rect 26092 15258 26116 15260
rect 26172 15258 26196 15260
rect 26034 15206 26036 15258
rect 26098 15206 26110 15258
rect 26172 15206 26174 15258
rect 26012 15204 26036 15206
rect 26092 15204 26116 15206
rect 26172 15204 26196 15206
rect 25956 15184 26252 15204
rect 26344 14278 26372 15943
rect 26436 14550 26464 15982
rect 26608 15496 26660 15502
rect 26608 15438 26660 15444
rect 26516 15360 26568 15366
rect 26516 15302 26568 15308
rect 26528 14958 26556 15302
rect 26516 14952 26568 14958
rect 26516 14894 26568 14900
rect 26528 14618 26556 14894
rect 26620 14822 26648 15438
rect 26608 14816 26660 14822
rect 26608 14758 26660 14764
rect 26516 14612 26568 14618
rect 26516 14554 26568 14560
rect 26424 14544 26476 14550
rect 26424 14486 26476 14492
rect 25872 14272 25924 14278
rect 25872 14214 25924 14220
rect 26332 14272 26384 14278
rect 26332 14214 26384 14220
rect 25884 13870 25912 14214
rect 25956 14172 26252 14192
rect 26012 14170 26036 14172
rect 26092 14170 26116 14172
rect 26172 14170 26196 14172
rect 26034 14118 26036 14170
rect 26098 14118 26110 14170
rect 26172 14118 26174 14170
rect 26012 14116 26036 14118
rect 26092 14116 26116 14118
rect 26172 14116 26196 14118
rect 25956 14096 26252 14116
rect 26514 14104 26570 14113
rect 26514 14039 26570 14048
rect 25872 13864 25924 13870
rect 25872 13806 25924 13812
rect 25884 13530 25912 13806
rect 26528 13569 26556 14039
rect 26514 13560 26570 13569
rect 25872 13524 25924 13530
rect 26514 13495 26570 13504
rect 25872 13466 25924 13472
rect 25872 13320 25924 13326
rect 25872 13262 25924 13268
rect 25884 12918 25912 13262
rect 26424 13252 26476 13258
rect 26424 13194 26476 13200
rect 26332 13184 26384 13190
rect 26332 13126 26384 13132
rect 25956 13084 26252 13104
rect 26012 13082 26036 13084
rect 26092 13082 26116 13084
rect 26172 13082 26196 13084
rect 26034 13030 26036 13082
rect 26098 13030 26110 13082
rect 26172 13030 26174 13082
rect 26012 13028 26036 13030
rect 26092 13028 26116 13030
rect 26172 13028 26196 13030
rect 25956 13008 26252 13028
rect 25872 12912 25924 12918
rect 25872 12854 25924 12860
rect 26148 12776 26200 12782
rect 26148 12718 26200 12724
rect 26160 12374 26188 12718
rect 26148 12368 26200 12374
rect 26148 12310 26200 12316
rect 25872 12096 25924 12102
rect 25872 12038 25924 12044
rect 25884 11694 25912 12038
rect 25956 11996 26252 12016
rect 26012 11994 26036 11996
rect 26092 11994 26116 11996
rect 26172 11994 26196 11996
rect 26034 11942 26036 11994
rect 26098 11942 26110 11994
rect 26172 11942 26174 11994
rect 26012 11940 26036 11942
rect 26092 11940 26116 11942
rect 26172 11940 26196 11942
rect 25956 11920 26252 11940
rect 25872 11688 25924 11694
rect 25872 11630 25924 11636
rect 26344 11354 26372 13126
rect 26436 12782 26464 13194
rect 26424 12776 26476 12782
rect 26424 12718 26476 12724
rect 26422 12608 26478 12617
rect 26422 12543 26478 12552
rect 26332 11348 26384 11354
rect 26332 11290 26384 11296
rect 25956 10908 26252 10928
rect 26012 10906 26036 10908
rect 26092 10906 26116 10908
rect 26172 10906 26196 10908
rect 26034 10854 26036 10906
rect 26098 10854 26110 10906
rect 26172 10854 26174 10906
rect 26012 10852 26036 10854
rect 26092 10852 26116 10854
rect 26172 10852 26196 10854
rect 25956 10832 26252 10852
rect 26436 10810 26464 12543
rect 26528 12442 26556 13495
rect 26620 12481 26648 14758
rect 26712 14362 26740 20198
rect 27526 20088 27582 20097
rect 27526 20023 27582 20032
rect 27252 19916 27304 19922
rect 27252 19858 27304 19864
rect 26976 19848 27028 19854
rect 26976 19790 27028 19796
rect 26988 18873 27016 19790
rect 27264 19174 27292 19858
rect 27436 19848 27488 19854
rect 27436 19790 27488 19796
rect 27448 19310 27476 19790
rect 27436 19304 27488 19310
rect 27436 19246 27488 19252
rect 27540 19258 27568 20023
rect 27252 19168 27304 19174
rect 27252 19110 27304 19116
rect 26974 18864 27030 18873
rect 26974 18799 27030 18808
rect 27264 18057 27292 19110
rect 27344 18624 27396 18630
rect 27344 18566 27396 18572
rect 27356 18086 27384 18566
rect 27344 18080 27396 18086
rect 27250 18048 27306 18057
rect 27344 18022 27396 18028
rect 27250 17983 27306 17992
rect 27448 17678 27476 19246
rect 27540 19230 27660 19258
rect 27632 19174 27660 19230
rect 27620 19168 27672 19174
rect 27620 19110 27672 19116
rect 27632 18873 27660 19110
rect 27618 18864 27674 18873
rect 27618 18799 27674 18808
rect 27528 18080 27580 18086
rect 27528 18022 27580 18028
rect 27436 17672 27488 17678
rect 27436 17614 27488 17620
rect 27448 17338 27476 17614
rect 27540 17524 27568 18022
rect 27620 17536 27672 17542
rect 27540 17496 27620 17524
rect 27620 17478 27672 17484
rect 27436 17332 27488 17338
rect 27436 17274 27488 17280
rect 27632 17241 27660 17478
rect 27618 17232 27674 17241
rect 27618 17167 27674 17176
rect 27528 16992 27580 16998
rect 27528 16934 27580 16940
rect 26884 16652 26936 16658
rect 26884 16594 26936 16600
rect 26976 16652 27028 16658
rect 26976 16594 27028 16600
rect 26896 16561 26924 16594
rect 26882 16552 26938 16561
rect 26882 16487 26938 16496
rect 26988 16153 27016 16594
rect 26974 16144 27030 16153
rect 26974 16079 27030 16088
rect 27540 16046 27568 16934
rect 28078 16552 28134 16561
rect 28078 16487 28134 16496
rect 28092 16250 28120 16487
rect 28080 16244 28132 16250
rect 28080 16186 28132 16192
rect 27528 16040 27580 16046
rect 27528 15982 27580 15988
rect 27344 15904 27396 15910
rect 27344 15846 27396 15852
rect 27158 15600 27214 15609
rect 27158 15535 27214 15544
rect 26792 14816 26844 14822
rect 26792 14758 26844 14764
rect 26804 14521 26832 14758
rect 26790 14512 26846 14521
rect 26790 14447 26846 14456
rect 26884 14476 26936 14482
rect 26884 14418 26936 14424
rect 26896 14385 26924 14418
rect 26976 14408 27028 14414
rect 26882 14376 26938 14385
rect 26712 14334 26832 14362
rect 26698 13832 26754 13841
rect 26698 13767 26754 13776
rect 26606 12472 26662 12481
rect 26516 12436 26568 12442
rect 26606 12407 26662 12416
rect 26516 12378 26568 12384
rect 26516 12300 26568 12306
rect 26516 12242 26568 12248
rect 26528 11898 26556 12242
rect 26516 11892 26568 11898
rect 26516 11834 26568 11840
rect 26516 11620 26568 11626
rect 26516 11562 26568 11568
rect 26528 11354 26556 11562
rect 26516 11348 26568 11354
rect 26516 11290 26568 11296
rect 26424 10804 26476 10810
rect 26424 10746 26476 10752
rect 26712 10266 26740 13767
rect 26804 10606 26832 14334
rect 26976 14350 27028 14356
rect 26882 14311 26938 14320
rect 26884 14272 26936 14278
rect 26884 14214 26936 14220
rect 26896 10674 26924 14214
rect 26988 14006 27016 14350
rect 27172 14278 27200 15535
rect 27356 15026 27384 15846
rect 27540 15706 27568 15982
rect 27528 15700 27580 15706
rect 27528 15642 27580 15648
rect 27436 15564 27488 15570
rect 27436 15506 27488 15512
rect 27344 15020 27396 15026
rect 27344 14962 27396 14968
rect 27356 14929 27384 14962
rect 27342 14920 27398 14929
rect 27264 14878 27342 14906
rect 27264 14618 27292 14878
rect 27342 14855 27398 14864
rect 27344 14816 27396 14822
rect 27344 14758 27396 14764
rect 27252 14612 27304 14618
rect 27252 14554 27304 14560
rect 27160 14272 27212 14278
rect 27160 14214 27212 14220
rect 26976 14000 27028 14006
rect 26974 13968 26976 13977
rect 27028 13968 27030 13977
rect 26974 13903 27030 13912
rect 26988 13877 27016 13903
rect 27160 13728 27212 13734
rect 27160 13670 27212 13676
rect 27172 13326 27200 13670
rect 26976 13320 27028 13326
rect 26976 13262 27028 13268
rect 27160 13320 27212 13326
rect 27160 13262 27212 13268
rect 26988 12714 27016 13262
rect 27172 12986 27200 13262
rect 27160 12980 27212 12986
rect 27160 12922 27212 12928
rect 27264 12850 27292 14554
rect 27356 12889 27384 14758
rect 27448 14600 27476 15506
rect 27540 15502 27568 15642
rect 27528 15496 27580 15502
rect 27528 15438 27580 15444
rect 27620 14884 27672 14890
rect 27620 14826 27672 14832
rect 27632 14600 27660 14826
rect 27448 14572 27660 14600
rect 27342 12880 27398 12889
rect 27252 12844 27304 12850
rect 27342 12815 27398 12824
rect 27252 12786 27304 12792
rect 26976 12708 27028 12714
rect 26976 12650 27028 12656
rect 27252 12708 27304 12714
rect 27252 12650 27304 12656
rect 27160 12640 27212 12646
rect 27160 12582 27212 12588
rect 26976 12436 27028 12442
rect 26976 12378 27028 12384
rect 26988 11898 27016 12378
rect 27172 12238 27200 12582
rect 27160 12232 27212 12238
rect 27160 12174 27212 12180
rect 27172 11898 27200 12174
rect 26976 11892 27028 11898
rect 26976 11834 27028 11840
rect 27160 11892 27212 11898
rect 27160 11834 27212 11840
rect 27068 11824 27120 11830
rect 26974 11792 27030 11801
rect 27068 11766 27120 11772
rect 26974 11727 27030 11736
rect 26988 11694 27016 11727
rect 26976 11688 27028 11694
rect 26976 11630 27028 11636
rect 26884 10668 26936 10674
rect 26884 10610 26936 10616
rect 26792 10600 26844 10606
rect 26792 10542 26844 10548
rect 26974 10568 27030 10577
rect 26974 10503 27030 10512
rect 26988 10266 27016 10503
rect 26700 10260 26752 10266
rect 26700 10202 26752 10208
rect 26976 10260 27028 10266
rect 26976 10202 27028 10208
rect 26792 10124 26844 10130
rect 26792 10066 26844 10072
rect 25956 9820 26252 9840
rect 26012 9818 26036 9820
rect 26092 9818 26116 9820
rect 26172 9818 26196 9820
rect 26034 9766 26036 9818
rect 26098 9766 26110 9818
rect 26172 9766 26174 9818
rect 26012 9764 26036 9766
rect 26092 9764 26116 9766
rect 26172 9764 26196 9766
rect 25956 9744 26252 9764
rect 26804 9450 26832 10066
rect 26988 9722 27016 10202
rect 26976 9716 27028 9722
rect 26976 9658 27028 9664
rect 26792 9444 26844 9450
rect 26792 9386 26844 9392
rect 26884 9376 26936 9382
rect 26884 9318 26936 9324
rect 26422 9208 26478 9217
rect 26422 9143 26478 9152
rect 25872 8832 25924 8838
rect 25872 8774 25924 8780
rect 25780 8628 25832 8634
rect 25780 8570 25832 8576
rect 25792 8430 25820 8570
rect 25780 8424 25832 8430
rect 25780 8366 25832 8372
rect 25884 8242 25912 8774
rect 25956 8732 26252 8752
rect 26012 8730 26036 8732
rect 26092 8730 26116 8732
rect 26172 8730 26196 8732
rect 26034 8678 26036 8730
rect 26098 8678 26110 8730
rect 26172 8678 26174 8730
rect 26012 8676 26036 8678
rect 26092 8676 26116 8678
rect 26172 8676 26196 8678
rect 25956 8656 26252 8676
rect 26240 8560 26292 8566
rect 26240 8502 26292 8508
rect 25792 8214 25912 8242
rect 25792 4593 25820 8214
rect 26252 7954 26280 8502
rect 26436 8430 26464 9143
rect 26516 9036 26568 9042
rect 26516 8978 26568 8984
rect 26528 8945 26556 8978
rect 26514 8936 26570 8945
rect 26514 8871 26570 8880
rect 26528 8634 26556 8871
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 26608 8560 26660 8566
rect 26608 8502 26660 8508
rect 26424 8424 26476 8430
rect 26424 8366 26476 8372
rect 26240 7948 26292 7954
rect 26240 7890 26292 7896
rect 25956 7644 26252 7664
rect 26012 7642 26036 7644
rect 26092 7642 26116 7644
rect 26172 7642 26196 7644
rect 26034 7590 26036 7642
rect 26098 7590 26110 7642
rect 26172 7590 26174 7642
rect 26012 7588 26036 7590
rect 26092 7588 26116 7590
rect 26172 7588 26196 7590
rect 25956 7568 26252 7588
rect 26620 7449 26648 8502
rect 26792 7744 26844 7750
rect 26792 7686 26844 7692
rect 26606 7440 26662 7449
rect 26606 7375 26662 7384
rect 26514 7304 26570 7313
rect 26514 7239 26570 7248
rect 26332 7200 26384 7206
rect 26332 7142 26384 7148
rect 25956 6556 26252 6576
rect 26012 6554 26036 6556
rect 26092 6554 26116 6556
rect 26172 6554 26196 6556
rect 26034 6502 26036 6554
rect 26098 6502 26110 6554
rect 26172 6502 26174 6554
rect 26012 6500 26036 6502
rect 26092 6500 26116 6502
rect 26172 6500 26196 6502
rect 25956 6480 26252 6500
rect 25956 5468 26252 5488
rect 26012 5466 26036 5468
rect 26092 5466 26116 5468
rect 26172 5466 26196 5468
rect 26034 5414 26036 5466
rect 26098 5414 26110 5466
rect 26172 5414 26174 5466
rect 26012 5412 26036 5414
rect 26092 5412 26116 5414
rect 26172 5412 26196 5414
rect 25956 5392 26252 5412
rect 26344 4978 26372 7142
rect 26528 6866 26556 7239
rect 26516 6860 26568 6866
rect 26516 6802 26568 6808
rect 26528 6458 26556 6802
rect 26700 6656 26752 6662
rect 26700 6598 26752 6604
rect 26516 6452 26568 6458
rect 26516 6394 26568 6400
rect 26712 6361 26740 6598
rect 26698 6352 26754 6361
rect 26698 6287 26754 6296
rect 26422 5264 26478 5273
rect 26422 5199 26478 5208
rect 26436 5166 26464 5199
rect 26424 5160 26476 5166
rect 26424 5102 26476 5108
rect 26606 5128 26662 5137
rect 26606 5063 26662 5072
rect 26620 5030 26648 5063
rect 25884 4950 26372 4978
rect 26608 5024 26660 5030
rect 26608 4966 26660 4972
rect 25778 4584 25834 4593
rect 25778 4519 25834 4528
rect 25686 3904 25742 3913
rect 25686 3839 25742 3848
rect 25594 3496 25650 3505
rect 25594 3431 25650 3440
rect 25410 2408 25466 2417
rect 25410 2343 25466 2352
rect 24860 2032 24912 2038
rect 24860 1974 24912 1980
rect 25884 1465 25912 4950
rect 25956 4380 26252 4400
rect 26012 4378 26036 4380
rect 26092 4378 26116 4380
rect 26172 4378 26196 4380
rect 26034 4326 26036 4378
rect 26098 4326 26110 4378
rect 26172 4326 26174 4378
rect 26012 4324 26036 4326
rect 26092 4324 26116 4326
rect 26172 4324 26196 4326
rect 25956 4304 26252 4324
rect 26422 4040 26478 4049
rect 26422 3975 26478 3984
rect 25956 3292 26252 3312
rect 26012 3290 26036 3292
rect 26092 3290 26116 3292
rect 26172 3290 26196 3292
rect 26034 3238 26036 3290
rect 26098 3238 26110 3290
rect 26172 3238 26174 3290
rect 26012 3236 26036 3238
rect 26092 3236 26116 3238
rect 26172 3236 26196 3238
rect 25956 3216 26252 3236
rect 26436 2990 26464 3975
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 26608 2848 26660 2854
rect 26606 2816 26608 2825
rect 26660 2816 26662 2825
rect 26606 2751 26662 2760
rect 25956 2204 26252 2224
rect 26012 2202 26036 2204
rect 26092 2202 26116 2204
rect 26172 2202 26196 2204
rect 26034 2150 26036 2202
rect 26098 2150 26110 2202
rect 26172 2150 26174 2202
rect 26012 2148 26036 2150
rect 26092 2148 26116 2150
rect 26172 2148 26196 2150
rect 25956 2128 26252 2148
rect 26148 2032 26200 2038
rect 26148 1974 26200 1980
rect 25870 1456 25926 1465
rect 25870 1391 25926 1400
rect 26160 480 26188 1974
rect 4066 368 4122 377
rect 4066 303 4122 312
rect 11150 0 11206 480
rect 18694 0 18750 480
rect 26146 0 26202 480
rect 26804 377 26832 7686
rect 26896 921 26924 9318
rect 26976 7948 27028 7954
rect 26976 7890 27028 7896
rect 26988 7546 27016 7890
rect 26976 7540 27028 7546
rect 26976 7482 27028 7488
rect 27080 7342 27108 11766
rect 27172 11150 27200 11834
rect 27160 11144 27212 11150
rect 27160 11086 27212 11092
rect 27160 10668 27212 10674
rect 27160 10610 27212 10616
rect 27172 10062 27200 10610
rect 27160 10056 27212 10062
rect 27160 9998 27212 10004
rect 27172 9178 27200 9998
rect 27264 9654 27292 12650
rect 27356 11642 27384 12815
rect 27448 12345 27476 14572
rect 27618 14376 27674 14385
rect 27618 14311 27674 14320
rect 27712 14340 27764 14346
rect 27632 13530 27660 14311
rect 27712 14282 27764 14288
rect 27724 14074 27752 14282
rect 27712 14068 27764 14074
rect 27712 14010 27764 14016
rect 27620 13524 27672 13530
rect 27620 13466 27672 13472
rect 27528 13388 27580 13394
rect 27528 13330 27580 13336
rect 27540 12889 27568 13330
rect 27526 12880 27582 12889
rect 27526 12815 27582 12824
rect 27528 12776 27580 12782
rect 27528 12718 27580 12724
rect 27434 12336 27490 12345
rect 27434 12271 27490 12280
rect 27356 11614 27476 11642
rect 27344 11552 27396 11558
rect 27344 11494 27396 11500
rect 27356 10713 27384 11494
rect 27342 10704 27398 10713
rect 27342 10639 27398 10648
rect 27342 10160 27398 10169
rect 27342 10095 27398 10104
rect 27252 9648 27304 9654
rect 27252 9590 27304 9596
rect 27160 9172 27212 9178
rect 27160 9114 27212 9120
rect 27356 8430 27384 10095
rect 27344 8424 27396 8430
rect 27344 8366 27396 8372
rect 27448 7478 27476 11614
rect 27540 10674 27568 12718
rect 27528 10668 27580 10674
rect 27528 10610 27580 10616
rect 27526 9616 27582 9625
rect 27526 9551 27582 9560
rect 27710 9616 27766 9625
rect 27710 9551 27766 9560
rect 27540 9518 27568 9551
rect 27528 9512 27580 9518
rect 27528 9454 27580 9460
rect 27724 8634 27752 9551
rect 27804 9376 27856 9382
rect 27804 9318 27856 9324
rect 27712 8628 27764 8634
rect 27712 8570 27764 8576
rect 27436 7472 27488 7478
rect 27436 7414 27488 7420
rect 27068 7336 27120 7342
rect 27068 7278 27120 7284
rect 27712 7200 27764 7206
rect 27712 7142 27764 7148
rect 27724 7041 27752 7142
rect 27710 7032 27766 7041
rect 27710 6967 27766 6976
rect 27816 5681 27844 9318
rect 27802 5672 27858 5681
rect 27802 5607 27858 5616
rect 26882 912 26938 921
rect 26882 847 26938 856
rect 26790 368 26846 377
rect 26790 303 26846 312
<< via2 >>
rect 3514 23568 3570 23624
rect 3422 23024 3478 23080
rect 25042 23568 25098 23624
rect 3238 22344 3294 22400
rect 2962 20576 3018 20632
rect 1766 15680 1822 15736
rect 1674 14456 1730 14512
rect 2042 15408 2098 15464
rect 1582 13368 1638 13424
rect 570 12824 626 12880
rect 1490 12144 1546 12200
rect 2410 19488 2466 19544
rect 2042 12144 2098 12200
rect 1950 10512 2006 10568
rect 1490 7384 1546 7440
rect 1582 6296 1638 6352
rect 1398 5772 1454 5808
rect 1398 5752 1400 5772
rect 1400 5752 1452 5772
rect 1452 5752 1454 5772
rect 1674 5616 1730 5672
rect 570 3304 626 3360
rect 3054 17720 3110 17776
rect 2686 14340 2742 14376
rect 2686 14320 2688 14340
rect 2688 14320 2740 14340
rect 2740 14320 2742 14340
rect 3146 15952 3202 16008
rect 2778 12960 2834 13016
rect 2962 12824 3018 12880
rect 2410 11600 2466 11656
rect 1950 9444 2006 9480
rect 1950 9424 1952 9444
rect 1952 9424 2004 9444
rect 2004 9424 2006 9444
rect 2962 11736 3018 11792
rect 2686 11192 2742 11248
rect 3790 21800 3846 21856
rect 4066 21256 4122 21312
rect 3698 19216 3754 19272
rect 3882 19116 3884 19136
rect 3884 19116 3936 19136
rect 3936 19116 3938 19136
rect 3882 19080 3938 19116
rect 3790 18808 3846 18864
rect 3514 18264 3570 18320
rect 3698 18264 3754 18320
rect 3330 17856 3386 17912
rect 3514 16632 3570 16688
rect 3514 15036 3516 15056
rect 3516 15036 3568 15056
rect 3568 15036 3570 15056
rect 3514 15000 3570 15036
rect 4434 20052 4490 20088
rect 4434 20032 4436 20052
rect 4436 20032 4488 20052
rect 4488 20032 4490 20052
rect 5956 21786 6012 21788
rect 6036 21786 6092 21788
rect 6116 21786 6172 21788
rect 6196 21786 6252 21788
rect 5956 21734 5982 21786
rect 5982 21734 6012 21786
rect 6036 21734 6046 21786
rect 6046 21734 6092 21786
rect 6116 21734 6162 21786
rect 6162 21734 6172 21786
rect 6196 21734 6226 21786
rect 6226 21734 6252 21786
rect 5956 21732 6012 21734
rect 6036 21732 6092 21734
rect 6116 21732 6172 21734
rect 6196 21732 6252 21734
rect 4618 19488 4674 19544
rect 4250 17856 4306 17912
rect 4434 17720 4490 17776
rect 4158 16768 4214 16824
rect 3790 15952 3846 16008
rect 3790 15816 3846 15872
rect 3606 14456 3662 14512
rect 3238 10648 3294 10704
rect 3146 10240 3202 10296
rect 2042 7268 2098 7304
rect 2042 7248 2044 7268
rect 2044 7248 2096 7268
rect 2096 7248 2098 7268
rect 2502 8608 2558 8664
rect 2410 6976 2466 7032
rect 2410 6316 2466 6352
rect 2410 6296 2412 6316
rect 2412 6296 2464 6316
rect 2464 6296 2466 6316
rect 2778 8336 2834 8392
rect 2686 6840 2742 6896
rect 2226 5072 2282 5128
rect 1858 4392 1914 4448
rect 2042 3984 2098 4040
rect 1582 2624 1638 2680
rect 1490 1400 1546 1456
rect 3146 9988 3202 10024
rect 3146 9968 3148 9988
rect 3148 9968 3200 9988
rect 3200 9968 3202 9988
rect 3238 9424 3294 9480
rect 3422 9560 3478 9616
rect 3882 15544 3938 15600
rect 4066 15272 4122 15328
rect 3698 13912 3754 13968
rect 4066 13640 4122 13696
rect 3790 13232 3846 13288
rect 4066 12280 4122 12336
rect 5956 20698 6012 20700
rect 6036 20698 6092 20700
rect 6116 20698 6172 20700
rect 6196 20698 6252 20700
rect 5956 20646 5982 20698
rect 5982 20646 6012 20698
rect 6036 20646 6046 20698
rect 6046 20646 6092 20698
rect 6116 20646 6162 20698
rect 6162 20646 6172 20698
rect 6196 20646 6226 20698
rect 6226 20646 6252 20698
rect 5956 20644 6012 20646
rect 6036 20644 6092 20646
rect 6116 20644 6172 20646
rect 6196 20644 6252 20646
rect 7378 20204 7380 20224
rect 7380 20204 7432 20224
rect 7432 20204 7434 20224
rect 7378 20168 7434 20204
rect 6550 20032 6606 20088
rect 5078 18944 5134 19000
rect 4618 15816 4674 15872
rect 4526 15700 4582 15736
rect 4526 15680 4528 15700
rect 4528 15680 4580 15700
rect 4580 15680 4582 15700
rect 4434 15000 4490 15056
rect 4710 14864 4766 14920
rect 4526 14048 4582 14104
rect 3882 11736 3938 11792
rect 4250 11056 4306 11112
rect 4066 10376 4122 10432
rect 3790 9832 3846 9888
rect 3606 8064 3662 8120
rect 4250 9424 4306 9480
rect 3514 6976 3570 7032
rect 3698 3440 3754 3496
rect 2778 2080 2834 2136
rect 2686 856 2742 912
rect 4618 10240 4674 10296
rect 4434 9016 4490 9072
rect 5956 19610 6012 19612
rect 6036 19610 6092 19612
rect 6116 19610 6172 19612
rect 6196 19610 6252 19612
rect 5956 19558 5982 19610
rect 5982 19558 6012 19610
rect 6036 19558 6046 19610
rect 6046 19558 6092 19610
rect 6116 19558 6162 19610
rect 6162 19558 6172 19610
rect 6196 19558 6226 19610
rect 6226 19558 6252 19610
rect 5956 19556 6012 19558
rect 6036 19556 6092 19558
rect 6116 19556 6172 19558
rect 6196 19556 6252 19558
rect 6090 19216 6146 19272
rect 5078 17584 5134 17640
rect 5262 17584 5318 17640
rect 5446 16360 5502 16416
rect 5956 18522 6012 18524
rect 6036 18522 6092 18524
rect 6116 18522 6172 18524
rect 6196 18522 6252 18524
rect 5956 18470 5982 18522
rect 5982 18470 6012 18522
rect 6036 18470 6046 18522
rect 6046 18470 6092 18522
rect 6116 18470 6162 18522
rect 6162 18470 6172 18522
rect 6196 18470 6226 18522
rect 6226 18470 6252 18522
rect 5956 18468 6012 18470
rect 6036 18468 6092 18470
rect 6116 18468 6172 18470
rect 6196 18468 6252 18470
rect 5956 17434 6012 17436
rect 6036 17434 6092 17436
rect 6116 17434 6172 17436
rect 6196 17434 6252 17436
rect 5956 17382 5982 17434
rect 5982 17382 6012 17434
rect 6036 17382 6046 17434
rect 6046 17382 6092 17434
rect 6116 17382 6162 17434
rect 6162 17382 6172 17434
rect 6196 17382 6226 17434
rect 6226 17382 6252 17434
rect 5956 17380 6012 17382
rect 6036 17380 6092 17382
rect 6116 17380 6172 17382
rect 6196 17380 6252 17382
rect 6642 17332 6698 17368
rect 6642 17312 6644 17332
rect 6644 17312 6696 17332
rect 6696 17312 6698 17332
rect 5814 17040 5870 17096
rect 5722 16088 5778 16144
rect 5078 15952 5134 16008
rect 5354 15680 5410 15736
rect 5170 11500 5172 11520
rect 5172 11500 5224 11520
rect 5224 11500 5226 11520
rect 5170 11464 5226 11500
rect 5446 14764 5448 14784
rect 5448 14764 5500 14784
rect 5500 14764 5502 14784
rect 5446 14728 5502 14764
rect 5538 12980 5594 13016
rect 5538 12960 5540 12980
rect 5540 12960 5592 12980
rect 5592 12960 5594 12980
rect 5956 16346 6012 16348
rect 6036 16346 6092 16348
rect 6116 16346 6172 16348
rect 6196 16346 6252 16348
rect 5956 16294 5982 16346
rect 5982 16294 6012 16346
rect 6036 16294 6046 16346
rect 6046 16294 6092 16346
rect 6116 16294 6162 16346
rect 6162 16294 6172 16346
rect 6196 16294 6226 16346
rect 6226 16294 6252 16346
rect 5956 16292 6012 16294
rect 6036 16292 6092 16294
rect 6116 16292 6172 16294
rect 6196 16292 6252 16294
rect 6090 15408 6146 15464
rect 5956 15258 6012 15260
rect 6036 15258 6092 15260
rect 6116 15258 6172 15260
rect 6196 15258 6252 15260
rect 5956 15206 5982 15258
rect 5982 15206 6012 15258
rect 6036 15206 6046 15258
rect 6046 15206 6092 15258
rect 6116 15206 6162 15258
rect 6162 15206 6172 15258
rect 6196 15206 6226 15258
rect 6226 15206 6252 15258
rect 5956 15204 6012 15206
rect 6036 15204 6092 15206
rect 6116 15204 6172 15206
rect 6196 15204 6252 15206
rect 5956 14170 6012 14172
rect 6036 14170 6092 14172
rect 6116 14170 6172 14172
rect 6196 14170 6252 14172
rect 5956 14118 5982 14170
rect 5982 14118 6012 14170
rect 6036 14118 6046 14170
rect 6046 14118 6092 14170
rect 6116 14118 6162 14170
rect 6162 14118 6172 14170
rect 6196 14118 6226 14170
rect 6226 14118 6252 14170
rect 5956 14116 6012 14118
rect 6036 14116 6092 14118
rect 6116 14116 6172 14118
rect 6196 14116 6252 14118
rect 5906 13368 5962 13424
rect 5956 13082 6012 13084
rect 6036 13082 6092 13084
rect 6116 13082 6172 13084
rect 6196 13082 6252 13084
rect 5956 13030 5982 13082
rect 5982 13030 6012 13082
rect 6036 13030 6046 13082
rect 6046 13030 6092 13082
rect 6116 13030 6162 13082
rect 6162 13030 6172 13082
rect 6196 13030 6226 13082
rect 6226 13030 6252 13082
rect 5956 13028 6012 13030
rect 6036 13028 6092 13030
rect 6116 13028 6172 13030
rect 6196 13028 6252 13030
rect 5814 12824 5870 12880
rect 6182 12860 6184 12880
rect 6184 12860 6236 12880
rect 6236 12860 6238 12880
rect 6182 12824 6238 12860
rect 5538 11328 5594 11384
rect 5630 10260 5686 10296
rect 5630 10240 5632 10260
rect 5632 10240 5684 10260
rect 5684 10240 5686 10260
rect 6550 14592 6606 14648
rect 6458 13640 6514 13696
rect 5906 12180 5908 12200
rect 5908 12180 5960 12200
rect 5960 12180 5962 12200
rect 5906 12144 5962 12180
rect 6274 12144 6330 12200
rect 5956 11994 6012 11996
rect 6036 11994 6092 11996
rect 6116 11994 6172 11996
rect 6196 11994 6252 11996
rect 5956 11942 5982 11994
rect 5982 11942 6012 11994
rect 6036 11942 6046 11994
rect 6046 11942 6092 11994
rect 6116 11942 6162 11994
rect 6162 11942 6172 11994
rect 6196 11942 6226 11994
rect 6226 11942 6252 11994
rect 5956 11940 6012 11942
rect 6036 11940 6092 11942
rect 6116 11940 6172 11942
rect 6196 11940 6252 11942
rect 6366 11892 6422 11928
rect 6366 11872 6368 11892
rect 6368 11872 6420 11892
rect 6420 11872 6422 11892
rect 5956 10906 6012 10908
rect 6036 10906 6092 10908
rect 6116 10906 6172 10908
rect 6196 10906 6252 10908
rect 5956 10854 5982 10906
rect 5982 10854 6012 10906
rect 6036 10854 6046 10906
rect 6046 10854 6092 10906
rect 6116 10854 6162 10906
rect 6162 10854 6172 10906
rect 6196 10854 6226 10906
rect 6226 10854 6252 10906
rect 5956 10852 6012 10854
rect 6036 10852 6092 10854
rect 6116 10852 6172 10854
rect 6196 10852 6252 10854
rect 5998 10260 6054 10296
rect 5998 10240 6000 10260
rect 6000 10240 6052 10260
rect 6052 10240 6054 10260
rect 6090 10140 6092 10160
rect 6092 10140 6144 10160
rect 6144 10140 6146 10160
rect 6090 10104 6146 10140
rect 5956 9818 6012 9820
rect 6036 9818 6092 9820
rect 6116 9818 6172 9820
rect 6196 9818 6252 9820
rect 5956 9766 5982 9818
rect 5982 9766 6012 9818
rect 6036 9766 6046 9818
rect 6046 9766 6092 9818
rect 6116 9766 6162 9818
rect 6162 9766 6172 9818
rect 6196 9766 6226 9818
rect 6226 9766 6252 9818
rect 5956 9764 6012 9766
rect 6036 9764 6092 9766
rect 6116 9764 6172 9766
rect 6196 9764 6252 9766
rect 5814 9324 5816 9344
rect 5816 9324 5868 9344
rect 5868 9324 5870 9344
rect 5814 9288 5870 9324
rect 4894 9016 4950 9072
rect 5956 8730 6012 8732
rect 6036 8730 6092 8732
rect 6116 8730 6172 8732
rect 6196 8730 6252 8732
rect 5956 8678 5982 8730
rect 5982 8678 6012 8730
rect 6036 8678 6046 8730
rect 6046 8678 6092 8730
rect 6116 8678 6162 8730
rect 6162 8678 6172 8730
rect 6196 8678 6226 8730
rect 6226 8678 6252 8730
rect 5956 8676 6012 8678
rect 6036 8676 6092 8678
rect 6116 8676 6172 8678
rect 6196 8676 6252 8678
rect 5538 8336 5594 8392
rect 5354 7792 5410 7848
rect 5956 7642 6012 7644
rect 6036 7642 6092 7644
rect 6116 7642 6172 7644
rect 6196 7642 6252 7644
rect 5956 7590 5982 7642
rect 5982 7590 6012 7642
rect 6036 7590 6046 7642
rect 6046 7590 6092 7642
rect 6116 7590 6162 7642
rect 6162 7590 6172 7642
rect 6196 7590 6226 7642
rect 6226 7590 6252 7642
rect 5956 7588 6012 7590
rect 6036 7588 6092 7590
rect 6116 7588 6172 7590
rect 6196 7588 6252 7590
rect 6366 10104 6422 10160
rect 7194 19080 7250 19136
rect 6826 18264 6882 18320
rect 7010 18672 7066 18728
rect 6734 14456 6790 14512
rect 7102 16224 7158 16280
rect 9310 20168 9366 20224
rect 7654 18964 7710 19000
rect 7654 18944 7656 18964
rect 7656 18944 7708 18964
rect 7708 18944 7710 18964
rect 7470 17720 7526 17776
rect 7194 15544 7250 15600
rect 7286 15020 7342 15056
rect 7286 15000 7288 15020
rect 7288 15000 7340 15020
rect 7340 15000 7342 15020
rect 6918 12688 6974 12744
rect 6826 11736 6882 11792
rect 9034 19216 9090 19272
rect 8942 18536 8998 18592
rect 8298 17720 8354 17776
rect 8022 17040 8078 17096
rect 7930 16768 7986 16824
rect 7654 16632 7710 16688
rect 8390 17312 8446 17368
rect 7562 14320 7618 14376
rect 8942 17992 8998 18048
rect 7562 14048 7618 14104
rect 7286 11736 7342 11792
rect 7654 13368 7710 13424
rect 7838 13368 7894 13424
rect 7746 12960 7802 13016
rect 7470 12416 7526 12472
rect 7562 12300 7618 12336
rect 7562 12280 7564 12300
rect 7564 12280 7616 12300
rect 7616 12280 7618 12300
rect 7562 12008 7618 12064
rect 5956 6554 6012 6556
rect 6036 6554 6092 6556
rect 6116 6554 6172 6556
rect 6196 6554 6252 6556
rect 5956 6502 5982 6554
rect 5982 6502 6012 6554
rect 6036 6502 6046 6554
rect 6046 6502 6092 6554
rect 6116 6502 6162 6554
rect 6162 6502 6172 6554
rect 6196 6502 6226 6554
rect 6226 6502 6252 6554
rect 5956 6500 6012 6502
rect 6036 6500 6092 6502
rect 6116 6500 6172 6502
rect 6196 6500 6252 6502
rect 5956 5466 6012 5468
rect 6036 5466 6092 5468
rect 6116 5466 6172 5468
rect 6196 5466 6252 5468
rect 5956 5414 5982 5466
rect 5982 5414 6012 5466
rect 6036 5414 6046 5466
rect 6046 5414 6092 5466
rect 6116 5414 6162 5466
rect 6162 5414 6172 5466
rect 6196 5414 6226 5466
rect 6226 5414 6252 5466
rect 5956 5412 6012 5414
rect 6036 5412 6092 5414
rect 6116 5412 6172 5414
rect 6196 5412 6252 5414
rect 5956 4378 6012 4380
rect 6036 4378 6092 4380
rect 6116 4378 6172 4380
rect 6196 4378 6252 4380
rect 5956 4326 5982 4378
rect 5982 4326 6012 4378
rect 6036 4326 6046 4378
rect 6046 4326 6092 4378
rect 6116 4326 6162 4378
rect 6162 4326 6172 4378
rect 6196 4326 6226 4378
rect 6226 4326 6252 4378
rect 5956 4324 6012 4326
rect 6036 4324 6092 4326
rect 6116 4324 6172 4326
rect 6196 4324 6252 4326
rect 4342 3848 4398 3904
rect 5956 3290 6012 3292
rect 6036 3290 6092 3292
rect 6116 3290 6172 3292
rect 6196 3290 6252 3292
rect 5956 3238 5982 3290
rect 5982 3238 6012 3290
rect 6036 3238 6046 3290
rect 6046 3238 6092 3290
rect 6116 3238 6162 3290
rect 6162 3238 6172 3290
rect 6196 3238 6226 3290
rect 6226 3238 6252 3290
rect 5956 3236 6012 3238
rect 6036 3236 6092 3238
rect 6116 3236 6172 3238
rect 6196 3236 6252 3238
rect 7194 9988 7250 10024
rect 7194 9968 7196 9988
rect 7196 9968 7248 9988
rect 7248 9968 7250 9988
rect 7194 8372 7196 8392
rect 7196 8372 7248 8392
rect 7248 8372 7250 8392
rect 7194 8336 7250 8372
rect 7378 7792 7434 7848
rect 8390 11600 8446 11656
rect 8298 11212 8354 11248
rect 8298 11192 8300 11212
rect 8300 11192 8352 11212
rect 8352 11192 8354 11212
rect 8390 10240 8446 10296
rect 8298 9560 8354 9616
rect 7930 6976 7986 7032
rect 6918 5752 6974 5808
rect 8390 7792 8446 7848
rect 8114 3984 8170 4040
rect 8850 11500 8852 11520
rect 8852 11500 8904 11520
rect 8904 11500 8906 11520
rect 8850 11464 8906 11500
rect 9586 19488 9642 19544
rect 9586 19352 9642 19408
rect 9586 18164 9588 18184
rect 9588 18164 9640 18184
rect 9640 18164 9642 18184
rect 9586 18128 9642 18164
rect 9402 17176 9458 17232
rect 9494 16632 9550 16688
rect 10956 21242 11012 21244
rect 11036 21242 11092 21244
rect 11116 21242 11172 21244
rect 11196 21242 11252 21244
rect 10956 21190 10982 21242
rect 10982 21190 11012 21242
rect 11036 21190 11046 21242
rect 11046 21190 11092 21242
rect 11116 21190 11162 21242
rect 11162 21190 11172 21242
rect 11196 21190 11226 21242
rect 11226 21190 11252 21242
rect 10956 21188 11012 21190
rect 11036 21188 11092 21190
rect 11116 21188 11172 21190
rect 11196 21188 11252 21190
rect 10956 20154 11012 20156
rect 11036 20154 11092 20156
rect 11116 20154 11172 20156
rect 11196 20154 11252 20156
rect 10956 20102 10982 20154
rect 10982 20102 11012 20154
rect 11036 20102 11046 20154
rect 11046 20102 11092 20154
rect 11116 20102 11162 20154
rect 11162 20102 11172 20154
rect 11196 20102 11226 20154
rect 11226 20102 11252 20154
rect 10956 20100 11012 20102
rect 11036 20100 11092 20102
rect 11116 20100 11172 20102
rect 11196 20100 11252 20102
rect 10956 19066 11012 19068
rect 11036 19066 11092 19068
rect 11116 19066 11172 19068
rect 11196 19066 11252 19068
rect 10956 19014 10982 19066
rect 10982 19014 11012 19066
rect 11036 19014 11046 19066
rect 11046 19014 11092 19066
rect 11116 19014 11162 19066
rect 11162 19014 11172 19066
rect 11196 19014 11226 19066
rect 11226 19014 11252 19066
rect 10956 19012 11012 19014
rect 11036 19012 11092 19014
rect 11116 19012 11172 19014
rect 11196 19012 11252 19014
rect 15956 21786 16012 21788
rect 16036 21786 16092 21788
rect 16116 21786 16172 21788
rect 16196 21786 16252 21788
rect 15956 21734 15982 21786
rect 15982 21734 16012 21786
rect 16036 21734 16046 21786
rect 16046 21734 16092 21786
rect 16116 21734 16162 21786
rect 16162 21734 16172 21786
rect 16196 21734 16226 21786
rect 16226 21734 16252 21786
rect 15956 21732 16012 21734
rect 16036 21732 16092 21734
rect 16116 21732 16172 21734
rect 16196 21732 16252 21734
rect 15956 20698 16012 20700
rect 16036 20698 16092 20700
rect 16116 20698 16172 20700
rect 16196 20698 16252 20700
rect 15956 20646 15982 20698
rect 15982 20646 16012 20698
rect 16036 20646 16046 20698
rect 16046 20646 16092 20698
rect 16116 20646 16162 20698
rect 16162 20646 16172 20698
rect 16196 20646 16226 20698
rect 16226 20646 16252 20698
rect 15956 20644 16012 20646
rect 16036 20644 16092 20646
rect 16116 20644 16172 20646
rect 16196 20644 16252 20646
rect 10782 18808 10838 18864
rect 9954 15952 10010 16008
rect 9402 12144 9458 12200
rect 10506 16224 10562 16280
rect 10414 14728 10470 14784
rect 10414 14184 10470 14240
rect 10414 13776 10470 13832
rect 10230 11736 10286 11792
rect 11150 18264 11206 18320
rect 11702 18808 11758 18864
rect 11794 18672 11850 18728
rect 11702 18536 11758 18592
rect 11794 18400 11850 18456
rect 12070 19216 12126 19272
rect 10782 18028 10784 18048
rect 10784 18028 10836 18048
rect 10836 18028 10838 18048
rect 10782 17992 10838 18028
rect 10956 17978 11012 17980
rect 11036 17978 11092 17980
rect 11116 17978 11172 17980
rect 11196 17978 11252 17980
rect 10956 17926 10982 17978
rect 10982 17926 11012 17978
rect 11036 17926 11046 17978
rect 11046 17926 11092 17978
rect 11116 17926 11162 17978
rect 11162 17926 11172 17978
rect 11196 17926 11226 17978
rect 11226 17926 11252 17978
rect 10956 17924 11012 17926
rect 11036 17924 11092 17926
rect 11116 17924 11172 17926
rect 11196 17924 11252 17926
rect 11150 17176 11206 17232
rect 11794 17584 11850 17640
rect 11242 17060 11298 17096
rect 11242 17040 11244 17060
rect 11244 17040 11296 17060
rect 11296 17040 11298 17060
rect 10956 16890 11012 16892
rect 11036 16890 11092 16892
rect 11116 16890 11172 16892
rect 11196 16890 11252 16892
rect 10956 16838 10982 16890
rect 10982 16838 11012 16890
rect 11036 16838 11046 16890
rect 11046 16838 11092 16890
rect 11116 16838 11162 16890
rect 11162 16838 11172 16890
rect 11196 16838 11226 16890
rect 11226 16838 11252 16890
rect 10956 16836 11012 16838
rect 11036 16836 11092 16838
rect 11116 16836 11172 16838
rect 11196 16836 11252 16838
rect 11334 16632 11390 16688
rect 11610 17040 11666 17096
rect 10690 15816 10746 15872
rect 10598 15680 10654 15736
rect 10598 13948 10600 13968
rect 10600 13948 10652 13968
rect 10652 13948 10654 13968
rect 10598 13912 10654 13948
rect 8942 10512 8998 10568
rect 9310 11348 9366 11384
rect 9310 11328 9312 11348
rect 9312 11328 9364 11348
rect 9364 11328 9366 11348
rect 10956 15802 11012 15804
rect 11036 15802 11092 15804
rect 11116 15802 11172 15804
rect 11196 15802 11252 15804
rect 10956 15750 10982 15802
rect 10982 15750 11012 15802
rect 11036 15750 11046 15802
rect 11046 15750 11092 15802
rect 11116 15750 11162 15802
rect 11162 15750 11172 15802
rect 11196 15750 11226 15802
rect 11226 15750 11252 15802
rect 10956 15748 11012 15750
rect 11036 15748 11092 15750
rect 11116 15748 11172 15750
rect 11196 15748 11252 15750
rect 10956 14714 11012 14716
rect 11036 14714 11092 14716
rect 11116 14714 11172 14716
rect 11196 14714 11252 14716
rect 10956 14662 10982 14714
rect 10982 14662 11012 14714
rect 11036 14662 11046 14714
rect 11046 14662 11092 14714
rect 11116 14662 11162 14714
rect 11162 14662 11172 14714
rect 11196 14662 11226 14714
rect 11226 14662 11252 14714
rect 10956 14660 11012 14662
rect 11036 14660 11092 14662
rect 11116 14660 11172 14662
rect 11196 14660 11252 14662
rect 10956 13626 11012 13628
rect 11036 13626 11092 13628
rect 11116 13626 11172 13628
rect 11196 13626 11252 13628
rect 10956 13574 10982 13626
rect 10982 13574 11012 13626
rect 11036 13574 11046 13626
rect 11046 13574 11092 13626
rect 11116 13574 11162 13626
rect 11162 13574 11172 13626
rect 11196 13574 11226 13626
rect 11226 13574 11252 13626
rect 10956 13572 11012 13574
rect 11036 13572 11092 13574
rect 11116 13572 11172 13574
rect 11196 13572 11252 13574
rect 11794 16244 11850 16280
rect 11794 16224 11796 16244
rect 11796 16224 11848 16244
rect 11848 16224 11850 16244
rect 11702 15952 11758 16008
rect 10782 12688 10838 12744
rect 10956 12538 11012 12540
rect 11036 12538 11092 12540
rect 11116 12538 11172 12540
rect 11196 12538 11252 12540
rect 10956 12486 10982 12538
rect 10982 12486 11012 12538
rect 11036 12486 11046 12538
rect 11046 12486 11092 12538
rect 11116 12486 11162 12538
rect 11162 12486 11172 12538
rect 11196 12486 11226 12538
rect 11226 12486 11252 12538
rect 10956 12484 11012 12486
rect 11036 12484 11092 12486
rect 11116 12484 11172 12486
rect 11196 12484 11252 12486
rect 10956 11450 11012 11452
rect 11036 11450 11092 11452
rect 11116 11450 11172 11452
rect 11196 11450 11252 11452
rect 10956 11398 10982 11450
rect 10982 11398 11012 11450
rect 11036 11398 11046 11450
rect 11046 11398 11092 11450
rect 11116 11398 11162 11450
rect 11162 11398 11172 11450
rect 11196 11398 11226 11450
rect 11226 11398 11252 11450
rect 10956 11396 11012 11398
rect 11036 11396 11092 11398
rect 11116 11396 11172 11398
rect 11196 11396 11252 11398
rect 11702 15408 11758 15464
rect 11794 14456 11850 14512
rect 11610 12960 11666 13016
rect 10598 10784 10654 10840
rect 10956 10362 11012 10364
rect 11036 10362 11092 10364
rect 11116 10362 11172 10364
rect 11196 10362 11252 10364
rect 10956 10310 10982 10362
rect 10982 10310 11012 10362
rect 11036 10310 11046 10362
rect 11046 10310 11092 10362
rect 11116 10310 11162 10362
rect 11162 10310 11172 10362
rect 11196 10310 11226 10362
rect 11226 10310 11252 10362
rect 10956 10308 11012 10310
rect 11036 10308 11092 10310
rect 11116 10308 11172 10310
rect 11196 10308 11252 10310
rect 10322 10004 10324 10024
rect 10324 10004 10376 10024
rect 10376 10004 10378 10024
rect 10322 9968 10378 10004
rect 8758 9696 8814 9752
rect 10956 9274 11012 9276
rect 11036 9274 11092 9276
rect 11116 9274 11172 9276
rect 11196 9274 11252 9276
rect 10956 9222 10982 9274
rect 10982 9222 11012 9274
rect 11036 9222 11046 9274
rect 11046 9222 11092 9274
rect 11116 9222 11162 9274
rect 11162 9222 11172 9274
rect 11196 9222 11226 9274
rect 11226 9222 11252 9274
rect 10956 9220 11012 9222
rect 11036 9220 11092 9222
rect 11116 9220 11172 9222
rect 11196 9220 11252 9222
rect 8850 8472 8906 8528
rect 10956 8186 11012 8188
rect 11036 8186 11092 8188
rect 11116 8186 11172 8188
rect 11196 8186 11252 8188
rect 10956 8134 10982 8186
rect 10982 8134 11012 8186
rect 11036 8134 11046 8186
rect 11046 8134 11092 8186
rect 11116 8134 11162 8186
rect 11162 8134 11172 8186
rect 11196 8134 11226 8186
rect 11226 8134 11252 8186
rect 10956 8132 11012 8134
rect 11036 8132 11092 8134
rect 11116 8132 11172 8134
rect 11196 8132 11252 8134
rect 11978 13268 11980 13288
rect 11980 13268 12032 13288
rect 12032 13268 12034 13288
rect 11978 13232 12034 13268
rect 20956 21242 21012 21244
rect 21036 21242 21092 21244
rect 21116 21242 21172 21244
rect 21196 21242 21252 21244
rect 20956 21190 20982 21242
rect 20982 21190 21012 21242
rect 21036 21190 21046 21242
rect 21046 21190 21092 21242
rect 21116 21190 21162 21242
rect 21162 21190 21172 21242
rect 21196 21190 21226 21242
rect 21226 21190 21252 21242
rect 20956 21188 21012 21190
rect 21036 21188 21092 21190
rect 21116 21188 21172 21190
rect 21196 21188 21252 21190
rect 17774 20340 17776 20360
rect 17776 20340 17828 20360
rect 17828 20340 17830 20360
rect 17774 20304 17830 20340
rect 15382 19760 15438 19816
rect 14278 19624 14334 19680
rect 13266 17176 13322 17232
rect 12990 16632 13046 16688
rect 12346 15972 12402 16008
rect 12346 15952 12348 15972
rect 12348 15952 12400 15972
rect 12400 15952 12402 15972
rect 12898 15852 12900 15872
rect 12900 15852 12952 15872
rect 12952 15852 12954 15872
rect 12898 15816 12954 15852
rect 12162 12860 12164 12880
rect 12164 12860 12216 12880
rect 12216 12860 12218 12880
rect 12162 12824 12218 12860
rect 11794 11620 11850 11656
rect 11794 11600 11796 11620
rect 11796 11600 11848 11620
rect 11848 11600 11850 11620
rect 13818 16788 13874 16824
rect 13818 16768 13820 16788
rect 13820 16768 13872 16788
rect 13872 16768 13874 16788
rect 14002 16768 14058 16824
rect 14830 18808 14886 18864
rect 15014 17992 15070 18048
rect 15198 14864 15254 14920
rect 14830 14592 14886 14648
rect 13266 14048 13322 14104
rect 13818 13776 13874 13832
rect 13634 12824 13690 12880
rect 13910 12724 13912 12744
rect 13912 12724 13964 12744
rect 13964 12724 13966 12744
rect 13910 12688 13966 12724
rect 14738 14184 14794 14240
rect 14094 13524 14150 13560
rect 14094 13504 14096 13524
rect 14096 13504 14148 13524
rect 14148 13504 14150 13524
rect 14922 13404 14924 13424
rect 14924 13404 14976 13424
rect 14976 13404 14978 13424
rect 14922 13368 14978 13404
rect 14094 12980 14150 13016
rect 14094 12960 14096 12980
rect 14096 12960 14148 12980
rect 14148 12960 14150 12980
rect 15956 19610 16012 19612
rect 16036 19610 16092 19612
rect 16116 19610 16172 19612
rect 16196 19610 16252 19612
rect 15956 19558 15982 19610
rect 15982 19558 16012 19610
rect 16036 19558 16046 19610
rect 16046 19558 16092 19610
rect 16116 19558 16162 19610
rect 16162 19558 16172 19610
rect 16196 19558 16226 19610
rect 16226 19558 16252 19610
rect 15956 19556 16012 19558
rect 16036 19556 16092 19558
rect 16116 19556 16172 19558
rect 16196 19556 16252 19558
rect 16394 18536 16450 18592
rect 15956 18522 16012 18524
rect 16036 18522 16092 18524
rect 16116 18522 16172 18524
rect 16196 18522 16252 18524
rect 15956 18470 15982 18522
rect 15982 18470 16012 18522
rect 16036 18470 16046 18522
rect 16046 18470 16092 18522
rect 16116 18470 16162 18522
rect 16162 18470 16172 18522
rect 16196 18470 16226 18522
rect 16226 18470 16252 18522
rect 15956 18468 16012 18470
rect 16036 18468 16092 18470
rect 16116 18468 16172 18470
rect 16196 18468 16252 18470
rect 15658 17720 15714 17776
rect 16670 17992 16726 18048
rect 15956 17434 16012 17436
rect 16036 17434 16092 17436
rect 16116 17434 16172 17436
rect 16196 17434 16252 17436
rect 15956 17382 15982 17434
rect 15982 17382 16012 17434
rect 16036 17382 16046 17434
rect 16046 17382 16092 17434
rect 16116 17382 16162 17434
rect 16162 17382 16172 17434
rect 16196 17382 16226 17434
rect 16226 17382 16252 17434
rect 15956 17380 16012 17382
rect 16036 17380 16092 17382
rect 16116 17380 16172 17382
rect 16196 17380 16252 17382
rect 16578 17448 16634 17504
rect 16302 16496 16358 16552
rect 15956 16346 16012 16348
rect 16036 16346 16092 16348
rect 16116 16346 16172 16348
rect 16196 16346 16252 16348
rect 15956 16294 15982 16346
rect 15982 16294 16012 16346
rect 16036 16294 16046 16346
rect 16046 16294 16092 16346
rect 16116 16294 16162 16346
rect 16162 16294 16172 16346
rect 16196 16294 16226 16346
rect 16226 16294 16252 16346
rect 15956 16292 16012 16294
rect 16036 16292 16092 16294
rect 16116 16292 16172 16294
rect 16196 16292 16252 16294
rect 16854 16768 16910 16824
rect 15956 15258 16012 15260
rect 16036 15258 16092 15260
rect 16116 15258 16172 15260
rect 16196 15258 16252 15260
rect 15956 15206 15982 15258
rect 15982 15206 16012 15258
rect 16036 15206 16046 15258
rect 16046 15206 16092 15258
rect 16116 15206 16162 15258
rect 16162 15206 16172 15258
rect 16196 15206 16226 15258
rect 16226 15206 16252 15258
rect 15956 15204 16012 15206
rect 16036 15204 16092 15206
rect 16116 15204 16172 15206
rect 16196 15204 16252 15206
rect 15566 13676 15568 13696
rect 15568 13676 15620 13696
rect 15620 13676 15622 13696
rect 15566 13640 15622 13676
rect 15290 13096 15346 13152
rect 15198 12552 15254 12608
rect 15474 12824 15530 12880
rect 15290 12144 15346 12200
rect 14738 12008 14794 12064
rect 12898 11872 12954 11928
rect 11978 10104 12034 10160
rect 11518 7248 11574 7304
rect 10956 7098 11012 7100
rect 11036 7098 11092 7100
rect 11116 7098 11172 7100
rect 11196 7098 11252 7100
rect 10956 7046 10982 7098
rect 10982 7046 11012 7098
rect 11036 7046 11046 7098
rect 11046 7046 11092 7098
rect 11116 7046 11162 7098
rect 11162 7046 11172 7098
rect 11196 7046 11226 7098
rect 11226 7046 11252 7098
rect 10956 7044 11012 7046
rect 11036 7044 11092 7046
rect 11116 7044 11172 7046
rect 11196 7044 11252 7046
rect 10956 6010 11012 6012
rect 11036 6010 11092 6012
rect 11116 6010 11172 6012
rect 11196 6010 11252 6012
rect 10956 5958 10982 6010
rect 10982 5958 11012 6010
rect 11036 5958 11046 6010
rect 11046 5958 11092 6010
rect 11116 5958 11162 6010
rect 11162 5958 11172 6010
rect 11196 5958 11226 6010
rect 11226 5958 11252 6010
rect 10956 5956 11012 5958
rect 11036 5956 11092 5958
rect 11116 5956 11172 5958
rect 11196 5956 11252 5958
rect 14278 11736 14334 11792
rect 14278 10784 14334 10840
rect 15956 14170 16012 14172
rect 16036 14170 16092 14172
rect 16116 14170 16172 14172
rect 16196 14170 16252 14172
rect 15956 14118 15982 14170
rect 15982 14118 16012 14170
rect 16036 14118 16046 14170
rect 16046 14118 16092 14170
rect 16116 14118 16162 14170
rect 16162 14118 16172 14170
rect 16196 14118 16226 14170
rect 16226 14118 16252 14170
rect 15956 14116 16012 14118
rect 16036 14116 16092 14118
rect 16116 14116 16172 14118
rect 16196 14116 16252 14118
rect 16026 13504 16082 13560
rect 15956 13082 16012 13084
rect 16036 13082 16092 13084
rect 16116 13082 16172 13084
rect 16196 13082 16252 13084
rect 15956 13030 15982 13082
rect 15982 13030 16012 13082
rect 16036 13030 16046 13082
rect 16046 13030 16092 13082
rect 16116 13030 16162 13082
rect 16162 13030 16172 13082
rect 16196 13030 16226 13082
rect 16226 13030 16252 13082
rect 15956 13028 16012 13030
rect 16036 13028 16092 13030
rect 16116 13028 16172 13030
rect 16196 13028 16252 13030
rect 16210 12824 16266 12880
rect 15658 12688 15714 12744
rect 15842 12552 15898 12608
rect 15934 12300 15990 12336
rect 15934 12280 15936 12300
rect 15936 12280 15988 12300
rect 15988 12280 15990 12300
rect 15956 11994 16012 11996
rect 16036 11994 16092 11996
rect 16116 11994 16172 11996
rect 16196 11994 16252 11996
rect 15956 11942 15982 11994
rect 15982 11942 16012 11994
rect 16036 11942 16046 11994
rect 16046 11942 16092 11994
rect 16116 11942 16162 11994
rect 16162 11942 16172 11994
rect 16196 11942 16226 11994
rect 16226 11942 16252 11994
rect 15956 11940 16012 11942
rect 16036 11940 16092 11942
rect 16116 11940 16172 11942
rect 16196 11940 16252 11942
rect 17958 19896 18014 19952
rect 17498 16632 17554 16688
rect 20350 20596 20406 20632
rect 20350 20576 20352 20596
rect 20352 20576 20404 20596
rect 20404 20576 20406 20596
rect 19154 19252 19156 19272
rect 19156 19252 19208 19272
rect 19208 19252 19210 19272
rect 19154 19216 19210 19252
rect 19430 18808 19486 18864
rect 19062 18148 19118 18184
rect 19062 18128 19064 18148
rect 19064 18128 19116 18148
rect 19116 18128 19118 18148
rect 19430 18028 19432 18048
rect 19432 18028 19484 18048
rect 19484 18028 19486 18048
rect 19430 17992 19486 18028
rect 19154 17720 19210 17776
rect 17498 13776 17554 13832
rect 16486 12688 16542 12744
rect 16578 12280 16634 12336
rect 16670 12008 16726 12064
rect 15956 10906 16012 10908
rect 16036 10906 16092 10908
rect 16116 10906 16172 10908
rect 16196 10906 16252 10908
rect 15956 10854 15982 10906
rect 15982 10854 16012 10906
rect 16036 10854 16046 10906
rect 16046 10854 16092 10906
rect 16116 10854 16162 10906
rect 16162 10854 16172 10906
rect 16196 10854 16226 10906
rect 16226 10854 16252 10906
rect 15956 10852 16012 10854
rect 16036 10852 16092 10854
rect 16116 10852 16172 10854
rect 16196 10852 16252 10854
rect 15956 9818 16012 9820
rect 16036 9818 16092 9820
rect 16116 9818 16172 9820
rect 16196 9818 16252 9820
rect 15956 9766 15982 9818
rect 15982 9766 16012 9818
rect 16036 9766 16046 9818
rect 16046 9766 16092 9818
rect 16116 9766 16162 9818
rect 16162 9766 16172 9818
rect 16196 9766 16226 9818
rect 16226 9766 16252 9818
rect 15956 9764 16012 9766
rect 16036 9764 16092 9766
rect 16116 9764 16172 9766
rect 16196 9764 16252 9766
rect 15750 9696 15806 9752
rect 15934 9424 15990 9480
rect 15956 8730 16012 8732
rect 16036 8730 16092 8732
rect 16116 8730 16172 8732
rect 16196 8730 16252 8732
rect 15956 8678 15982 8730
rect 15982 8678 16012 8730
rect 16036 8678 16046 8730
rect 16046 8678 16092 8730
rect 16116 8678 16162 8730
rect 16162 8678 16172 8730
rect 16196 8678 16226 8730
rect 16226 8678 16252 8730
rect 15956 8676 16012 8678
rect 16036 8676 16092 8678
rect 16116 8676 16172 8678
rect 16196 8676 16252 8678
rect 16486 9288 16542 9344
rect 16578 9152 16634 9208
rect 15956 7642 16012 7644
rect 16036 7642 16092 7644
rect 16116 7642 16172 7644
rect 16196 7642 16252 7644
rect 15956 7590 15982 7642
rect 15982 7590 16012 7642
rect 16036 7590 16046 7642
rect 16046 7590 16092 7642
rect 16116 7590 16162 7642
rect 16162 7590 16172 7642
rect 16196 7590 16226 7642
rect 16226 7590 16252 7642
rect 15956 7588 16012 7590
rect 16036 7588 16092 7590
rect 16116 7588 16172 7590
rect 16196 7588 16252 7590
rect 12898 5208 12954 5264
rect 10956 4922 11012 4924
rect 11036 4922 11092 4924
rect 11116 4922 11172 4924
rect 11196 4922 11252 4924
rect 10956 4870 10982 4922
rect 10982 4870 11012 4922
rect 11036 4870 11046 4922
rect 11046 4870 11092 4922
rect 11116 4870 11162 4922
rect 11162 4870 11172 4922
rect 11196 4870 11226 4922
rect 11226 4870 11252 4922
rect 10956 4868 11012 4870
rect 11036 4868 11092 4870
rect 11116 4868 11172 4870
rect 11196 4868 11252 4870
rect 10956 3834 11012 3836
rect 11036 3834 11092 3836
rect 11116 3834 11172 3836
rect 11196 3834 11252 3836
rect 10956 3782 10982 3834
rect 10982 3782 11012 3834
rect 11036 3782 11046 3834
rect 11046 3782 11092 3834
rect 11116 3782 11162 3834
rect 11162 3782 11172 3834
rect 11196 3782 11226 3834
rect 11226 3782 11252 3834
rect 10956 3780 11012 3782
rect 11036 3780 11092 3782
rect 11116 3780 11172 3782
rect 11196 3780 11252 3782
rect 15956 6554 16012 6556
rect 16036 6554 16092 6556
rect 16116 6554 16172 6556
rect 16196 6554 16252 6556
rect 15956 6502 15982 6554
rect 15982 6502 16012 6554
rect 16036 6502 16046 6554
rect 16046 6502 16092 6554
rect 16116 6502 16162 6554
rect 16162 6502 16172 6554
rect 16196 6502 16226 6554
rect 16226 6502 16252 6554
rect 15956 6500 16012 6502
rect 16036 6500 16092 6502
rect 16116 6500 16172 6502
rect 16196 6500 16252 6502
rect 18142 15000 18198 15056
rect 19338 17312 19394 17368
rect 19154 17040 19210 17096
rect 20956 20154 21012 20156
rect 21036 20154 21092 20156
rect 21116 20154 21172 20156
rect 21196 20154 21252 20156
rect 20956 20102 20982 20154
rect 20982 20102 21012 20154
rect 21036 20102 21046 20154
rect 21046 20102 21092 20154
rect 21116 20102 21162 20154
rect 21162 20102 21172 20154
rect 21196 20102 21226 20154
rect 21226 20102 21252 20154
rect 20956 20100 21012 20102
rect 21036 20100 21092 20102
rect 21116 20100 21172 20102
rect 21196 20100 21252 20102
rect 20718 19216 20774 19272
rect 20956 19066 21012 19068
rect 21036 19066 21092 19068
rect 21116 19066 21172 19068
rect 21196 19066 21252 19068
rect 20956 19014 20982 19066
rect 20982 19014 21012 19066
rect 21036 19014 21046 19066
rect 21046 19014 21092 19066
rect 21116 19014 21162 19066
rect 21162 19014 21172 19066
rect 21196 19014 21226 19066
rect 21226 19014 21252 19066
rect 20956 19012 21012 19014
rect 21036 19012 21092 19014
rect 21116 19012 21172 19014
rect 21196 19012 21252 19014
rect 19982 18300 19984 18320
rect 19984 18300 20036 18320
rect 20036 18300 20038 18320
rect 19982 18264 20038 18300
rect 18786 15816 18842 15872
rect 18970 15816 19026 15872
rect 18694 15136 18750 15192
rect 18602 15000 18658 15056
rect 18510 13640 18566 13696
rect 17130 10512 17186 10568
rect 17222 10104 17278 10160
rect 17406 10124 17462 10160
rect 17406 10104 17408 10124
rect 17408 10104 17460 10124
rect 17460 10104 17462 10124
rect 17222 9696 17278 9752
rect 16854 9580 16910 9616
rect 16854 9560 16856 9580
rect 16856 9560 16908 9580
rect 16908 9560 16910 9580
rect 18418 11328 18474 11384
rect 17406 9016 17462 9072
rect 18510 9288 18566 9344
rect 19338 16088 19394 16144
rect 19982 15852 19984 15872
rect 19984 15852 20036 15872
rect 20036 15852 20038 15872
rect 19982 15816 20038 15852
rect 19338 15544 19394 15600
rect 19154 14864 19210 14920
rect 19246 13912 19302 13968
rect 19430 13776 19486 13832
rect 19890 14592 19946 14648
rect 19706 14476 19762 14512
rect 19706 14456 19708 14476
rect 19708 14456 19760 14476
rect 19760 14456 19762 14476
rect 20074 14068 20130 14104
rect 20074 14048 20076 14068
rect 20076 14048 20128 14068
rect 20128 14048 20130 14068
rect 19614 13640 19670 13696
rect 21546 20576 21602 20632
rect 20956 17978 21012 17980
rect 21036 17978 21092 17980
rect 21116 17978 21172 17980
rect 21196 17978 21252 17980
rect 20956 17926 20982 17978
rect 20982 17926 21012 17978
rect 21036 17926 21046 17978
rect 21046 17926 21092 17978
rect 21116 17926 21162 17978
rect 21162 17926 21172 17978
rect 21196 17926 21226 17978
rect 21226 17926 21252 17978
rect 20956 17924 21012 17926
rect 21036 17924 21092 17926
rect 21116 17924 21172 17926
rect 21196 17924 21252 17926
rect 20956 16890 21012 16892
rect 21036 16890 21092 16892
rect 21116 16890 21172 16892
rect 21196 16890 21252 16892
rect 20956 16838 20982 16890
rect 20982 16838 21012 16890
rect 21036 16838 21046 16890
rect 21046 16838 21092 16890
rect 21116 16838 21162 16890
rect 21162 16838 21172 16890
rect 21196 16838 21226 16890
rect 21226 16838 21252 16890
rect 20956 16836 21012 16838
rect 21036 16836 21092 16838
rect 21116 16836 21172 16838
rect 21196 16836 21252 16838
rect 20718 15408 20774 15464
rect 20350 14184 20406 14240
rect 19614 12960 19670 13016
rect 19706 12824 19762 12880
rect 18602 8336 18658 8392
rect 19246 8608 19302 8664
rect 19246 8336 19302 8392
rect 19062 7828 19064 7848
rect 19064 7828 19116 7848
rect 19116 7828 19118 7848
rect 19062 7792 19118 7828
rect 19522 8744 19578 8800
rect 19522 7792 19578 7848
rect 16762 6296 16818 6352
rect 15956 5466 16012 5468
rect 16036 5466 16092 5468
rect 16116 5466 16172 5468
rect 16196 5466 16252 5468
rect 15956 5414 15982 5466
rect 15982 5414 16012 5466
rect 16036 5414 16046 5466
rect 16046 5414 16092 5466
rect 16116 5414 16162 5466
rect 16162 5414 16172 5466
rect 16196 5414 16226 5466
rect 16226 5414 16252 5466
rect 15956 5412 16012 5414
rect 16036 5412 16092 5414
rect 16116 5412 16172 5414
rect 16196 5412 16252 5414
rect 15956 4378 16012 4380
rect 16036 4378 16092 4380
rect 16116 4378 16172 4380
rect 16196 4378 16252 4380
rect 15956 4326 15982 4378
rect 15982 4326 16012 4378
rect 16036 4326 16046 4378
rect 16046 4326 16092 4378
rect 16116 4326 16162 4378
rect 16162 4326 16172 4378
rect 16196 4326 16226 4378
rect 16226 4326 16252 4378
rect 15956 4324 16012 4326
rect 16036 4324 16092 4326
rect 16116 4324 16172 4326
rect 16196 4324 16252 4326
rect 15566 3440 15622 3496
rect 15956 3290 16012 3292
rect 16036 3290 16092 3292
rect 16116 3290 16172 3292
rect 16196 3290 16252 3292
rect 15956 3238 15982 3290
rect 15982 3238 16012 3290
rect 16036 3238 16046 3290
rect 16046 3238 16092 3290
rect 16116 3238 16162 3290
rect 16162 3238 16172 3290
rect 16196 3238 16226 3290
rect 16226 3238 16252 3290
rect 15956 3236 16012 3238
rect 16036 3236 16092 3238
rect 16116 3236 16172 3238
rect 16196 3236 16252 3238
rect 10956 2746 11012 2748
rect 11036 2746 11092 2748
rect 11116 2746 11172 2748
rect 11196 2746 11252 2748
rect 10956 2694 10982 2746
rect 10982 2694 11012 2746
rect 11036 2694 11046 2746
rect 11046 2694 11092 2746
rect 11116 2694 11162 2746
rect 11162 2694 11172 2746
rect 11196 2694 11226 2746
rect 11226 2694 11252 2746
rect 10956 2692 11012 2694
rect 11036 2692 11092 2694
rect 11116 2692 11172 2694
rect 11196 2692 11252 2694
rect 7470 2352 7526 2408
rect 11150 2352 11206 2408
rect 5956 2202 6012 2204
rect 6036 2202 6092 2204
rect 6116 2202 6172 2204
rect 6196 2202 6252 2204
rect 5956 2150 5982 2202
rect 5982 2150 6012 2202
rect 6036 2150 6046 2202
rect 6046 2150 6092 2202
rect 6116 2150 6162 2202
rect 6162 2150 6172 2202
rect 6196 2150 6226 2202
rect 6226 2150 6252 2202
rect 5956 2148 6012 2150
rect 6036 2148 6092 2150
rect 6116 2148 6172 2150
rect 6196 2148 6252 2150
rect 15956 2202 16012 2204
rect 16036 2202 16092 2204
rect 16116 2202 16172 2204
rect 16196 2202 16252 2204
rect 15956 2150 15982 2202
rect 15982 2150 16012 2202
rect 16036 2150 16046 2202
rect 16046 2150 16092 2202
rect 16116 2150 16162 2202
rect 16162 2150 16172 2202
rect 16196 2150 16226 2202
rect 16226 2150 16252 2202
rect 15956 2148 16012 2150
rect 16036 2148 16092 2150
rect 16116 2148 16172 2150
rect 16196 2148 16252 2150
rect 19246 7248 19302 7304
rect 20074 10920 20130 10976
rect 20626 13504 20682 13560
rect 20956 15802 21012 15804
rect 21036 15802 21092 15804
rect 21116 15802 21172 15804
rect 21196 15802 21252 15804
rect 20956 15750 20982 15802
rect 20982 15750 21012 15802
rect 21036 15750 21046 15802
rect 21046 15750 21092 15802
rect 21116 15750 21162 15802
rect 21162 15750 21172 15802
rect 21196 15750 21226 15802
rect 21226 15750 21252 15802
rect 20956 15748 21012 15750
rect 21036 15748 21092 15750
rect 21116 15748 21172 15750
rect 21196 15748 21252 15750
rect 21454 16224 21510 16280
rect 21362 15408 21418 15464
rect 20956 14714 21012 14716
rect 21036 14714 21092 14716
rect 21116 14714 21172 14716
rect 21196 14714 21252 14716
rect 20956 14662 20982 14714
rect 20982 14662 21012 14714
rect 21036 14662 21046 14714
rect 21046 14662 21092 14714
rect 21116 14662 21162 14714
rect 21162 14662 21172 14714
rect 21196 14662 21226 14714
rect 21226 14662 21252 14714
rect 20956 14660 21012 14662
rect 21036 14660 21092 14662
rect 21116 14660 21172 14662
rect 21196 14660 21252 14662
rect 20534 13368 20590 13424
rect 20718 13096 20774 13152
rect 20956 13626 21012 13628
rect 21036 13626 21092 13628
rect 21116 13626 21172 13628
rect 21196 13626 21252 13628
rect 20956 13574 20982 13626
rect 20982 13574 21012 13626
rect 21036 13574 21046 13626
rect 21046 13574 21092 13626
rect 21116 13574 21162 13626
rect 21162 13574 21172 13626
rect 21196 13574 21226 13626
rect 21226 13574 21252 13626
rect 20956 13572 21012 13574
rect 21036 13572 21092 13574
rect 21116 13572 21172 13574
rect 21196 13572 21252 13574
rect 21454 13504 21510 13560
rect 21546 13096 21602 13152
rect 21454 12688 21510 12744
rect 20956 12538 21012 12540
rect 21036 12538 21092 12540
rect 21116 12538 21172 12540
rect 21196 12538 21252 12540
rect 20956 12486 20982 12538
rect 20982 12486 21012 12538
rect 21036 12486 21046 12538
rect 21046 12486 21092 12538
rect 21116 12486 21162 12538
rect 21162 12486 21172 12538
rect 21196 12486 21226 12538
rect 21226 12486 21252 12538
rect 20956 12484 21012 12486
rect 21036 12484 21092 12486
rect 21116 12484 21172 12486
rect 21196 12484 21252 12486
rect 20994 12280 21050 12336
rect 20442 10784 20498 10840
rect 19706 8492 19762 8528
rect 20956 11450 21012 11452
rect 21036 11450 21092 11452
rect 21116 11450 21172 11452
rect 21196 11450 21252 11452
rect 20956 11398 20982 11450
rect 20982 11398 21012 11450
rect 21036 11398 21046 11450
rect 21046 11398 21092 11450
rect 21116 11398 21162 11450
rect 21162 11398 21172 11450
rect 21196 11398 21226 11450
rect 21226 11398 21252 11450
rect 20956 11396 21012 11398
rect 21036 11396 21092 11398
rect 21116 11396 21172 11398
rect 21196 11396 21252 11398
rect 20810 11328 20866 11384
rect 20956 10362 21012 10364
rect 21036 10362 21092 10364
rect 21116 10362 21172 10364
rect 21196 10362 21252 10364
rect 20956 10310 20982 10362
rect 20982 10310 21012 10362
rect 21036 10310 21046 10362
rect 21046 10310 21092 10362
rect 21116 10310 21162 10362
rect 21162 10310 21172 10362
rect 21196 10310 21226 10362
rect 21226 10310 21252 10362
rect 20956 10308 21012 10310
rect 21036 10308 21092 10310
rect 21116 10308 21172 10310
rect 21196 10308 21252 10310
rect 21546 12416 21602 12472
rect 21270 9560 21326 9616
rect 20956 9274 21012 9276
rect 21036 9274 21092 9276
rect 21116 9274 21172 9276
rect 21196 9274 21252 9276
rect 20956 9222 20982 9274
rect 20982 9222 21012 9274
rect 21036 9222 21046 9274
rect 21046 9222 21092 9274
rect 21116 9222 21162 9274
rect 21162 9222 21172 9274
rect 21196 9222 21226 9274
rect 21226 9222 21252 9274
rect 20956 9220 21012 9222
rect 21036 9220 21092 9222
rect 21116 9220 21172 9222
rect 21196 9220 21252 9222
rect 19706 8472 19708 8492
rect 19708 8472 19760 8492
rect 19760 8472 19762 8492
rect 21454 9560 21510 9616
rect 20956 8186 21012 8188
rect 21036 8186 21092 8188
rect 21116 8186 21172 8188
rect 21196 8186 21252 8188
rect 20956 8134 20982 8186
rect 20982 8134 21012 8186
rect 21036 8134 21046 8186
rect 21046 8134 21092 8186
rect 21116 8134 21162 8186
rect 21162 8134 21172 8186
rect 21196 8134 21226 8186
rect 21226 8134 21252 8186
rect 20956 8132 21012 8134
rect 21036 8132 21092 8134
rect 21116 8132 21172 8134
rect 21196 8132 21252 8134
rect 21914 19216 21970 19272
rect 21914 17484 21916 17504
rect 21916 17484 21968 17504
rect 21968 17484 21970 17504
rect 21914 17448 21970 17484
rect 23846 18672 23902 18728
rect 23110 18128 23166 18184
rect 22650 17584 22706 17640
rect 22098 17040 22154 17096
rect 22006 16632 22062 16688
rect 22006 12144 22062 12200
rect 22926 15136 22982 15192
rect 22926 13776 22982 13832
rect 22742 13368 22798 13424
rect 22650 13232 22706 13288
rect 22742 12280 22798 12336
rect 23570 16652 23626 16688
rect 23570 16632 23572 16652
rect 23572 16632 23624 16652
rect 23624 16632 23626 16652
rect 23386 15952 23442 16008
rect 23202 15020 23258 15056
rect 23202 15000 23204 15020
rect 23204 15000 23256 15020
rect 23256 15000 23258 15020
rect 23202 13524 23258 13560
rect 23202 13504 23204 13524
rect 23204 13504 23256 13524
rect 23256 13504 23258 13524
rect 23018 12008 23074 12064
rect 23662 15000 23718 15056
rect 23754 14864 23810 14920
rect 23938 16496 23994 16552
rect 23478 14068 23534 14104
rect 23478 14048 23480 14068
rect 23480 14048 23532 14068
rect 23532 14048 23534 14068
rect 22650 11600 22706 11656
rect 22466 10104 22522 10160
rect 23202 10784 23258 10840
rect 23846 10920 23902 10976
rect 25594 23024 25650 23080
rect 25870 22344 25926 22400
rect 25686 21528 25742 21584
rect 25778 21256 25834 21312
rect 25226 19896 25282 19952
rect 24490 18264 24546 18320
rect 25042 18264 25098 18320
rect 24214 17856 24270 17912
rect 23938 10784 23994 10840
rect 24214 14320 24270 14376
rect 24398 14884 24454 14920
rect 24398 14864 24400 14884
rect 24400 14864 24452 14884
rect 24452 14864 24454 14884
rect 24582 17176 24638 17232
rect 25410 20476 25412 20496
rect 25412 20476 25464 20496
rect 25464 20476 25466 20496
rect 25410 20440 25466 20476
rect 25956 21786 26012 21788
rect 26036 21786 26092 21788
rect 26116 21786 26172 21788
rect 26196 21786 26252 21788
rect 25956 21734 25982 21786
rect 25982 21734 26012 21786
rect 26036 21734 26046 21786
rect 26046 21734 26092 21786
rect 26116 21734 26162 21786
rect 26162 21734 26172 21786
rect 26196 21734 26226 21786
rect 26226 21734 26252 21786
rect 25956 21732 26012 21734
rect 26036 21732 26092 21734
rect 26116 21732 26172 21734
rect 26196 21732 26252 21734
rect 25956 20698 26012 20700
rect 26036 20698 26092 20700
rect 26116 20698 26172 20700
rect 26196 20698 26252 20700
rect 25956 20646 25982 20698
rect 25982 20646 26012 20698
rect 26036 20646 26046 20698
rect 26046 20646 26092 20698
rect 26116 20646 26162 20698
rect 26162 20646 26172 20698
rect 26196 20646 26226 20698
rect 26226 20646 26252 20698
rect 25956 20644 26012 20646
rect 26036 20644 26092 20646
rect 26116 20644 26172 20646
rect 26196 20644 26252 20646
rect 27158 20440 27214 20496
rect 25318 18536 25374 18592
rect 25502 18264 25558 18320
rect 24950 15680 25006 15736
rect 24674 15564 24730 15600
rect 24674 15544 24676 15564
rect 24676 15544 24728 15564
rect 24728 15544 24730 15564
rect 24858 15408 24914 15464
rect 24766 15000 24822 15056
rect 24674 13812 24676 13832
rect 24676 13812 24728 13832
rect 24728 13812 24730 13832
rect 24674 13776 24730 13812
rect 24582 12552 24638 12608
rect 24582 12144 24638 12200
rect 24122 10648 24178 10704
rect 24398 10376 24454 10432
rect 25410 15544 25466 15600
rect 25042 14592 25098 14648
rect 24950 13504 25006 13560
rect 24858 11736 24914 11792
rect 24950 10920 25006 10976
rect 24950 10512 25006 10568
rect 24582 9560 24638 9616
rect 24214 9460 24216 9480
rect 24216 9460 24268 9480
rect 24268 9460 24270 9480
rect 24214 9424 24270 9460
rect 24398 9324 24400 9344
rect 24400 9324 24452 9344
rect 24452 9324 24454 9344
rect 24398 9288 24454 9324
rect 23202 9152 23258 9208
rect 20956 7098 21012 7100
rect 21036 7098 21092 7100
rect 21116 7098 21172 7100
rect 21196 7098 21252 7100
rect 20956 7046 20982 7098
rect 20982 7046 21012 7098
rect 21036 7046 21046 7098
rect 21046 7046 21092 7098
rect 21116 7046 21162 7098
rect 21162 7046 21172 7098
rect 21196 7046 21226 7098
rect 21226 7046 21252 7098
rect 20956 7044 21012 7046
rect 21036 7044 21092 7046
rect 21116 7044 21172 7046
rect 21196 7044 21252 7046
rect 20956 6010 21012 6012
rect 21036 6010 21092 6012
rect 21116 6010 21172 6012
rect 21196 6010 21252 6012
rect 20956 5958 20982 6010
rect 20982 5958 21012 6010
rect 21036 5958 21046 6010
rect 21046 5958 21092 6010
rect 21116 5958 21162 6010
rect 21162 5958 21172 6010
rect 21196 5958 21226 6010
rect 21226 5958 21252 6010
rect 20956 5956 21012 5958
rect 21036 5956 21092 5958
rect 21116 5956 21172 5958
rect 21196 5956 21252 5958
rect 20956 4922 21012 4924
rect 21036 4922 21092 4924
rect 21116 4922 21172 4924
rect 21196 4922 21252 4924
rect 20956 4870 20982 4922
rect 20982 4870 21012 4922
rect 21036 4870 21046 4922
rect 21046 4870 21092 4922
rect 21116 4870 21162 4922
rect 21162 4870 21172 4922
rect 21196 4870 21226 4922
rect 21226 4870 21252 4922
rect 20956 4868 21012 4870
rect 21036 4868 21092 4870
rect 21116 4868 21172 4870
rect 21196 4868 21252 4870
rect 19890 3984 19946 4040
rect 20956 3834 21012 3836
rect 21036 3834 21092 3836
rect 21116 3834 21172 3836
rect 21196 3834 21252 3836
rect 20956 3782 20982 3834
rect 20982 3782 21012 3834
rect 21036 3782 21046 3834
rect 21046 3782 21092 3834
rect 21116 3782 21162 3834
rect 21162 3782 21172 3834
rect 21196 3782 21226 3834
rect 21226 3782 21252 3834
rect 20956 3780 21012 3782
rect 21036 3780 21092 3782
rect 21116 3780 21172 3782
rect 21196 3780 21252 3782
rect 20956 2746 21012 2748
rect 21036 2746 21092 2748
rect 21116 2746 21172 2748
rect 21196 2746 21252 2748
rect 20956 2694 20982 2746
rect 20982 2694 21012 2746
rect 21036 2694 21046 2746
rect 21046 2694 21092 2746
rect 21116 2694 21162 2746
rect 21162 2694 21172 2746
rect 21196 2694 21226 2746
rect 21226 2694 21252 2746
rect 20956 2692 21012 2694
rect 21036 2692 21092 2694
rect 21116 2692 21172 2694
rect 21196 2692 21252 2694
rect 25594 17756 25596 17776
rect 25596 17756 25648 17776
rect 25648 17756 25650 17776
rect 25594 17720 25650 17756
rect 25956 19610 26012 19612
rect 26036 19610 26092 19612
rect 26116 19610 26172 19612
rect 26196 19610 26252 19612
rect 25956 19558 25982 19610
rect 25982 19558 26012 19610
rect 26036 19558 26046 19610
rect 26046 19558 26092 19610
rect 26116 19558 26162 19610
rect 26162 19558 26172 19610
rect 26196 19558 26226 19610
rect 26226 19558 26252 19610
rect 25956 19556 26012 19558
rect 26036 19556 26092 19558
rect 26116 19556 26172 19558
rect 26196 19556 26252 19558
rect 25956 18522 26012 18524
rect 26036 18522 26092 18524
rect 26116 18522 26172 18524
rect 26196 18522 26252 18524
rect 25956 18470 25982 18522
rect 25982 18470 26012 18522
rect 26036 18470 26046 18522
rect 26046 18470 26092 18522
rect 26116 18470 26162 18522
rect 26162 18470 26172 18522
rect 26196 18470 26226 18522
rect 26226 18470 26252 18522
rect 25956 18468 26012 18470
rect 26036 18468 26092 18470
rect 26116 18468 26172 18470
rect 26196 18468 26252 18470
rect 25956 17434 26012 17436
rect 26036 17434 26092 17436
rect 26116 17434 26172 17436
rect 26196 17434 26252 17436
rect 25956 17382 25982 17434
rect 25982 17382 26012 17434
rect 26036 17382 26046 17434
rect 26046 17382 26092 17434
rect 26116 17382 26162 17434
rect 26162 17382 26172 17434
rect 26196 17382 26226 17434
rect 26226 17382 26252 17434
rect 25956 17380 26012 17382
rect 26036 17380 26092 17382
rect 26116 17380 26172 17382
rect 26196 17380 26252 17382
rect 25778 15952 25834 16008
rect 25686 13640 25742 13696
rect 25594 13504 25650 13560
rect 25502 11056 25558 11112
rect 25226 10920 25282 10976
rect 25226 10784 25282 10840
rect 25318 9968 25374 10024
rect 25318 9036 25374 9072
rect 25318 9016 25320 9036
rect 25320 9016 25372 9036
rect 25372 9016 25374 9036
rect 25042 8744 25098 8800
rect 25686 10648 25742 10704
rect 25502 8472 25558 8528
rect 25502 8064 25558 8120
rect 25956 16346 26012 16348
rect 26036 16346 26092 16348
rect 26116 16346 26172 16348
rect 26196 16346 26252 16348
rect 25956 16294 25982 16346
rect 25982 16294 26012 16346
rect 26036 16294 26046 16346
rect 26046 16294 26092 16346
rect 26116 16294 26162 16346
rect 26162 16294 26172 16346
rect 26196 16294 26226 16346
rect 26226 16294 26252 16346
rect 25956 16292 26012 16294
rect 26036 16292 26092 16294
rect 26116 16292 26172 16294
rect 26196 16292 26252 16294
rect 25962 16124 25964 16144
rect 25964 16124 26016 16144
rect 26016 16124 26018 16144
rect 25962 16088 26018 16124
rect 26330 15952 26386 16008
rect 25956 15258 26012 15260
rect 26036 15258 26092 15260
rect 26116 15258 26172 15260
rect 26196 15258 26252 15260
rect 25956 15206 25982 15258
rect 25982 15206 26012 15258
rect 26036 15206 26046 15258
rect 26046 15206 26092 15258
rect 26116 15206 26162 15258
rect 26162 15206 26172 15258
rect 26196 15206 26226 15258
rect 26226 15206 26252 15258
rect 25956 15204 26012 15206
rect 26036 15204 26092 15206
rect 26116 15204 26172 15206
rect 26196 15204 26252 15206
rect 25956 14170 26012 14172
rect 26036 14170 26092 14172
rect 26116 14170 26172 14172
rect 26196 14170 26252 14172
rect 25956 14118 25982 14170
rect 25982 14118 26012 14170
rect 26036 14118 26046 14170
rect 26046 14118 26092 14170
rect 26116 14118 26162 14170
rect 26162 14118 26172 14170
rect 26196 14118 26226 14170
rect 26226 14118 26252 14170
rect 25956 14116 26012 14118
rect 26036 14116 26092 14118
rect 26116 14116 26172 14118
rect 26196 14116 26252 14118
rect 26514 14048 26570 14104
rect 26514 13504 26570 13560
rect 25956 13082 26012 13084
rect 26036 13082 26092 13084
rect 26116 13082 26172 13084
rect 26196 13082 26252 13084
rect 25956 13030 25982 13082
rect 25982 13030 26012 13082
rect 26036 13030 26046 13082
rect 26046 13030 26092 13082
rect 26116 13030 26162 13082
rect 26162 13030 26172 13082
rect 26196 13030 26226 13082
rect 26226 13030 26252 13082
rect 25956 13028 26012 13030
rect 26036 13028 26092 13030
rect 26116 13028 26172 13030
rect 26196 13028 26252 13030
rect 25956 11994 26012 11996
rect 26036 11994 26092 11996
rect 26116 11994 26172 11996
rect 26196 11994 26252 11996
rect 25956 11942 25982 11994
rect 25982 11942 26012 11994
rect 26036 11942 26046 11994
rect 26046 11942 26092 11994
rect 26116 11942 26162 11994
rect 26162 11942 26172 11994
rect 26196 11942 26226 11994
rect 26226 11942 26252 11994
rect 25956 11940 26012 11942
rect 26036 11940 26092 11942
rect 26116 11940 26172 11942
rect 26196 11940 26252 11942
rect 26422 12552 26478 12608
rect 25956 10906 26012 10908
rect 26036 10906 26092 10908
rect 26116 10906 26172 10908
rect 26196 10906 26252 10908
rect 25956 10854 25982 10906
rect 25982 10854 26012 10906
rect 26036 10854 26046 10906
rect 26046 10854 26092 10906
rect 26116 10854 26162 10906
rect 26162 10854 26172 10906
rect 26196 10854 26226 10906
rect 26226 10854 26252 10906
rect 25956 10852 26012 10854
rect 26036 10852 26092 10854
rect 26116 10852 26172 10854
rect 26196 10852 26252 10854
rect 27526 20032 27582 20088
rect 26974 18808 27030 18864
rect 27250 17992 27306 18048
rect 27618 18808 27674 18864
rect 27618 17176 27674 17232
rect 26882 16496 26938 16552
rect 26974 16088 27030 16144
rect 28078 16496 28134 16552
rect 27158 15544 27214 15600
rect 26790 14456 26846 14512
rect 26698 13776 26754 13832
rect 26606 12416 26662 12472
rect 26882 14320 26938 14376
rect 27342 14864 27398 14920
rect 26974 13948 26976 13968
rect 26976 13948 27028 13968
rect 27028 13948 27030 13968
rect 26974 13912 27030 13948
rect 27342 12824 27398 12880
rect 26974 11736 27030 11792
rect 26974 10512 27030 10568
rect 25956 9818 26012 9820
rect 26036 9818 26092 9820
rect 26116 9818 26172 9820
rect 26196 9818 26252 9820
rect 25956 9766 25982 9818
rect 25982 9766 26012 9818
rect 26036 9766 26046 9818
rect 26046 9766 26092 9818
rect 26116 9766 26162 9818
rect 26162 9766 26172 9818
rect 26196 9766 26226 9818
rect 26226 9766 26252 9818
rect 25956 9764 26012 9766
rect 26036 9764 26092 9766
rect 26116 9764 26172 9766
rect 26196 9764 26252 9766
rect 26422 9152 26478 9208
rect 25956 8730 26012 8732
rect 26036 8730 26092 8732
rect 26116 8730 26172 8732
rect 26196 8730 26252 8732
rect 25956 8678 25982 8730
rect 25982 8678 26012 8730
rect 26036 8678 26046 8730
rect 26046 8678 26092 8730
rect 26116 8678 26162 8730
rect 26162 8678 26172 8730
rect 26196 8678 26226 8730
rect 26226 8678 26252 8730
rect 25956 8676 26012 8678
rect 26036 8676 26092 8678
rect 26116 8676 26172 8678
rect 26196 8676 26252 8678
rect 26514 8880 26570 8936
rect 25956 7642 26012 7644
rect 26036 7642 26092 7644
rect 26116 7642 26172 7644
rect 26196 7642 26252 7644
rect 25956 7590 25982 7642
rect 25982 7590 26012 7642
rect 26036 7590 26046 7642
rect 26046 7590 26092 7642
rect 26116 7590 26162 7642
rect 26162 7590 26172 7642
rect 26196 7590 26226 7642
rect 26226 7590 26252 7642
rect 25956 7588 26012 7590
rect 26036 7588 26092 7590
rect 26116 7588 26172 7590
rect 26196 7588 26252 7590
rect 26606 7384 26662 7440
rect 26514 7248 26570 7304
rect 25956 6554 26012 6556
rect 26036 6554 26092 6556
rect 26116 6554 26172 6556
rect 26196 6554 26252 6556
rect 25956 6502 25982 6554
rect 25982 6502 26012 6554
rect 26036 6502 26046 6554
rect 26046 6502 26092 6554
rect 26116 6502 26162 6554
rect 26162 6502 26172 6554
rect 26196 6502 26226 6554
rect 26226 6502 26252 6554
rect 25956 6500 26012 6502
rect 26036 6500 26092 6502
rect 26116 6500 26172 6502
rect 26196 6500 26252 6502
rect 25956 5466 26012 5468
rect 26036 5466 26092 5468
rect 26116 5466 26172 5468
rect 26196 5466 26252 5468
rect 25956 5414 25982 5466
rect 25982 5414 26012 5466
rect 26036 5414 26046 5466
rect 26046 5414 26092 5466
rect 26116 5414 26162 5466
rect 26162 5414 26172 5466
rect 26196 5414 26226 5466
rect 26226 5414 26252 5466
rect 25956 5412 26012 5414
rect 26036 5412 26092 5414
rect 26116 5412 26172 5414
rect 26196 5412 26252 5414
rect 26698 6296 26754 6352
rect 26422 5208 26478 5264
rect 26606 5072 26662 5128
rect 25778 4528 25834 4584
rect 25686 3848 25742 3904
rect 25594 3440 25650 3496
rect 25410 2352 25466 2408
rect 25956 4378 26012 4380
rect 26036 4378 26092 4380
rect 26116 4378 26172 4380
rect 26196 4378 26252 4380
rect 25956 4326 25982 4378
rect 25982 4326 26012 4378
rect 26036 4326 26046 4378
rect 26046 4326 26092 4378
rect 26116 4326 26162 4378
rect 26162 4326 26172 4378
rect 26196 4326 26226 4378
rect 26226 4326 26252 4378
rect 25956 4324 26012 4326
rect 26036 4324 26092 4326
rect 26116 4324 26172 4326
rect 26196 4324 26252 4326
rect 26422 3984 26478 4040
rect 25956 3290 26012 3292
rect 26036 3290 26092 3292
rect 26116 3290 26172 3292
rect 26196 3290 26252 3292
rect 25956 3238 25982 3290
rect 25982 3238 26012 3290
rect 26036 3238 26046 3290
rect 26046 3238 26092 3290
rect 26116 3238 26162 3290
rect 26162 3238 26172 3290
rect 26196 3238 26226 3290
rect 26226 3238 26252 3290
rect 25956 3236 26012 3238
rect 26036 3236 26092 3238
rect 26116 3236 26172 3238
rect 26196 3236 26252 3238
rect 26606 2796 26608 2816
rect 26608 2796 26660 2816
rect 26660 2796 26662 2816
rect 26606 2760 26662 2796
rect 25956 2202 26012 2204
rect 26036 2202 26092 2204
rect 26116 2202 26172 2204
rect 26196 2202 26252 2204
rect 25956 2150 25982 2202
rect 25982 2150 26012 2202
rect 26036 2150 26046 2202
rect 26046 2150 26092 2202
rect 26116 2150 26162 2202
rect 26162 2150 26172 2202
rect 26196 2150 26226 2202
rect 26226 2150 26252 2202
rect 25956 2148 26012 2150
rect 26036 2148 26092 2150
rect 26116 2148 26172 2150
rect 26196 2148 26252 2150
rect 25870 1400 25926 1456
rect 4066 312 4122 368
rect 27618 14320 27674 14376
rect 27526 12824 27582 12880
rect 27434 12280 27490 12336
rect 27342 10648 27398 10704
rect 27342 10104 27398 10160
rect 27526 9560 27582 9616
rect 27710 9560 27766 9616
rect 27710 6976 27766 7032
rect 27802 5616 27858 5672
rect 26882 856 26938 912
rect 26790 312 26846 368
<< metal3 >>
rect 0 23626 480 23656
rect 3509 23626 3575 23629
rect 0 23624 3575 23626
rect 0 23568 3514 23624
rect 3570 23568 3575 23624
rect 0 23566 3575 23568
rect 0 23536 480 23566
rect 3509 23563 3575 23566
rect 25037 23626 25103 23629
rect 29520 23626 30000 23656
rect 25037 23624 30000 23626
rect 25037 23568 25042 23624
rect 25098 23568 30000 23624
rect 25037 23566 30000 23568
rect 25037 23563 25103 23566
rect 29520 23536 30000 23566
rect 0 23082 480 23112
rect 3417 23082 3483 23085
rect 0 23080 3483 23082
rect 0 23024 3422 23080
rect 3478 23024 3483 23080
rect 0 23022 3483 23024
rect 0 22992 480 23022
rect 3417 23019 3483 23022
rect 25589 23082 25655 23085
rect 29520 23082 30000 23112
rect 25589 23080 30000 23082
rect 25589 23024 25594 23080
rect 25650 23024 30000 23080
rect 25589 23022 30000 23024
rect 25589 23019 25655 23022
rect 29520 22992 30000 23022
rect 0 22402 480 22432
rect 3233 22402 3299 22405
rect 0 22400 3299 22402
rect 0 22344 3238 22400
rect 3294 22344 3299 22400
rect 0 22342 3299 22344
rect 0 22312 480 22342
rect 3233 22339 3299 22342
rect 25865 22402 25931 22405
rect 29520 22402 30000 22432
rect 25865 22400 30000 22402
rect 25865 22344 25870 22400
rect 25926 22344 30000 22400
rect 25865 22342 30000 22344
rect 25865 22339 25931 22342
rect 29520 22312 30000 22342
rect 0 21858 480 21888
rect 3785 21858 3851 21861
rect 29520 21858 30000 21888
rect 0 21856 3851 21858
rect 0 21800 3790 21856
rect 3846 21800 3851 21856
rect 0 21798 3851 21800
rect 0 21768 480 21798
rect 3785 21795 3851 21798
rect 26374 21798 30000 21858
rect 5944 21792 6264 21793
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 21727 6264 21728
rect 15944 21792 16264 21793
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 21727 16264 21728
rect 25944 21792 26264 21793
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 21727 26264 21728
rect 25681 21586 25747 21589
rect 26374 21586 26434 21798
rect 29520 21768 30000 21798
rect 25681 21584 26434 21586
rect 25681 21528 25686 21584
rect 25742 21528 26434 21584
rect 25681 21526 26434 21528
rect 25681 21523 25747 21526
rect 0 21314 480 21344
rect 4061 21314 4127 21317
rect 0 21312 4127 21314
rect 0 21256 4066 21312
rect 4122 21256 4127 21312
rect 0 21254 4127 21256
rect 0 21224 480 21254
rect 4061 21251 4127 21254
rect 25773 21314 25839 21317
rect 29520 21314 30000 21344
rect 25773 21312 30000 21314
rect 25773 21256 25778 21312
rect 25834 21256 30000 21312
rect 25773 21254 30000 21256
rect 25773 21251 25839 21254
rect 10944 21248 11264 21249
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 21183 11264 21184
rect 20944 21248 21264 21249
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 29520 21224 30000 21254
rect 20944 21183 21264 21184
rect 5944 20704 6264 20705
rect 0 20634 480 20664
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 20639 6264 20640
rect 15944 20704 16264 20705
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 20639 16264 20640
rect 25944 20704 26264 20705
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 20639 26264 20640
rect 2957 20634 3023 20637
rect 0 20632 3023 20634
rect 0 20576 2962 20632
rect 3018 20576 3023 20632
rect 0 20574 3023 20576
rect 0 20544 480 20574
rect 2957 20571 3023 20574
rect 20345 20634 20411 20637
rect 21541 20634 21607 20637
rect 29520 20634 30000 20664
rect 20345 20632 21607 20634
rect 20345 20576 20350 20632
rect 20406 20576 21546 20632
rect 21602 20576 21607 20632
rect 20345 20574 21607 20576
rect 20345 20571 20411 20574
rect 21541 20571 21607 20574
rect 27294 20574 30000 20634
rect 25405 20498 25471 20501
rect 27153 20498 27219 20501
rect 25405 20496 27219 20498
rect 25405 20440 25410 20496
rect 25466 20440 27158 20496
rect 27214 20440 27219 20496
rect 25405 20438 27219 20440
rect 25405 20435 25471 20438
rect 27153 20435 27219 20438
rect 17769 20362 17835 20365
rect 614 20360 17835 20362
rect 614 20304 17774 20360
rect 17830 20304 17835 20360
rect 614 20302 17835 20304
rect 0 20090 480 20120
rect 614 20090 674 20302
rect 17769 20299 17835 20302
rect 7373 20226 7439 20229
rect 9305 20226 9371 20229
rect 7373 20224 9371 20226
rect 7373 20168 7378 20224
rect 7434 20168 9310 20224
rect 9366 20168 9371 20224
rect 7373 20166 9371 20168
rect 7373 20163 7439 20166
rect 9305 20163 9371 20166
rect 10944 20160 11264 20161
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 20095 11264 20096
rect 20944 20160 21264 20161
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 20095 21264 20096
rect 0 20030 674 20090
rect 4429 20090 4495 20093
rect 6545 20090 6611 20093
rect 4429 20088 6611 20090
rect 4429 20032 4434 20088
rect 4490 20032 6550 20088
rect 6606 20032 6611 20088
rect 4429 20030 6611 20032
rect 0 20000 480 20030
rect 4429 20027 4495 20030
rect 6545 20027 6611 20030
rect 17953 19954 18019 19957
rect 25221 19954 25287 19957
rect 17953 19952 25287 19954
rect 17953 19896 17958 19952
rect 18014 19896 25226 19952
rect 25282 19896 25287 19952
rect 17953 19894 25287 19896
rect 17953 19891 18019 19894
rect 25221 19891 25287 19894
rect 15377 19818 15443 19821
rect 27294 19818 27354 20574
rect 29520 20544 30000 20574
rect 27521 20090 27587 20093
rect 29520 20090 30000 20120
rect 27521 20088 30000 20090
rect 27521 20032 27526 20088
rect 27582 20032 30000 20088
rect 27521 20030 30000 20032
rect 27521 20027 27587 20030
rect 29520 20000 30000 20030
rect 15377 19816 27354 19818
rect 15377 19760 15382 19816
rect 15438 19760 27354 19816
rect 15377 19758 27354 19760
rect 15377 19755 15443 19758
rect 9622 19620 9628 19684
rect 9692 19682 9698 19684
rect 14273 19682 14339 19685
rect 9692 19680 14339 19682
rect 9692 19624 14278 19680
rect 14334 19624 14339 19680
rect 9692 19622 14339 19624
rect 9692 19620 9698 19622
rect 14273 19619 14339 19622
rect 5944 19616 6264 19617
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 19551 6264 19552
rect 15944 19616 16264 19617
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 19551 16264 19552
rect 25944 19616 26264 19617
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 19551 26264 19552
rect 2405 19546 2471 19549
rect 4613 19546 4679 19549
rect 9581 19546 9647 19549
rect 2405 19544 4679 19546
rect 2405 19488 2410 19544
rect 2466 19488 4618 19544
rect 4674 19488 4679 19544
rect 2405 19486 4679 19488
rect 2405 19483 2471 19486
rect 4613 19483 4679 19486
rect 6502 19544 9647 19546
rect 6502 19488 9586 19544
rect 9642 19488 9647 19544
rect 6502 19486 9647 19488
rect 0 19410 480 19440
rect 6502 19410 6562 19486
rect 9581 19483 9647 19486
rect 0 19350 6562 19410
rect 9581 19412 9647 19413
rect 9581 19408 9628 19412
rect 9692 19410 9698 19412
rect 29520 19410 30000 19440
rect 9581 19352 9586 19408
rect 0 19320 480 19350
rect 9581 19348 9628 19352
rect 9692 19350 9774 19410
rect 25822 19350 30000 19410
rect 9692 19348 9698 19350
rect 9581 19347 9647 19348
rect 3693 19274 3759 19277
rect 6085 19274 6151 19277
rect 3693 19272 6151 19274
rect 3693 19216 3698 19272
rect 3754 19216 6090 19272
rect 6146 19216 6151 19272
rect 3693 19214 6151 19216
rect 3693 19211 3759 19214
rect 6085 19211 6151 19214
rect 9029 19274 9095 19277
rect 12065 19274 12131 19277
rect 9029 19272 12131 19274
rect 9029 19216 9034 19272
rect 9090 19216 12070 19272
rect 12126 19216 12131 19272
rect 9029 19214 12131 19216
rect 9029 19211 9095 19214
rect 12065 19211 12131 19214
rect 19149 19274 19215 19277
rect 20713 19274 20779 19277
rect 19149 19272 20779 19274
rect 19149 19216 19154 19272
rect 19210 19216 20718 19272
rect 20774 19216 20779 19272
rect 19149 19214 20779 19216
rect 19149 19211 19215 19214
rect 20713 19211 20779 19214
rect 21909 19274 21975 19277
rect 25822 19274 25882 19350
rect 29520 19320 30000 19350
rect 21909 19272 25882 19274
rect 21909 19216 21914 19272
rect 21970 19216 25882 19272
rect 21909 19214 25882 19216
rect 21909 19211 21975 19214
rect 3877 19138 3943 19141
rect 7189 19138 7255 19141
rect 3877 19136 7255 19138
rect 3877 19080 3882 19136
rect 3938 19080 7194 19136
rect 7250 19080 7255 19136
rect 3877 19078 7255 19080
rect 3877 19075 3943 19078
rect 7189 19075 7255 19078
rect 10944 19072 11264 19073
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 19007 11264 19008
rect 20944 19072 21264 19073
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 19007 21264 19008
rect 5073 19002 5139 19005
rect 7649 19002 7715 19005
rect 5073 19000 7715 19002
rect 5073 18944 5078 19000
rect 5134 18944 7654 19000
rect 7710 18944 7715 19000
rect 5073 18942 7715 18944
rect 5073 18939 5139 18942
rect 7649 18939 7715 18942
rect 11470 18942 17234 19002
rect 0 18866 480 18896
rect 3785 18866 3851 18869
rect 0 18864 3851 18866
rect 0 18808 3790 18864
rect 3846 18808 3851 18864
rect 0 18806 3851 18808
rect 0 18776 480 18806
rect 3785 18803 3851 18806
rect 10777 18866 10843 18869
rect 11470 18866 11530 18942
rect 10777 18864 11530 18866
rect 10777 18808 10782 18864
rect 10838 18808 11530 18864
rect 10777 18806 11530 18808
rect 11697 18866 11763 18869
rect 14825 18866 14891 18869
rect 11697 18864 14891 18866
rect 11697 18808 11702 18864
rect 11758 18808 14830 18864
rect 14886 18808 14891 18864
rect 11697 18806 14891 18808
rect 10777 18803 10843 18806
rect 11697 18803 11763 18806
rect 14825 18803 14891 18806
rect 7005 18730 7071 18733
rect 11789 18730 11855 18733
rect 7005 18728 11855 18730
rect 7005 18672 7010 18728
rect 7066 18672 11794 18728
rect 11850 18672 11855 18728
rect 7005 18670 11855 18672
rect 17174 18730 17234 18942
rect 19425 18866 19491 18869
rect 26969 18866 27035 18869
rect 27613 18866 27679 18869
rect 29520 18866 30000 18896
rect 19425 18864 27679 18866
rect 19425 18808 19430 18864
rect 19486 18808 26974 18864
rect 27030 18808 27618 18864
rect 27674 18808 27679 18864
rect 19425 18806 27679 18808
rect 19425 18803 19491 18806
rect 26969 18803 27035 18806
rect 27613 18803 27679 18806
rect 27846 18806 30000 18866
rect 23841 18730 23907 18733
rect 27846 18730 27906 18806
rect 29520 18776 30000 18806
rect 17174 18728 27906 18730
rect 17174 18672 23846 18728
rect 23902 18672 27906 18728
rect 17174 18670 27906 18672
rect 7005 18667 7071 18670
rect 11789 18667 11855 18670
rect 23841 18667 23907 18670
rect 8937 18594 9003 18597
rect 11697 18594 11763 18597
rect 8937 18592 11763 18594
rect 8937 18536 8942 18592
rect 8998 18536 11702 18592
rect 11758 18536 11763 18592
rect 8937 18534 11763 18536
rect 8937 18531 9003 18534
rect 11697 18531 11763 18534
rect 16389 18594 16455 18597
rect 25313 18594 25379 18597
rect 16389 18592 25379 18594
rect 16389 18536 16394 18592
rect 16450 18536 25318 18592
rect 25374 18536 25379 18592
rect 16389 18534 25379 18536
rect 16389 18531 16455 18534
rect 25313 18531 25379 18534
rect 5944 18528 6264 18529
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 18463 6264 18464
rect 15944 18528 16264 18529
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 18463 16264 18464
rect 25944 18528 26264 18529
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 18463 26264 18464
rect 11789 18458 11855 18461
rect 11789 18456 15716 18458
rect 11789 18400 11794 18456
rect 11850 18400 15716 18456
rect 11789 18398 15716 18400
rect 11789 18395 11855 18398
rect 0 18322 480 18352
rect 3509 18322 3575 18325
rect 0 18320 3575 18322
rect 0 18264 3514 18320
rect 3570 18264 3575 18320
rect 0 18262 3575 18264
rect 0 18232 480 18262
rect 3509 18259 3575 18262
rect 3693 18322 3759 18325
rect 6821 18322 6887 18325
rect 3693 18320 6887 18322
rect 3693 18264 3698 18320
rect 3754 18264 6826 18320
rect 6882 18264 6887 18320
rect 3693 18262 6887 18264
rect 3693 18259 3759 18262
rect 6821 18259 6887 18262
rect 11145 18322 11211 18325
rect 15656 18322 15716 18398
rect 19977 18322 20043 18325
rect 24485 18322 24551 18325
rect 25037 18322 25103 18325
rect 11145 18320 15578 18322
rect 11145 18264 11150 18320
rect 11206 18264 15578 18320
rect 11145 18262 15578 18264
rect 15656 18320 25103 18322
rect 15656 18264 19982 18320
rect 20038 18264 24490 18320
rect 24546 18264 25042 18320
rect 25098 18264 25103 18320
rect 15656 18262 25103 18264
rect 11145 18259 11211 18262
rect 9581 18186 9647 18189
rect 15518 18186 15578 18262
rect 19977 18259 20043 18262
rect 24485 18259 24551 18262
rect 25037 18259 25103 18262
rect 25497 18322 25563 18325
rect 29520 18322 30000 18352
rect 25497 18320 30000 18322
rect 25497 18264 25502 18320
rect 25558 18264 30000 18320
rect 25497 18262 30000 18264
rect 25497 18259 25563 18262
rect 29520 18232 30000 18262
rect 19057 18186 19123 18189
rect 23105 18186 23171 18189
rect 9581 18184 14474 18186
rect 9581 18128 9586 18184
rect 9642 18128 14474 18184
rect 9581 18126 14474 18128
rect 15518 18184 23171 18186
rect 15518 18128 19062 18184
rect 19118 18128 23110 18184
rect 23166 18128 23171 18184
rect 15518 18126 23171 18128
rect 9581 18123 9647 18126
rect 8937 18050 9003 18053
rect 10777 18050 10843 18053
rect 8937 18048 10843 18050
rect 8937 17992 8942 18048
rect 8998 17992 10782 18048
rect 10838 17992 10843 18048
rect 8937 17990 10843 17992
rect 8937 17987 9003 17990
rect 10777 17987 10843 17990
rect 10944 17984 11264 17985
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 17919 11264 17920
rect 3325 17914 3391 17917
rect 4245 17914 4311 17917
rect 3325 17912 4311 17914
rect 3325 17856 3330 17912
rect 3386 17856 4250 17912
rect 4306 17856 4311 17912
rect 3325 17854 4311 17856
rect 14414 17914 14474 18126
rect 19057 18123 19123 18126
rect 23105 18123 23171 18126
rect 15009 18050 15075 18053
rect 16665 18050 16731 18053
rect 19425 18050 19491 18053
rect 27245 18050 27311 18053
rect 15009 18048 16731 18050
rect 15009 17992 15014 18048
rect 15070 17992 16670 18048
rect 16726 17992 16731 18048
rect 15009 17990 16731 17992
rect 15009 17987 15075 17990
rect 16665 17987 16731 17990
rect 16806 18048 19491 18050
rect 16806 17992 19430 18048
rect 19486 17992 19491 18048
rect 16806 17990 19491 17992
rect 16806 17914 16866 17990
rect 19425 17987 19491 17990
rect 26006 18048 27311 18050
rect 26006 17992 27250 18048
rect 27306 17992 27311 18048
rect 26006 17990 27311 17992
rect 20944 17984 21264 17985
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 17919 21264 17920
rect 14414 17854 16866 17914
rect 24209 17914 24275 17917
rect 26006 17914 26066 17990
rect 27245 17987 27311 17990
rect 24209 17912 26066 17914
rect 24209 17856 24214 17912
rect 24270 17856 26066 17912
rect 24209 17854 26066 17856
rect 3325 17851 3391 17854
rect 4245 17851 4311 17854
rect 24209 17851 24275 17854
rect 3049 17778 3115 17781
rect 4429 17778 4495 17781
rect 3049 17776 4495 17778
rect 3049 17720 3054 17776
rect 3110 17720 4434 17776
rect 4490 17720 4495 17776
rect 3049 17718 4495 17720
rect 3049 17715 3115 17718
rect 4429 17715 4495 17718
rect 7465 17778 7531 17781
rect 8293 17778 8359 17781
rect 15653 17778 15719 17781
rect 7465 17776 15719 17778
rect 7465 17720 7470 17776
rect 7526 17720 8298 17776
rect 8354 17720 15658 17776
rect 15714 17720 15719 17776
rect 7465 17718 15719 17720
rect 7465 17715 7531 17718
rect 8293 17715 8359 17718
rect 15653 17715 15719 17718
rect 19149 17778 19215 17781
rect 25589 17778 25655 17781
rect 19149 17776 25655 17778
rect 19149 17720 19154 17776
rect 19210 17720 25594 17776
rect 25650 17720 25655 17776
rect 19149 17718 25655 17720
rect 19149 17715 19215 17718
rect 25589 17715 25655 17718
rect 0 17642 480 17672
rect 5073 17642 5139 17645
rect 0 17640 5139 17642
rect 0 17584 5078 17640
rect 5134 17584 5139 17640
rect 0 17582 5139 17584
rect 0 17552 480 17582
rect 5073 17579 5139 17582
rect 5257 17642 5323 17645
rect 11789 17642 11855 17645
rect 5257 17640 11855 17642
rect 5257 17584 5262 17640
rect 5318 17584 11794 17640
rect 11850 17584 11855 17640
rect 5257 17582 11855 17584
rect 5257 17579 5323 17582
rect 11789 17579 11855 17582
rect 22645 17642 22711 17645
rect 29520 17642 30000 17672
rect 22645 17640 30000 17642
rect 22645 17584 22650 17640
rect 22706 17584 30000 17640
rect 22645 17582 30000 17584
rect 22645 17579 22711 17582
rect 29520 17552 30000 17582
rect 16573 17506 16639 17509
rect 21909 17506 21975 17509
rect 16573 17504 21975 17506
rect 16573 17448 16578 17504
rect 16634 17448 21914 17504
rect 21970 17448 21975 17504
rect 16573 17446 21975 17448
rect 16573 17443 16639 17446
rect 21909 17443 21975 17446
rect 5944 17440 6264 17441
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 17375 6264 17376
rect 15944 17440 16264 17441
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 17375 16264 17376
rect 25944 17440 26264 17441
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 17375 26264 17376
rect 6637 17370 6703 17373
rect 8385 17370 8451 17373
rect 19333 17370 19399 17373
rect 6637 17368 8451 17370
rect 6637 17312 6642 17368
rect 6698 17312 8390 17368
rect 8446 17312 8451 17368
rect 6637 17310 8451 17312
rect 6637 17307 6703 17310
rect 8385 17307 8451 17310
rect 16392 17368 19399 17370
rect 16392 17312 19338 17368
rect 19394 17312 19399 17368
rect 16392 17310 19399 17312
rect 9397 17234 9463 17237
rect 11145 17234 11211 17237
rect 9397 17232 11211 17234
rect 9397 17176 9402 17232
rect 9458 17176 11150 17232
rect 11206 17176 11211 17232
rect 9397 17174 11211 17176
rect 9397 17171 9463 17174
rect 11145 17171 11211 17174
rect 13261 17234 13327 17237
rect 16392 17234 16452 17310
rect 19333 17307 19399 17310
rect 13261 17232 16452 17234
rect 13261 17176 13266 17232
rect 13322 17176 16452 17232
rect 13261 17174 16452 17176
rect 24577 17234 24643 17237
rect 27613 17234 27679 17237
rect 24577 17232 27679 17234
rect 24577 17176 24582 17232
rect 24638 17176 27618 17232
rect 27674 17176 27679 17232
rect 24577 17174 27679 17176
rect 13261 17171 13327 17174
rect 24577 17171 24643 17174
rect 27613 17171 27679 17174
rect 0 17098 480 17128
rect 5809 17098 5875 17101
rect 0 17096 5875 17098
rect 0 17040 5814 17096
rect 5870 17040 5875 17096
rect 0 17038 5875 17040
rect 0 17008 480 17038
rect 5809 17035 5875 17038
rect 8017 17098 8083 17101
rect 11237 17098 11303 17101
rect 8017 17096 11303 17098
rect 8017 17040 8022 17096
rect 8078 17040 11242 17096
rect 11298 17040 11303 17096
rect 8017 17038 11303 17040
rect 8017 17035 8083 17038
rect 11237 17035 11303 17038
rect 11605 17098 11671 17101
rect 19149 17098 19215 17101
rect 11605 17096 19215 17098
rect 11605 17040 11610 17096
rect 11666 17040 19154 17096
rect 19210 17040 19215 17096
rect 11605 17038 19215 17040
rect 11605 17035 11671 17038
rect 19149 17035 19215 17038
rect 22093 17098 22159 17101
rect 29520 17098 30000 17128
rect 22093 17096 30000 17098
rect 22093 17040 22098 17096
rect 22154 17040 30000 17096
rect 22093 17038 30000 17040
rect 22093 17035 22159 17038
rect 29520 17008 30000 17038
rect 10944 16896 11264 16897
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 16831 11264 16832
rect 20944 16896 21264 16897
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 16831 21264 16832
rect 4153 16826 4219 16829
rect 7925 16826 7991 16829
rect 4153 16824 7991 16826
rect 4153 16768 4158 16824
rect 4214 16768 7930 16824
rect 7986 16768 7991 16824
rect 4153 16766 7991 16768
rect 4153 16763 4219 16766
rect 7925 16763 7991 16766
rect 13813 16826 13879 16829
rect 13997 16826 14063 16829
rect 16849 16826 16915 16829
rect 13813 16824 16915 16826
rect 13813 16768 13818 16824
rect 13874 16768 14002 16824
rect 14058 16768 16854 16824
rect 16910 16768 16915 16824
rect 13813 16766 16915 16768
rect 13813 16763 13879 16766
rect 13997 16763 14063 16766
rect 16849 16763 16915 16766
rect 3509 16690 3575 16693
rect 7649 16690 7715 16693
rect 3509 16688 7715 16690
rect 3509 16632 3514 16688
rect 3570 16632 7654 16688
rect 7710 16632 7715 16688
rect 3509 16630 7715 16632
rect 3509 16627 3575 16630
rect 7649 16627 7715 16630
rect 9489 16690 9555 16693
rect 11329 16690 11395 16693
rect 9489 16688 11395 16690
rect 9489 16632 9494 16688
rect 9550 16632 11334 16688
rect 11390 16632 11395 16688
rect 9489 16630 11395 16632
rect 9489 16627 9555 16630
rect 11329 16627 11395 16630
rect 12985 16690 13051 16693
rect 17493 16690 17559 16693
rect 12985 16688 17559 16690
rect 12985 16632 12990 16688
rect 13046 16632 17498 16688
rect 17554 16632 17559 16688
rect 12985 16630 17559 16632
rect 12985 16627 13051 16630
rect 17493 16627 17559 16630
rect 22001 16690 22067 16693
rect 23565 16690 23631 16693
rect 22001 16688 23631 16690
rect 22001 16632 22006 16688
rect 22062 16632 23570 16688
rect 23626 16632 23631 16688
rect 22001 16630 23631 16632
rect 22001 16627 22067 16630
rect 23565 16627 23631 16630
rect 16297 16554 16363 16557
rect 23933 16554 23999 16557
rect 26877 16554 26943 16557
rect 28073 16554 28139 16557
rect 16297 16552 23999 16554
rect 16297 16496 16302 16552
rect 16358 16496 23938 16552
rect 23994 16496 23999 16552
rect 16297 16494 23999 16496
rect 16297 16491 16363 16494
rect 23933 16491 23999 16494
rect 25822 16552 28274 16554
rect 25822 16496 26882 16552
rect 26938 16496 28078 16552
rect 28134 16496 28274 16552
rect 25822 16494 28274 16496
rect 0 16418 480 16448
rect 5441 16418 5507 16421
rect 0 16416 5507 16418
rect 0 16360 5446 16416
rect 5502 16360 5507 16416
rect 0 16358 5507 16360
rect 0 16328 480 16358
rect 5441 16355 5507 16358
rect 5944 16352 6264 16353
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 16287 6264 16288
rect 15944 16352 16264 16353
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 16287 16264 16288
rect 7097 16282 7163 16285
rect 10501 16282 10567 16285
rect 11789 16282 11855 16285
rect 21449 16282 21515 16285
rect 25822 16282 25882 16494
rect 26877 16491 26943 16494
rect 28073 16491 28139 16494
rect 28214 16418 28274 16494
rect 29520 16418 30000 16448
rect 28214 16358 30000 16418
rect 25944 16352 26264 16353
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 29520 16328 30000 16358
rect 25944 16287 26264 16288
rect 7097 16280 11855 16282
rect 7097 16224 7102 16280
rect 7158 16224 10506 16280
rect 10562 16224 11794 16280
rect 11850 16224 11855 16280
rect 7097 16222 11855 16224
rect 7097 16219 7163 16222
rect 10501 16219 10567 16222
rect 11789 16219 11855 16222
rect 18462 16280 25882 16282
rect 18462 16224 21454 16280
rect 21510 16224 25882 16280
rect 18462 16222 25882 16224
rect 5717 16146 5783 16149
rect 18462 16146 18522 16222
rect 21449 16219 21515 16222
rect 5717 16144 18522 16146
rect 5717 16088 5722 16144
rect 5778 16088 18522 16144
rect 5717 16086 18522 16088
rect 19333 16146 19399 16149
rect 25957 16146 26023 16149
rect 26969 16146 27035 16149
rect 19333 16144 27035 16146
rect 19333 16088 19338 16144
rect 19394 16088 25962 16144
rect 26018 16088 26974 16144
rect 27030 16088 27035 16144
rect 19333 16086 27035 16088
rect 5717 16083 5783 16086
rect 19333 16083 19399 16086
rect 25957 16083 26023 16086
rect 26969 16083 27035 16086
rect 3141 16010 3207 16013
rect 3785 16010 3851 16013
rect 3141 16008 3851 16010
rect 3141 15952 3146 16008
rect 3202 15952 3790 16008
rect 3846 15952 3851 16008
rect 3141 15950 3851 15952
rect 3141 15947 3207 15950
rect 3785 15947 3851 15950
rect 5073 16010 5139 16013
rect 9949 16010 10015 16013
rect 11697 16010 11763 16013
rect 12341 16010 12407 16013
rect 23381 16010 23447 16013
rect 5073 16008 11530 16010
rect 5073 15952 5078 16008
rect 5134 15952 9954 16008
rect 10010 15952 11530 16008
rect 5073 15950 11530 15952
rect 5073 15947 5139 15950
rect 9949 15947 10015 15950
rect 0 15874 480 15904
rect 3785 15874 3851 15877
rect 0 15872 3851 15874
rect 0 15816 3790 15872
rect 3846 15816 3851 15872
rect 0 15814 3851 15816
rect 0 15784 480 15814
rect 3785 15811 3851 15814
rect 4613 15874 4679 15877
rect 10685 15874 10751 15877
rect 4613 15872 10751 15874
rect 4613 15816 4618 15872
rect 4674 15816 10690 15872
rect 10746 15816 10751 15872
rect 4613 15814 10751 15816
rect 4613 15811 4679 15814
rect 10685 15811 10751 15814
rect 10944 15808 11264 15809
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 15743 11264 15744
rect 1761 15738 1827 15741
rect 4521 15738 4587 15741
rect 1761 15736 4587 15738
rect 1761 15680 1766 15736
rect 1822 15680 4526 15736
rect 4582 15680 4587 15736
rect 1761 15678 4587 15680
rect 1761 15675 1827 15678
rect 4521 15675 4587 15678
rect 5349 15738 5415 15741
rect 10593 15738 10659 15741
rect 5349 15736 10659 15738
rect 5349 15680 5354 15736
rect 5410 15680 10598 15736
rect 10654 15680 10659 15736
rect 5349 15678 10659 15680
rect 11470 15738 11530 15950
rect 11697 16008 23447 16010
rect 11697 15952 11702 16008
rect 11758 15952 12346 16008
rect 12402 15952 23386 16008
rect 23442 15952 23447 16008
rect 11697 15950 23447 15952
rect 11697 15947 11763 15950
rect 12341 15947 12407 15950
rect 23381 15947 23447 15950
rect 25773 16010 25839 16013
rect 26325 16010 26391 16013
rect 25773 16008 26391 16010
rect 25773 15952 25778 16008
rect 25834 15952 26330 16008
rect 26386 15952 26391 16008
rect 25773 15950 26391 15952
rect 25773 15947 25839 15950
rect 26325 15947 26391 15950
rect 12893 15874 12959 15877
rect 18781 15874 18847 15877
rect 18965 15874 19031 15877
rect 19977 15874 20043 15877
rect 29520 15874 30000 15904
rect 12893 15872 20178 15874
rect 12893 15816 12898 15872
rect 12954 15816 18786 15872
rect 18842 15816 18970 15872
rect 19026 15816 19982 15872
rect 20038 15816 20178 15872
rect 12893 15814 20178 15816
rect 12893 15811 12959 15814
rect 18781 15811 18847 15814
rect 18965 15811 19031 15814
rect 19977 15811 20043 15814
rect 11470 15678 19994 15738
rect 5349 15675 5415 15678
rect 10593 15675 10659 15678
rect 3877 15602 3943 15605
rect 7189 15602 7255 15605
rect 19333 15602 19399 15605
rect 3877 15600 7114 15602
rect 3877 15544 3882 15600
rect 3938 15544 7114 15600
rect 3877 15542 7114 15544
rect 3877 15539 3943 15542
rect 2037 15466 2103 15469
rect 6085 15466 6151 15469
rect 2037 15464 6151 15466
rect 2037 15408 2042 15464
rect 2098 15408 6090 15464
rect 6146 15408 6151 15464
rect 2037 15406 6151 15408
rect 7054 15466 7114 15542
rect 7189 15600 19399 15602
rect 7189 15544 7194 15600
rect 7250 15544 19338 15600
rect 19394 15544 19399 15600
rect 7189 15542 19399 15544
rect 7189 15539 7255 15542
rect 19333 15539 19399 15542
rect 11697 15466 11763 15469
rect 7054 15464 11763 15466
rect 7054 15408 11702 15464
rect 11758 15408 11763 15464
rect 7054 15406 11763 15408
rect 19934 15466 19994 15678
rect 20118 15602 20178 15814
rect 27294 15814 30000 15874
rect 20944 15808 21264 15809
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 20944 15743 21264 15744
rect 24945 15738 25011 15741
rect 27294 15738 27354 15814
rect 29520 15784 30000 15814
rect 24945 15736 27354 15738
rect 24945 15680 24950 15736
rect 25006 15680 27354 15736
rect 24945 15678 27354 15680
rect 24945 15675 25011 15678
rect 24669 15602 24735 15605
rect 20118 15600 24735 15602
rect 20118 15544 24674 15600
rect 24730 15544 24735 15600
rect 20118 15542 24735 15544
rect 24669 15539 24735 15542
rect 25405 15602 25471 15605
rect 27153 15602 27219 15605
rect 25405 15600 27219 15602
rect 25405 15544 25410 15600
rect 25466 15544 27158 15600
rect 27214 15544 27219 15600
rect 25405 15542 27219 15544
rect 25405 15539 25471 15542
rect 27153 15539 27219 15542
rect 20713 15466 20779 15469
rect 21357 15466 21423 15469
rect 19934 15464 21423 15466
rect 19934 15408 20718 15464
rect 20774 15408 21362 15464
rect 21418 15408 21423 15464
rect 19934 15406 21423 15408
rect 2037 15403 2103 15406
rect 6085 15403 6151 15406
rect 11697 15403 11763 15406
rect 20713 15403 20779 15406
rect 21357 15403 21423 15406
rect 24853 15466 24919 15469
rect 24853 15464 26802 15466
rect 24853 15408 24858 15464
rect 24914 15408 26802 15464
rect 24853 15406 26802 15408
rect 24853 15403 24919 15406
rect 0 15330 480 15360
rect 4061 15330 4127 15333
rect 0 15328 4127 15330
rect 0 15272 4066 15328
rect 4122 15272 4127 15328
rect 0 15270 4127 15272
rect 26742 15330 26802 15406
rect 29520 15330 30000 15360
rect 26742 15270 30000 15330
rect 0 15240 480 15270
rect 4061 15267 4127 15270
rect 5944 15264 6264 15265
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 15199 6264 15200
rect 15944 15264 16264 15265
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 15199 16264 15200
rect 25944 15264 26264 15265
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 29520 15240 30000 15270
rect 25944 15199 26264 15200
rect 18689 15194 18755 15197
rect 22921 15194 22987 15197
rect 18689 15192 22987 15194
rect 18689 15136 18694 15192
rect 18750 15136 22926 15192
rect 22982 15136 22987 15192
rect 18689 15134 22987 15136
rect 18689 15131 18755 15134
rect 22921 15131 22987 15134
rect 3509 15058 3575 15061
rect 4429 15058 4495 15061
rect 7281 15058 7347 15061
rect 3509 15056 7347 15058
rect 3509 15000 3514 15056
rect 3570 15000 4434 15056
rect 4490 15000 7286 15056
rect 7342 15000 7347 15056
rect 3509 14998 7347 15000
rect 3509 14995 3575 14998
rect 4429 14995 4495 14998
rect 7281 14995 7347 14998
rect 18137 15058 18203 15061
rect 18597 15058 18663 15061
rect 23197 15058 23263 15061
rect 23657 15058 23723 15061
rect 24761 15058 24827 15061
rect 18137 15056 24827 15058
rect 18137 15000 18142 15056
rect 18198 15000 18602 15056
rect 18658 15000 23202 15056
rect 23258 15000 23662 15056
rect 23718 15000 24766 15056
rect 24822 15000 24827 15056
rect 18137 14998 24827 15000
rect 18137 14995 18203 14998
rect 18597 14995 18663 14998
rect 23197 14995 23263 14998
rect 23657 14995 23723 14998
rect 24761 14995 24827 14998
rect 4705 14922 4771 14925
rect 15193 14922 15259 14925
rect 4705 14920 15259 14922
rect 4705 14864 4710 14920
rect 4766 14864 15198 14920
rect 15254 14864 15259 14920
rect 4705 14862 15259 14864
rect 4705 14859 4771 14862
rect 15193 14859 15259 14862
rect 19149 14922 19215 14925
rect 23749 14922 23815 14925
rect 24393 14922 24459 14925
rect 27337 14922 27403 14925
rect 19149 14920 27403 14922
rect 19149 14864 19154 14920
rect 19210 14864 23754 14920
rect 23810 14864 24398 14920
rect 24454 14864 27342 14920
rect 27398 14864 27403 14920
rect 19149 14862 27403 14864
rect 19149 14859 19215 14862
rect 23749 14859 23815 14862
rect 24393 14859 24459 14862
rect 27337 14859 27403 14862
rect 5441 14786 5507 14789
rect 10409 14786 10475 14789
rect 5441 14784 10475 14786
rect 5441 14728 5446 14784
rect 5502 14728 10414 14784
rect 10470 14728 10475 14784
rect 5441 14726 10475 14728
rect 5441 14723 5507 14726
rect 10409 14723 10475 14726
rect 10944 14720 11264 14721
rect 0 14650 480 14680
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 14655 11264 14656
rect 20944 14720 21264 14721
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 14655 21264 14656
rect 6545 14650 6611 14653
rect 0 14648 6611 14650
rect 0 14592 6550 14648
rect 6606 14592 6611 14648
rect 0 14590 6611 14592
rect 0 14560 480 14590
rect 6545 14587 6611 14590
rect 14825 14650 14891 14653
rect 19885 14650 19951 14653
rect 14825 14648 19951 14650
rect 14825 14592 14830 14648
rect 14886 14592 19890 14648
rect 19946 14592 19951 14648
rect 14825 14590 19951 14592
rect 14825 14587 14891 14590
rect 19885 14587 19951 14590
rect 25037 14650 25103 14653
rect 29520 14650 30000 14680
rect 25037 14648 30000 14650
rect 25037 14592 25042 14648
rect 25098 14592 30000 14648
rect 25037 14590 30000 14592
rect 25037 14587 25103 14590
rect 29520 14560 30000 14590
rect 1669 14514 1735 14517
rect 3601 14514 3667 14517
rect 1669 14512 3667 14514
rect 1669 14456 1674 14512
rect 1730 14456 3606 14512
rect 3662 14456 3667 14512
rect 1669 14454 3667 14456
rect 1669 14451 1735 14454
rect 3601 14451 3667 14454
rect 6729 14514 6795 14517
rect 11789 14514 11855 14517
rect 6729 14512 11855 14514
rect 6729 14456 6734 14512
rect 6790 14456 11794 14512
rect 11850 14456 11855 14512
rect 6729 14454 11855 14456
rect 6729 14451 6795 14454
rect 11789 14451 11855 14454
rect 19701 14514 19767 14517
rect 26785 14514 26851 14517
rect 19701 14512 26851 14514
rect 19701 14456 19706 14512
rect 19762 14456 26790 14512
rect 26846 14456 26851 14512
rect 19701 14454 26851 14456
rect 19701 14451 19767 14454
rect 26785 14451 26851 14454
rect 2681 14378 2747 14381
rect 7557 14378 7623 14381
rect 2681 14376 7623 14378
rect 2681 14320 2686 14376
rect 2742 14320 7562 14376
rect 7618 14320 7623 14376
rect 2681 14318 7623 14320
rect 2681 14315 2747 14318
rect 7557 14315 7623 14318
rect 24209 14378 24275 14381
rect 26877 14378 26943 14381
rect 27613 14378 27679 14381
rect 24209 14376 27679 14378
rect 24209 14320 24214 14376
rect 24270 14320 26882 14376
rect 26938 14320 27618 14376
rect 27674 14320 27679 14376
rect 24209 14318 27679 14320
rect 24209 14315 24275 14318
rect 26877 14315 26943 14318
rect 27613 14315 27679 14318
rect 10409 14242 10475 14245
rect 14733 14242 14799 14245
rect 20345 14242 20411 14245
rect 10409 14240 14799 14242
rect 10409 14184 10414 14240
rect 10470 14184 14738 14240
rect 14794 14184 14799 14240
rect 10409 14182 14799 14184
rect 10409 14179 10475 14182
rect 14733 14179 14799 14182
rect 18646 14240 20411 14242
rect 18646 14184 20350 14240
rect 20406 14184 20411 14240
rect 18646 14182 20411 14184
rect 5944 14176 6264 14177
rect 0 14106 480 14136
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 14111 6264 14112
rect 15944 14176 16264 14177
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 14111 16264 14112
rect 4521 14106 4587 14109
rect 0 14104 4587 14106
rect 0 14048 4526 14104
rect 4582 14048 4587 14104
rect 0 14046 4587 14048
rect 0 14016 480 14046
rect 4521 14043 4587 14046
rect 7557 14106 7623 14109
rect 13261 14106 13327 14109
rect 7557 14104 13327 14106
rect 7557 14048 7562 14104
rect 7618 14048 13266 14104
rect 13322 14048 13327 14104
rect 7557 14046 13327 14048
rect 7557 14043 7623 14046
rect 13261 14043 13327 14046
rect 3693 13970 3759 13973
rect 10593 13970 10659 13973
rect 18646 13970 18706 14182
rect 20345 14179 20411 14182
rect 25944 14176 26264 14177
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 14111 26264 14112
rect 20069 14106 20135 14109
rect 23473 14106 23539 14109
rect 20069 14104 23539 14106
rect 20069 14048 20074 14104
rect 20130 14048 23478 14104
rect 23534 14048 23539 14104
rect 20069 14046 23539 14048
rect 20069 14043 20135 14046
rect 23473 14043 23539 14046
rect 26509 14106 26575 14109
rect 29520 14106 30000 14136
rect 26509 14104 30000 14106
rect 26509 14048 26514 14104
rect 26570 14048 30000 14104
rect 26509 14046 30000 14048
rect 26509 14043 26575 14046
rect 29520 14016 30000 14046
rect 3693 13968 18706 13970
rect 3693 13912 3698 13968
rect 3754 13912 10598 13968
rect 10654 13912 18706 13968
rect 3693 13910 18706 13912
rect 19241 13970 19307 13973
rect 26969 13970 27035 13973
rect 19241 13968 27035 13970
rect 19241 13912 19246 13968
rect 19302 13912 26974 13968
rect 27030 13912 27035 13968
rect 19241 13910 27035 13912
rect 3693 13907 3759 13910
rect 10593 13907 10659 13910
rect 19241 13907 19307 13910
rect 26969 13907 27035 13910
rect 10409 13834 10475 13837
rect 13813 13834 13879 13837
rect 10409 13832 13879 13834
rect 10409 13776 10414 13832
rect 10470 13776 13818 13832
rect 13874 13776 13879 13832
rect 10409 13774 13879 13776
rect 10409 13771 10475 13774
rect 13813 13771 13879 13774
rect 17493 13834 17559 13837
rect 19425 13834 19491 13837
rect 17493 13832 19491 13834
rect 17493 13776 17498 13832
rect 17554 13776 19430 13832
rect 19486 13776 19491 13832
rect 17493 13774 19491 13776
rect 17493 13771 17559 13774
rect 19425 13771 19491 13774
rect 22921 13834 22987 13837
rect 24669 13834 24735 13837
rect 26693 13834 26759 13837
rect 22921 13832 23490 13834
rect 22921 13776 22926 13832
rect 22982 13776 23490 13832
rect 22921 13774 23490 13776
rect 22921 13771 22987 13774
rect 4061 13698 4127 13701
rect 6453 13698 6519 13701
rect 4061 13696 6519 13698
rect 4061 13640 4066 13696
rect 4122 13640 6458 13696
rect 6514 13640 6519 13696
rect 4061 13638 6519 13640
rect 4061 13635 4127 13638
rect 6453 13635 6519 13638
rect 15561 13698 15627 13701
rect 18505 13698 18571 13701
rect 19609 13698 19675 13701
rect 15561 13696 19675 13698
rect 15561 13640 15566 13696
rect 15622 13640 18510 13696
rect 18566 13640 19614 13696
rect 19670 13640 19675 13696
rect 15561 13638 19675 13640
rect 23430 13698 23490 13774
rect 24669 13832 26759 13834
rect 24669 13776 24674 13832
rect 24730 13776 26698 13832
rect 26754 13776 26759 13832
rect 24669 13774 26759 13776
rect 24669 13771 24735 13774
rect 26693 13771 26759 13774
rect 25681 13698 25747 13701
rect 23430 13696 25747 13698
rect 23430 13640 25686 13696
rect 25742 13640 25747 13696
rect 23430 13638 25747 13640
rect 15561 13635 15627 13638
rect 18505 13635 18571 13638
rect 19609 13635 19675 13638
rect 25681 13635 25747 13638
rect 10944 13632 11264 13633
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 13567 11264 13568
rect 20944 13632 21264 13633
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 13567 21264 13568
rect 14089 13562 14155 13565
rect 16021 13562 16087 13565
rect 20621 13562 20687 13565
rect 14089 13560 20687 13562
rect 14089 13504 14094 13560
rect 14150 13504 16026 13560
rect 16082 13504 20626 13560
rect 20682 13504 20687 13560
rect 14089 13502 20687 13504
rect 14089 13499 14155 13502
rect 16021 13499 16087 13502
rect 20621 13499 20687 13502
rect 21449 13562 21515 13565
rect 23197 13562 23263 13565
rect 24945 13562 25011 13565
rect 21449 13560 25011 13562
rect 21449 13504 21454 13560
rect 21510 13504 23202 13560
rect 23258 13504 24950 13560
rect 25006 13504 25011 13560
rect 21449 13502 25011 13504
rect 21449 13499 21515 13502
rect 23197 13499 23263 13502
rect 24945 13499 25011 13502
rect 25589 13562 25655 13565
rect 26509 13562 26575 13565
rect 25589 13560 26575 13562
rect 25589 13504 25594 13560
rect 25650 13504 26514 13560
rect 26570 13504 26575 13560
rect 25589 13502 26575 13504
rect 25589 13499 25655 13502
rect 26509 13499 26575 13502
rect 0 13426 480 13456
rect 1577 13426 1643 13429
rect 0 13424 1643 13426
rect 0 13368 1582 13424
rect 1638 13368 1643 13424
rect 0 13366 1643 13368
rect 0 13336 480 13366
rect 1577 13363 1643 13366
rect 5901 13426 5967 13429
rect 7649 13426 7715 13429
rect 5901 13424 7715 13426
rect 5901 13368 5906 13424
rect 5962 13368 7654 13424
rect 7710 13368 7715 13424
rect 5901 13366 7715 13368
rect 5901 13363 5967 13366
rect 7649 13363 7715 13366
rect 7833 13426 7899 13429
rect 14917 13426 14983 13429
rect 7833 13424 14983 13426
rect 7833 13368 7838 13424
rect 7894 13368 14922 13424
rect 14978 13368 14983 13424
rect 7833 13366 14983 13368
rect 7833 13363 7899 13366
rect 14917 13363 14983 13366
rect 20529 13426 20595 13429
rect 22737 13426 22803 13429
rect 29520 13426 30000 13456
rect 20529 13424 22803 13426
rect 20529 13368 20534 13424
rect 20590 13368 22742 13424
rect 22798 13368 22803 13424
rect 20529 13366 22803 13368
rect 20529 13363 20595 13366
rect 22737 13363 22803 13366
rect 25822 13366 30000 13426
rect 3785 13290 3851 13293
rect 11973 13290 12039 13293
rect 22645 13290 22711 13293
rect 3785 13288 6562 13290
rect 3785 13232 3790 13288
rect 3846 13232 6562 13288
rect 3785 13230 6562 13232
rect 3785 13227 3851 13230
rect 6502 13154 6562 13230
rect 11973 13288 22711 13290
rect 11973 13232 11978 13288
rect 12034 13232 22650 13288
rect 22706 13232 22711 13288
rect 11973 13230 22711 13232
rect 11973 13227 12039 13230
rect 22645 13227 22711 13230
rect 15285 13154 15351 13157
rect 6502 13152 15351 13154
rect 6502 13096 15290 13152
rect 15346 13096 15351 13152
rect 6502 13094 15351 13096
rect 15285 13091 15351 13094
rect 20713 13154 20779 13157
rect 21541 13154 21607 13157
rect 20713 13152 21607 13154
rect 20713 13096 20718 13152
rect 20774 13096 21546 13152
rect 21602 13096 21607 13152
rect 20713 13094 21607 13096
rect 20713 13091 20779 13094
rect 21541 13091 21607 13094
rect 5944 13088 6264 13089
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 13023 6264 13024
rect 15944 13088 16264 13089
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 13023 16264 13024
rect 2773 13018 2839 13021
rect 5533 13018 5599 13021
rect 2773 13016 5599 13018
rect 2773 12960 2778 13016
rect 2834 12960 5538 13016
rect 5594 12960 5599 13016
rect 2773 12958 5599 12960
rect 2773 12955 2839 12958
rect 5533 12955 5599 12958
rect 7741 13018 7807 13021
rect 11605 13018 11671 13021
rect 14089 13018 14155 13021
rect 7741 13016 14155 13018
rect 7741 12960 7746 13016
rect 7802 12960 11610 13016
rect 11666 12960 14094 13016
rect 14150 12960 14155 13016
rect 7741 12958 14155 12960
rect 7741 12955 7807 12958
rect 11605 12955 11671 12958
rect 14089 12955 14155 12958
rect 19609 13018 19675 13021
rect 25822 13018 25882 13366
rect 29520 13336 30000 13366
rect 25944 13088 26264 13089
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 13023 26264 13024
rect 19609 13016 25882 13018
rect 19609 12960 19614 13016
rect 19670 12960 25882 13016
rect 19609 12958 25882 12960
rect 19609 12955 19675 12958
rect 0 12882 480 12912
rect 565 12882 631 12885
rect 0 12880 631 12882
rect 0 12824 570 12880
rect 626 12824 631 12880
rect 0 12822 631 12824
rect 0 12792 480 12822
rect 565 12819 631 12822
rect 2957 12882 3023 12885
rect 5809 12882 5875 12885
rect 2957 12880 5875 12882
rect 2957 12824 2962 12880
rect 3018 12824 5814 12880
rect 5870 12824 5875 12880
rect 2957 12822 5875 12824
rect 2957 12819 3023 12822
rect 5809 12819 5875 12822
rect 6177 12882 6243 12885
rect 12157 12882 12223 12885
rect 6177 12880 12223 12882
rect 6177 12824 6182 12880
rect 6238 12824 12162 12880
rect 12218 12824 12223 12880
rect 6177 12822 12223 12824
rect 6177 12819 6243 12822
rect 12157 12819 12223 12822
rect 13629 12882 13695 12885
rect 15469 12882 15535 12885
rect 13629 12880 15535 12882
rect 13629 12824 13634 12880
rect 13690 12824 15474 12880
rect 15530 12824 15535 12880
rect 13629 12822 15535 12824
rect 13629 12819 13695 12822
rect 15469 12819 15535 12822
rect 16205 12882 16271 12885
rect 19701 12882 19767 12885
rect 27337 12882 27403 12885
rect 16205 12880 27403 12882
rect 16205 12824 16210 12880
rect 16266 12824 19706 12880
rect 19762 12824 27342 12880
rect 27398 12824 27403 12880
rect 16205 12822 27403 12824
rect 16205 12819 16271 12822
rect 19701 12819 19767 12822
rect 27337 12819 27403 12822
rect 27521 12882 27587 12885
rect 29520 12882 30000 12912
rect 27521 12880 30000 12882
rect 27521 12824 27526 12880
rect 27582 12824 30000 12880
rect 27521 12822 30000 12824
rect 27521 12819 27587 12822
rect 29520 12792 30000 12822
rect 6913 12746 6979 12749
rect 10777 12746 10843 12749
rect 13905 12746 13971 12749
rect 6913 12744 13971 12746
rect 6913 12688 6918 12744
rect 6974 12688 10782 12744
rect 10838 12688 13910 12744
rect 13966 12688 13971 12744
rect 6913 12686 13971 12688
rect 6913 12683 6979 12686
rect 10777 12683 10843 12686
rect 13905 12683 13971 12686
rect 15653 12746 15719 12749
rect 16481 12746 16547 12749
rect 21449 12746 21515 12749
rect 15653 12744 16547 12746
rect 15653 12688 15658 12744
rect 15714 12688 16486 12744
rect 16542 12688 16547 12744
rect 15653 12686 16547 12688
rect 15653 12683 15719 12686
rect 16481 12683 16547 12686
rect 20670 12744 21515 12746
rect 20670 12688 21454 12744
rect 21510 12688 21515 12744
rect 20670 12686 21515 12688
rect 15193 12610 15259 12613
rect 15837 12610 15903 12613
rect 20670 12610 20730 12686
rect 21449 12683 21515 12686
rect 15193 12608 20730 12610
rect 15193 12552 15198 12608
rect 15254 12552 15842 12608
rect 15898 12552 20730 12608
rect 15193 12550 20730 12552
rect 24577 12610 24643 12613
rect 26417 12610 26483 12613
rect 24577 12608 26483 12610
rect 24577 12552 24582 12608
rect 24638 12552 26422 12608
rect 26478 12552 26483 12608
rect 24577 12550 26483 12552
rect 15193 12547 15259 12550
rect 15837 12547 15903 12550
rect 24577 12547 24643 12550
rect 26417 12547 26483 12550
rect 10944 12544 11264 12545
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 12479 11264 12480
rect 20944 12544 21264 12545
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 12479 21264 12480
rect 7465 12474 7531 12477
rect 21541 12474 21607 12477
rect 26601 12474 26667 12477
rect 7465 12472 8402 12474
rect 7465 12416 7470 12472
rect 7526 12416 8402 12472
rect 7465 12414 8402 12416
rect 7465 12411 7531 12414
rect 0 12338 480 12368
rect 4061 12338 4127 12341
rect 7557 12338 7623 12341
rect 0 12336 4127 12338
rect 0 12280 4066 12336
rect 4122 12280 4127 12336
rect 0 12278 4127 12280
rect 0 12248 480 12278
rect 4061 12275 4127 12278
rect 5766 12336 7623 12338
rect 5766 12280 7562 12336
rect 7618 12280 7623 12336
rect 5766 12278 7623 12280
rect 8342 12338 8402 12414
rect 21541 12472 26667 12474
rect 21541 12416 21546 12472
rect 21602 12416 26606 12472
rect 26662 12416 26667 12472
rect 21541 12414 26667 12416
rect 21541 12411 21607 12414
rect 26601 12411 26667 12414
rect 15929 12338 15995 12341
rect 8342 12336 15995 12338
rect 8342 12280 15934 12336
rect 15990 12280 15995 12336
rect 8342 12278 15995 12280
rect 1485 12202 1551 12205
rect 2037 12202 2103 12205
rect 5766 12202 5826 12278
rect 7557 12275 7623 12278
rect 15929 12275 15995 12278
rect 16573 12338 16639 12341
rect 20989 12338 21055 12341
rect 16573 12336 21055 12338
rect 16573 12280 16578 12336
rect 16634 12280 20994 12336
rect 21050 12280 21055 12336
rect 16573 12278 21055 12280
rect 16573 12275 16639 12278
rect 20989 12275 21055 12278
rect 22737 12338 22803 12341
rect 27429 12338 27495 12341
rect 29520 12338 30000 12368
rect 22737 12336 30000 12338
rect 22737 12280 22742 12336
rect 22798 12280 27434 12336
rect 27490 12280 30000 12336
rect 22737 12278 30000 12280
rect 22737 12275 22803 12278
rect 27429 12275 27495 12278
rect 29520 12248 30000 12278
rect 1485 12200 5826 12202
rect 1485 12144 1490 12200
rect 1546 12144 2042 12200
rect 2098 12144 5826 12200
rect 1485 12142 5826 12144
rect 5901 12202 5967 12205
rect 6269 12202 6335 12205
rect 9397 12202 9463 12205
rect 5901 12200 9463 12202
rect 5901 12144 5906 12200
rect 5962 12144 6274 12200
rect 6330 12144 9402 12200
rect 9458 12144 9463 12200
rect 5901 12142 9463 12144
rect 1485 12139 1551 12142
rect 2037 12139 2103 12142
rect 5901 12139 5967 12142
rect 6269 12139 6335 12142
rect 9397 12139 9463 12142
rect 15285 12202 15351 12205
rect 22001 12202 22067 12205
rect 24577 12202 24643 12205
rect 15285 12200 16498 12202
rect 15285 12144 15290 12200
rect 15346 12144 16498 12200
rect 15285 12142 16498 12144
rect 15285 12139 15351 12142
rect 7557 12066 7623 12069
rect 14733 12066 14799 12069
rect 7557 12064 14799 12066
rect 7557 12008 7562 12064
rect 7618 12008 14738 12064
rect 14794 12008 14799 12064
rect 7557 12006 14799 12008
rect 16438 12066 16498 12142
rect 22001 12200 24643 12202
rect 22001 12144 22006 12200
rect 22062 12144 24582 12200
rect 24638 12144 24643 12200
rect 22001 12142 24643 12144
rect 22001 12139 22067 12142
rect 24577 12139 24643 12142
rect 16665 12066 16731 12069
rect 23013 12066 23079 12069
rect 16438 12064 25882 12066
rect 16438 12008 16670 12064
rect 16726 12008 23018 12064
rect 23074 12008 25882 12064
rect 16438 12006 25882 12008
rect 7557 12003 7623 12006
rect 14733 12003 14799 12006
rect 16665 12003 16731 12006
rect 23013 12003 23079 12006
rect 5944 12000 6264 12001
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 11935 6264 11936
rect 15944 12000 16264 12001
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 11935 16264 11936
rect 6361 11930 6427 11933
rect 6494 11930 6500 11932
rect 6361 11928 6500 11930
rect 6361 11872 6366 11928
rect 6422 11872 6500 11928
rect 6361 11870 6500 11872
rect 6361 11867 6427 11870
rect 6494 11868 6500 11870
rect 6564 11868 6570 11932
rect 12750 11868 12756 11932
rect 12820 11930 12826 11932
rect 12893 11930 12959 11933
rect 12820 11928 12959 11930
rect 12820 11872 12898 11928
rect 12954 11872 12959 11928
rect 12820 11870 12959 11872
rect 12820 11868 12826 11870
rect 12893 11867 12959 11870
rect 2957 11794 3023 11797
rect 1350 11792 3023 11794
rect 1350 11736 2962 11792
rect 3018 11736 3023 11792
rect 1350 11734 3023 11736
rect 0 11658 480 11688
rect 1350 11658 1410 11734
rect 2957 11731 3023 11734
rect 3877 11794 3943 11797
rect 6821 11794 6887 11797
rect 3877 11792 6887 11794
rect 3877 11736 3882 11792
rect 3938 11736 6826 11792
rect 6882 11736 6887 11792
rect 3877 11734 6887 11736
rect 3877 11731 3943 11734
rect 6821 11731 6887 11734
rect 7281 11794 7347 11797
rect 10225 11794 10291 11797
rect 7281 11792 10291 11794
rect 7281 11736 7286 11792
rect 7342 11736 10230 11792
rect 10286 11736 10291 11792
rect 7281 11734 10291 11736
rect 7281 11731 7347 11734
rect 10225 11731 10291 11734
rect 14273 11794 14339 11797
rect 24853 11794 24919 11797
rect 14273 11792 24919 11794
rect 14273 11736 14278 11792
rect 14334 11736 24858 11792
rect 24914 11736 24919 11792
rect 14273 11734 24919 11736
rect 25822 11794 25882 12006
rect 25944 12000 26264 12001
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 11935 26264 11936
rect 26969 11794 27035 11797
rect 25822 11792 27035 11794
rect 25822 11736 26974 11792
rect 27030 11736 27035 11792
rect 25822 11734 27035 11736
rect 14273 11731 14339 11734
rect 24853 11731 24919 11734
rect 26969 11731 27035 11734
rect 0 11598 1410 11658
rect 2405 11658 2471 11661
rect 8385 11658 8451 11661
rect 11789 11658 11855 11661
rect 2405 11656 8451 11658
rect 2405 11600 2410 11656
rect 2466 11600 8390 11656
rect 8446 11600 8451 11656
rect 2405 11598 8451 11600
rect 0 11568 480 11598
rect 2405 11595 2471 11598
rect 8385 11595 8451 11598
rect 8894 11656 11855 11658
rect 8894 11600 11794 11656
rect 11850 11600 11855 11656
rect 8894 11598 11855 11600
rect 8894 11525 8954 11598
rect 11789 11595 11855 11598
rect 22645 11658 22711 11661
rect 29520 11658 30000 11688
rect 22645 11656 30000 11658
rect 22645 11600 22650 11656
rect 22706 11600 30000 11656
rect 22645 11598 30000 11600
rect 22645 11595 22711 11598
rect 29520 11568 30000 11598
rect 5165 11522 5231 11525
rect 8845 11522 8954 11525
rect 5165 11520 8954 11522
rect 5165 11464 5170 11520
rect 5226 11464 8850 11520
rect 8906 11464 8954 11520
rect 5165 11462 8954 11464
rect 5165 11459 5231 11462
rect 8845 11459 8911 11462
rect 10944 11456 11264 11457
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 11391 11264 11392
rect 20944 11456 21264 11457
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 11391 21264 11392
rect 5533 11386 5599 11389
rect 9305 11386 9371 11389
rect 5533 11384 9371 11386
rect 5533 11328 5538 11384
rect 5594 11328 9310 11384
rect 9366 11328 9371 11384
rect 5533 11326 9371 11328
rect 5533 11323 5599 11326
rect 9305 11323 9371 11326
rect 18413 11386 18479 11389
rect 20805 11386 20871 11389
rect 18413 11384 20871 11386
rect 18413 11328 18418 11384
rect 18474 11328 20810 11384
rect 20866 11328 20871 11384
rect 18413 11326 20871 11328
rect 18413 11323 18479 11326
rect 20805 11323 20871 11326
rect 2681 11250 2747 11253
rect 8293 11250 8359 11253
rect 2681 11248 8359 11250
rect 2681 11192 2686 11248
rect 2742 11192 8298 11248
rect 8354 11192 8359 11248
rect 2681 11190 8359 11192
rect 2681 11187 2747 11190
rect 8293 11187 8359 11190
rect 0 11114 480 11144
rect 4245 11114 4311 11117
rect 0 11112 4311 11114
rect 0 11056 4250 11112
rect 4306 11056 4311 11112
rect 0 11054 4311 11056
rect 0 11024 480 11054
rect 4245 11051 4311 11054
rect 25497 11114 25563 11117
rect 29520 11114 30000 11144
rect 25497 11112 30000 11114
rect 25497 11056 25502 11112
rect 25558 11056 30000 11112
rect 25497 11054 30000 11056
rect 25497 11051 25563 11054
rect 29520 11024 30000 11054
rect 20069 10978 20135 10981
rect 23841 10978 23907 10981
rect 20069 10976 23907 10978
rect 20069 10920 20074 10976
rect 20130 10920 23846 10976
rect 23902 10920 23907 10976
rect 20069 10918 23907 10920
rect 20069 10915 20135 10918
rect 23841 10915 23907 10918
rect 24945 10978 25011 10981
rect 25221 10978 25287 10981
rect 24945 10976 25287 10978
rect 24945 10920 24950 10976
rect 25006 10920 25226 10976
rect 25282 10920 25287 10976
rect 24945 10918 25287 10920
rect 24945 10915 25011 10918
rect 25221 10915 25287 10918
rect 5944 10912 6264 10913
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 10847 6264 10848
rect 15944 10912 16264 10913
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 10847 16264 10848
rect 25944 10912 26264 10913
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 10847 26264 10848
rect 10593 10842 10659 10845
rect 14273 10842 14339 10845
rect 10593 10840 14339 10842
rect 10593 10784 10598 10840
rect 10654 10784 14278 10840
rect 14334 10784 14339 10840
rect 10593 10782 14339 10784
rect 10593 10779 10659 10782
rect 14273 10779 14339 10782
rect 20437 10842 20503 10845
rect 23197 10842 23263 10845
rect 20437 10840 23263 10842
rect 20437 10784 20442 10840
rect 20498 10784 23202 10840
rect 23258 10784 23263 10840
rect 20437 10782 23263 10784
rect 20437 10779 20503 10782
rect 23197 10779 23263 10782
rect 23933 10842 23999 10845
rect 25221 10842 25287 10845
rect 23933 10840 25287 10842
rect 23933 10784 23938 10840
rect 23994 10784 25226 10840
rect 25282 10784 25287 10840
rect 23933 10782 25287 10784
rect 23933 10779 23999 10782
rect 25221 10779 25287 10782
rect 3233 10706 3299 10709
rect 24117 10706 24183 10709
rect 3233 10704 24183 10706
rect 3233 10648 3238 10704
rect 3294 10648 24122 10704
rect 24178 10648 24183 10704
rect 3233 10646 24183 10648
rect 3233 10643 3299 10646
rect 24117 10643 24183 10646
rect 25681 10706 25747 10709
rect 27337 10706 27403 10709
rect 25681 10704 27403 10706
rect 25681 10648 25686 10704
rect 25742 10648 27342 10704
rect 27398 10648 27403 10704
rect 25681 10646 27403 10648
rect 25681 10643 25747 10646
rect 27337 10643 27403 10646
rect 1945 10570 2011 10573
rect 8937 10570 9003 10573
rect 1945 10568 9003 10570
rect 1945 10512 1950 10568
rect 2006 10512 8942 10568
rect 8998 10512 9003 10568
rect 1945 10510 9003 10512
rect 1945 10507 2011 10510
rect 8937 10507 9003 10510
rect 17125 10570 17191 10573
rect 24945 10570 25011 10573
rect 26969 10570 27035 10573
rect 17125 10568 27035 10570
rect 17125 10512 17130 10568
rect 17186 10512 24950 10568
rect 25006 10512 26974 10568
rect 27030 10512 27035 10568
rect 17125 10510 27035 10512
rect 17125 10507 17191 10510
rect 24945 10507 25011 10510
rect 26969 10507 27035 10510
rect 0 10434 480 10464
rect 4061 10434 4127 10437
rect 0 10432 4127 10434
rect 0 10376 4066 10432
rect 4122 10376 4127 10432
rect 0 10374 4127 10376
rect 0 10344 480 10374
rect 4061 10371 4127 10374
rect 24393 10434 24459 10437
rect 29520 10434 30000 10464
rect 24393 10432 30000 10434
rect 24393 10376 24398 10432
rect 24454 10376 30000 10432
rect 24393 10374 30000 10376
rect 24393 10371 24459 10374
rect 10944 10368 11264 10369
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 10303 11264 10304
rect 20944 10368 21264 10369
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 29520 10344 30000 10374
rect 20944 10303 21264 10304
rect 3141 10298 3207 10301
rect 4613 10298 4679 10301
rect 5625 10298 5691 10301
rect 3141 10296 5691 10298
rect 3141 10240 3146 10296
rect 3202 10240 4618 10296
rect 4674 10240 5630 10296
rect 5686 10240 5691 10296
rect 3141 10238 5691 10240
rect 3141 10235 3207 10238
rect 4613 10235 4679 10238
rect 5625 10235 5691 10238
rect 5993 10298 6059 10301
rect 8385 10298 8451 10301
rect 5993 10296 8451 10298
rect 5993 10240 5998 10296
rect 6054 10240 8390 10296
rect 8446 10240 8451 10296
rect 5993 10238 8451 10240
rect 5993 10235 6059 10238
rect 8385 10235 8451 10238
rect 6085 10162 6151 10165
rect 6361 10162 6427 10165
rect 11973 10162 12039 10165
rect 17217 10162 17283 10165
rect 6085 10160 8770 10162
rect 6085 10104 6090 10160
rect 6146 10104 6366 10160
rect 6422 10104 8770 10160
rect 6085 10102 8770 10104
rect 6085 10099 6151 10102
rect 6361 10099 6427 10102
rect 3141 10026 3207 10029
rect 7189 10026 7255 10029
rect 3141 10024 7255 10026
rect 3141 9968 3146 10024
rect 3202 9968 7194 10024
rect 7250 9968 7255 10024
rect 3141 9966 7255 9968
rect 8710 10026 8770 10102
rect 11973 10160 17283 10162
rect 11973 10104 11978 10160
rect 12034 10104 17222 10160
rect 17278 10104 17283 10160
rect 11973 10102 17283 10104
rect 11973 10099 12039 10102
rect 17217 10099 17283 10102
rect 17401 10162 17467 10165
rect 22461 10162 22527 10165
rect 27337 10162 27403 10165
rect 17401 10160 27403 10162
rect 17401 10104 17406 10160
rect 17462 10104 22466 10160
rect 22522 10104 27342 10160
rect 27398 10104 27403 10160
rect 17401 10102 27403 10104
rect 17401 10099 17467 10102
rect 22461 10099 22527 10102
rect 27337 10099 27403 10102
rect 10317 10026 10383 10029
rect 25313 10026 25379 10029
rect 8710 10024 25379 10026
rect 8710 9968 10322 10024
rect 10378 9968 25318 10024
rect 25374 9968 25379 10024
rect 8710 9966 25379 9968
rect 3141 9963 3207 9966
rect 7189 9963 7255 9966
rect 10317 9963 10383 9966
rect 25313 9963 25379 9966
rect 0 9890 480 9920
rect 3785 9890 3851 9893
rect 29520 9890 30000 9920
rect 0 9888 3851 9890
rect 0 9832 3790 9888
rect 3846 9832 3851 9888
rect 0 9830 3851 9832
rect 0 9800 480 9830
rect 3785 9827 3851 9830
rect 27846 9830 30000 9890
rect 5944 9824 6264 9825
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 9759 6264 9760
rect 15944 9824 16264 9825
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 9759 16264 9760
rect 25944 9824 26264 9825
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 25944 9759 26264 9760
rect 8753 9754 8819 9757
rect 15745 9754 15811 9757
rect 8753 9752 15811 9754
rect 8753 9696 8758 9752
rect 8814 9696 15750 9752
rect 15806 9696 15811 9752
rect 8753 9694 15811 9696
rect 8753 9691 8819 9694
rect 15745 9691 15811 9694
rect 17217 9754 17283 9757
rect 17217 9752 22202 9754
rect 17217 9696 17222 9752
rect 17278 9696 22202 9752
rect 17217 9694 22202 9696
rect 17217 9691 17283 9694
rect 21452 9621 21512 9694
rect 3417 9618 3483 9621
rect 8293 9618 8359 9621
rect 3417 9616 8359 9618
rect 3417 9560 3422 9616
rect 3478 9560 8298 9616
rect 8354 9560 8359 9616
rect 3417 9558 8359 9560
rect 3417 9555 3483 9558
rect 8293 9555 8359 9558
rect 16849 9618 16915 9621
rect 21265 9618 21331 9621
rect 16849 9616 21331 9618
rect 16849 9560 16854 9616
rect 16910 9560 21270 9616
rect 21326 9560 21331 9616
rect 16849 9558 21331 9560
rect 16849 9555 16915 9558
rect 21265 9555 21331 9558
rect 21449 9616 21515 9621
rect 21449 9560 21454 9616
rect 21510 9560 21515 9616
rect 21449 9555 21515 9560
rect 1945 9482 2011 9485
rect 3233 9482 3299 9485
rect 1945 9480 3299 9482
rect 1945 9424 1950 9480
rect 2006 9424 3238 9480
rect 3294 9424 3299 9480
rect 1945 9422 3299 9424
rect 1945 9419 2011 9422
rect 3233 9419 3299 9422
rect 4245 9482 4311 9485
rect 15929 9482 15995 9485
rect 4245 9480 15995 9482
rect 4245 9424 4250 9480
rect 4306 9424 15934 9480
rect 15990 9424 15995 9480
rect 4245 9422 15995 9424
rect 22142 9482 22202 9694
rect 24577 9618 24643 9621
rect 27521 9618 27587 9621
rect 24577 9616 27587 9618
rect 24577 9560 24582 9616
rect 24638 9560 27526 9616
rect 27582 9560 27587 9616
rect 24577 9558 27587 9560
rect 24577 9555 24643 9558
rect 27521 9555 27587 9558
rect 27705 9618 27771 9621
rect 27846 9618 27906 9830
rect 29520 9800 30000 9830
rect 27705 9616 27906 9618
rect 27705 9560 27710 9616
rect 27766 9560 27906 9616
rect 27705 9558 27906 9560
rect 27705 9555 27771 9558
rect 24209 9482 24275 9485
rect 22142 9480 24275 9482
rect 22142 9424 24214 9480
rect 24270 9424 24275 9480
rect 22142 9422 24275 9424
rect 4245 9419 4311 9422
rect 15929 9419 15995 9422
rect 24209 9419 24275 9422
rect 0 9346 480 9376
rect 5809 9346 5875 9349
rect 0 9344 5875 9346
rect 0 9288 5814 9344
rect 5870 9288 5875 9344
rect 0 9286 5875 9288
rect 0 9256 480 9286
rect 5809 9283 5875 9286
rect 16481 9346 16547 9349
rect 18505 9346 18571 9349
rect 16481 9344 18571 9346
rect 16481 9288 16486 9344
rect 16542 9288 18510 9344
rect 18566 9288 18571 9344
rect 16481 9286 18571 9288
rect 16481 9283 16547 9286
rect 18505 9283 18571 9286
rect 24393 9346 24459 9349
rect 29520 9346 30000 9376
rect 24393 9344 30000 9346
rect 24393 9288 24398 9344
rect 24454 9288 30000 9344
rect 24393 9286 30000 9288
rect 24393 9283 24459 9286
rect 10944 9280 11264 9281
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 9215 11264 9216
rect 20944 9280 21264 9281
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 29520 9256 30000 9286
rect 20944 9215 21264 9216
rect 16573 9210 16639 9213
rect 23197 9210 23263 9213
rect 26417 9210 26483 9213
rect 16573 9208 17602 9210
rect 16573 9152 16578 9208
rect 16634 9152 17602 9208
rect 16573 9150 17602 9152
rect 16573 9147 16639 9150
rect 4429 9074 4495 9077
rect 4889 9074 4955 9077
rect 17401 9074 17467 9077
rect 4429 9072 17467 9074
rect 4429 9016 4434 9072
rect 4490 9016 4894 9072
rect 4950 9016 17406 9072
rect 17462 9016 17467 9072
rect 4429 9014 17467 9016
rect 17542 9074 17602 9150
rect 23197 9208 26483 9210
rect 23197 9152 23202 9208
rect 23258 9152 26422 9208
rect 26478 9152 26483 9208
rect 23197 9150 26483 9152
rect 23197 9147 23263 9150
rect 26417 9147 26483 9150
rect 25313 9074 25379 9077
rect 17542 9072 25379 9074
rect 17542 9016 25318 9072
rect 25374 9016 25379 9072
rect 17542 9014 25379 9016
rect 4429 9011 4495 9014
rect 4889 9011 4955 9014
rect 17401 9011 17467 9014
rect 25313 9011 25379 9014
rect 26509 8938 26575 8941
rect 25822 8936 26575 8938
rect 25822 8880 26514 8936
rect 26570 8880 26575 8936
rect 25822 8878 26575 8880
rect 19517 8802 19583 8805
rect 25037 8802 25103 8805
rect 19517 8800 25103 8802
rect 19517 8744 19522 8800
rect 19578 8744 25042 8800
rect 25098 8744 25103 8800
rect 19517 8742 25103 8744
rect 19517 8739 19583 8742
rect 25037 8739 25103 8742
rect 5944 8736 6264 8737
rect 0 8666 480 8696
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 8671 6264 8672
rect 15944 8736 16264 8737
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 8671 16264 8672
rect 2497 8666 2563 8669
rect 0 8664 2563 8666
rect 0 8608 2502 8664
rect 2558 8608 2563 8664
rect 0 8606 2563 8608
rect 0 8576 480 8606
rect 2497 8603 2563 8606
rect 19241 8666 19307 8669
rect 25822 8666 25882 8878
rect 26509 8875 26575 8878
rect 25944 8736 26264 8737
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 8671 26264 8672
rect 29520 8666 30000 8696
rect 19241 8664 25882 8666
rect 19241 8608 19246 8664
rect 19302 8608 25882 8664
rect 19241 8606 25882 8608
rect 26374 8606 30000 8666
rect 19241 8603 19307 8606
rect 8845 8530 8911 8533
rect 19701 8530 19767 8533
rect 8845 8528 19767 8530
rect 8845 8472 8850 8528
rect 8906 8472 19706 8528
rect 19762 8472 19767 8528
rect 8845 8470 19767 8472
rect 8845 8467 8911 8470
rect 19701 8467 19767 8470
rect 25497 8530 25563 8533
rect 26374 8530 26434 8606
rect 29520 8576 30000 8606
rect 25497 8528 26434 8530
rect 25497 8472 25502 8528
rect 25558 8472 26434 8528
rect 25497 8470 26434 8472
rect 25497 8467 25563 8470
rect 2773 8394 2839 8397
rect 5533 8394 5599 8397
rect 2773 8392 5599 8394
rect 2773 8336 2778 8392
rect 2834 8336 5538 8392
rect 5594 8336 5599 8392
rect 2773 8334 5599 8336
rect 2773 8331 2839 8334
rect 5533 8331 5599 8334
rect 7189 8394 7255 8397
rect 18597 8394 18663 8397
rect 19241 8394 19307 8397
rect 7189 8392 19307 8394
rect 7189 8336 7194 8392
rect 7250 8336 18602 8392
rect 18658 8336 19246 8392
rect 19302 8336 19307 8392
rect 7189 8334 19307 8336
rect 7189 8331 7255 8334
rect 18597 8331 18663 8334
rect 19241 8331 19307 8334
rect 10944 8192 11264 8193
rect 0 8122 480 8152
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 8127 11264 8128
rect 20944 8192 21264 8193
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 8127 21264 8128
rect 3601 8122 3667 8125
rect 0 8120 3667 8122
rect 0 8064 3606 8120
rect 3662 8064 3667 8120
rect 0 8062 3667 8064
rect 0 8032 480 8062
rect 3601 8059 3667 8062
rect 25497 8122 25563 8125
rect 29520 8122 30000 8152
rect 25497 8120 30000 8122
rect 25497 8064 25502 8120
rect 25558 8064 30000 8120
rect 25497 8062 30000 8064
rect 25497 8059 25563 8062
rect 29520 8032 30000 8062
rect 5349 7850 5415 7853
rect 7373 7850 7439 7853
rect 5349 7848 7439 7850
rect 5349 7792 5354 7848
rect 5410 7792 7378 7848
rect 7434 7792 7439 7848
rect 5349 7790 7439 7792
rect 5349 7787 5415 7790
rect 7373 7787 7439 7790
rect 8385 7850 8451 7853
rect 19057 7850 19123 7853
rect 19517 7850 19583 7853
rect 8385 7848 19583 7850
rect 8385 7792 8390 7848
rect 8446 7792 19062 7848
rect 19118 7792 19522 7848
rect 19578 7792 19583 7848
rect 8385 7790 19583 7792
rect 8385 7787 8451 7790
rect 19057 7787 19123 7790
rect 19517 7787 19583 7790
rect 5944 7648 6264 7649
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 7583 6264 7584
rect 15944 7648 16264 7649
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 7583 16264 7584
rect 25944 7648 26264 7649
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 7583 26264 7584
rect 0 7442 480 7472
rect 1485 7442 1551 7445
rect 0 7440 1551 7442
rect 0 7384 1490 7440
rect 1546 7384 1551 7440
rect 0 7382 1551 7384
rect 0 7352 480 7382
rect 1485 7379 1551 7382
rect 26601 7442 26667 7445
rect 29520 7442 30000 7472
rect 26601 7440 30000 7442
rect 26601 7384 26606 7440
rect 26662 7384 30000 7440
rect 26601 7382 30000 7384
rect 26601 7379 26667 7382
rect 29520 7352 30000 7382
rect 2037 7306 2103 7309
rect 11513 7306 11579 7309
rect 2037 7304 11579 7306
rect 2037 7248 2042 7304
rect 2098 7248 11518 7304
rect 11574 7248 11579 7304
rect 2037 7246 11579 7248
rect 2037 7243 2103 7246
rect 11513 7243 11579 7246
rect 19241 7306 19307 7309
rect 26509 7306 26575 7309
rect 19241 7304 26575 7306
rect 19241 7248 19246 7304
rect 19302 7248 26514 7304
rect 26570 7248 26575 7304
rect 19241 7246 26575 7248
rect 19241 7243 19307 7246
rect 26509 7243 26575 7246
rect 10944 7104 11264 7105
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 7039 11264 7040
rect 20944 7104 21264 7105
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 7039 21264 7040
rect 2405 7034 2471 7037
rect 3509 7034 3575 7037
rect 7925 7034 7991 7037
rect 2405 7032 7991 7034
rect 2405 6976 2410 7032
rect 2466 6976 3514 7032
rect 3570 6976 7930 7032
rect 7986 6976 7991 7032
rect 2405 6974 7991 6976
rect 2405 6971 2471 6974
rect 3509 6971 3575 6974
rect 7925 6971 7991 6974
rect 27705 7034 27771 7037
rect 27705 7032 27906 7034
rect 27705 6976 27710 7032
rect 27766 6976 27906 7032
rect 27705 6974 27906 6976
rect 27705 6971 27771 6974
rect 0 6898 480 6928
rect 2681 6898 2747 6901
rect 0 6896 2747 6898
rect 0 6840 2686 6896
rect 2742 6840 2747 6896
rect 0 6838 2747 6840
rect 27846 6898 27906 6974
rect 29520 6898 30000 6928
rect 27846 6838 30000 6898
rect 0 6808 480 6838
rect 2681 6835 2747 6838
rect 29520 6808 30000 6838
rect 5944 6560 6264 6561
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 6495 6264 6496
rect 15944 6560 16264 6561
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 6495 16264 6496
rect 25944 6560 26264 6561
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 6495 26264 6496
rect 0 6354 480 6384
rect 1577 6354 1643 6357
rect 0 6352 1643 6354
rect 0 6296 1582 6352
rect 1638 6296 1643 6352
rect 0 6294 1643 6296
rect 0 6264 480 6294
rect 1577 6291 1643 6294
rect 2405 6354 2471 6357
rect 16757 6354 16823 6357
rect 2405 6352 16823 6354
rect 2405 6296 2410 6352
rect 2466 6296 16762 6352
rect 16818 6296 16823 6352
rect 2405 6294 16823 6296
rect 2405 6291 2471 6294
rect 16757 6291 16823 6294
rect 26693 6354 26759 6357
rect 29520 6354 30000 6384
rect 26693 6352 30000 6354
rect 26693 6296 26698 6352
rect 26754 6296 30000 6352
rect 26693 6294 30000 6296
rect 26693 6291 26759 6294
rect 29520 6264 30000 6294
rect 10944 6016 11264 6017
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 5951 11264 5952
rect 20944 6016 21264 6017
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 5951 21264 5952
rect 1393 5810 1459 5813
rect 6913 5810 6979 5813
rect 1393 5808 6979 5810
rect 1393 5752 1398 5808
rect 1454 5752 6918 5808
rect 6974 5752 6979 5808
rect 1393 5750 6979 5752
rect 1393 5747 1459 5750
rect 6913 5747 6979 5750
rect 0 5674 480 5704
rect 1669 5674 1735 5677
rect 0 5672 1735 5674
rect 0 5616 1674 5672
rect 1730 5616 1735 5672
rect 0 5614 1735 5616
rect 0 5584 480 5614
rect 1669 5611 1735 5614
rect 27797 5674 27863 5677
rect 29520 5674 30000 5704
rect 27797 5672 30000 5674
rect 27797 5616 27802 5672
rect 27858 5616 30000 5672
rect 27797 5614 30000 5616
rect 27797 5611 27863 5614
rect 29520 5584 30000 5614
rect 5944 5472 6264 5473
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 5407 6264 5408
rect 15944 5472 16264 5473
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 5407 16264 5408
rect 25944 5472 26264 5473
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 5407 26264 5408
rect 12893 5266 12959 5269
rect 26417 5266 26483 5269
rect 12893 5264 26483 5266
rect 12893 5208 12898 5264
rect 12954 5208 26422 5264
rect 26478 5208 26483 5264
rect 12893 5206 26483 5208
rect 12893 5203 12959 5206
rect 26417 5203 26483 5206
rect 0 5130 480 5160
rect 2221 5130 2287 5133
rect 0 5128 2287 5130
rect 0 5072 2226 5128
rect 2282 5072 2287 5128
rect 0 5070 2287 5072
rect 0 5040 480 5070
rect 2221 5067 2287 5070
rect 26601 5130 26667 5133
rect 29520 5130 30000 5160
rect 26601 5128 30000 5130
rect 26601 5072 26606 5128
rect 26662 5072 30000 5128
rect 26601 5070 30000 5072
rect 26601 5067 26667 5070
rect 29520 5040 30000 5070
rect 10944 4928 11264 4929
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 4863 11264 4864
rect 20944 4928 21264 4929
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 4863 21264 4864
rect 25773 4586 25839 4589
rect 25773 4584 26434 4586
rect 25773 4528 25778 4584
rect 25834 4528 26434 4584
rect 25773 4526 26434 4528
rect 25773 4523 25839 4526
rect 0 4450 480 4480
rect 1853 4450 1919 4453
rect 0 4448 1919 4450
rect 0 4392 1858 4448
rect 1914 4392 1919 4448
rect 0 4390 1919 4392
rect 26374 4450 26434 4526
rect 29520 4450 30000 4480
rect 26374 4390 30000 4450
rect 0 4360 480 4390
rect 1853 4387 1919 4390
rect 5944 4384 6264 4385
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 4319 6264 4320
rect 15944 4384 16264 4385
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 4319 16264 4320
rect 25944 4384 26264 4385
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 29520 4360 30000 4390
rect 25944 4319 26264 4320
rect 2037 4042 2103 4045
rect 8109 4042 8175 4045
rect 2037 4040 8175 4042
rect 2037 3984 2042 4040
rect 2098 3984 8114 4040
rect 8170 3984 8175 4040
rect 2037 3982 8175 3984
rect 2037 3979 2103 3982
rect 8109 3979 8175 3982
rect 19885 4042 19951 4045
rect 26417 4042 26483 4045
rect 19885 4040 26483 4042
rect 19885 3984 19890 4040
rect 19946 3984 26422 4040
rect 26478 3984 26483 4040
rect 19885 3982 26483 3984
rect 19885 3979 19951 3982
rect 26417 3979 26483 3982
rect 0 3906 480 3936
rect 4337 3906 4403 3909
rect 0 3904 4403 3906
rect 0 3848 4342 3904
rect 4398 3848 4403 3904
rect 0 3846 4403 3848
rect 0 3816 480 3846
rect 4337 3843 4403 3846
rect 25681 3906 25747 3909
rect 29520 3906 30000 3936
rect 25681 3904 30000 3906
rect 25681 3848 25686 3904
rect 25742 3848 30000 3904
rect 25681 3846 30000 3848
rect 25681 3843 25747 3846
rect 10944 3840 11264 3841
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 3775 11264 3776
rect 20944 3840 21264 3841
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 29520 3816 30000 3846
rect 20944 3775 21264 3776
rect 3693 3498 3759 3501
rect 15561 3498 15627 3501
rect 3693 3496 15627 3498
rect 3693 3440 3698 3496
rect 3754 3440 15566 3496
rect 15622 3440 15627 3496
rect 3693 3438 15627 3440
rect 3693 3435 3759 3438
rect 15561 3435 15627 3438
rect 25589 3498 25655 3501
rect 25589 3496 26434 3498
rect 25589 3440 25594 3496
rect 25650 3440 26434 3496
rect 25589 3438 26434 3440
rect 25589 3435 25655 3438
rect 0 3362 480 3392
rect 565 3362 631 3365
rect 0 3360 631 3362
rect 0 3304 570 3360
rect 626 3304 631 3360
rect 0 3302 631 3304
rect 26374 3362 26434 3438
rect 29520 3362 30000 3392
rect 26374 3302 30000 3362
rect 0 3272 480 3302
rect 565 3299 631 3302
rect 5944 3296 6264 3297
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 3231 6264 3232
rect 15944 3296 16264 3297
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 3231 16264 3232
rect 25944 3296 26264 3297
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 29520 3272 30000 3302
rect 25944 3231 26264 3232
rect 26601 2818 26667 2821
rect 26601 2816 26802 2818
rect 26601 2760 26606 2816
rect 26662 2760 26802 2816
rect 26601 2758 26802 2760
rect 26601 2755 26667 2758
rect 10944 2752 11264 2753
rect 0 2682 480 2712
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2687 11264 2688
rect 20944 2752 21264 2753
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2687 21264 2688
rect 1577 2682 1643 2685
rect 0 2680 1643 2682
rect 0 2624 1582 2680
rect 1638 2624 1643 2680
rect 0 2622 1643 2624
rect 26742 2682 26802 2758
rect 29520 2682 30000 2712
rect 26742 2622 30000 2682
rect 0 2592 480 2622
rect 1577 2619 1643 2622
rect 29520 2592 30000 2622
rect 7465 2410 7531 2413
rect 11145 2410 11211 2413
rect 7465 2408 11211 2410
rect 7465 2352 7470 2408
rect 7526 2352 11150 2408
rect 11206 2352 11211 2408
rect 7465 2350 11211 2352
rect 7465 2347 7531 2350
rect 11145 2347 11211 2350
rect 25405 2410 25471 2413
rect 25405 2408 27906 2410
rect 25405 2352 25410 2408
rect 25466 2352 27906 2408
rect 25405 2350 27906 2352
rect 25405 2347 25471 2350
rect 5944 2208 6264 2209
rect 0 2138 480 2168
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2143 6264 2144
rect 15944 2208 16264 2209
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2143 16264 2144
rect 25944 2208 26264 2209
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2143 26264 2144
rect 2773 2138 2839 2141
rect 0 2136 2839 2138
rect 0 2080 2778 2136
rect 2834 2080 2839 2136
rect 0 2078 2839 2080
rect 27846 2138 27906 2350
rect 29520 2138 30000 2168
rect 27846 2078 30000 2138
rect 0 2048 480 2078
rect 2773 2075 2839 2078
rect 29520 2048 30000 2078
rect 0 1458 480 1488
rect 1485 1458 1551 1461
rect 0 1456 1551 1458
rect 0 1400 1490 1456
rect 1546 1400 1551 1456
rect 0 1398 1551 1400
rect 0 1368 480 1398
rect 1485 1395 1551 1398
rect 25865 1458 25931 1461
rect 29520 1458 30000 1488
rect 25865 1456 30000 1458
rect 25865 1400 25870 1456
rect 25926 1400 30000 1456
rect 25865 1398 30000 1400
rect 25865 1395 25931 1398
rect 29520 1368 30000 1398
rect 0 914 480 944
rect 2681 914 2747 917
rect 0 912 2747 914
rect 0 856 2686 912
rect 2742 856 2747 912
rect 0 854 2747 856
rect 0 824 480 854
rect 2681 851 2747 854
rect 26877 914 26943 917
rect 29520 914 30000 944
rect 26877 912 30000 914
rect 26877 856 26882 912
rect 26938 856 30000 912
rect 26877 854 30000 856
rect 26877 851 26943 854
rect 29520 824 30000 854
rect 0 370 480 400
rect 4061 370 4127 373
rect 0 368 4127 370
rect 0 312 4066 368
rect 4122 312 4127 368
rect 0 310 4127 312
rect 0 280 480 310
rect 4061 307 4127 310
rect 26785 370 26851 373
rect 29520 370 30000 400
rect 26785 368 30000 370
rect 26785 312 26790 368
rect 26846 312 30000 368
rect 26785 310 30000 312
rect 26785 307 26851 310
rect 29520 280 30000 310
<< via3 >>
rect 5952 21788 6016 21792
rect 5952 21732 5956 21788
rect 5956 21732 6012 21788
rect 6012 21732 6016 21788
rect 5952 21728 6016 21732
rect 6032 21788 6096 21792
rect 6032 21732 6036 21788
rect 6036 21732 6092 21788
rect 6092 21732 6096 21788
rect 6032 21728 6096 21732
rect 6112 21788 6176 21792
rect 6112 21732 6116 21788
rect 6116 21732 6172 21788
rect 6172 21732 6176 21788
rect 6112 21728 6176 21732
rect 6192 21788 6256 21792
rect 6192 21732 6196 21788
rect 6196 21732 6252 21788
rect 6252 21732 6256 21788
rect 6192 21728 6256 21732
rect 15952 21788 16016 21792
rect 15952 21732 15956 21788
rect 15956 21732 16012 21788
rect 16012 21732 16016 21788
rect 15952 21728 16016 21732
rect 16032 21788 16096 21792
rect 16032 21732 16036 21788
rect 16036 21732 16092 21788
rect 16092 21732 16096 21788
rect 16032 21728 16096 21732
rect 16112 21788 16176 21792
rect 16112 21732 16116 21788
rect 16116 21732 16172 21788
rect 16172 21732 16176 21788
rect 16112 21728 16176 21732
rect 16192 21788 16256 21792
rect 16192 21732 16196 21788
rect 16196 21732 16252 21788
rect 16252 21732 16256 21788
rect 16192 21728 16256 21732
rect 25952 21788 26016 21792
rect 25952 21732 25956 21788
rect 25956 21732 26012 21788
rect 26012 21732 26016 21788
rect 25952 21728 26016 21732
rect 26032 21788 26096 21792
rect 26032 21732 26036 21788
rect 26036 21732 26092 21788
rect 26092 21732 26096 21788
rect 26032 21728 26096 21732
rect 26112 21788 26176 21792
rect 26112 21732 26116 21788
rect 26116 21732 26172 21788
rect 26172 21732 26176 21788
rect 26112 21728 26176 21732
rect 26192 21788 26256 21792
rect 26192 21732 26196 21788
rect 26196 21732 26252 21788
rect 26252 21732 26256 21788
rect 26192 21728 26256 21732
rect 10952 21244 11016 21248
rect 10952 21188 10956 21244
rect 10956 21188 11012 21244
rect 11012 21188 11016 21244
rect 10952 21184 11016 21188
rect 11032 21244 11096 21248
rect 11032 21188 11036 21244
rect 11036 21188 11092 21244
rect 11092 21188 11096 21244
rect 11032 21184 11096 21188
rect 11112 21244 11176 21248
rect 11112 21188 11116 21244
rect 11116 21188 11172 21244
rect 11172 21188 11176 21244
rect 11112 21184 11176 21188
rect 11192 21244 11256 21248
rect 11192 21188 11196 21244
rect 11196 21188 11252 21244
rect 11252 21188 11256 21244
rect 11192 21184 11256 21188
rect 20952 21244 21016 21248
rect 20952 21188 20956 21244
rect 20956 21188 21012 21244
rect 21012 21188 21016 21244
rect 20952 21184 21016 21188
rect 21032 21244 21096 21248
rect 21032 21188 21036 21244
rect 21036 21188 21092 21244
rect 21092 21188 21096 21244
rect 21032 21184 21096 21188
rect 21112 21244 21176 21248
rect 21112 21188 21116 21244
rect 21116 21188 21172 21244
rect 21172 21188 21176 21244
rect 21112 21184 21176 21188
rect 21192 21244 21256 21248
rect 21192 21188 21196 21244
rect 21196 21188 21252 21244
rect 21252 21188 21256 21244
rect 21192 21184 21256 21188
rect 5952 20700 6016 20704
rect 5952 20644 5956 20700
rect 5956 20644 6012 20700
rect 6012 20644 6016 20700
rect 5952 20640 6016 20644
rect 6032 20700 6096 20704
rect 6032 20644 6036 20700
rect 6036 20644 6092 20700
rect 6092 20644 6096 20700
rect 6032 20640 6096 20644
rect 6112 20700 6176 20704
rect 6112 20644 6116 20700
rect 6116 20644 6172 20700
rect 6172 20644 6176 20700
rect 6112 20640 6176 20644
rect 6192 20700 6256 20704
rect 6192 20644 6196 20700
rect 6196 20644 6252 20700
rect 6252 20644 6256 20700
rect 6192 20640 6256 20644
rect 15952 20700 16016 20704
rect 15952 20644 15956 20700
rect 15956 20644 16012 20700
rect 16012 20644 16016 20700
rect 15952 20640 16016 20644
rect 16032 20700 16096 20704
rect 16032 20644 16036 20700
rect 16036 20644 16092 20700
rect 16092 20644 16096 20700
rect 16032 20640 16096 20644
rect 16112 20700 16176 20704
rect 16112 20644 16116 20700
rect 16116 20644 16172 20700
rect 16172 20644 16176 20700
rect 16112 20640 16176 20644
rect 16192 20700 16256 20704
rect 16192 20644 16196 20700
rect 16196 20644 16252 20700
rect 16252 20644 16256 20700
rect 16192 20640 16256 20644
rect 25952 20700 26016 20704
rect 25952 20644 25956 20700
rect 25956 20644 26012 20700
rect 26012 20644 26016 20700
rect 25952 20640 26016 20644
rect 26032 20700 26096 20704
rect 26032 20644 26036 20700
rect 26036 20644 26092 20700
rect 26092 20644 26096 20700
rect 26032 20640 26096 20644
rect 26112 20700 26176 20704
rect 26112 20644 26116 20700
rect 26116 20644 26172 20700
rect 26172 20644 26176 20700
rect 26112 20640 26176 20644
rect 26192 20700 26256 20704
rect 26192 20644 26196 20700
rect 26196 20644 26252 20700
rect 26252 20644 26256 20700
rect 26192 20640 26256 20644
rect 10952 20156 11016 20160
rect 10952 20100 10956 20156
rect 10956 20100 11012 20156
rect 11012 20100 11016 20156
rect 10952 20096 11016 20100
rect 11032 20156 11096 20160
rect 11032 20100 11036 20156
rect 11036 20100 11092 20156
rect 11092 20100 11096 20156
rect 11032 20096 11096 20100
rect 11112 20156 11176 20160
rect 11112 20100 11116 20156
rect 11116 20100 11172 20156
rect 11172 20100 11176 20156
rect 11112 20096 11176 20100
rect 11192 20156 11256 20160
rect 11192 20100 11196 20156
rect 11196 20100 11252 20156
rect 11252 20100 11256 20156
rect 11192 20096 11256 20100
rect 20952 20156 21016 20160
rect 20952 20100 20956 20156
rect 20956 20100 21012 20156
rect 21012 20100 21016 20156
rect 20952 20096 21016 20100
rect 21032 20156 21096 20160
rect 21032 20100 21036 20156
rect 21036 20100 21092 20156
rect 21092 20100 21096 20156
rect 21032 20096 21096 20100
rect 21112 20156 21176 20160
rect 21112 20100 21116 20156
rect 21116 20100 21172 20156
rect 21172 20100 21176 20156
rect 21112 20096 21176 20100
rect 21192 20156 21256 20160
rect 21192 20100 21196 20156
rect 21196 20100 21252 20156
rect 21252 20100 21256 20156
rect 21192 20096 21256 20100
rect 9628 19620 9692 19684
rect 5952 19612 6016 19616
rect 5952 19556 5956 19612
rect 5956 19556 6012 19612
rect 6012 19556 6016 19612
rect 5952 19552 6016 19556
rect 6032 19612 6096 19616
rect 6032 19556 6036 19612
rect 6036 19556 6092 19612
rect 6092 19556 6096 19612
rect 6032 19552 6096 19556
rect 6112 19612 6176 19616
rect 6112 19556 6116 19612
rect 6116 19556 6172 19612
rect 6172 19556 6176 19612
rect 6112 19552 6176 19556
rect 6192 19612 6256 19616
rect 6192 19556 6196 19612
rect 6196 19556 6252 19612
rect 6252 19556 6256 19612
rect 6192 19552 6256 19556
rect 15952 19612 16016 19616
rect 15952 19556 15956 19612
rect 15956 19556 16012 19612
rect 16012 19556 16016 19612
rect 15952 19552 16016 19556
rect 16032 19612 16096 19616
rect 16032 19556 16036 19612
rect 16036 19556 16092 19612
rect 16092 19556 16096 19612
rect 16032 19552 16096 19556
rect 16112 19612 16176 19616
rect 16112 19556 16116 19612
rect 16116 19556 16172 19612
rect 16172 19556 16176 19612
rect 16112 19552 16176 19556
rect 16192 19612 16256 19616
rect 16192 19556 16196 19612
rect 16196 19556 16252 19612
rect 16252 19556 16256 19612
rect 16192 19552 16256 19556
rect 25952 19612 26016 19616
rect 25952 19556 25956 19612
rect 25956 19556 26012 19612
rect 26012 19556 26016 19612
rect 25952 19552 26016 19556
rect 26032 19612 26096 19616
rect 26032 19556 26036 19612
rect 26036 19556 26092 19612
rect 26092 19556 26096 19612
rect 26032 19552 26096 19556
rect 26112 19612 26176 19616
rect 26112 19556 26116 19612
rect 26116 19556 26172 19612
rect 26172 19556 26176 19612
rect 26112 19552 26176 19556
rect 26192 19612 26256 19616
rect 26192 19556 26196 19612
rect 26196 19556 26252 19612
rect 26252 19556 26256 19612
rect 26192 19552 26256 19556
rect 9628 19408 9692 19412
rect 9628 19352 9642 19408
rect 9642 19352 9692 19408
rect 9628 19348 9692 19352
rect 10952 19068 11016 19072
rect 10952 19012 10956 19068
rect 10956 19012 11012 19068
rect 11012 19012 11016 19068
rect 10952 19008 11016 19012
rect 11032 19068 11096 19072
rect 11032 19012 11036 19068
rect 11036 19012 11092 19068
rect 11092 19012 11096 19068
rect 11032 19008 11096 19012
rect 11112 19068 11176 19072
rect 11112 19012 11116 19068
rect 11116 19012 11172 19068
rect 11172 19012 11176 19068
rect 11112 19008 11176 19012
rect 11192 19068 11256 19072
rect 11192 19012 11196 19068
rect 11196 19012 11252 19068
rect 11252 19012 11256 19068
rect 11192 19008 11256 19012
rect 20952 19068 21016 19072
rect 20952 19012 20956 19068
rect 20956 19012 21012 19068
rect 21012 19012 21016 19068
rect 20952 19008 21016 19012
rect 21032 19068 21096 19072
rect 21032 19012 21036 19068
rect 21036 19012 21092 19068
rect 21092 19012 21096 19068
rect 21032 19008 21096 19012
rect 21112 19068 21176 19072
rect 21112 19012 21116 19068
rect 21116 19012 21172 19068
rect 21172 19012 21176 19068
rect 21112 19008 21176 19012
rect 21192 19068 21256 19072
rect 21192 19012 21196 19068
rect 21196 19012 21252 19068
rect 21252 19012 21256 19068
rect 21192 19008 21256 19012
rect 5952 18524 6016 18528
rect 5952 18468 5956 18524
rect 5956 18468 6012 18524
rect 6012 18468 6016 18524
rect 5952 18464 6016 18468
rect 6032 18524 6096 18528
rect 6032 18468 6036 18524
rect 6036 18468 6092 18524
rect 6092 18468 6096 18524
rect 6032 18464 6096 18468
rect 6112 18524 6176 18528
rect 6112 18468 6116 18524
rect 6116 18468 6172 18524
rect 6172 18468 6176 18524
rect 6112 18464 6176 18468
rect 6192 18524 6256 18528
rect 6192 18468 6196 18524
rect 6196 18468 6252 18524
rect 6252 18468 6256 18524
rect 6192 18464 6256 18468
rect 15952 18524 16016 18528
rect 15952 18468 15956 18524
rect 15956 18468 16012 18524
rect 16012 18468 16016 18524
rect 15952 18464 16016 18468
rect 16032 18524 16096 18528
rect 16032 18468 16036 18524
rect 16036 18468 16092 18524
rect 16092 18468 16096 18524
rect 16032 18464 16096 18468
rect 16112 18524 16176 18528
rect 16112 18468 16116 18524
rect 16116 18468 16172 18524
rect 16172 18468 16176 18524
rect 16112 18464 16176 18468
rect 16192 18524 16256 18528
rect 16192 18468 16196 18524
rect 16196 18468 16252 18524
rect 16252 18468 16256 18524
rect 16192 18464 16256 18468
rect 25952 18524 26016 18528
rect 25952 18468 25956 18524
rect 25956 18468 26012 18524
rect 26012 18468 26016 18524
rect 25952 18464 26016 18468
rect 26032 18524 26096 18528
rect 26032 18468 26036 18524
rect 26036 18468 26092 18524
rect 26092 18468 26096 18524
rect 26032 18464 26096 18468
rect 26112 18524 26176 18528
rect 26112 18468 26116 18524
rect 26116 18468 26172 18524
rect 26172 18468 26176 18524
rect 26112 18464 26176 18468
rect 26192 18524 26256 18528
rect 26192 18468 26196 18524
rect 26196 18468 26252 18524
rect 26252 18468 26256 18524
rect 26192 18464 26256 18468
rect 10952 17980 11016 17984
rect 10952 17924 10956 17980
rect 10956 17924 11012 17980
rect 11012 17924 11016 17980
rect 10952 17920 11016 17924
rect 11032 17980 11096 17984
rect 11032 17924 11036 17980
rect 11036 17924 11092 17980
rect 11092 17924 11096 17980
rect 11032 17920 11096 17924
rect 11112 17980 11176 17984
rect 11112 17924 11116 17980
rect 11116 17924 11172 17980
rect 11172 17924 11176 17980
rect 11112 17920 11176 17924
rect 11192 17980 11256 17984
rect 11192 17924 11196 17980
rect 11196 17924 11252 17980
rect 11252 17924 11256 17980
rect 11192 17920 11256 17924
rect 20952 17980 21016 17984
rect 20952 17924 20956 17980
rect 20956 17924 21012 17980
rect 21012 17924 21016 17980
rect 20952 17920 21016 17924
rect 21032 17980 21096 17984
rect 21032 17924 21036 17980
rect 21036 17924 21092 17980
rect 21092 17924 21096 17980
rect 21032 17920 21096 17924
rect 21112 17980 21176 17984
rect 21112 17924 21116 17980
rect 21116 17924 21172 17980
rect 21172 17924 21176 17980
rect 21112 17920 21176 17924
rect 21192 17980 21256 17984
rect 21192 17924 21196 17980
rect 21196 17924 21252 17980
rect 21252 17924 21256 17980
rect 21192 17920 21256 17924
rect 5952 17436 6016 17440
rect 5952 17380 5956 17436
rect 5956 17380 6012 17436
rect 6012 17380 6016 17436
rect 5952 17376 6016 17380
rect 6032 17436 6096 17440
rect 6032 17380 6036 17436
rect 6036 17380 6092 17436
rect 6092 17380 6096 17436
rect 6032 17376 6096 17380
rect 6112 17436 6176 17440
rect 6112 17380 6116 17436
rect 6116 17380 6172 17436
rect 6172 17380 6176 17436
rect 6112 17376 6176 17380
rect 6192 17436 6256 17440
rect 6192 17380 6196 17436
rect 6196 17380 6252 17436
rect 6252 17380 6256 17436
rect 6192 17376 6256 17380
rect 15952 17436 16016 17440
rect 15952 17380 15956 17436
rect 15956 17380 16012 17436
rect 16012 17380 16016 17436
rect 15952 17376 16016 17380
rect 16032 17436 16096 17440
rect 16032 17380 16036 17436
rect 16036 17380 16092 17436
rect 16092 17380 16096 17436
rect 16032 17376 16096 17380
rect 16112 17436 16176 17440
rect 16112 17380 16116 17436
rect 16116 17380 16172 17436
rect 16172 17380 16176 17436
rect 16112 17376 16176 17380
rect 16192 17436 16256 17440
rect 16192 17380 16196 17436
rect 16196 17380 16252 17436
rect 16252 17380 16256 17436
rect 16192 17376 16256 17380
rect 25952 17436 26016 17440
rect 25952 17380 25956 17436
rect 25956 17380 26012 17436
rect 26012 17380 26016 17436
rect 25952 17376 26016 17380
rect 26032 17436 26096 17440
rect 26032 17380 26036 17436
rect 26036 17380 26092 17436
rect 26092 17380 26096 17436
rect 26032 17376 26096 17380
rect 26112 17436 26176 17440
rect 26112 17380 26116 17436
rect 26116 17380 26172 17436
rect 26172 17380 26176 17436
rect 26112 17376 26176 17380
rect 26192 17436 26256 17440
rect 26192 17380 26196 17436
rect 26196 17380 26252 17436
rect 26252 17380 26256 17436
rect 26192 17376 26256 17380
rect 10952 16892 11016 16896
rect 10952 16836 10956 16892
rect 10956 16836 11012 16892
rect 11012 16836 11016 16892
rect 10952 16832 11016 16836
rect 11032 16892 11096 16896
rect 11032 16836 11036 16892
rect 11036 16836 11092 16892
rect 11092 16836 11096 16892
rect 11032 16832 11096 16836
rect 11112 16892 11176 16896
rect 11112 16836 11116 16892
rect 11116 16836 11172 16892
rect 11172 16836 11176 16892
rect 11112 16832 11176 16836
rect 11192 16892 11256 16896
rect 11192 16836 11196 16892
rect 11196 16836 11252 16892
rect 11252 16836 11256 16892
rect 11192 16832 11256 16836
rect 20952 16892 21016 16896
rect 20952 16836 20956 16892
rect 20956 16836 21012 16892
rect 21012 16836 21016 16892
rect 20952 16832 21016 16836
rect 21032 16892 21096 16896
rect 21032 16836 21036 16892
rect 21036 16836 21092 16892
rect 21092 16836 21096 16892
rect 21032 16832 21096 16836
rect 21112 16892 21176 16896
rect 21112 16836 21116 16892
rect 21116 16836 21172 16892
rect 21172 16836 21176 16892
rect 21112 16832 21176 16836
rect 21192 16892 21256 16896
rect 21192 16836 21196 16892
rect 21196 16836 21252 16892
rect 21252 16836 21256 16892
rect 21192 16832 21256 16836
rect 5952 16348 6016 16352
rect 5952 16292 5956 16348
rect 5956 16292 6012 16348
rect 6012 16292 6016 16348
rect 5952 16288 6016 16292
rect 6032 16348 6096 16352
rect 6032 16292 6036 16348
rect 6036 16292 6092 16348
rect 6092 16292 6096 16348
rect 6032 16288 6096 16292
rect 6112 16348 6176 16352
rect 6112 16292 6116 16348
rect 6116 16292 6172 16348
rect 6172 16292 6176 16348
rect 6112 16288 6176 16292
rect 6192 16348 6256 16352
rect 6192 16292 6196 16348
rect 6196 16292 6252 16348
rect 6252 16292 6256 16348
rect 6192 16288 6256 16292
rect 15952 16348 16016 16352
rect 15952 16292 15956 16348
rect 15956 16292 16012 16348
rect 16012 16292 16016 16348
rect 15952 16288 16016 16292
rect 16032 16348 16096 16352
rect 16032 16292 16036 16348
rect 16036 16292 16092 16348
rect 16092 16292 16096 16348
rect 16032 16288 16096 16292
rect 16112 16348 16176 16352
rect 16112 16292 16116 16348
rect 16116 16292 16172 16348
rect 16172 16292 16176 16348
rect 16112 16288 16176 16292
rect 16192 16348 16256 16352
rect 16192 16292 16196 16348
rect 16196 16292 16252 16348
rect 16252 16292 16256 16348
rect 16192 16288 16256 16292
rect 25952 16348 26016 16352
rect 25952 16292 25956 16348
rect 25956 16292 26012 16348
rect 26012 16292 26016 16348
rect 25952 16288 26016 16292
rect 26032 16348 26096 16352
rect 26032 16292 26036 16348
rect 26036 16292 26092 16348
rect 26092 16292 26096 16348
rect 26032 16288 26096 16292
rect 26112 16348 26176 16352
rect 26112 16292 26116 16348
rect 26116 16292 26172 16348
rect 26172 16292 26176 16348
rect 26112 16288 26176 16292
rect 26192 16348 26256 16352
rect 26192 16292 26196 16348
rect 26196 16292 26252 16348
rect 26252 16292 26256 16348
rect 26192 16288 26256 16292
rect 10952 15804 11016 15808
rect 10952 15748 10956 15804
rect 10956 15748 11012 15804
rect 11012 15748 11016 15804
rect 10952 15744 11016 15748
rect 11032 15804 11096 15808
rect 11032 15748 11036 15804
rect 11036 15748 11092 15804
rect 11092 15748 11096 15804
rect 11032 15744 11096 15748
rect 11112 15804 11176 15808
rect 11112 15748 11116 15804
rect 11116 15748 11172 15804
rect 11172 15748 11176 15804
rect 11112 15744 11176 15748
rect 11192 15804 11256 15808
rect 11192 15748 11196 15804
rect 11196 15748 11252 15804
rect 11252 15748 11256 15804
rect 11192 15744 11256 15748
rect 20952 15804 21016 15808
rect 20952 15748 20956 15804
rect 20956 15748 21012 15804
rect 21012 15748 21016 15804
rect 20952 15744 21016 15748
rect 21032 15804 21096 15808
rect 21032 15748 21036 15804
rect 21036 15748 21092 15804
rect 21092 15748 21096 15804
rect 21032 15744 21096 15748
rect 21112 15804 21176 15808
rect 21112 15748 21116 15804
rect 21116 15748 21172 15804
rect 21172 15748 21176 15804
rect 21112 15744 21176 15748
rect 21192 15804 21256 15808
rect 21192 15748 21196 15804
rect 21196 15748 21252 15804
rect 21252 15748 21256 15804
rect 21192 15744 21256 15748
rect 5952 15260 6016 15264
rect 5952 15204 5956 15260
rect 5956 15204 6012 15260
rect 6012 15204 6016 15260
rect 5952 15200 6016 15204
rect 6032 15260 6096 15264
rect 6032 15204 6036 15260
rect 6036 15204 6092 15260
rect 6092 15204 6096 15260
rect 6032 15200 6096 15204
rect 6112 15260 6176 15264
rect 6112 15204 6116 15260
rect 6116 15204 6172 15260
rect 6172 15204 6176 15260
rect 6112 15200 6176 15204
rect 6192 15260 6256 15264
rect 6192 15204 6196 15260
rect 6196 15204 6252 15260
rect 6252 15204 6256 15260
rect 6192 15200 6256 15204
rect 15952 15260 16016 15264
rect 15952 15204 15956 15260
rect 15956 15204 16012 15260
rect 16012 15204 16016 15260
rect 15952 15200 16016 15204
rect 16032 15260 16096 15264
rect 16032 15204 16036 15260
rect 16036 15204 16092 15260
rect 16092 15204 16096 15260
rect 16032 15200 16096 15204
rect 16112 15260 16176 15264
rect 16112 15204 16116 15260
rect 16116 15204 16172 15260
rect 16172 15204 16176 15260
rect 16112 15200 16176 15204
rect 16192 15260 16256 15264
rect 16192 15204 16196 15260
rect 16196 15204 16252 15260
rect 16252 15204 16256 15260
rect 16192 15200 16256 15204
rect 25952 15260 26016 15264
rect 25952 15204 25956 15260
rect 25956 15204 26012 15260
rect 26012 15204 26016 15260
rect 25952 15200 26016 15204
rect 26032 15260 26096 15264
rect 26032 15204 26036 15260
rect 26036 15204 26092 15260
rect 26092 15204 26096 15260
rect 26032 15200 26096 15204
rect 26112 15260 26176 15264
rect 26112 15204 26116 15260
rect 26116 15204 26172 15260
rect 26172 15204 26176 15260
rect 26112 15200 26176 15204
rect 26192 15260 26256 15264
rect 26192 15204 26196 15260
rect 26196 15204 26252 15260
rect 26252 15204 26256 15260
rect 26192 15200 26256 15204
rect 10952 14716 11016 14720
rect 10952 14660 10956 14716
rect 10956 14660 11012 14716
rect 11012 14660 11016 14716
rect 10952 14656 11016 14660
rect 11032 14716 11096 14720
rect 11032 14660 11036 14716
rect 11036 14660 11092 14716
rect 11092 14660 11096 14716
rect 11032 14656 11096 14660
rect 11112 14716 11176 14720
rect 11112 14660 11116 14716
rect 11116 14660 11172 14716
rect 11172 14660 11176 14716
rect 11112 14656 11176 14660
rect 11192 14716 11256 14720
rect 11192 14660 11196 14716
rect 11196 14660 11252 14716
rect 11252 14660 11256 14716
rect 11192 14656 11256 14660
rect 20952 14716 21016 14720
rect 20952 14660 20956 14716
rect 20956 14660 21012 14716
rect 21012 14660 21016 14716
rect 20952 14656 21016 14660
rect 21032 14716 21096 14720
rect 21032 14660 21036 14716
rect 21036 14660 21092 14716
rect 21092 14660 21096 14716
rect 21032 14656 21096 14660
rect 21112 14716 21176 14720
rect 21112 14660 21116 14716
rect 21116 14660 21172 14716
rect 21172 14660 21176 14716
rect 21112 14656 21176 14660
rect 21192 14716 21256 14720
rect 21192 14660 21196 14716
rect 21196 14660 21252 14716
rect 21252 14660 21256 14716
rect 21192 14656 21256 14660
rect 5952 14172 6016 14176
rect 5952 14116 5956 14172
rect 5956 14116 6012 14172
rect 6012 14116 6016 14172
rect 5952 14112 6016 14116
rect 6032 14172 6096 14176
rect 6032 14116 6036 14172
rect 6036 14116 6092 14172
rect 6092 14116 6096 14172
rect 6032 14112 6096 14116
rect 6112 14172 6176 14176
rect 6112 14116 6116 14172
rect 6116 14116 6172 14172
rect 6172 14116 6176 14172
rect 6112 14112 6176 14116
rect 6192 14172 6256 14176
rect 6192 14116 6196 14172
rect 6196 14116 6252 14172
rect 6252 14116 6256 14172
rect 6192 14112 6256 14116
rect 15952 14172 16016 14176
rect 15952 14116 15956 14172
rect 15956 14116 16012 14172
rect 16012 14116 16016 14172
rect 15952 14112 16016 14116
rect 16032 14172 16096 14176
rect 16032 14116 16036 14172
rect 16036 14116 16092 14172
rect 16092 14116 16096 14172
rect 16032 14112 16096 14116
rect 16112 14172 16176 14176
rect 16112 14116 16116 14172
rect 16116 14116 16172 14172
rect 16172 14116 16176 14172
rect 16112 14112 16176 14116
rect 16192 14172 16256 14176
rect 16192 14116 16196 14172
rect 16196 14116 16252 14172
rect 16252 14116 16256 14172
rect 16192 14112 16256 14116
rect 25952 14172 26016 14176
rect 25952 14116 25956 14172
rect 25956 14116 26012 14172
rect 26012 14116 26016 14172
rect 25952 14112 26016 14116
rect 26032 14172 26096 14176
rect 26032 14116 26036 14172
rect 26036 14116 26092 14172
rect 26092 14116 26096 14172
rect 26032 14112 26096 14116
rect 26112 14172 26176 14176
rect 26112 14116 26116 14172
rect 26116 14116 26172 14172
rect 26172 14116 26176 14172
rect 26112 14112 26176 14116
rect 26192 14172 26256 14176
rect 26192 14116 26196 14172
rect 26196 14116 26252 14172
rect 26252 14116 26256 14172
rect 26192 14112 26256 14116
rect 10952 13628 11016 13632
rect 10952 13572 10956 13628
rect 10956 13572 11012 13628
rect 11012 13572 11016 13628
rect 10952 13568 11016 13572
rect 11032 13628 11096 13632
rect 11032 13572 11036 13628
rect 11036 13572 11092 13628
rect 11092 13572 11096 13628
rect 11032 13568 11096 13572
rect 11112 13628 11176 13632
rect 11112 13572 11116 13628
rect 11116 13572 11172 13628
rect 11172 13572 11176 13628
rect 11112 13568 11176 13572
rect 11192 13628 11256 13632
rect 11192 13572 11196 13628
rect 11196 13572 11252 13628
rect 11252 13572 11256 13628
rect 11192 13568 11256 13572
rect 20952 13628 21016 13632
rect 20952 13572 20956 13628
rect 20956 13572 21012 13628
rect 21012 13572 21016 13628
rect 20952 13568 21016 13572
rect 21032 13628 21096 13632
rect 21032 13572 21036 13628
rect 21036 13572 21092 13628
rect 21092 13572 21096 13628
rect 21032 13568 21096 13572
rect 21112 13628 21176 13632
rect 21112 13572 21116 13628
rect 21116 13572 21172 13628
rect 21172 13572 21176 13628
rect 21112 13568 21176 13572
rect 21192 13628 21256 13632
rect 21192 13572 21196 13628
rect 21196 13572 21252 13628
rect 21252 13572 21256 13628
rect 21192 13568 21256 13572
rect 5952 13084 6016 13088
rect 5952 13028 5956 13084
rect 5956 13028 6012 13084
rect 6012 13028 6016 13084
rect 5952 13024 6016 13028
rect 6032 13084 6096 13088
rect 6032 13028 6036 13084
rect 6036 13028 6092 13084
rect 6092 13028 6096 13084
rect 6032 13024 6096 13028
rect 6112 13084 6176 13088
rect 6112 13028 6116 13084
rect 6116 13028 6172 13084
rect 6172 13028 6176 13084
rect 6112 13024 6176 13028
rect 6192 13084 6256 13088
rect 6192 13028 6196 13084
rect 6196 13028 6252 13084
rect 6252 13028 6256 13084
rect 6192 13024 6256 13028
rect 15952 13084 16016 13088
rect 15952 13028 15956 13084
rect 15956 13028 16012 13084
rect 16012 13028 16016 13084
rect 15952 13024 16016 13028
rect 16032 13084 16096 13088
rect 16032 13028 16036 13084
rect 16036 13028 16092 13084
rect 16092 13028 16096 13084
rect 16032 13024 16096 13028
rect 16112 13084 16176 13088
rect 16112 13028 16116 13084
rect 16116 13028 16172 13084
rect 16172 13028 16176 13084
rect 16112 13024 16176 13028
rect 16192 13084 16256 13088
rect 16192 13028 16196 13084
rect 16196 13028 16252 13084
rect 16252 13028 16256 13084
rect 16192 13024 16256 13028
rect 25952 13084 26016 13088
rect 25952 13028 25956 13084
rect 25956 13028 26012 13084
rect 26012 13028 26016 13084
rect 25952 13024 26016 13028
rect 26032 13084 26096 13088
rect 26032 13028 26036 13084
rect 26036 13028 26092 13084
rect 26092 13028 26096 13084
rect 26032 13024 26096 13028
rect 26112 13084 26176 13088
rect 26112 13028 26116 13084
rect 26116 13028 26172 13084
rect 26172 13028 26176 13084
rect 26112 13024 26176 13028
rect 26192 13084 26256 13088
rect 26192 13028 26196 13084
rect 26196 13028 26252 13084
rect 26252 13028 26256 13084
rect 26192 13024 26256 13028
rect 10952 12540 11016 12544
rect 10952 12484 10956 12540
rect 10956 12484 11012 12540
rect 11012 12484 11016 12540
rect 10952 12480 11016 12484
rect 11032 12540 11096 12544
rect 11032 12484 11036 12540
rect 11036 12484 11092 12540
rect 11092 12484 11096 12540
rect 11032 12480 11096 12484
rect 11112 12540 11176 12544
rect 11112 12484 11116 12540
rect 11116 12484 11172 12540
rect 11172 12484 11176 12540
rect 11112 12480 11176 12484
rect 11192 12540 11256 12544
rect 11192 12484 11196 12540
rect 11196 12484 11252 12540
rect 11252 12484 11256 12540
rect 11192 12480 11256 12484
rect 20952 12540 21016 12544
rect 20952 12484 20956 12540
rect 20956 12484 21012 12540
rect 21012 12484 21016 12540
rect 20952 12480 21016 12484
rect 21032 12540 21096 12544
rect 21032 12484 21036 12540
rect 21036 12484 21092 12540
rect 21092 12484 21096 12540
rect 21032 12480 21096 12484
rect 21112 12540 21176 12544
rect 21112 12484 21116 12540
rect 21116 12484 21172 12540
rect 21172 12484 21176 12540
rect 21112 12480 21176 12484
rect 21192 12540 21256 12544
rect 21192 12484 21196 12540
rect 21196 12484 21252 12540
rect 21252 12484 21256 12540
rect 21192 12480 21256 12484
rect 5952 11996 6016 12000
rect 5952 11940 5956 11996
rect 5956 11940 6012 11996
rect 6012 11940 6016 11996
rect 5952 11936 6016 11940
rect 6032 11996 6096 12000
rect 6032 11940 6036 11996
rect 6036 11940 6092 11996
rect 6092 11940 6096 11996
rect 6032 11936 6096 11940
rect 6112 11996 6176 12000
rect 6112 11940 6116 11996
rect 6116 11940 6172 11996
rect 6172 11940 6176 11996
rect 6112 11936 6176 11940
rect 6192 11996 6256 12000
rect 6192 11940 6196 11996
rect 6196 11940 6252 11996
rect 6252 11940 6256 11996
rect 6192 11936 6256 11940
rect 15952 11996 16016 12000
rect 15952 11940 15956 11996
rect 15956 11940 16012 11996
rect 16012 11940 16016 11996
rect 15952 11936 16016 11940
rect 16032 11996 16096 12000
rect 16032 11940 16036 11996
rect 16036 11940 16092 11996
rect 16092 11940 16096 11996
rect 16032 11936 16096 11940
rect 16112 11996 16176 12000
rect 16112 11940 16116 11996
rect 16116 11940 16172 11996
rect 16172 11940 16176 11996
rect 16112 11936 16176 11940
rect 16192 11996 16256 12000
rect 16192 11940 16196 11996
rect 16196 11940 16252 11996
rect 16252 11940 16256 11996
rect 16192 11936 16256 11940
rect 6500 11868 6564 11932
rect 12756 11868 12820 11932
rect 25952 11996 26016 12000
rect 25952 11940 25956 11996
rect 25956 11940 26012 11996
rect 26012 11940 26016 11996
rect 25952 11936 26016 11940
rect 26032 11996 26096 12000
rect 26032 11940 26036 11996
rect 26036 11940 26092 11996
rect 26092 11940 26096 11996
rect 26032 11936 26096 11940
rect 26112 11996 26176 12000
rect 26112 11940 26116 11996
rect 26116 11940 26172 11996
rect 26172 11940 26176 11996
rect 26112 11936 26176 11940
rect 26192 11996 26256 12000
rect 26192 11940 26196 11996
rect 26196 11940 26252 11996
rect 26252 11940 26256 11996
rect 26192 11936 26256 11940
rect 10952 11452 11016 11456
rect 10952 11396 10956 11452
rect 10956 11396 11012 11452
rect 11012 11396 11016 11452
rect 10952 11392 11016 11396
rect 11032 11452 11096 11456
rect 11032 11396 11036 11452
rect 11036 11396 11092 11452
rect 11092 11396 11096 11452
rect 11032 11392 11096 11396
rect 11112 11452 11176 11456
rect 11112 11396 11116 11452
rect 11116 11396 11172 11452
rect 11172 11396 11176 11452
rect 11112 11392 11176 11396
rect 11192 11452 11256 11456
rect 11192 11396 11196 11452
rect 11196 11396 11252 11452
rect 11252 11396 11256 11452
rect 11192 11392 11256 11396
rect 20952 11452 21016 11456
rect 20952 11396 20956 11452
rect 20956 11396 21012 11452
rect 21012 11396 21016 11452
rect 20952 11392 21016 11396
rect 21032 11452 21096 11456
rect 21032 11396 21036 11452
rect 21036 11396 21092 11452
rect 21092 11396 21096 11452
rect 21032 11392 21096 11396
rect 21112 11452 21176 11456
rect 21112 11396 21116 11452
rect 21116 11396 21172 11452
rect 21172 11396 21176 11452
rect 21112 11392 21176 11396
rect 21192 11452 21256 11456
rect 21192 11396 21196 11452
rect 21196 11396 21252 11452
rect 21252 11396 21256 11452
rect 21192 11392 21256 11396
rect 5952 10908 6016 10912
rect 5952 10852 5956 10908
rect 5956 10852 6012 10908
rect 6012 10852 6016 10908
rect 5952 10848 6016 10852
rect 6032 10908 6096 10912
rect 6032 10852 6036 10908
rect 6036 10852 6092 10908
rect 6092 10852 6096 10908
rect 6032 10848 6096 10852
rect 6112 10908 6176 10912
rect 6112 10852 6116 10908
rect 6116 10852 6172 10908
rect 6172 10852 6176 10908
rect 6112 10848 6176 10852
rect 6192 10908 6256 10912
rect 6192 10852 6196 10908
rect 6196 10852 6252 10908
rect 6252 10852 6256 10908
rect 6192 10848 6256 10852
rect 15952 10908 16016 10912
rect 15952 10852 15956 10908
rect 15956 10852 16012 10908
rect 16012 10852 16016 10908
rect 15952 10848 16016 10852
rect 16032 10908 16096 10912
rect 16032 10852 16036 10908
rect 16036 10852 16092 10908
rect 16092 10852 16096 10908
rect 16032 10848 16096 10852
rect 16112 10908 16176 10912
rect 16112 10852 16116 10908
rect 16116 10852 16172 10908
rect 16172 10852 16176 10908
rect 16112 10848 16176 10852
rect 16192 10908 16256 10912
rect 16192 10852 16196 10908
rect 16196 10852 16252 10908
rect 16252 10852 16256 10908
rect 16192 10848 16256 10852
rect 25952 10908 26016 10912
rect 25952 10852 25956 10908
rect 25956 10852 26012 10908
rect 26012 10852 26016 10908
rect 25952 10848 26016 10852
rect 26032 10908 26096 10912
rect 26032 10852 26036 10908
rect 26036 10852 26092 10908
rect 26092 10852 26096 10908
rect 26032 10848 26096 10852
rect 26112 10908 26176 10912
rect 26112 10852 26116 10908
rect 26116 10852 26172 10908
rect 26172 10852 26176 10908
rect 26112 10848 26176 10852
rect 26192 10908 26256 10912
rect 26192 10852 26196 10908
rect 26196 10852 26252 10908
rect 26252 10852 26256 10908
rect 26192 10848 26256 10852
rect 10952 10364 11016 10368
rect 10952 10308 10956 10364
rect 10956 10308 11012 10364
rect 11012 10308 11016 10364
rect 10952 10304 11016 10308
rect 11032 10364 11096 10368
rect 11032 10308 11036 10364
rect 11036 10308 11092 10364
rect 11092 10308 11096 10364
rect 11032 10304 11096 10308
rect 11112 10364 11176 10368
rect 11112 10308 11116 10364
rect 11116 10308 11172 10364
rect 11172 10308 11176 10364
rect 11112 10304 11176 10308
rect 11192 10364 11256 10368
rect 11192 10308 11196 10364
rect 11196 10308 11252 10364
rect 11252 10308 11256 10364
rect 11192 10304 11256 10308
rect 20952 10364 21016 10368
rect 20952 10308 20956 10364
rect 20956 10308 21012 10364
rect 21012 10308 21016 10364
rect 20952 10304 21016 10308
rect 21032 10364 21096 10368
rect 21032 10308 21036 10364
rect 21036 10308 21092 10364
rect 21092 10308 21096 10364
rect 21032 10304 21096 10308
rect 21112 10364 21176 10368
rect 21112 10308 21116 10364
rect 21116 10308 21172 10364
rect 21172 10308 21176 10364
rect 21112 10304 21176 10308
rect 21192 10364 21256 10368
rect 21192 10308 21196 10364
rect 21196 10308 21252 10364
rect 21252 10308 21256 10364
rect 21192 10304 21256 10308
rect 5952 9820 6016 9824
rect 5952 9764 5956 9820
rect 5956 9764 6012 9820
rect 6012 9764 6016 9820
rect 5952 9760 6016 9764
rect 6032 9820 6096 9824
rect 6032 9764 6036 9820
rect 6036 9764 6092 9820
rect 6092 9764 6096 9820
rect 6032 9760 6096 9764
rect 6112 9820 6176 9824
rect 6112 9764 6116 9820
rect 6116 9764 6172 9820
rect 6172 9764 6176 9820
rect 6112 9760 6176 9764
rect 6192 9820 6256 9824
rect 6192 9764 6196 9820
rect 6196 9764 6252 9820
rect 6252 9764 6256 9820
rect 6192 9760 6256 9764
rect 15952 9820 16016 9824
rect 15952 9764 15956 9820
rect 15956 9764 16012 9820
rect 16012 9764 16016 9820
rect 15952 9760 16016 9764
rect 16032 9820 16096 9824
rect 16032 9764 16036 9820
rect 16036 9764 16092 9820
rect 16092 9764 16096 9820
rect 16032 9760 16096 9764
rect 16112 9820 16176 9824
rect 16112 9764 16116 9820
rect 16116 9764 16172 9820
rect 16172 9764 16176 9820
rect 16112 9760 16176 9764
rect 16192 9820 16256 9824
rect 16192 9764 16196 9820
rect 16196 9764 16252 9820
rect 16252 9764 16256 9820
rect 16192 9760 16256 9764
rect 25952 9820 26016 9824
rect 25952 9764 25956 9820
rect 25956 9764 26012 9820
rect 26012 9764 26016 9820
rect 25952 9760 26016 9764
rect 26032 9820 26096 9824
rect 26032 9764 26036 9820
rect 26036 9764 26092 9820
rect 26092 9764 26096 9820
rect 26032 9760 26096 9764
rect 26112 9820 26176 9824
rect 26112 9764 26116 9820
rect 26116 9764 26172 9820
rect 26172 9764 26176 9820
rect 26112 9760 26176 9764
rect 26192 9820 26256 9824
rect 26192 9764 26196 9820
rect 26196 9764 26252 9820
rect 26252 9764 26256 9820
rect 26192 9760 26256 9764
rect 10952 9276 11016 9280
rect 10952 9220 10956 9276
rect 10956 9220 11012 9276
rect 11012 9220 11016 9276
rect 10952 9216 11016 9220
rect 11032 9276 11096 9280
rect 11032 9220 11036 9276
rect 11036 9220 11092 9276
rect 11092 9220 11096 9276
rect 11032 9216 11096 9220
rect 11112 9276 11176 9280
rect 11112 9220 11116 9276
rect 11116 9220 11172 9276
rect 11172 9220 11176 9276
rect 11112 9216 11176 9220
rect 11192 9276 11256 9280
rect 11192 9220 11196 9276
rect 11196 9220 11252 9276
rect 11252 9220 11256 9276
rect 11192 9216 11256 9220
rect 20952 9276 21016 9280
rect 20952 9220 20956 9276
rect 20956 9220 21012 9276
rect 21012 9220 21016 9276
rect 20952 9216 21016 9220
rect 21032 9276 21096 9280
rect 21032 9220 21036 9276
rect 21036 9220 21092 9276
rect 21092 9220 21096 9276
rect 21032 9216 21096 9220
rect 21112 9276 21176 9280
rect 21112 9220 21116 9276
rect 21116 9220 21172 9276
rect 21172 9220 21176 9276
rect 21112 9216 21176 9220
rect 21192 9276 21256 9280
rect 21192 9220 21196 9276
rect 21196 9220 21252 9276
rect 21252 9220 21256 9276
rect 21192 9216 21256 9220
rect 5952 8732 6016 8736
rect 5952 8676 5956 8732
rect 5956 8676 6012 8732
rect 6012 8676 6016 8732
rect 5952 8672 6016 8676
rect 6032 8732 6096 8736
rect 6032 8676 6036 8732
rect 6036 8676 6092 8732
rect 6092 8676 6096 8732
rect 6032 8672 6096 8676
rect 6112 8732 6176 8736
rect 6112 8676 6116 8732
rect 6116 8676 6172 8732
rect 6172 8676 6176 8732
rect 6112 8672 6176 8676
rect 6192 8732 6256 8736
rect 6192 8676 6196 8732
rect 6196 8676 6252 8732
rect 6252 8676 6256 8732
rect 6192 8672 6256 8676
rect 15952 8732 16016 8736
rect 15952 8676 15956 8732
rect 15956 8676 16012 8732
rect 16012 8676 16016 8732
rect 15952 8672 16016 8676
rect 16032 8732 16096 8736
rect 16032 8676 16036 8732
rect 16036 8676 16092 8732
rect 16092 8676 16096 8732
rect 16032 8672 16096 8676
rect 16112 8732 16176 8736
rect 16112 8676 16116 8732
rect 16116 8676 16172 8732
rect 16172 8676 16176 8732
rect 16112 8672 16176 8676
rect 16192 8732 16256 8736
rect 16192 8676 16196 8732
rect 16196 8676 16252 8732
rect 16252 8676 16256 8732
rect 16192 8672 16256 8676
rect 25952 8732 26016 8736
rect 25952 8676 25956 8732
rect 25956 8676 26012 8732
rect 26012 8676 26016 8732
rect 25952 8672 26016 8676
rect 26032 8732 26096 8736
rect 26032 8676 26036 8732
rect 26036 8676 26092 8732
rect 26092 8676 26096 8732
rect 26032 8672 26096 8676
rect 26112 8732 26176 8736
rect 26112 8676 26116 8732
rect 26116 8676 26172 8732
rect 26172 8676 26176 8732
rect 26112 8672 26176 8676
rect 26192 8732 26256 8736
rect 26192 8676 26196 8732
rect 26196 8676 26252 8732
rect 26252 8676 26256 8732
rect 26192 8672 26256 8676
rect 10952 8188 11016 8192
rect 10952 8132 10956 8188
rect 10956 8132 11012 8188
rect 11012 8132 11016 8188
rect 10952 8128 11016 8132
rect 11032 8188 11096 8192
rect 11032 8132 11036 8188
rect 11036 8132 11092 8188
rect 11092 8132 11096 8188
rect 11032 8128 11096 8132
rect 11112 8188 11176 8192
rect 11112 8132 11116 8188
rect 11116 8132 11172 8188
rect 11172 8132 11176 8188
rect 11112 8128 11176 8132
rect 11192 8188 11256 8192
rect 11192 8132 11196 8188
rect 11196 8132 11252 8188
rect 11252 8132 11256 8188
rect 11192 8128 11256 8132
rect 20952 8188 21016 8192
rect 20952 8132 20956 8188
rect 20956 8132 21012 8188
rect 21012 8132 21016 8188
rect 20952 8128 21016 8132
rect 21032 8188 21096 8192
rect 21032 8132 21036 8188
rect 21036 8132 21092 8188
rect 21092 8132 21096 8188
rect 21032 8128 21096 8132
rect 21112 8188 21176 8192
rect 21112 8132 21116 8188
rect 21116 8132 21172 8188
rect 21172 8132 21176 8188
rect 21112 8128 21176 8132
rect 21192 8188 21256 8192
rect 21192 8132 21196 8188
rect 21196 8132 21252 8188
rect 21252 8132 21256 8188
rect 21192 8128 21256 8132
rect 5952 7644 6016 7648
rect 5952 7588 5956 7644
rect 5956 7588 6012 7644
rect 6012 7588 6016 7644
rect 5952 7584 6016 7588
rect 6032 7644 6096 7648
rect 6032 7588 6036 7644
rect 6036 7588 6092 7644
rect 6092 7588 6096 7644
rect 6032 7584 6096 7588
rect 6112 7644 6176 7648
rect 6112 7588 6116 7644
rect 6116 7588 6172 7644
rect 6172 7588 6176 7644
rect 6112 7584 6176 7588
rect 6192 7644 6256 7648
rect 6192 7588 6196 7644
rect 6196 7588 6252 7644
rect 6252 7588 6256 7644
rect 6192 7584 6256 7588
rect 15952 7644 16016 7648
rect 15952 7588 15956 7644
rect 15956 7588 16012 7644
rect 16012 7588 16016 7644
rect 15952 7584 16016 7588
rect 16032 7644 16096 7648
rect 16032 7588 16036 7644
rect 16036 7588 16092 7644
rect 16092 7588 16096 7644
rect 16032 7584 16096 7588
rect 16112 7644 16176 7648
rect 16112 7588 16116 7644
rect 16116 7588 16172 7644
rect 16172 7588 16176 7644
rect 16112 7584 16176 7588
rect 16192 7644 16256 7648
rect 16192 7588 16196 7644
rect 16196 7588 16252 7644
rect 16252 7588 16256 7644
rect 16192 7584 16256 7588
rect 25952 7644 26016 7648
rect 25952 7588 25956 7644
rect 25956 7588 26012 7644
rect 26012 7588 26016 7644
rect 25952 7584 26016 7588
rect 26032 7644 26096 7648
rect 26032 7588 26036 7644
rect 26036 7588 26092 7644
rect 26092 7588 26096 7644
rect 26032 7584 26096 7588
rect 26112 7644 26176 7648
rect 26112 7588 26116 7644
rect 26116 7588 26172 7644
rect 26172 7588 26176 7644
rect 26112 7584 26176 7588
rect 26192 7644 26256 7648
rect 26192 7588 26196 7644
rect 26196 7588 26252 7644
rect 26252 7588 26256 7644
rect 26192 7584 26256 7588
rect 10952 7100 11016 7104
rect 10952 7044 10956 7100
rect 10956 7044 11012 7100
rect 11012 7044 11016 7100
rect 10952 7040 11016 7044
rect 11032 7100 11096 7104
rect 11032 7044 11036 7100
rect 11036 7044 11092 7100
rect 11092 7044 11096 7100
rect 11032 7040 11096 7044
rect 11112 7100 11176 7104
rect 11112 7044 11116 7100
rect 11116 7044 11172 7100
rect 11172 7044 11176 7100
rect 11112 7040 11176 7044
rect 11192 7100 11256 7104
rect 11192 7044 11196 7100
rect 11196 7044 11252 7100
rect 11252 7044 11256 7100
rect 11192 7040 11256 7044
rect 20952 7100 21016 7104
rect 20952 7044 20956 7100
rect 20956 7044 21012 7100
rect 21012 7044 21016 7100
rect 20952 7040 21016 7044
rect 21032 7100 21096 7104
rect 21032 7044 21036 7100
rect 21036 7044 21092 7100
rect 21092 7044 21096 7100
rect 21032 7040 21096 7044
rect 21112 7100 21176 7104
rect 21112 7044 21116 7100
rect 21116 7044 21172 7100
rect 21172 7044 21176 7100
rect 21112 7040 21176 7044
rect 21192 7100 21256 7104
rect 21192 7044 21196 7100
rect 21196 7044 21252 7100
rect 21252 7044 21256 7100
rect 21192 7040 21256 7044
rect 5952 6556 6016 6560
rect 5952 6500 5956 6556
rect 5956 6500 6012 6556
rect 6012 6500 6016 6556
rect 5952 6496 6016 6500
rect 6032 6556 6096 6560
rect 6032 6500 6036 6556
rect 6036 6500 6092 6556
rect 6092 6500 6096 6556
rect 6032 6496 6096 6500
rect 6112 6556 6176 6560
rect 6112 6500 6116 6556
rect 6116 6500 6172 6556
rect 6172 6500 6176 6556
rect 6112 6496 6176 6500
rect 6192 6556 6256 6560
rect 6192 6500 6196 6556
rect 6196 6500 6252 6556
rect 6252 6500 6256 6556
rect 6192 6496 6256 6500
rect 15952 6556 16016 6560
rect 15952 6500 15956 6556
rect 15956 6500 16012 6556
rect 16012 6500 16016 6556
rect 15952 6496 16016 6500
rect 16032 6556 16096 6560
rect 16032 6500 16036 6556
rect 16036 6500 16092 6556
rect 16092 6500 16096 6556
rect 16032 6496 16096 6500
rect 16112 6556 16176 6560
rect 16112 6500 16116 6556
rect 16116 6500 16172 6556
rect 16172 6500 16176 6556
rect 16112 6496 16176 6500
rect 16192 6556 16256 6560
rect 16192 6500 16196 6556
rect 16196 6500 16252 6556
rect 16252 6500 16256 6556
rect 16192 6496 16256 6500
rect 25952 6556 26016 6560
rect 25952 6500 25956 6556
rect 25956 6500 26012 6556
rect 26012 6500 26016 6556
rect 25952 6496 26016 6500
rect 26032 6556 26096 6560
rect 26032 6500 26036 6556
rect 26036 6500 26092 6556
rect 26092 6500 26096 6556
rect 26032 6496 26096 6500
rect 26112 6556 26176 6560
rect 26112 6500 26116 6556
rect 26116 6500 26172 6556
rect 26172 6500 26176 6556
rect 26112 6496 26176 6500
rect 26192 6556 26256 6560
rect 26192 6500 26196 6556
rect 26196 6500 26252 6556
rect 26252 6500 26256 6556
rect 26192 6496 26256 6500
rect 10952 6012 11016 6016
rect 10952 5956 10956 6012
rect 10956 5956 11012 6012
rect 11012 5956 11016 6012
rect 10952 5952 11016 5956
rect 11032 6012 11096 6016
rect 11032 5956 11036 6012
rect 11036 5956 11092 6012
rect 11092 5956 11096 6012
rect 11032 5952 11096 5956
rect 11112 6012 11176 6016
rect 11112 5956 11116 6012
rect 11116 5956 11172 6012
rect 11172 5956 11176 6012
rect 11112 5952 11176 5956
rect 11192 6012 11256 6016
rect 11192 5956 11196 6012
rect 11196 5956 11252 6012
rect 11252 5956 11256 6012
rect 11192 5952 11256 5956
rect 20952 6012 21016 6016
rect 20952 5956 20956 6012
rect 20956 5956 21012 6012
rect 21012 5956 21016 6012
rect 20952 5952 21016 5956
rect 21032 6012 21096 6016
rect 21032 5956 21036 6012
rect 21036 5956 21092 6012
rect 21092 5956 21096 6012
rect 21032 5952 21096 5956
rect 21112 6012 21176 6016
rect 21112 5956 21116 6012
rect 21116 5956 21172 6012
rect 21172 5956 21176 6012
rect 21112 5952 21176 5956
rect 21192 6012 21256 6016
rect 21192 5956 21196 6012
rect 21196 5956 21252 6012
rect 21252 5956 21256 6012
rect 21192 5952 21256 5956
rect 5952 5468 6016 5472
rect 5952 5412 5956 5468
rect 5956 5412 6012 5468
rect 6012 5412 6016 5468
rect 5952 5408 6016 5412
rect 6032 5468 6096 5472
rect 6032 5412 6036 5468
rect 6036 5412 6092 5468
rect 6092 5412 6096 5468
rect 6032 5408 6096 5412
rect 6112 5468 6176 5472
rect 6112 5412 6116 5468
rect 6116 5412 6172 5468
rect 6172 5412 6176 5468
rect 6112 5408 6176 5412
rect 6192 5468 6256 5472
rect 6192 5412 6196 5468
rect 6196 5412 6252 5468
rect 6252 5412 6256 5468
rect 6192 5408 6256 5412
rect 15952 5468 16016 5472
rect 15952 5412 15956 5468
rect 15956 5412 16012 5468
rect 16012 5412 16016 5468
rect 15952 5408 16016 5412
rect 16032 5468 16096 5472
rect 16032 5412 16036 5468
rect 16036 5412 16092 5468
rect 16092 5412 16096 5468
rect 16032 5408 16096 5412
rect 16112 5468 16176 5472
rect 16112 5412 16116 5468
rect 16116 5412 16172 5468
rect 16172 5412 16176 5468
rect 16112 5408 16176 5412
rect 16192 5468 16256 5472
rect 16192 5412 16196 5468
rect 16196 5412 16252 5468
rect 16252 5412 16256 5468
rect 16192 5408 16256 5412
rect 25952 5468 26016 5472
rect 25952 5412 25956 5468
rect 25956 5412 26012 5468
rect 26012 5412 26016 5468
rect 25952 5408 26016 5412
rect 26032 5468 26096 5472
rect 26032 5412 26036 5468
rect 26036 5412 26092 5468
rect 26092 5412 26096 5468
rect 26032 5408 26096 5412
rect 26112 5468 26176 5472
rect 26112 5412 26116 5468
rect 26116 5412 26172 5468
rect 26172 5412 26176 5468
rect 26112 5408 26176 5412
rect 26192 5468 26256 5472
rect 26192 5412 26196 5468
rect 26196 5412 26252 5468
rect 26252 5412 26256 5468
rect 26192 5408 26256 5412
rect 10952 4924 11016 4928
rect 10952 4868 10956 4924
rect 10956 4868 11012 4924
rect 11012 4868 11016 4924
rect 10952 4864 11016 4868
rect 11032 4924 11096 4928
rect 11032 4868 11036 4924
rect 11036 4868 11092 4924
rect 11092 4868 11096 4924
rect 11032 4864 11096 4868
rect 11112 4924 11176 4928
rect 11112 4868 11116 4924
rect 11116 4868 11172 4924
rect 11172 4868 11176 4924
rect 11112 4864 11176 4868
rect 11192 4924 11256 4928
rect 11192 4868 11196 4924
rect 11196 4868 11252 4924
rect 11252 4868 11256 4924
rect 11192 4864 11256 4868
rect 20952 4924 21016 4928
rect 20952 4868 20956 4924
rect 20956 4868 21012 4924
rect 21012 4868 21016 4924
rect 20952 4864 21016 4868
rect 21032 4924 21096 4928
rect 21032 4868 21036 4924
rect 21036 4868 21092 4924
rect 21092 4868 21096 4924
rect 21032 4864 21096 4868
rect 21112 4924 21176 4928
rect 21112 4868 21116 4924
rect 21116 4868 21172 4924
rect 21172 4868 21176 4924
rect 21112 4864 21176 4868
rect 21192 4924 21256 4928
rect 21192 4868 21196 4924
rect 21196 4868 21252 4924
rect 21252 4868 21256 4924
rect 21192 4864 21256 4868
rect 5952 4380 6016 4384
rect 5952 4324 5956 4380
rect 5956 4324 6012 4380
rect 6012 4324 6016 4380
rect 5952 4320 6016 4324
rect 6032 4380 6096 4384
rect 6032 4324 6036 4380
rect 6036 4324 6092 4380
rect 6092 4324 6096 4380
rect 6032 4320 6096 4324
rect 6112 4380 6176 4384
rect 6112 4324 6116 4380
rect 6116 4324 6172 4380
rect 6172 4324 6176 4380
rect 6112 4320 6176 4324
rect 6192 4380 6256 4384
rect 6192 4324 6196 4380
rect 6196 4324 6252 4380
rect 6252 4324 6256 4380
rect 6192 4320 6256 4324
rect 15952 4380 16016 4384
rect 15952 4324 15956 4380
rect 15956 4324 16012 4380
rect 16012 4324 16016 4380
rect 15952 4320 16016 4324
rect 16032 4380 16096 4384
rect 16032 4324 16036 4380
rect 16036 4324 16092 4380
rect 16092 4324 16096 4380
rect 16032 4320 16096 4324
rect 16112 4380 16176 4384
rect 16112 4324 16116 4380
rect 16116 4324 16172 4380
rect 16172 4324 16176 4380
rect 16112 4320 16176 4324
rect 16192 4380 16256 4384
rect 16192 4324 16196 4380
rect 16196 4324 16252 4380
rect 16252 4324 16256 4380
rect 16192 4320 16256 4324
rect 25952 4380 26016 4384
rect 25952 4324 25956 4380
rect 25956 4324 26012 4380
rect 26012 4324 26016 4380
rect 25952 4320 26016 4324
rect 26032 4380 26096 4384
rect 26032 4324 26036 4380
rect 26036 4324 26092 4380
rect 26092 4324 26096 4380
rect 26032 4320 26096 4324
rect 26112 4380 26176 4384
rect 26112 4324 26116 4380
rect 26116 4324 26172 4380
rect 26172 4324 26176 4380
rect 26112 4320 26176 4324
rect 26192 4380 26256 4384
rect 26192 4324 26196 4380
rect 26196 4324 26252 4380
rect 26252 4324 26256 4380
rect 26192 4320 26256 4324
rect 10952 3836 11016 3840
rect 10952 3780 10956 3836
rect 10956 3780 11012 3836
rect 11012 3780 11016 3836
rect 10952 3776 11016 3780
rect 11032 3836 11096 3840
rect 11032 3780 11036 3836
rect 11036 3780 11092 3836
rect 11092 3780 11096 3836
rect 11032 3776 11096 3780
rect 11112 3836 11176 3840
rect 11112 3780 11116 3836
rect 11116 3780 11172 3836
rect 11172 3780 11176 3836
rect 11112 3776 11176 3780
rect 11192 3836 11256 3840
rect 11192 3780 11196 3836
rect 11196 3780 11252 3836
rect 11252 3780 11256 3836
rect 11192 3776 11256 3780
rect 20952 3836 21016 3840
rect 20952 3780 20956 3836
rect 20956 3780 21012 3836
rect 21012 3780 21016 3836
rect 20952 3776 21016 3780
rect 21032 3836 21096 3840
rect 21032 3780 21036 3836
rect 21036 3780 21092 3836
rect 21092 3780 21096 3836
rect 21032 3776 21096 3780
rect 21112 3836 21176 3840
rect 21112 3780 21116 3836
rect 21116 3780 21172 3836
rect 21172 3780 21176 3836
rect 21112 3776 21176 3780
rect 21192 3836 21256 3840
rect 21192 3780 21196 3836
rect 21196 3780 21252 3836
rect 21252 3780 21256 3836
rect 21192 3776 21256 3780
rect 5952 3292 6016 3296
rect 5952 3236 5956 3292
rect 5956 3236 6012 3292
rect 6012 3236 6016 3292
rect 5952 3232 6016 3236
rect 6032 3292 6096 3296
rect 6032 3236 6036 3292
rect 6036 3236 6092 3292
rect 6092 3236 6096 3292
rect 6032 3232 6096 3236
rect 6112 3292 6176 3296
rect 6112 3236 6116 3292
rect 6116 3236 6172 3292
rect 6172 3236 6176 3292
rect 6112 3232 6176 3236
rect 6192 3292 6256 3296
rect 6192 3236 6196 3292
rect 6196 3236 6252 3292
rect 6252 3236 6256 3292
rect 6192 3232 6256 3236
rect 15952 3292 16016 3296
rect 15952 3236 15956 3292
rect 15956 3236 16012 3292
rect 16012 3236 16016 3292
rect 15952 3232 16016 3236
rect 16032 3292 16096 3296
rect 16032 3236 16036 3292
rect 16036 3236 16092 3292
rect 16092 3236 16096 3292
rect 16032 3232 16096 3236
rect 16112 3292 16176 3296
rect 16112 3236 16116 3292
rect 16116 3236 16172 3292
rect 16172 3236 16176 3292
rect 16112 3232 16176 3236
rect 16192 3292 16256 3296
rect 16192 3236 16196 3292
rect 16196 3236 16252 3292
rect 16252 3236 16256 3292
rect 16192 3232 16256 3236
rect 25952 3292 26016 3296
rect 25952 3236 25956 3292
rect 25956 3236 26012 3292
rect 26012 3236 26016 3292
rect 25952 3232 26016 3236
rect 26032 3292 26096 3296
rect 26032 3236 26036 3292
rect 26036 3236 26092 3292
rect 26092 3236 26096 3292
rect 26032 3232 26096 3236
rect 26112 3292 26176 3296
rect 26112 3236 26116 3292
rect 26116 3236 26172 3292
rect 26172 3236 26176 3292
rect 26112 3232 26176 3236
rect 26192 3292 26256 3296
rect 26192 3236 26196 3292
rect 26196 3236 26252 3292
rect 26252 3236 26256 3292
rect 26192 3232 26256 3236
rect 10952 2748 11016 2752
rect 10952 2692 10956 2748
rect 10956 2692 11012 2748
rect 11012 2692 11016 2748
rect 10952 2688 11016 2692
rect 11032 2748 11096 2752
rect 11032 2692 11036 2748
rect 11036 2692 11092 2748
rect 11092 2692 11096 2748
rect 11032 2688 11096 2692
rect 11112 2748 11176 2752
rect 11112 2692 11116 2748
rect 11116 2692 11172 2748
rect 11172 2692 11176 2748
rect 11112 2688 11176 2692
rect 11192 2748 11256 2752
rect 11192 2692 11196 2748
rect 11196 2692 11252 2748
rect 11252 2692 11256 2748
rect 11192 2688 11256 2692
rect 20952 2748 21016 2752
rect 20952 2692 20956 2748
rect 20956 2692 21012 2748
rect 21012 2692 21016 2748
rect 20952 2688 21016 2692
rect 21032 2748 21096 2752
rect 21032 2692 21036 2748
rect 21036 2692 21092 2748
rect 21092 2692 21096 2748
rect 21032 2688 21096 2692
rect 21112 2748 21176 2752
rect 21112 2692 21116 2748
rect 21116 2692 21172 2748
rect 21172 2692 21176 2748
rect 21112 2688 21176 2692
rect 21192 2748 21256 2752
rect 21192 2692 21196 2748
rect 21196 2692 21252 2748
rect 21252 2692 21256 2748
rect 21192 2688 21256 2692
rect 5952 2204 6016 2208
rect 5952 2148 5956 2204
rect 5956 2148 6012 2204
rect 6012 2148 6016 2204
rect 5952 2144 6016 2148
rect 6032 2204 6096 2208
rect 6032 2148 6036 2204
rect 6036 2148 6092 2204
rect 6092 2148 6096 2204
rect 6032 2144 6096 2148
rect 6112 2204 6176 2208
rect 6112 2148 6116 2204
rect 6116 2148 6172 2204
rect 6172 2148 6176 2204
rect 6112 2144 6176 2148
rect 6192 2204 6256 2208
rect 6192 2148 6196 2204
rect 6196 2148 6252 2204
rect 6252 2148 6256 2204
rect 6192 2144 6256 2148
rect 15952 2204 16016 2208
rect 15952 2148 15956 2204
rect 15956 2148 16012 2204
rect 16012 2148 16016 2204
rect 15952 2144 16016 2148
rect 16032 2204 16096 2208
rect 16032 2148 16036 2204
rect 16036 2148 16092 2204
rect 16092 2148 16096 2204
rect 16032 2144 16096 2148
rect 16112 2204 16176 2208
rect 16112 2148 16116 2204
rect 16116 2148 16172 2204
rect 16172 2148 16176 2204
rect 16112 2144 16176 2148
rect 16192 2204 16256 2208
rect 16192 2148 16196 2204
rect 16196 2148 16252 2204
rect 16252 2148 16256 2204
rect 16192 2144 16256 2148
rect 25952 2204 26016 2208
rect 25952 2148 25956 2204
rect 25956 2148 26012 2204
rect 26012 2148 26016 2204
rect 25952 2144 26016 2148
rect 26032 2204 26096 2208
rect 26032 2148 26036 2204
rect 26036 2148 26092 2204
rect 26092 2148 26096 2204
rect 26032 2144 26096 2148
rect 26112 2204 26176 2208
rect 26112 2148 26116 2204
rect 26116 2148 26172 2204
rect 26172 2148 26176 2204
rect 26112 2144 26176 2148
rect 26192 2204 26256 2208
rect 26192 2148 26196 2204
rect 26196 2148 26252 2204
rect 26252 2148 26256 2204
rect 26192 2144 26256 2148
<< metal4 >>
rect 5944 21792 6264 21808
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 20704 6264 21728
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 19616 6264 20640
rect 10944 21248 11264 21808
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 20160 11264 21184
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 9627 19684 9693 19685
rect 9627 19620 9628 19684
rect 9692 19620 9693 19684
rect 9627 19619 9693 19620
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 18528 6264 19552
rect 9630 19413 9690 19619
rect 9627 19412 9693 19413
rect 9627 19348 9628 19412
rect 9692 19348 9693 19412
rect 9627 19347 9693 19348
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 17440 6264 18464
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 16352 6264 17376
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 15264 6264 16288
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 14176 6264 15200
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 13088 6264 14112
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 12000 6264 13024
rect 10944 19072 11264 20096
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 17984 11264 19008
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 16896 11264 17920
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 15808 11264 16832
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 14720 11264 15744
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 13632 11264 14656
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 12544 11264 13568
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 10912 6264 11936
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 9824 6264 10848
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 8736 6264 9760
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 7648 6264 8672
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 6560 6264 7584
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 5472 6264 6496
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 4384 6264 5408
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 3296 6264 4320
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 2208 6264 3232
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2128 6264 2144
rect 10944 11456 11264 12480
rect 15944 21792 16264 21808
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 20704 16264 21728
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 19616 16264 20640
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 18528 16264 19552
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 17440 16264 18464
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 16352 16264 17376
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 15264 16264 16288
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 14176 16264 15200
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 13088 16264 14112
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 12000 16264 13024
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 10368 11264 11392
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 9280 11264 10304
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 8192 11264 9216
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 7104 11264 8128
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 6016 11264 7040
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 4928 11264 5952
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 3840 11264 4864
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 2752 11264 3776
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2128 11264 2688
rect 15944 10912 16264 11936
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 9824 16264 10848
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 8736 16264 9760
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 7648 16264 8672
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 6560 16264 7584
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 5472 16264 6496
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 4384 16264 5408
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 3296 16264 4320
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 2208 16264 3232
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2128 16264 2144
rect 20944 21248 21264 21808
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 20944 20160 21264 21184
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 19072 21264 20096
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 17984 21264 19008
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 16896 21264 17920
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 15808 21264 16832
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 20944 14720 21264 15744
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 13632 21264 14656
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 12544 21264 13568
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 11456 21264 12480
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 10368 21264 11392
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 20944 9280 21264 10304
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 20944 8192 21264 9216
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 7104 21264 8128
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 6016 21264 7040
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 4928 21264 5952
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 3840 21264 4864
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 20944 2752 21264 3776
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2128 21264 2688
rect 25944 21792 26264 21808
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 20704 26264 21728
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 19616 26264 20640
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 18528 26264 19552
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 17440 26264 18464
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 16352 26264 17376
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 15264 26264 16288
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 25944 14176 26264 15200
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 13088 26264 14112
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 12000 26264 13024
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 10912 26264 11936
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 9824 26264 10848
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 25944 8736 26264 9760
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 7648 26264 8672
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 6560 26264 7584
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 5472 26264 6496
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 4384 26264 5408
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 25944 3296 26264 4320
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 25944 2208 26264 3232
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2128 26264 2144
<< via4 >>
rect 6414 11932 6650 12018
rect 6414 11868 6500 11932
rect 6500 11868 6564 11932
rect 6564 11868 6650 11932
rect 6414 11782 6650 11868
rect 12670 11932 12906 12018
rect 12670 11868 12756 11932
rect 12756 11868 12820 11932
rect 12820 11868 12906 11932
rect 12670 11782 12906 11868
<< metal5 >>
rect 6372 12018 12948 12060
rect 6372 11782 6414 12018
rect 6650 11782 12670 12018
rect 12906 11782 12948 12018
rect 6372 11740 12948 11782
use scs8hd_buf_2  _49_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__49__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_11
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_72 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_23
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_35
timestamp 1586364061
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_47
timestamp 1586364061
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7176 0 -1 2720
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_85 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_118 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _69_
timestamp 1586364061
transform 1 0 26404 0 1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_6  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__69__A
timestamp 1586364061
transform 1 0 26956 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_280
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_292
timestamp 1586364061
transform 1 0 27968 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_279
timestamp 1586364061
transform 1 0 26772 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_283
timestamp 1586364061
transform 1 0 27140 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_295
timestamp 1586364061
transform 1 0 28244 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 28888 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 28888 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_298 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 28520 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_288
timestamp 1586364061
transform 1 0 27600 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_296
timestamp 1586364061
transform 1 0 28336 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 28888 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_281
timestamp 1586364061
transform 1 0 26956 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_3_293
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 590 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 28888 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_288
timestamp 1586364061
transform 1 0 27600 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_296
timestamp 1586364061
transform 1 0 28336 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 28888 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 1564 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_19
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_31
timestamp 1586364061
transform 1 0 3956 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_43
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_5_55
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _65_
timestamp 1586364061
transform 1 0 26404 0 1 4896
box -38 -48 406 592
use scs8hd_decap_6  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__65__A
timestamp 1586364061
transform 1 0 26956 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_279
timestamp 1586364061
transform 1 0 26772 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_283
timestamp 1586364061
transform 1 0 27140 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_5_295
timestamp 1586364061
transform 1 0 28244 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 28888 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_7
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 1932 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _51_
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use scs8hd_buf_2  _41_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_19
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_11
timestamp 1586364061
transform 1 0 2116 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _52_
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_17
timestamp 1586364061
transform 1 0 2668 0 -1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_29
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_23
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_35
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_47
timestamp 1586364061
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_157
timestamp 1586364061
transform 1 0 15548 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_169
timestamp 1586364061
transform 1 0 16652 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_181
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__63__A
timestamp 1586364061
transform 1 0 26496 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_275
timestamp 1586364061
transform 1 0 26404 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_288
timestamp 1586364061
transform 1 0 27600 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_296
timestamp 1586364061
transform 1 0 28336 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_278
timestamp 1586364061
transform 1 0 26680 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_290
timestamp 1586364061
transform 1 0 27784 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 28888 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 28888 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_298
timestamp 1586364061
transform 1 0 28520 0 1 5984
box -38 -48 130 592
use scs8hd_buf_2  _39_
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 406 592
use scs8hd_buf_2  _43_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 2300 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_11
timestamp 1586364061
transform 1 0 2116 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_19
timestamp 1586364061
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 3036 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_36
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_48
timestamp 1586364061
transform 1 0 5520 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_59
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_65
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_77
timestamp 1586364061
transform 1 0 8188 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_89
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_1  mux_top_ipin_0.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15364 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_158
timestamp 1586364061
transform 1 0 15640 0 -1 7072
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_168
timestamp 1586364061
transform 1 0 16560 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_172
timestamp 1586364061
transform 1 0 16928 0 -1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_184
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_8_196
timestamp 1586364061
transform 1 0 19136 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_200
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_204
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_212
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _63_
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_280
timestamp 1586364061
transform 1 0 26864 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_8_292
timestamp 1586364061
transform 1 0 27968 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 28888 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_298
timestamp 1586364061
transform 1 0 28520 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  _42_
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 406 592
use scs8hd_buf_2  _44_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_11
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_19
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _37_
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 406 592
use scs8hd_buf_2  _53_
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 5244 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_43
timestamp 1586364061
transform 1 0 5060 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_47
timestamp 1586364061
transform 1 0 5428 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l1_in_1_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6900 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_72
timestamp 1586364061
transform 1 0 7728 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_76
timestamp 1586364061
transform 1 0 8096 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_88
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_100
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_112
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_120
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use scs8hd_mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_162
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_194
timestamp 1586364061
transform 1 0 18952 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_190
timestamp 1586364061
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18768 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 19320 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 20332 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_207
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_211
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_223
timestamp 1586364061
transform 1 0 21620 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_235
timestamp 1586364061
transform 1 0 22724 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_243
timestamp 1586364061
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _71_
timestamp 1586364061
transform 1 0 26404 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__71__A
timestamp 1586364061
transform 1 0 26220 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 406 592
use scs8hd_buf_2  _62_
timestamp 1586364061
transform 1 0 27508 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__73__A
timestamp 1586364061
transform 1 0 26956 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__62__A
timestamp 1586364061
transform 1 0 28060 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_279
timestamp 1586364061
transform 1 0 26772 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_283
timestamp 1586364061
transform 1 0 27140 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_291
timestamp 1586364061
transform 1 0 27876 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_295
timestamp 1586364061
transform 1 0 28244 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 28888 0 1 7072
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l4_in_0_
timestamp 1586364061
transform 1 0 1932 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_18
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_22
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_26
timestamp 1586364061
transform 1 0 3496 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6164 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_10_53
timestamp 1586364061
transform 1 0 5980 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_66
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_70
timestamp 1586364061
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_74
timestamp 1586364061
transform 1 0 7912 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_78
timestamp 1586364061
transform 1 0 8280 0 -1 8160
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_81
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_89
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_top_ipin_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 16744 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_162
timestamp 1586364061
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_165
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_169
timestamp 1586364061
transform 1 0 16652 0 -1 8160
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_189
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_193
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21160 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 20240 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_210
timestamp 1586364061
transform 1 0 20424 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_3  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 21528 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_220
timestamp 1586364061
transform 1 0 21344 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_224
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_228
timestamp 1586364061
transform 1 0 22080 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_240
timestamp 1586364061
transform 1 0 23184 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_252
timestamp 1586364061
transform 1 0 24288 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_2  _73_
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_264
timestamp 1586364061
transform 1 0 25392 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_272
timestamp 1586364061
transform 1 0 26128 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_280
timestamp 1586364061
transform 1 0 26864 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_10_292
timestamp 1586364061
transform 1 0 27968 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 28888 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_298
timestamp 1586364061
transform 1 0 28520 0 -1 8160
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l3_in_1_
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_16
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_20
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_24
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_38
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _50_
timestamp 1586364061
transform 1 0 5336 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_42
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_50
timestamp 1586364061
transform 1 0 5704 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_54
timestamp 1586364061
transform 1 0 6072 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_58
timestamp 1586364061
transform 1 0 6440 0 1 8160
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_75
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_88
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_92
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_104
timestamp 1586364061
transform 1 0 10672 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_11_116
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_11_155
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_158
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_162
timestamp 1586364061
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_199
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_210
timestamp 1586364061
transform 1 0 20424 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_214
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_227
timestamp 1586364061
transform 1 0 21988 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_231
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_243
timestamp 1586364061
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 406 592
use scs8hd_buf_2  _60_
timestamp 1586364061
transform 1 0 25300 0 1 8160
box -38 -48 406 592
use scs8hd_buf_2  _61_
timestamp 1586364061
transform 1 0 26404 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__60__A
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__59__A
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_267
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_271
timestamp 1586364061
transform 1 0 26036 0 1 8160
box -38 -48 406 592
use scs8hd_buf_2  _57_
timestamp 1586364061
transform 1 0 27508 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__61__A
timestamp 1586364061
transform 1 0 26956 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__57__A
timestamp 1586364061
transform 1 0 28060 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__66__A
timestamp 1586364061
transform 1 0 27324 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_279
timestamp 1586364061
transform 1 0 26772 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_283
timestamp 1586364061
transform 1 0 27140 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_291
timestamp 1586364061
transform 1 0 27876 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_295
timestamp 1586364061
transform 1 0 28244 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 28888 0 1 8160
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l2_in_3_
timestamp 1586364061
transform 1 0 1932 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_18
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4692 0 -1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3128 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_24
timestamp 1586364061
transform 1 0 3312 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_28
timestamp 1586364061
transform 1 0 3680 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_58
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7176 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_62
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_65
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_75
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_81
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_89
timestamp 1586364061
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_conb_1  _20_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15456 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_ipin_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_159
timestamp 1586364061
transform 1 0 15732 0 -1 9248
box -38 -48 590 592
use scs8hd_mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 19228 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 18676 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_193
timestamp 1586364061
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_11.mux_l2_in_2_
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_236
timestamp 1586364061
transform 1 0 22816 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_248
timestamp 1586364061
transform 1 0 23920 0 -1 9248
box -38 -48 1142 592
use scs8hd_buf_2  _59_
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 406 592
use scs8hd_buf_2  _66_
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_260
timestamp 1586364061
transform 1 0 25024 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_267
timestamp 1586364061
transform 1 0 25668 0 -1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 27048 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_280
timestamp 1586364061
transform 1 0 26864 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_284
timestamp 1586364061
transform 1 0 27232 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_12_296
timestamp 1586364061
transform 1 0 28336 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 28888 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l2_in_2_
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 866 592
use scs8hd_conb_1  _21_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_18
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_14
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 5060 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_41
timestamp 1586364061
transform 1 0 4876 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_2  _38_
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_45
timestamp 1586364061
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_45
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_14_58
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6900 0 1 9248
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_64
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_75
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_79
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_87
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_83
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_82
timestamp 1586364061
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_14_91
timestamp 1586364061
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 10212 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 10580 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_101
timestamp 1586364061
transform 1 0 10396 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_155
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_158
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_168
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_164
timestamp 1586364061
transform 1 0 16192 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_162
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16008 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 16652 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17664 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_182
timestamp 1586364061
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_186
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_194
timestamp 1586364061
transform 1 0 18952 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_194
timestamp 1586364061
transform 1 0 18952 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_190
timestamp 1586364061
transform 1 0 18584 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 19044 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 18768 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_11.mux_l2_in_1_
timestamp 1586364061
transform 1 0 19228 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_ipin_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19320 0 1 9248
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_ipin_11.mux_l2_in_3_
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_206
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_210
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 21988 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 23000 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_221
timestamp 1586364061
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_225
timestamp 1586364061
transform 1 0 21804 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_229
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_236
timestamp 1586364061
transform 1 0 22816 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_243
timestamp 1586364061
transform 1 0 23460 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_13_241
timestamp 1586364061
transform 1 0 23276 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 23644 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_conb_1  _28_
timestamp 1586364061
transform 1 0 23184 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_255
timestamp 1586364061
transform 1 0 24564 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_247
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_255
timestamp 1586364061
transform 1 0 24564 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 24012 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__56__A
timestamp 1586364061
transform 1 0 24012 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _58_
timestamp 1586364061
transform 1 0 24196 0 1 9248
box -38 -48 406 592
use scs8hd_buf_2  _56_
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__58__A
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_267
timestamp 1586364061
transform 1 0 25668 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_267
timestamp 1586364061
transform 1 0 25668 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_259
timestamp 1586364061
transform 1 0 24932 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__68__A
timestamp 1586364061
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _68_
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 406 592
use scs8hd_buf_2  _55_
timestamp 1586364061
transform 1 0 25300 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_271
timestamp 1586364061
transform 1 0 26036 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__72__A
timestamp 1586364061
transform 1 0 26220 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_14.mux_l2_in_2_
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 866 592
use scs8hd_buf_2  _72_
timestamp 1586364061
transform 1 0 26404 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_283
timestamp 1586364061
transform 1 0 27140 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_279
timestamp 1586364061
transform 1 0 26772 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 27324 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 26956 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _64_
timestamp 1586364061
transform 1 0 27508 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_297
timestamp 1586364061
transform 1 0 28428 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_295
timestamp 1586364061
transform 1 0 28244 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_291
timestamp 1586364061
transform 1 0 27876 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__A
timestamp 1586364061
transform 1 0 28060 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_285
timestamp 1586364061
transform 1 0 27324 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 28888 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 28888 0 -1 10336
box -38 -48 314 592
use scs8hd_buf_2  _46_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2668 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_13
timestamp 1586364061
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_26
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_30
timestamp 1586364061
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _48_
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_83
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_87
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_91
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_95
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_108
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_112
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12604 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_127
timestamp 1586364061
transform 1 0 12788 0 1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_139
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_15_151
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_157
timestamp 1586364061
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_10.mux_l2_in_1_
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_161
timestamp 1586364061
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_165
timestamp 1586364061
transform 1 0 16284 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_11.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_ipin_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_199
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 21712 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 22080 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_222
timestamp 1586364061
transform 1 0 21528 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_226
timestamp 1586364061
transform 1 0 21896 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_230
timestamp 1586364061
transform 1 0 22264 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_234
timestamp 1586364061
transform 1 0 22632 0 1 10336
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_15.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_14.mux_l2_in_3_
timestamp 1586364061
transform 1 0 26404 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 26220 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__70__A
timestamp 1586364061
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_264
timestamp 1586364061
transform 1 0 25392 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_268
timestamp 1586364061
transform 1 0 25760 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_272
timestamp 1586364061
transform 1 0 26128 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 27416 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 27784 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 28152 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_284
timestamp 1586364061
transform 1 0 27232 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_288
timestamp 1586364061
transform 1 0 27600 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_292
timestamp 1586364061
transform 1 0 27968 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_296
timestamp 1586364061
transform 1 0 28336 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 28888 0 1 10336
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_11
timestamp 1586364061
transform 1 0 2116 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_2  _36_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4600 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_36
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4968 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_40
timestamp 1586364061
transform 1 0 4784 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_66
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_70
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 8924 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_83
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_87
timestamp 1586364061
transform 1 0 9108 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_91
timestamp 1586364061
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 11776 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_108
timestamp 1586364061
transform 1 0 11040 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_112
timestamp 1586364061
transform 1 0 11408 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_137
timestamp 1586364061
transform 1 0 13708 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 15548 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_149
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_10.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 15916 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_159
timestamp 1586364061
transform 1 0 15732 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_172
timestamp 1586364061
transform 1 0 16928 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_176
timestamp 1586364061
transform 1 0 17296 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_11.mux_l2_in_0_
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_ipin_11.mux_l3_in_1_
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_189
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_193
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_11.mux_l4_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use scs8hd_conb_1  _24_
timestamp 1586364061
transform 1 0 22448 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_228
timestamp 1586364061
transform 1 0 22080 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_6  FILLER_16_235
timestamp 1586364061
transform 1 0 22724 0 -1 11424
box -38 -48 590 592
use scs8hd_mux2_1  mux_bottom_ipin_15.mux_l3_in_1_
timestamp 1586364061
transform 1 0 23552 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 23368 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 24564 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_241
timestamp 1586364061
transform 1 0 23276 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_253
timestamp 1586364061
transform 1 0 24380 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_257
timestamp 1586364061
transform 1 0 24748 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  _70_
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_15.mux_l2_in_0_
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 26220 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 24932 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_261
timestamp 1586364061
transform 1 0 25116 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_267
timestamp 1586364061
transform 1 0 25668 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_285
timestamp 1586364061
transform 1 0 27324 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_16_297
timestamp 1586364061
transform 1 0 28428 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 28888 0 -1 11424
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 1786 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__35__A
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_30
timestamp 1586364061
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_34
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_40
timestamp 1586364061
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l3_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l4_in_0_
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_88
timestamp 1586364061
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_92
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_106
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_17_155
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_10.mux_l3_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_163
timestamp 1586364061
transform 1 0 16100 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_11.mux_l3_in_0_
timestamp 1586364061
transform 1 0 18400 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_11.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_201
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _54_
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21896 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_224
timestamp 1586364061
transform 1 0 21712 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_228
timestamp 1586364061
transform 1 0 22080 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_236
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_15.mux_l4_in_0_
timestamp 1586364061
transform 1 0 24012 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 23828 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_15.mux_l3_in_0_
timestamp 1586364061
transform 1 0 25576 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 26588 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 25392 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_258
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_262
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_275
timestamp 1586364061
transform 1 0 26404 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _67_
timestamp 1586364061
transform 1 0 27140 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__67__A
timestamp 1586364061
transform 1 0 27692 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 26956 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 28060 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_279
timestamp 1586364061
transform 1 0 26772 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_287
timestamp 1586364061
transform 1 0 27508 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_291
timestamp 1586364061
transform 1 0 27876 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_295
timestamp 1586364061
transform 1 0 28244 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 28888 0 1 11424
box -38 -48 314 592
use scs8hd_conb_1  _22_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _35_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_36
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 6532 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_40
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_46
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l2_in_3_
timestamp 1586364061
transform 1 0 7084 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 6900 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 8096 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_61
timestamp 1586364061
transform 1 0 6716 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_74
timestamp 1586364061
transform 1 0 7912 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_78
timestamp 1586364061
transform 1 0 8280 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_82
timestamp 1586364061
transform 1 0 8648 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_85
timestamp 1586364061
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_89
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_97
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 10212 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10580 0 -1 12512
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_18_101
timestamp 1586364061
transform 1 0 10396 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_122
timestamp 1586364061
transform 1 0 12328 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_126
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_134
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_138
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_10.mux_l2_in_2_
timestamp 1586364061
transform 1 0 15548 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_142
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_148
timestamp 1586364061
transform 1 0 14720 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_151
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_11.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 17112 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 16560 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 16928 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_170
timestamp 1586364061
transform 1 0 16744 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_193
timestamp 1586364061
transform 1 0 18860 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_203
timestamp 1586364061
transform 1 0 19780 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_199
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 19596 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_207
timestamp 1586364061
transform 1 0 20148 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 19964 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_211
timestamp 1586364061
transform 1 0 20516 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21160 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21436 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 22724 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_220
timestamp 1586364061
transform 1 0 21344 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_230
timestamp 1586364061
transform 1 0 22264 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_234
timestamp 1586364061
transform 1 0 22632 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_237
timestamp 1586364061
transform 1 0 22908 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_15.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 23368 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_241
timestamp 1586364061
transform 1 0 23276 0 -1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_15.mux_l2_in_1_
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 26128 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 25668 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_261
timestamp 1586364061
transform 1 0 25116 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_265
timestamp 1586364061
transform 1 0 25484 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_269
timestamp 1586364061
transform 1 0 25852 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_274
timestamp 1586364061
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_285
timestamp 1586364061
transform 1 0 27324 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_18_297
timestamp 1586364061
transform 1 0 28428 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 28888 0 -1 12512
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_1.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 1472 0 -1 13600
box -38 -48 1786 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_29
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_25
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_38
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_34
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_46
timestamp 1586364061
transform 1 0 5336 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_42
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_buf_2  _34_
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_20_57
timestamp 1586364061
transform 1 0 6348 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_53
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__34__A
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_64
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_61
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l2_in_2_
timestamp 1586364061
transform 1 0 7084 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_19_78
timestamp 1586364061
transform 1 0 8280 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 8096 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_4.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_107
timestamp 1586364061
transform 1 0 10948 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_107
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_102
timestamp 1586364061
transform 1 0 10488 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11132 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_111
timestamp 1586364061
transform 1 0 11316 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l2_in_2_
timestamp 1586364061
transform 1 0 11500 0 -1 13600
box -38 -48 866 592
use scs8hd_conb_1  _32_
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_126
timestamp 1586364061
transform 1 0 12696 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_122
timestamp 1586364061
transform 1 0 12328 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_130
timestamp 1586364061
transform 1 0 13064 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_138
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_10.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_146
timestamp 1586364061
transform 1 0 14536 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_142
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_158
timestamp 1586364061
transform 1 0 15640 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_152
timestamp 1586364061
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_158
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 14904 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_10.mux_l2_in_3_
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_162
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 15916 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_10.mux_l3_in_1_
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_10.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 16468 0 -1 13600
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_20_186
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18400 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_194
timestamp 1586364061
transform 1 0 18952 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l1_in_1_
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_11.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_207
timestamp 1586364061
transform 1 0 20148 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_203
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 19964 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_210
timestamp 1586364061
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_212
timestamp 1586364061
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_11.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 20976 0 1 12512
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l1_in_2_
timestamp 1586364061
transform 1 0 22724 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 22908 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 22172 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 22540 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_235
timestamp 1586364061
transform 1 0 22724 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_231
timestamp 1586364061
transform 1 0 22356 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_244
timestamp 1586364061
transform 1 0 23552 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_239
timestamp 1586364061
transform 1 0 23092 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 23736 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_15.mux_l2_in_2_
timestamp 1586364061
transform 1 0 23736 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_248
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_255
timestamp 1586364061
transform 1 0 24564 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 24104 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_15.mux_l2_in_3_
timestamp 1586364061
transform 1 0 24288 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_265
timestamp 1586364061
transform 1 0 25484 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_261
timestamp 1586364061
transform 1 0 25116 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_263
timestamp 1586364061
transform 1 0 25300 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_259
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 25576 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_274
timestamp 1586364061
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_270
timestamp 1586364061
transform 1 0 25944 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_268
timestamp 1586364061
transform 1 0 25760 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 26128 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 25760 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 25944 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_15.mux_l1_in_0_
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_15.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 26128 0 1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 28060 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 27508 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_291
timestamp 1586364061
transform 1 0 27876 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_295
timestamp 1586364061
transform 1 0 28244 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_285
timestamp 1586364061
transform 1 0 27324 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_289
timestamp 1586364061
transform 1 0 27692 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_297
timestamp 1586364061
transform 1 0 28428 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 28888 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 28888 0 -1 13600
box -38 -48 314 592
use scs8hd_buf_2  _45_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 1786 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_11
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__47__A
timestamp 1586364061
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_35
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_75
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_79
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l3_in_1_
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_83
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_97
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l2_in_3_
timestamp 1586364061
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_101
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l1_in_1_
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_142
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_146
timestamp 1586364061
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use scs8hd_conb_1  _23_
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_163
timestamp 1586364061
transform 1 0 16100 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_168
timestamp 1586364061
transform 1 0 16560 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_10.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_12.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 21068 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 19964 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_203
timestamp 1586364061
transform 1 0 19780 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_207
timestamp 1586364061
transform 1 0 20148 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_213
timestamp 1586364061
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_14.mux_l3_in_1_
timestamp 1586364061
transform 1 0 24196 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 23920 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_21_250
timestamp 1586364061
transform 1 0 24104 0 1 13600
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_15.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 25760 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 25576 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 25208 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_260
timestamp 1586364061
transform 1 0 25024 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_264
timestamp 1586364061
transform 1 0 25392 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 27692 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 28060 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_287
timestamp 1586364061
transform 1 0 27508 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_291
timestamp 1586364061
transform 1 0 27876 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_295
timestamp 1586364061
transform 1 0 28244 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 28888 0 1 13600
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_2.mux_l2_in_2_
timestamp 1586364061
transform 1 0 1932 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_18
timestamp 1586364061
transform 1 0 2760 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_2  _47_
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3496 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 2944 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4600 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_22
timestamp 1586364061
transform 1 0 3128 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  FILLER_22_28
timestamp 1586364061
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_36
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 5428 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_40
timestamp 1586364061
transform 1 0 4784 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_46
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_6.mux_l3_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_66
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_70
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 10212 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_97
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_6.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_101
timestamp 1586364061
transform 1 0 10396 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_107
timestamp 1586364061
transform 1 0 10948 0 -1 14688
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 13340 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_127
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_131
timestamp 1586364061
transform 1 0 13156 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_135
timestamp 1586364061
transform 1 0 13524 0 -1 14688
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 14904 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_152
timestamp 1586364061
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_10.mux_l4_in_0_
timestamp 1586364061
transform 1 0 17112 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16652 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_167
timestamp 1586364061
transform 1 0 16468 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_171
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_14.mux_l3_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 18492 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 18124 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 18860 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_183
timestamp 1586364061
transform 1 0 17940 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_187
timestamp 1586364061
transform 1 0 18308 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_191
timestamp 1586364061
transform 1 0 18676 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_195
timestamp 1586364061
transform 1 0 19044 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 21068 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_210
timestamp 1586364061
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_12.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 21436 0 -1 14688
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_22_219
timestamp 1586364061
transform 1 0 21252 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_14.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 23920 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 23368 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 23736 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_240
timestamp 1586364061
transform 1 0 23184 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_244
timestamp 1586364061
transform 1 0 23552 0 -1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_14.mux_l4_in_0_
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 26220 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 25852 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_267
timestamp 1586364061
transform 1 0 25668 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_271
timestamp 1586364061
transform 1 0 26036 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 27508 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_285
timestamp 1586364061
transform 1 0 27324 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_289
timestamp 1586364061
transform 1 0 27692 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_297
timestamp 1586364061
transform 1 0 28428 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 28888 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_2.mux_l2_in_3_
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_18
timestamp 1586364061
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_22
timestamp 1586364061
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_35
timestamp 1586364061
transform 1 0 4324 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _31_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_6.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 7268 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_65
timestamp 1586364061
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_69
timestamp 1586364061
transform 1 0 7452 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_5.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 9384 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 8832 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_82
timestamp 1586364061
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_109
timestamp 1586364061
transform 1 0 11132 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l1_in_2_
timestamp 1586364061
transform 1 0 12880 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 12696 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_137
timestamp 1586364061
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_141
timestamp 1586364061
transform 1 0 14076 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_154
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_158
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17020 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_14.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18492 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_198
timestamp 1586364061
transform 1 0 19320 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l2_in_1_
timestamp 1586364061
transform 1 0 20056 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 19872 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 21068 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 19504 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_202
timestamp 1586364061
transform 1 0 19688 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_215
timestamp 1586364061
transform 1 0 20884 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l2_in_3_
timestamp 1586364061
transform 1 0 21620 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_219
timestamp 1586364061
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_238
timestamp 1586364061
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_14.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 24288 0 1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 24104 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_242
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_249
timestamp 1586364061
transform 1 0 24012 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 26496 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_271
timestamp 1586364061
transform 1 0 26036 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_275
timestamp 1586364061
transform 1 0 26404 0 1 14688
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_14.mux_l2_in_0_
timestamp 1586364061
transform 1 0 26772 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 27784 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 28152 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_278
timestamp 1586364061
transform 1 0 26680 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_288
timestamp 1586364061
transform 1 0 27600 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_292
timestamp 1586364061
transform 1 0 27968 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_296
timestamp 1586364061
transform 1 0 28336 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 28888 0 1 14688
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 1472 0 -1 15776
box -38 -48 1786 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5704 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5520 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_41
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_46
timestamp 1586364061
transform 1 0 5336 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 8188 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_69
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_75
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_79
timestamp 1586364061
transform 1 0 8372 0 -1 15776
box -38 -48 222 592
use scs8hd_conb_1  _33_
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l4_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_6.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11776 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11408 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_24_107
timestamp 1586364061
transform 1 0 10948 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_111
timestamp 1586364061
transform 1 0 11316 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_114
timestamp 1586364061
transform 1 0 11592 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 13708 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_135
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_139
timestamp 1586364061
transform 1 0 13892 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_6  FILLER_24_147
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 17204 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_173
timestamp 1586364061
transform 1 0 17020 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_177
timestamp 1586364061
transform 1 0 17388 0 -1 15776
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_10.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18216 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 17664 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_182
timestamp 1586364061
transform 1 0 17848 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l3_in_0_
timestamp 1586364061
transform 1 0 21068 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 20148 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_205
timestamp 1586364061
transform 1 0 19964 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_209
timestamp 1586364061
transform 1 0 20332 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 22080 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_226
timestamp 1586364061
transform 1 0 21896 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_230
timestamp 1586364061
transform 1 0 22264 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_238
timestamp 1586364061
transform 1 0 23000 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23184 0 -1 15776
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l1_in_1_
timestamp 1586364061
transform 1 0 24748 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 24564 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_249
timestamp 1586364061
transform 1 0 24012 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_253
timestamp 1586364061
transform 1 0 24380 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_14.mux_l1_in_0_
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 26128 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 25760 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_266
timestamp 1586364061
transform 1 0 25576 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_270
timestamp 1586364061
transform 1 0 25944 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_274
timestamp 1586364061
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 27508 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_285
timestamp 1586364061
transform 1 0 27324 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_289
timestamp 1586364061
transform 1 0 27692 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_297
timestamp 1586364061
transform 1 0 28428 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 28888 0 -1 15776
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 1564 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_16
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 3312 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_20
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 5336 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_43
timestamp 1586364061
transform 1 0 5060 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_48
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_52
timestamp 1586364061
transform 1 0 5888 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_56
timestamp 1586364061
transform 1 0 6256 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_69
timestamp 1586364061
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_66
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_60
timestamp 1586364061
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_73
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_6.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_96
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_6.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_100
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_7.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_136
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 16100 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 16468 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_161
timestamp 1586364061
transform 1 0 15916 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_165
timestamp 1586364061
transform 1 0 16284 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_169
timestamp 1586364061
transform 1 0 16652 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_173
timestamp 1586364061
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_177
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_10.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 19964 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 20700 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_203
timestamp 1586364061
transform 1 0 19780 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_207
timestamp 1586364061
transform 1 0 20148 0 1 15776
box -38 -48 590 592
use scs8hd_fill_2  FILLER_25_215
timestamp 1586364061
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l3_in_1_
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 22356 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 22724 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_219
timestamp 1586364061
transform 1 0 21252 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_229
timestamp 1586364061
transform 1 0 22172 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_233
timestamp 1586364061
transform 1 0 22540 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_237
timestamp 1586364061
transform 1 0 22908 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l2_in_0_
timestamp 1586364061
transform 1 0 24564 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 23092 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 24012 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_241
timestamp 1586364061
transform 1 0 23276 0 1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_251
timestamp 1586364061
transform 1 0 24196 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_14.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 26128 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 25944 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_264
timestamp 1586364061
transform 1 0 25392 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_268
timestamp 1586364061
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 28060 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_291
timestamp 1586364061
transform 1 0 27876 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_295
timestamp 1586364061
transform 1 0 28244 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 28888 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_2.mux_l3_in_1_
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_2.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_27_26
timestamp 1586364061
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_26
timestamp 1586364061
transform 1 0 3496 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 3680 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3312 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_30
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_39
timestamp 1586364061
transform 1 0 4692 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_35
timestamp 1586364061
transform 1 0 4324 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_30
timestamp 1586364061
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 4508 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_conb_1  _29_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 5336 0 -1 16864
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 4968 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_66
timestamp 1586364061
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_65
timestamp 1586364061
transform 1 0 7084 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 6992 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_70
timestamp 1586364061
transform 1 0 7544 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_71
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 7728 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 8096 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_6.mux_l2_in_2_
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_6.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 8280 0 1 16864
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_ipin_6.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_97
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_101
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_107
timestamp 1586364061
transform 1 0 10948 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_6.mux_l3_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_111
timestamp 1586364061
transform 1 0 11316 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_7.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11408 0 -1 16864
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_7.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_138
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_26_138
timestamp 1586364061
transform 1 0 13800 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_135
timestamp 1586364061
transform 1 0 13524 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_131
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_143
timestamp 1586364061
transform 1 0 14260 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_144
timestamp 1586364061
transform 1 0 14352 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 14444 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use scs8hd_conb_1  _18_
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_150
timestamp 1586364061
transform 1 0 14904 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 14812 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l2_in_2_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_8.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 14996 0 1 16864
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l3_in_1_
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16928 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 16652 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_167
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_170
timestamp 1586364061
transform 1 0 16744 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_174
timestamp 1586364061
transform 1 0 17112 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_186
timestamp 1586364061
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_180
timestamp 1586364061
transform 1 0 17664 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18400 0 -1 16864
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18308 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_197
timestamp 1586364061
transform 1 0 19228 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19320 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_204
timestamp 1586364061
transform 1 0 19872 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_200
timestamp 1586364061
transform 1 0 19504 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_205
timestamp 1586364061
transform 1 0 19964 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19688 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 20148 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_213
timestamp 1586364061
transform 1 0 20700 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_209
timestamp 1586364061
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_210
timestamp 1586364061
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 20516 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_12.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 21068 0 1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_12.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 21068 0 -1 16864
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23000 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_236
timestamp 1586364061
transform 1 0 22816 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_236
timestamp 1586364061
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_247
timestamp 1586364061
transform 1 0 23828 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_240
timestamp 1586364061
transform 1 0 23184 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23368 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_conb_1  _25_
timestamp 1586364061
transform 1 0 23552 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_257
timestamp 1586364061
transform 1 0 24748 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 24564 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 24012 0 -1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_13.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_27_264
timestamp 1586364061
transform 1 0 25392 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_267
timestamp 1586364061
transform 1 0 25668 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 25576 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l2_in_1_
timestamp 1586364061
transform 1 0 24840 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_268
timestamp 1586364061
transform 1 0 25760 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_274
timestamp 1586364061
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_271
timestamp 1586364061
transform 1 0 26036 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 26128 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 25944 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l1_in_2_
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_14.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 26128 0 1 16864
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 28060 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_285
timestamp 1586364061
transform 1 0 27324 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_26_297
timestamp 1586364061
transform 1 0 28428 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_291
timestamp 1586364061
transform 1 0 27876 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_295
timestamp 1586364061
transform 1 0 28244 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 28888 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 28888 0 1 16864
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_2.mux_l4_in_0_
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 2760 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_16
timestamp 1586364061
transform 1 0 2576 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 4692 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 3312 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_20
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_4  FILLER_28_26
timestamp 1586364061
transform 1 0 3496 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_30
timestamp 1586364061
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_36
timestamp 1586364061
transform 1 0 4416 0 -1 17952
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4968 0 -1 17952
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_28_41
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_6.mux_l4_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6900 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_61
timestamp 1586364061
transform 1 0 6716 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_65
timestamp 1586364061
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_69
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_73
timestamp 1586364061
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_7.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11592 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 11960 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_112
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_116
timestamp 1586364061
transform 1 0 11776 0 -1 17952
box -38 -48 222 592
use scs8hd_conb_1  _17_
timestamp 1586364061
transform 1 0 12144 0 -1 17952
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l4_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_123
timestamp 1586364061
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_127
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_131
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_135
timestamp 1586364061
transform 1 0 13524 0 -1 17952
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_6  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_bottom_ipin_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15824 0 -1 17952
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18308 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18124 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_179
timestamp 1586364061
transform 1 0 17572 0 -1 17952
box -38 -48 590 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l4_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_210
timestamp 1586364061
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_13.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 22448 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 21896 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_224
timestamp 1586364061
transform 1 0 21712 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_228
timestamp 1586364061
transform 1 0 22080 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 24472 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_256
timestamp 1586364061
transform 1 0 24656 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_267
timestamp 1586364061
transform 1 0 25668 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_260
timestamp 1586364061
transform 1 0 25024 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25208 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 24840 0 -1 17952
box -38 -48 222 592
use scs8hd_conb_1  _26_
timestamp 1586364061
transform 1 0 25392 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_274
timestamp 1586364061
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_271
timestamp 1586364061
transform 1 0 26036 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 26128 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l2_in_3_
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 27508 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_285
timestamp 1586364061
transform 1 0 27324 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_289
timestamp 1586364061
transform 1 0 27692 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_297
timestamp 1586364061
transform 1 0 28428 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 28888 0 -1 17952
box -38 -48 314 592
use scs8hd_buf_2  _40_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_11
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_19
timestamp 1586364061
transform 1 0 2852 0 1 17952
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_3.mux_l2_in_3_
timestamp 1586364061
transform 1 0 3312 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_33
timestamp 1586364061
transform 1 0 4140 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_37
timestamp 1586364061
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4876 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5888 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_50
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_54
timestamp 1586364061
transform 1 0 6072 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_58
timestamp 1586364061
transform 1 0 6440 0 1 17952
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_75
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_6.mux_l2_in_3_
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_89
timestamp 1586364061
transform 1 0 9292 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_93
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_96
timestamp 1586364061
transform 1 0 9936 0 1 17952
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_7.mux_l2_in_2_
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_101
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_7.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 16468 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_161
timestamp 1586364061
transform 1 0 15916 0 1 17952
box -38 -48 590 592
use scs8hd_fill_2  FILLER_29_169
timestamp 1586364061
transform 1 0 16652 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_173
timestamp 1586364061
transform 1 0 17020 0 1 17952
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_197
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l2_in_3_
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_210
timestamp 1586364061
transform 1 0 20424 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_214
timestamp 1586364061
transform 1 0 20792 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_217
timestamp 1586364061
transform 1 0 21068 0 1 17952
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l2_in_2_
timestamp 1586364061
transform 1 0 21528 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 22540 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22908 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_231
timestamp 1586364061
transform 1 0 22356 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_235
timestamp 1586364061
transform 1 0 22724 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_13.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 24472 0 1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 24288 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 23920 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_239
timestamp 1586364061
transform 1 0 23092 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_243
timestamp 1586364061
transform 1 0 23460 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_250
timestamp 1586364061
transform 1 0 24104 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 26496 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_273
timestamp 1586364061
transform 1 0 26220 0 1 17952
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l3_in_0_
timestamp 1586364061
transform 1 0 26956 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 27968 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_278
timestamp 1586364061
transform 1 0 26680 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_290
timestamp 1586364061
transform 1 0 27784 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_294
timestamp 1586364061
transform 1 0 28152 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 28888 0 1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_29_298
timestamp 1586364061
transform 1 0 28520 0 1 17952
box -38 -48 130 592
use scs8hd_buf_1  mux_bottom_ipin_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2208 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2668 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_3  FILLER_30_9
timestamp 1586364061
transform 1 0 1932 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_19
timestamp 1586364061
transform 1 0 2852 0 -1 19040
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_3.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 4692 0 -1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 3312 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 4508 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_30_26
timestamp 1586364061
transform 1 0 3496 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_36
timestamp 1586364061
transform 1 0 4416 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_58
timestamp 1586364061
transform 1 0 6440 0 -1 19040
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 7176 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_64
timestamp 1586364061
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_75
timestamp 1586364061
transform 1 0 8004 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_79
timestamp 1586364061
transform 1 0 8372 0 -1 19040
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_7.mux_l3_in_1_
timestamp 1586364061
transform 1 0 9752 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_82
timestamp 1586364061
transform 1 0 8648 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_86
timestamp 1586364061
transform 1 0 9016 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_7.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11316 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_103
timestamp 1586364061
transform 1 0 10580 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_107
timestamp 1586364061
transform 1 0 10948 0 -1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 13248 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_130
timestamp 1586364061
transform 1 0 13064 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_134
timestamp 1586364061
transform 1 0 13432 0 -1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_144
timestamp 1586364061
transform 1 0 14352 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_150
timestamp 1586364061
transform 1 0 14904 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_bottom_ipin_9.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 16468 0 -1 19040
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l2_in_2_
timestamp 1586364061
transform 1 0 18952 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 18768 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 18400 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_186
timestamp 1586364061
transform 1 0 18216 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l1_in_2_
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 19964 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 20332 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_203
timestamp 1586364061
transform 1 0 19780 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_207
timestamp 1586364061
transform 1 0 20148 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_211
timestamp 1586364061
transform 1 0 20516 0 -1 19040
box -38 -48 314 592
use scs8hd_buf_1  mux_bottom_ipin_12.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22448 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 21896 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_224
timestamp 1586364061
transform 1 0 21712 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_228
timestamp 1586364061
transform 1 0 22080 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_235
timestamp 1586364061
transform 1 0 22724 0 -1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 24656 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_247
timestamp 1586364061
transform 1 0 23828 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_255
timestamp 1586364061
transform 1 0 24564 0 -1 19040
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l3_in_1_
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l4_in_0_
timestamp 1586364061
transform 1 0 24840 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 26220 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 25852 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_267
timestamp 1586364061
transform 1 0 25668 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_271
timestamp 1586364061
transform 1 0 26036 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 27508 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_285
timestamp 1586364061
transform 1 0 27324 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_289
timestamp 1586364061
transform 1 0 27692 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_297
timestamp 1586364061
transform 1 0 28428 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 28888 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_3.mux_l4_in_0_
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_21
timestamp 1586364061
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_34
timestamp 1586364061
transform 1 0 4232 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_38
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_55
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _30_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_65
timestamp 1586364061
transform 1 0 7084 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_31_77
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 590 592
use scs8hd_buf_1  mux_bottom_ipin_6.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 8832 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 9292 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_83
timestamp 1586364061
transform 1 0 8740 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_87
timestamp 1586364061
transform 1 0 9108 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_91
timestamp 1586364061
transform 1 0 9476 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_96
timestamp 1586364061
transform 1 0 9936 0 1 19040
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_7.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 11868 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_101
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_119
timestamp 1586364061
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_7.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 12512 0 1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l2_in_3_
timestamp 1586364061
transform 1 0 14996 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 14812 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_143
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 16468 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_160
timestamp 1586364061
transform 1 0 15824 0 1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_31_166
timestamp 1586364061
transform 1 0 16376 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_169
timestamp 1586364061
transform 1 0 16652 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_173
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_177
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 406 592
use scs8hd_conb_1  _19_
timestamp 1586364061
transform 1 0 18492 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 19320 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 18952 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 18308 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_192
timestamp 1586364061
transform 1 0 18768 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 19504 0 1 19040
box -38 -48 1786 592
use scs8hd_decap_12  FILLER_31_219
timestamp 1586364061
transform 1 0 21252 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_231
timestamp 1586364061
transform 1 0 22356 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_243
timestamp 1586364061
transform 1 0 23460 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_13.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 25300 0 1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 25116 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 27232 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 27600 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 27968 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_282
timestamp 1586364061
transform 1 0 27048 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_286
timestamp 1586364061
transform 1 0 27416 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_290
timestamp 1586364061
transform 1 0 27784 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_294
timestamp 1586364061
transform 1 0 28152 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 28888 0 1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_31_298
timestamp 1586364061
transform 1 0 28520 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 774 592
use scs8hd_buf_1  mux_bottom_ipin_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 4232 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_37
timestamp 1586364061
transform 1 0 4508 0 -1 20128
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_3.mux_l2_in_2_
timestamp 1586364061
transform 1 0 5244 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4968 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_41
timestamp 1586364061
transform 1 0 4876 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_54
timestamp 1586364061
transform 1 0 6072 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_58
timestamp 1586364061
transform 1 0 6440 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_70
timestamp 1586364061
transform 1 0 7544 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_82
timestamp 1586364061
transform 1 0 8648 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_90
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_mux2_1  mux_bottom_ipin_7.mux_l2_in_3_
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 11684 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 11316 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_107
timestamp 1586364061
transform 1 0 10948 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_113
timestamp 1586364061
transform 1 0 11500 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 12880 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_126
timestamp 1586364061
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_130
timestamp 1586364061
transform 1 0 13064 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_142
timestamp 1586364061
transform 1 0 14168 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_150
timestamp 1586364061
transform 1 0 14904 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l4_in_0_
timestamp 1586364061
transform 1 0 17204 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16652 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_171
timestamp 1586364061
transform 1 0 16836 0 -1 20128
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l3_in_1_
timestamp 1586364061
transform 1 0 18768 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 18216 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_184
timestamp 1586364061
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_188
timestamp 1586364061
transform 1 0 18400 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 19780 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_201
timestamp 1586364061
transform 1 0 19596 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_205
timestamp 1586364061
transform 1 0 19964 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_213
timestamp 1586364061
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l2_in_2_
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_265
timestamp 1586364061
transform 1 0 25484 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_273
timestamp 1586364061
transform 1 0 26220 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_285
timestamp 1586364061
transform 1 0 27324 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_32_297
timestamp 1586364061
transform 1 0 28428 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 28888 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_6
timestamp 1586364061
transform 1 0 1656 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1840 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_buf_1  mux_bottom_ipin_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_17
timestamp 1586364061
transform 1 0 2668 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_10
timestamp 1586364061
transform 1 0 2024 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2852 0 1 20128
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_ipin_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2392 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_21
timestamp 1586364061
transform 1 0 3036 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_33_33
timestamp 1586364061
transform 1 0 4140 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_38
timestamp 1586364061
transform 1 0 4600 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_8  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 774 592
use scs8hd_mux2_1  mux_bottom_ipin_3.mux_l3_in_1_
timestamp 1586364061
transform 1 0 4968 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 4784 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 4968 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_40
timestamp 1586364061
transform 1 0 4784 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_ipin_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 7268 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_65
timestamp 1586364061
transform 1 0 7084 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_69
timestamp 1586364061
transform 1 0 7452 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_ipin_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 9108 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 9568 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_81
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_90
timestamp 1586364061
transform 1 0 9384 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_94
timestamp 1586364061
transform 1 0 9752 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_106
timestamp 1586364061
transform 1 0 10856 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_7.mux_l4_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use scs8hd_buf_1  mux_bottom_ipin_7.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12144 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_132
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_34_123
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_127
timestamp 1586364061
transform 1 0 12788 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_ipin_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14444 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14904 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_144
timestamp 1586364061
transform 1 0 14352 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_148
timestamp 1586364061
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_152
timestamp 1586364061
transform 1 0 15088 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_139
timestamp 1586364061
transform 1 0 13892 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_34_151
timestamp 1586364061
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_33_164
timestamp 1586364061
transform 1 0 16192 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16468 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_174
timestamp 1586364061
transform 1 0 17112 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_176
timestamp 1586364061
transform 1 0 17296 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_172
timestamp 1586364061
transform 1 0 16928 0 1 20128
box -38 -48 406 592
use scs8hd_buf_1  mux_bottom_ipin_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16652 0 1 20128
box -38 -48 314 592
use scs8hd_buf_1  mux_bottom_ipin_10.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 17204 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18216 0 -1 21216
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18124 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_33_198
timestamp 1586364061
transform 1 0 19320 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_194
timestamp 1586364061
transform 1 0 18952 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_195
timestamp 1586364061
transform 1 0 19044 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_34_207
timestamp 1586364061
transform 1 0 20148 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_33_206
timestamp 1586364061
transform 1 0 20056 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_202
timestamp 1586364061
transform 1 0 19688 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 19504 0 1 20128
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_ipin_11.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20148 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_213
timestamp 1586364061
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_210
timestamp 1586364061
transform 1 0 20424 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20608 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_214
timestamp 1586364061
transform 1 0 20792 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_226
timestamp 1586364061
transform 1 0 21896 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_238
timestamp 1586364061
transform 1 0 23000 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_ipin_13.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24196 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24656 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_254
timestamp 1586364061
transform 1 0 24472 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_conb_1  _27_
timestamp 1586364061
transform 1 0 26404 0 1 20128
box -38 -48 314 592
use scs8hd_buf_1  mux_bottom_ipin_14.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 25208 0 1 20128
box -38 -48 314 592
use scs8hd_buf_1  mux_bottom_ipin_15.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25668 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_258
timestamp 1586364061
transform 1 0 24840 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_265
timestamp 1586364061
transform 1 0 25484 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 26864 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_278
timestamp 1586364061
transform 1 0 26680 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_282
timestamp 1586364061
transform 1 0 27048 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_33_294
timestamp 1586364061
transform 1 0 28152 0 1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_279
timestamp 1586364061
transform 1 0 26772 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_291
timestamp 1586364061
transform 1 0 27876 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 28888 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 28888 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_33_298
timestamp 1586364061
transform 1 0 28520 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_35_32
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_44
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_56
timestamp 1586364061
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_63
timestamp 1586364061
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_87
timestamp 1586364061
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_106
timestamp 1586364061
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_125
timestamp 1586364061
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_137
timestamp 1586364061
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_149
timestamp 1586364061
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_168
timestamp 1586364061
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_180
timestamp 1586364061
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_199
timestamp 1586364061
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_211
timestamp 1586364061
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_218
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_230
timestamp 1586364061
transform 1 0 22264 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23920 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_242
timestamp 1586364061
transform 1 0 23368 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_249
timestamp 1586364061
transform 1 0 24012 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_261
timestamp 1586364061
transform 1 0 25116 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_273
timestamp 1586364061
transform 1 0 26220 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 26772 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_280
timestamp 1586364061
transform 1 0 26864 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_292
timestamp 1586364061
transform 1 0 27968 0 1 21216
box -38 -48 590 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 28888 0 1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_35_298
timestamp 1586364061
transform 1 0 28520 0 1 21216
box -38 -48 130 592
<< labels >>
rlabel metal2 s 3698 0 3754 480 6 bottom_grid_pin_0_
port 0 nsew default tristate
rlabel metal2 s 11150 0 11206 480 6 ccff_head
port 1 nsew default input
rlabel metal2 s 18694 0 18750 480 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[0]
port 3 nsew default input
rlabel metal3 s 0 18232 480 18352 6 chanx_left_in[10]
port 4 nsew default input
rlabel metal3 s 0 18776 480 18896 6 chanx_left_in[11]
port 5 nsew default input
rlabel metal3 s 0 19320 480 19440 6 chanx_left_in[12]
port 6 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chanx_left_in[13]
port 7 nsew default input
rlabel metal3 s 0 20544 480 20664 6 chanx_left_in[14]
port 8 nsew default input
rlabel metal3 s 0 21224 480 21344 6 chanx_left_in[15]
port 9 nsew default input
rlabel metal3 s 0 21768 480 21888 6 chanx_left_in[16]
port 10 nsew default input
rlabel metal3 s 0 22312 480 22432 6 chanx_left_in[17]
port 11 nsew default input
rlabel metal3 s 0 22992 480 23112 6 chanx_left_in[18]
port 12 nsew default input
rlabel metal3 s 0 23536 480 23656 6 chanx_left_in[19]
port 13 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[1]
port 14 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[2]
port 15 nsew default input
rlabel metal3 s 0 14016 480 14136 6 chanx_left_in[3]
port 16 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[4]
port 17 nsew default input
rlabel metal3 s 0 15240 480 15360 6 chanx_left_in[5]
port 18 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[6]
port 19 nsew default input
rlabel metal3 s 0 16328 480 16448 6 chanx_left_in[7]
port 20 nsew default input
rlabel metal3 s 0 17008 480 17128 6 chanx_left_in[8]
port 21 nsew default input
rlabel metal3 s 0 17552 480 17672 6 chanx_left_in[9]
port 22 nsew default input
rlabel metal3 s 0 280 480 400 6 chanx_left_out[0]
port 23 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[10]
port 24 nsew default tristate
rlabel metal3 s 0 6808 480 6928 6 chanx_left_out[11]
port 25 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[12]
port 26 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 chanx_left_out[13]
port 27 nsew default tristate
rlabel metal3 s 0 8576 480 8696 6 chanx_left_out[14]
port 28 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[15]
port 29 nsew default tristate
rlabel metal3 s 0 9800 480 9920 6 chanx_left_out[16]
port 30 nsew default tristate
rlabel metal3 s 0 10344 480 10464 6 chanx_left_out[17]
port 31 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[18]
port 32 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 chanx_left_out[19]
port 33 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_out[1]
port 34 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[2]
port 35 nsew default tristate
rlabel metal3 s 0 2048 480 2168 6 chanx_left_out[3]
port 36 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[4]
port 37 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 chanx_left_out[5]
port 38 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_out[6]
port 39 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 chanx_left_out[7]
port 40 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[8]
port 41 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[9]
port 42 nsew default tristate
rlabel metal3 s 29520 12248 30000 12368 6 chanx_right_in[0]
port 43 nsew default input
rlabel metal3 s 29520 18232 30000 18352 6 chanx_right_in[10]
port 44 nsew default input
rlabel metal3 s 29520 18776 30000 18896 6 chanx_right_in[11]
port 45 nsew default input
rlabel metal3 s 29520 19320 30000 19440 6 chanx_right_in[12]
port 46 nsew default input
rlabel metal3 s 29520 20000 30000 20120 6 chanx_right_in[13]
port 47 nsew default input
rlabel metal3 s 29520 20544 30000 20664 6 chanx_right_in[14]
port 48 nsew default input
rlabel metal3 s 29520 21224 30000 21344 6 chanx_right_in[15]
port 49 nsew default input
rlabel metal3 s 29520 21768 30000 21888 6 chanx_right_in[16]
port 50 nsew default input
rlabel metal3 s 29520 22312 30000 22432 6 chanx_right_in[17]
port 51 nsew default input
rlabel metal3 s 29520 22992 30000 23112 6 chanx_right_in[18]
port 52 nsew default input
rlabel metal3 s 29520 23536 30000 23656 6 chanx_right_in[19]
port 53 nsew default input
rlabel metal3 s 29520 12792 30000 12912 6 chanx_right_in[1]
port 54 nsew default input
rlabel metal3 s 29520 13336 30000 13456 6 chanx_right_in[2]
port 55 nsew default input
rlabel metal3 s 29520 14016 30000 14136 6 chanx_right_in[3]
port 56 nsew default input
rlabel metal3 s 29520 14560 30000 14680 6 chanx_right_in[4]
port 57 nsew default input
rlabel metal3 s 29520 15240 30000 15360 6 chanx_right_in[5]
port 58 nsew default input
rlabel metal3 s 29520 15784 30000 15904 6 chanx_right_in[6]
port 59 nsew default input
rlabel metal3 s 29520 16328 30000 16448 6 chanx_right_in[7]
port 60 nsew default input
rlabel metal3 s 29520 17008 30000 17128 6 chanx_right_in[8]
port 61 nsew default input
rlabel metal3 s 29520 17552 30000 17672 6 chanx_right_in[9]
port 62 nsew default input
rlabel metal3 s 29520 280 30000 400 6 chanx_right_out[0]
port 63 nsew default tristate
rlabel metal3 s 29520 6264 30000 6384 6 chanx_right_out[10]
port 64 nsew default tristate
rlabel metal3 s 29520 6808 30000 6928 6 chanx_right_out[11]
port 65 nsew default tristate
rlabel metal3 s 29520 7352 30000 7472 6 chanx_right_out[12]
port 66 nsew default tristate
rlabel metal3 s 29520 8032 30000 8152 6 chanx_right_out[13]
port 67 nsew default tristate
rlabel metal3 s 29520 8576 30000 8696 6 chanx_right_out[14]
port 68 nsew default tristate
rlabel metal3 s 29520 9256 30000 9376 6 chanx_right_out[15]
port 69 nsew default tristate
rlabel metal3 s 29520 9800 30000 9920 6 chanx_right_out[16]
port 70 nsew default tristate
rlabel metal3 s 29520 10344 30000 10464 6 chanx_right_out[17]
port 71 nsew default tristate
rlabel metal3 s 29520 11024 30000 11144 6 chanx_right_out[18]
port 72 nsew default tristate
rlabel metal3 s 29520 11568 30000 11688 6 chanx_right_out[19]
port 73 nsew default tristate
rlabel metal3 s 29520 824 30000 944 6 chanx_right_out[1]
port 74 nsew default tristate
rlabel metal3 s 29520 1368 30000 1488 6 chanx_right_out[2]
port 75 nsew default tristate
rlabel metal3 s 29520 2048 30000 2168 6 chanx_right_out[3]
port 76 nsew default tristate
rlabel metal3 s 29520 2592 30000 2712 6 chanx_right_out[4]
port 77 nsew default tristate
rlabel metal3 s 29520 3272 30000 3392 6 chanx_right_out[5]
port 78 nsew default tristate
rlabel metal3 s 29520 3816 30000 3936 6 chanx_right_out[6]
port 79 nsew default tristate
rlabel metal3 s 29520 4360 30000 4480 6 chanx_right_out[7]
port 80 nsew default tristate
rlabel metal3 s 29520 5040 30000 5160 6 chanx_right_out[8]
port 81 nsew default tristate
rlabel metal3 s 29520 5584 30000 5704 6 chanx_right_out[9]
port 82 nsew default tristate
rlabel metal2 s 26146 0 26202 480 6 prog_clk
port 83 nsew default input
rlabel metal2 s 938 23520 994 24000 6 top_grid_pin_16_
port 84 nsew default tristate
rlabel metal2 s 2778 23520 2834 24000 6 top_grid_pin_17_
port 85 nsew default tristate
rlabel metal2 s 4618 23520 4674 24000 6 top_grid_pin_18_
port 86 nsew default tristate
rlabel metal2 s 6550 23520 6606 24000 6 top_grid_pin_19_
port 87 nsew default tristate
rlabel metal2 s 8390 23520 8446 24000 6 top_grid_pin_20_
port 88 nsew default tristate
rlabel metal2 s 10230 23520 10286 24000 6 top_grid_pin_21_
port 89 nsew default tristate
rlabel metal2 s 12162 23520 12218 24000 6 top_grid_pin_22_
port 90 nsew default tristate
rlabel metal2 s 14002 23520 14058 24000 6 top_grid_pin_23_
port 91 nsew default tristate
rlabel metal2 s 15934 23520 15990 24000 6 top_grid_pin_24_
port 92 nsew default tristate
rlabel metal2 s 17774 23520 17830 24000 6 top_grid_pin_25_
port 93 nsew default tristate
rlabel metal2 s 19614 23520 19670 24000 6 top_grid_pin_26_
port 94 nsew default tristate
rlabel metal2 s 21546 23520 21602 24000 6 top_grid_pin_27_
port 95 nsew default tristate
rlabel metal2 s 23386 23520 23442 24000 6 top_grid_pin_28_
port 96 nsew default tristate
rlabel metal2 s 25226 23520 25282 24000 6 top_grid_pin_29_
port 97 nsew default tristate
rlabel metal2 s 27158 23520 27214 24000 6 top_grid_pin_30_
port 98 nsew default tristate
rlabel metal2 s 28998 23520 29054 24000 6 top_grid_pin_31_
port 99 nsew default tristate
rlabel metal4 s 5944 2128 6264 21808 6 vpwr
port 100 nsew default input
rlabel metal4 s 10944 2128 11264 21808 6 vgnd
port 101 nsew default input
<< properties >>
string FIXED_BBOX 0 0 30000 24000
<< end >>
