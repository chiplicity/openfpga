* NGSPICE file created from sb_1__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand3_4 abstract view
.subckt scs8hd_nand3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

.subckt sb_1__0_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] chanx_left_in[0] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4]
+ chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_out[0]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_right_in[0] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ left_bottom_grid_pin_11_ left_bottom_grid_pin_13_ left_bottom_grid_pin_15_ left_bottom_grid_pin_1_
+ left_bottom_grid_pin_3_ left_bottom_grid_pin_5_ left_bottom_grid_pin_7_ left_bottom_grid_pin_9_
+ left_top_grid_pin_10_ right_bottom_grid_pin_11_ right_bottom_grid_pin_13_ right_bottom_grid_pin_15_
+ right_bottom_grid_pin_1_ right_bottom_grid_pin_3_ right_bottom_grid_pin_5_ right_bottom_grid_pin_7_
+ right_bottom_grid_pin_9_ right_top_grid_pin_10_ top_left_grid_pin_13_ top_right_grid_pin_11_
+ vpwr vgnd
XFILLER_22_199 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_41 vpwr vgnd scs8hd_fill_2
XFILLER_9_159 vpwr vgnd scs8hd_fill_2
XFILLER_13_188 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_12 vpwr vgnd scs8hd_fill_2
XANTENNA__113__B _112_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_214 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_107 vpwr vgnd scs8hd_fill_2
XFILLER_10_125 vpwr vgnd scs8hd_fill_2
XFILLER_12_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XFILLER_33_206 vgnd vpwr scs8hd_decap_8
XANTENNA__108__B _105_/X vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _074_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_173 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_3_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_206 vgnd vpwr scs8hd_decap_8
XFILLER_15_217 vgnd vpwr scs8hd_decap_12
XFILLER_23_20 vpwr vgnd scs8hd_fill_2
X_062_ _047_/Y address[2] address[0] _079_/A vgnd vpwr scs8hd_or3_4
X_131_ _131_/HI _131_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_31 vpwr vgnd scs8hd_fill_2
XFILLER_2_198 vgnd vpwr scs8hd_decap_4
XFILLER_2_165 vpwr vgnd scs8hd_fill_2
XFILLER_0_79 vgnd vpwr scs8hd_decap_8
XANTENNA__119__A _069_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_66 vpwr vgnd scs8hd_fill_2
XFILLER_12_209 vgnd vpwr scs8hd_decap_4
XFILLER_20_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_64 vpwr vgnd scs8hd_fill_2
X_045_ _045_/A _045_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__105__C address[6] vgnd vpwr scs8hd_diode_2
X_114_ _068_/A address[3] _112_/C _112_/D _114_/Y vgnd vpwr scs8hd_nor4_4
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_4_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__121__B _119_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_4_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_32 vgnd vpwr scs8hd_fill_1
XFILLER_20_87 vgnd vpwr scs8hd_decap_4
XFILLER_6_23 vpwr vgnd scs8hd_fill_2
XANTENNA__116__B _112_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_3
XFILLER_19_172 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_1_.latch data_in mem_right_track_8.LATCH_1_.latch/Q _073_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _131_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_219 vgnd vpwr scs8hd_decap_12
XANTENNA__042__A _042_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_109 vgnd vpwr scs8hd_decap_6
XFILLER_25_197 vgnd vpwr scs8hd_decap_8
XFILLER_15_54 vgnd vpwr scs8hd_fill_1
XFILLER_15_65 vpwr vgnd scs8hd_fill_2
XFILLER_31_75 vgnd vpwr scs8hd_decap_4
XFILLER_31_156 vgnd vpwr scs8hd_fill_1
XFILLER_31_123 vgnd vpwr scs8hd_fill_1
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB _092_/Y vgnd vpwr scs8hd_diode_2
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_134 vpwr vgnd scs8hd_fill_2
XFILLER_22_145 vpwr vgnd scs8hd_fill_2
XFILLER_26_75 vpwr vgnd scs8hd_fill_2
XFILLER_13_112 vpwr vgnd scs8hd_fill_2
XFILLER_13_123 vpwr vgnd scs8hd_fill_2
XFILLER_13_167 vpwr vgnd scs8hd_fill_2
XFILLER_9_138 vpwr vgnd scs8hd_fill_2
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XANTENNA__113__C _112_/C vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_5_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chanx_left_in[0] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A right_bottom_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_88 vpwr vgnd scs8hd_fill_2
XFILLER_33_218 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__124__B _119_/B vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _140_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_8.INVTX1_4_.scs8hd_inv_1 right_bottom_grid_pin_7_ mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__050__A enable vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_130_ _130_/HI _130_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_229 vgnd vpwr scs8hd_decap_4
X_061_ _063_/A _071_/A _061_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_177 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XFILLER_9_12 vpwr vgnd scs8hd_fill_2
XANTENNA__119__B _119_/B vgnd vpwr scs8hd_diode_2
XANTENNA__045__A _045_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_32 vpwr vgnd scs8hd_fill_2
X_113_ address[4] _112_/B _112_/C address[0] _113_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__105__D _083_/D vgnd vpwr scs8hd_diode_2
X_044_ _044_/A _044_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _089_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_7 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.INVTX1_6_.scs8hd_inv_1 left_bottom_grid_pin_5_ mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_20_11 vpwr vgnd scs8hd_fill_2
XFILLER_29_97 vpwr vgnd scs8hd_fill_2
XFILLER_28_195 vgnd vpwr scs8hd_decap_12
XFILLER_28_184 vpwr vgnd scs8hd_fill_2
XFILLER_28_151 vpwr vgnd scs8hd_fill_2
XFILLER_6_46 vpwr vgnd scs8hd_fill_2
XANTENNA__116__C _112_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _081_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_151 vgnd vpwr scs8hd_decap_3
XFILLER_19_195 vpwr vgnd scs8hd_fill_2
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_132 vpwr vgnd scs8hd_fill_2
XFILLER_15_11 vpwr vgnd scs8hd_fill_2
XFILLER_15_22 vpwr vgnd scs8hd_fill_2
XFILLER_15_44 vpwr vgnd scs8hd_fill_2
XFILLER_15_99 vpwr vgnd scs8hd_fill_2
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_168 vgnd vpwr scs8hd_decap_3
XFILLER_31_135 vpwr vgnd scs8hd_fill_2
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_198 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__143__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_22_102 vgnd vpwr scs8hd_decap_3
XFILLER_22_113 vgnd vpwr scs8hd_decap_8
XANTENNA__053__A address[3] vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _042_/Y mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_26_87 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_36 vpwr vgnd scs8hd_fill_2
XANTENNA__113__D address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__138__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_8_161 vpwr vgnd scs8hd_fill_2
XFILLER_8_172 vgnd vpwr scs8hd_decap_12
XANTENNA__048__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_12_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_153 vpwr vgnd scs8hd_fill_2
XFILLER_32_230 vgnd vpwr scs8hd_decap_3
XFILLER_24_219 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[4] mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_99 vgnd vpwr scs8hd_fill_1
X_060_ _047_/Y address[2] _112_/D _071_/A vgnd vpwr scs8hd_or3_4
XFILLER_2_112 vpwr vgnd scs8hd_fill_2
XFILLER_9_24 vgnd vpwr scs8hd_decap_3
XFILLER_9_46 vpwr vgnd scs8hd_fill_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XFILLER_9_79 vpwr vgnd scs8hd_fill_2
XANTENNA__151__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _042_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__061__A _063_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_22 vgnd vpwr scs8hd_decap_8
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _133_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_204 vpwr vgnd scs8hd_fill_2
XFILLER_7_215 vpwr vgnd scs8hd_fill_2
X_112_ address[4] _112_/B _112_/C _112_/D _112_/Y vgnd vpwr scs8hd_nor4_4
X_043_ _043_/A _043_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__146__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_1_80 vpwr vgnd scs8hd_fill_2
XANTENNA__056__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_4_218 vgnd vpwr scs8hd_decap_12
XFILLER_20_56 vgnd vpwr scs8hd_fill_1
XFILLER_29_76 vpwr vgnd scs8hd_fill_2
XFILLER_29_54 vgnd vpwr scs8hd_fill_1
XFILLER_6_69 vpwr vgnd scs8hd_fill_2
XANTENNA__116__D _112_/D vgnd vpwr scs8hd_diode_2
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_111 vgnd vpwr scs8hd_decap_4
XFILLER_15_34 vgnd vpwr scs8hd_fill_1
XFILLER_0_232 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _128_/HI mem_right_track_0.LATCH_2_.latch/Q
+ mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB _069_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_188 vgnd vpwr scs8hd_fill_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_180 vgnd vpwr scs8hd_decap_4
XFILLER_26_22 vgnd vpwr scs8hd_decap_6
XFILLER_9_107 vpwr vgnd scs8hd_fill_2
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_147 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _154_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_140 vgnd vpwr scs8hd_decap_6
XFILLER_8_184 vpwr vgnd scs8hd_fill_2
XFILLER_12_191 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_206 vgnd vpwr scs8hd_decap_8
XANTENNA__064__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _135_/HI vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_0.LATCH_0_.latch data_in mem_top_track_0.LATCH_0_.latch/Q _111_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A left_bottom_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__149__A _149_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_91 vgnd vpwr scs8hd_fill_1
XFILLER_23_231 vpwr vgnd scs8hd_fill_2
XANTENNA__059__A _063_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_27 vpwr vgnd scs8hd_fill_2
XFILLER_0_49 vpwr vgnd scs8hd_fill_2
XFILLER_14_231 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_3_.latch data_in mem_left_track_17.LATCH_3_.latch/Q _100_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__061__B _071_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XFILLER_11_212 vgnd vpwr scs8hd_decap_3
XFILLER_34_99 vgnd vpwr scs8hd_fill_1
X_111_ _074_/A _105_/X _111_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _065_/Y vgnd vpwr scs8hd_diode_2
X_042_ _042_/A _042_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _042_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__162__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_92 vgnd vpwr scs8hd_decap_4
XANTENNA__056__B _112_/B vgnd vpwr scs8hd_diode_2
XANTENNA__072__A _079_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_22 vgnd vpwr scs8hd_decap_12
XFILLER_29_11 vpwr vgnd scs8hd_fill_2
XFILLER_20_46 vpwr vgnd scs8hd_fill_2
XFILLER_20_68 vpwr vgnd scs8hd_fill_2
XFILLER_20_79 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_7 vpwr vgnd scs8hd_fill_2
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XANTENNA__157__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_178 vpwr vgnd scs8hd_fill_2
XFILLER_25_156 vgnd vpwr scs8hd_decap_3
XANTENNA__067__A _063_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_31_56 vgnd vpwr scs8hd_decap_3
XFILLER_31_12 vgnd vpwr scs8hd_decap_12
XFILLER_0_222 vpwr vgnd scs8hd_fill_2
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_3 vgnd vpwr scs8hd_decap_3
XFILLER_22_159 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_1_.latch data_in mem_left_track_1.LATCH_1_.latch/Q _088_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_56 vgnd vpwr scs8hd_decap_6
XFILLER_26_45 vgnd vpwr scs8hd_decap_8
XFILLER_3_16 vgnd vpwr scs8hd_decap_4
XFILLER_3_49 vpwr vgnd scs8hd_fill_2
XFILLER_8_152 vgnd vpwr scs8hd_fill_1
XFILLER_12_181 vgnd vpwr scs8hd_fill_1
Xmem_right_track_16.LATCH_2_.latch data_in mem_right_track_16.LATCH_2_.latch/Q _079_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__064__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_10_129 vgnd vpwr scs8hd_decap_4
XFILLER_12_36 vgnd vpwr scs8hd_decap_3
XANTENNA__080__A _073_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_177 vgnd vpwr scs8hd_decap_4
XFILLER_5_199 vpwr vgnd scs8hd_fill_2
XFILLER_32_210 vgnd vpwr scs8hd_decap_4
XANTENNA__059__B _077_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_79 vgnd vpwr scs8hd_decap_3
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XANTENNA__075__A _068_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_35 vgnd vpwr scs8hd_decap_3
XFILLER_2_169 vgnd vpwr scs8hd_decap_4
XFILLER_2_147 vgnd vpwr scs8hd_decap_6
XFILLER_2_125 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_68 vgnd vpwr scs8hd_decap_4
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
X_110_ _073_/A _105_/X _110_/Y vgnd vpwr scs8hd_nor2_4
X_041_ _041_/A _041_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__056__C _068_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__072__B _073_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_34 vgnd vpwr scs8hd_decap_3
XFILLER_28_154 vpwr vgnd scs8hd_fill_2
XFILLER_28_143 vgnd vpwr scs8hd_decap_8
XFILLER_6_16 vgnd vpwr scs8hd_decap_4
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_10_91 vgnd vpwr scs8hd_fill_1
XFILLER_19_176 vgnd vpwr scs8hd_decap_6
XFILLER_19_187 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
XFILLER_33_190 vpwr vgnd scs8hd_fill_2
XFILLER_31_24 vgnd vpwr scs8hd_decap_12
XANTENNA__067__B _074_/A vgnd vpwr scs8hd_diode_2
XANTENNA__083__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_15_69 vpwr vgnd scs8hd_fill_2
XFILLER_31_79 vgnd vpwr scs8hd_fill_1
XFILLER_31_149 vgnd vpwr scs8hd_decap_4
XFILLER_31_127 vpwr vgnd scs8hd_fill_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_124 vgnd vpwr scs8hd_decap_8
XFILLER_16_168 vgnd vpwr scs8hd_decap_12
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_138 vgnd vpwr scs8hd_decap_4
XFILLER_22_149 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_26_79 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_116 vgnd vpwr scs8hd_decap_4
XANTENNA__078__A _071_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_230 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_219 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__064__C _112_/D vgnd vpwr scs8hd_diode_2
XFILLER_10_108 vpwr vgnd scs8hd_fill_2
XANTENNA__080__B _077_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_9 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_219 vgnd vpwr scs8hd_decap_12
Xmem_right_track_0.LATCH_1_.latch data_in mem_right_track_0.LATCH_1_.latch/Q _065_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_112 vpwr vgnd scs8hd_fill_2
XFILLER_5_134 vpwr vgnd scs8hd_fill_2
Xmem_top_track_8.LATCH_1_.latch data_in _043_/A _114_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_60 vgnd vpwr scs8hd_decap_6
XANTENNA__075__B _112_/B vgnd vpwr scs8hd_diode_2
XANTENNA__091__A _069_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_137 vpwr vgnd scs8hd_fill_2
XFILLER_9_16 vgnd vpwr scs8hd_decap_8
XFILLER_1_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[0] mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_36 vgnd vpwr scs8hd_decap_4
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XANTENNA__086__A _071_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_3 vpwr vgnd scs8hd_fill_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_57 vpwr vgnd scs8hd_fill_2
XFILLER_29_46 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_188 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_199 vgnd vpwr scs8hd_fill_1
XFILLER_34_136 vgnd vpwr scs8hd_fill_1
XFILLER_25_136 vgnd vpwr scs8hd_decap_3
XFILLER_15_26 vpwr vgnd scs8hd_fill_2
XFILLER_15_48 vgnd vpwr scs8hd_decap_6
XFILLER_31_36 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__083__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_31_139 vgnd vpwr scs8hd_fill_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_track_0.LATCH_3_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_60 vgnd vpwr scs8hd_fill_1
XFILLER_7_82 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_2_.latch data_in mem_left_track_9.LATCH_2_.latch/Q _094_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__078__B _077_/B vgnd vpwr scs8hd_diode_2
XANTENNA__094__A _079_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_128 vpwr vgnd scs8hd_fill_2
Xmem_top_track_14.LATCH_0_.latch data_in _046_/A _117_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_154 vpwr vgnd scs8hd_fill_2
XFILLER_16_91 vgnd vpwr scs8hd_fill_1
XFILLER_8_165 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _041_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_27 vpwr vgnd scs8hd_fill_2
XANTENNA__089__A _074_/A vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_3_.latch data_in mem_top_track_16.LATCH_3_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.INVTX1_4_.scs8hd_inv_1 right_bottom_grid_pin_5_ mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_157 vgnd vpwr scs8hd_decap_4
Xmux_top_track_14.tap_buf4_0_.scs8hd_inv_1 mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _155_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_4_83 vpwr vgnd scs8hd_fill_2
XFILLER_23_223 vgnd vpwr scs8hd_decap_8
XFILLER_23_212 vgnd vpwr scs8hd_fill_1
XANTENNA__075__C _068_/C vgnd vpwr scs8hd_diode_2
XFILLER_3_7 vgnd vpwr scs8hd_decap_3
XANTENNA__091__B _090_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_70 vgnd vpwr scs8hd_decap_3
XFILLER_13_92 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A left_bottom_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__086__B _089_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_59 vgnd vpwr scs8hd_decap_3
XFILLER_7_208 vgnd vpwr scs8hd_decap_4
XFILLER_7_219 vpwr vgnd scs8hd_fill_2
XFILLER_24_80 vpwr vgnd scs8hd_fill_2
XFILLER_6_230 vgnd vpwr scs8hd_decap_3
X_099_ _077_/A _102_/B _099_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_3 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_51 vgnd vpwr scs8hd_decap_6
XFILLER_1_62 vpwr vgnd scs8hd_fill_2
XFILLER_1_84 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_5_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_167 vgnd vpwr scs8hd_decap_8
XANTENNA__097__A _068_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_71 vpwr vgnd scs8hd_fill_2
XFILLER_10_82 vgnd vpwr scs8hd_decap_6
XFILLER_10_93 vpwr vgnd scs8hd_fill_2
XFILLER_34_104 vgnd vpwr scs8hd_decap_12
XFILLER_19_101 vpwr vgnd scs8hd_fill_2
XFILLER_19_112 vpwr vgnd scs8hd_fill_2
XFILLER_19_134 vpwr vgnd scs8hd_fill_2
XFILLER_19_156 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB _072_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_115 vgnd vpwr scs8hd_fill_1
XFILLER_31_48 vgnd vpwr scs8hd_decap_8
XANTENNA__083__C _083_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_203 vgnd vpwr scs8hd_decap_3
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_170 vgnd vpwr scs8hd_decap_4
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_81 vpwr vgnd scs8hd_fill_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_22_107 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__094__B _090_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_162 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB _084_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_184 vgnd vpwr scs8hd_decap_12
XFILLER_32_91 vgnd vpwr scs8hd_fill_1
XFILLER_8_111 vgnd vpwr scs8hd_decap_4
XFILLER_8_122 vgnd vpwr scs8hd_fill_1
XFILLER_12_151 vpwr vgnd scs8hd_fill_2
XANTENNA__089__B _089_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_4_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmem_right_track_8.LATCH_2_.latch data_in mem_right_track_8.LATCH_2_.latch/Q _072_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB _076_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_180 vgnd vpwr scs8hd_decap_8
XFILLER_23_16 vpwr vgnd scs8hd_fill_2
XFILLER_23_27 vpwr vgnd scs8hd_fill_2
XFILLER_23_49 vgnd vpwr scs8hd_decap_6
Xmux_left_track_17.INVTX1_6_.scs8hd_inv_1 left_bottom_grid_pin_9_ mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_5_.scs8hd_inv_1 right_bottom_grid_pin_15_ mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_29 vpwr vgnd scs8hd_fill_2
XFILLER_14_213 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_5_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _131_/HI mem_top_track_0.LATCH_5_.latch/Q
+ mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_49 vgnd vpwr scs8hd_decap_8
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_098_ _069_/A _102_/B _098_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_96 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__097__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_3_223 vpwr vgnd scs8hd_fill_2
XFILLER_3_212 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _115_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB _100_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_116 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_168 vpwr vgnd scs8hd_fill_2
XFILLER_33_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__083__D _083_/D vgnd vpwr scs8hd_diode_2
XFILLER_0_226 vgnd vpwr scs8hd_decap_6
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_105 vgnd vpwr scs8hd_decap_8
XFILLER_16_149 vpwr vgnd scs8hd_fill_2
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_60 vgnd vpwr scs8hd_fill_1
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_160 vgnd vpwr scs8hd_decap_4
XFILLER_30_163 vpwr vgnd scs8hd_fill_2
XFILLER_30_152 vgnd vpwr scs8hd_fill_1
XFILLER_7_62 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A right_bottom_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_108 vpwr vgnd scs8hd_fill_2
XFILLER_21_196 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _126_/HI mem_left_track_17.LATCH_2_.latch/Q
+ mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_16_93 vgnd vpwr scs8hd_decap_3
XFILLER_12_130 vgnd vpwr scs8hd_decap_6
XFILLER_35_211 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_26_211 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_92 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _144_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_107 vgnd vpwr scs8hd_decap_3
Xmux_top_track_2.tap_buf4_0_.scs8hd_inv_1 mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _161_/A vgnd vpwr scs8hd_inv_1
XFILLER_13_50 vpwr vgnd scs8hd_fill_2
XFILLER_1_184 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XFILLER_11_217 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _127_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_097_ _068_/A address[3] _083_/C _083_/D _102_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_18 vgnd vpwr scs8hd_decap_12
XFILLER_28_125 vgnd vpwr scs8hd_decap_3
XFILLER_28_103 vgnd vpwr scs8hd_fill_1
XANTENNA__097__C _083_/C vgnd vpwr scs8hd_diode_2
XFILLER_19_71 vgnd vpwr scs8hd_decap_4
XFILLER_34_128 vgnd vpwr scs8hd_decap_8
X_149_ _149_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_32_3 vpwr vgnd scs8hd_fill_2
XFILLER_33_194 vgnd vpwr scs8hd_decap_12
XFILLER_15_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_216 vgnd vpwr scs8hd_fill_1
XFILLER_31_109 vgnd vpwr scs8hd_decap_12
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_72 vgnd vpwr scs8hd_decap_3
XFILLER_30_142 vpwr vgnd scs8hd_fill_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_150 vgnd vpwr scs8hd_decap_4
XFILLER_30_186 vgnd vpwr scs8hd_decap_12
XFILLER_7_52 vpwr vgnd scs8hd_fill_2
XFILLER_26_28 vgnd vpwr scs8hd_fill_1
XFILLER_21_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_72 vpwr vgnd scs8hd_fill_2
XFILLER_16_83 vgnd vpwr scs8hd_decap_8
XFILLER_32_93 vpwr vgnd scs8hd_fill_2
XFILLER_12_197 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_116 vgnd vpwr scs8hd_decap_4
XFILLER_5_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_71 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A right_bottom_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_62 vpwr vgnd scs8hd_fill_2
XFILLER_13_84 vgnd vpwr scs8hd_decap_8
XFILLER_13_95 vpwr vgnd scs8hd_fill_2
XFILLER_1_174 vgnd vpwr scs8hd_decap_3
XANTENNA__100__A _071_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_230 vgnd vpwr scs8hd_decap_3
XFILLER_11_229 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_7 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_200 vgnd vpwr scs8hd_decap_12
X_096_ _074_/A _090_/X _096_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_track_0.LATCH_1_.latch data_in mem_top_track_0.LATCH_1_.latch/Q _110_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_115 vgnd vpwr scs8hd_decap_8
XANTENNA__097__D _083_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.INVTX1_1_.scs8hd_inv_1 chanx_left_in[8] mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_181 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_148_ chanx_left_in[4] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
X_079_ _079_/A _077_/B _079_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_3 vgnd vpwr scs8hd_decap_4
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XFILLER_33_184 vgnd vpwr scs8hd_decap_3
Xmem_left_track_17.LATCH_4_.latch data_in mem_left_track_17.LATCH_4_.latch/Q _099_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_151 vpwr vgnd scs8hd_fill_2
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_21_62 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XPHY_4 vgnd vpwr scs8hd_decap_3
Xmux_left_track_9.INVTX1_5_.scs8hd_inv_1 left_bottom_grid_pin_1_ mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_184 vgnd vpwr scs8hd_decap_3
XFILLER_30_198 vgnd vpwr scs8hd_decap_12
XFILLER_7_86 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _042_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_125 vpwr vgnd scs8hd_fill_2
XFILLER_8_136 vpwr vgnd scs8hd_fill_2
XFILLER_12_165 vgnd vpwr scs8hd_decap_12
XFILLER_16_62 vgnd vpwr scs8hd_fill_1
XFILLER_32_83 vpwr vgnd scs8hd_fill_2
XFILLER_32_72 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A left_bottom_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__103__A _074_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_191 vpwr vgnd scs8hd_fill_2
XFILLER_4_43 vpwr vgnd scs8hd_fill_2
XFILLER_4_32 vpwr vgnd scs8hd_fill_2
XFILLER_4_87 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_153 vpwr vgnd scs8hd_fill_2
Xmem_left_track_1.LATCH_2_.latch data_in mem_left_track_1.LATCH_2_.latch/Q _087_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__100__B _102_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_219 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_16.LATCH_3_.latch data_in mem_right_track_16.LATCH_3_.latch/Q _078_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_84 vgnd vpwr scs8hd_decap_8
XFILLER_24_73 vgnd vpwr scs8hd_decap_4
X_095_ _073_/A _090_/X _095_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_212 vpwr vgnd scs8hd_fill_2
XFILLER_10_230 vgnd vpwr scs8hd_decap_3
XANTENNA__111__A _074_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_66 vgnd vpwr scs8hd_decap_3
XFILLER_1_99 vpwr vgnd scs8hd_fill_2
XFILLER_29_18 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_6_.scs8hd_inv_1 chanx_left_in[1] mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_97 vpwr vgnd scs8hd_fill_2
XFILLER_27_171 vgnd vpwr scs8hd_decap_4
XFILLER_19_40 vpwr vgnd scs8hd_fill_2
XFILLER_19_84 vpwr vgnd scs8hd_fill_2
XFILLER_19_105 vpwr vgnd scs8hd_fill_2
XFILLER_19_116 vgnd vpwr scs8hd_decap_4
XFILLER_19_138 vpwr vgnd scs8hd_fill_2
XFILLER_35_94 vgnd vpwr scs8hd_decap_12
X_147_ chanx_left_in[5] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA__106__A _069_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_078_ _071_/A _077_/B _078_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_185 vpwr vgnd scs8hd_fill_2
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_96 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_3_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB _087_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_130 vpwr vgnd scs8hd_fill_2
XFILLER_7_10 vgnd vpwr scs8hd_decap_4
XFILLER_21_100 vgnd vpwr scs8hd_decap_3
XFILLER_21_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_155 vgnd vpwr scs8hd_decap_4
XFILLER_16_30 vgnd vpwr scs8hd_fill_1
XFILLER_8_115 vgnd vpwr scs8hd_fill_1
XFILLER_8_148 vgnd vpwr scs8hd_decap_4
XFILLER_12_177 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_3_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__103__B _102_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB _079_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_203 vgnd vpwr scs8hd_decap_8
XFILLER_27_51 vpwr vgnd scs8hd_fill_2
XFILLER_17_214 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_2_.scs8hd_inv_1 chany_top_in[7] mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__114__A _068_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_198 vpwr vgnd scs8hd_fill_2
XANTENNA__109__A _079_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_209 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_094_ _079_/A _090_/X _094_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__111__B _105_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_34 vpwr vgnd scs8hd_fill_2
Xmem_right_track_0.LATCH_2_.latch data_in mem_right_track_0.LATCH_2_.latch/Q _063_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _103_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_139 vpwr vgnd scs8hd_fill_2
XFILLER_3_227 vgnd vpwr scs8hd_decap_6
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_27_194 vgnd vpwr scs8hd_decap_12
XFILLER_27_150 vpwr vgnd scs8hd_fill_2
X_077_ _077_/A _077_/B _077_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__106__B _105_/X vgnd vpwr scs8hd_diode_2
XANTENNA__122__A _079_/A vgnd vpwr scs8hd_diode_2
X_146_ chanx_left_in[6] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_33_142 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_208 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_24_120 vgnd vpwr scs8hd_decap_3
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_20 vpwr vgnd scs8hd_fill_2
XFILLER_21_53 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_175 vgnd vpwr scs8hd_decap_6
XFILLER_30_167 vgnd vpwr scs8hd_decap_4
XFILLER_7_66 vgnd vpwr scs8hd_fill_1
XANTENNA__117__A _068_/A vgnd vpwr scs8hd_diode_2
X_129_ _129_/HI _129_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_99 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_21_123 vgnd vpwr scs8hd_decap_3
Xmux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_145 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _130_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_182 vgnd vpwr scs8hd_fill_1
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_32_218 vgnd vpwr scs8hd_decap_12
XANTENNA__114__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_4_163 vpwr vgnd scs8hd_fill_2
XFILLER_4_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_54 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_3_.latch data_in mem_left_track_9.LATCH_3_.latch/Q _093_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_3 vpwr vgnd scs8hd_fill_2
XANTENNA__109__B _105_/X vgnd vpwr scs8hd_diode_2
Xmem_top_track_14.LATCH_1_.latch data_in _045_/A _116_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_24_42 vpwr vgnd scs8hd_fill_2
X_162_ _162_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
X_093_ _071_/A _090_/X _093_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_13 vgnd vpwr scs8hd_fill_1
Xmem_top_track_16.LATCH_4_.latch data_in mem_top_track_16.LATCH_4_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_217 vgnd vpwr scs8hd_decap_3
XFILLER_10_44 vgnd vpwr scs8hd_fill_1
XFILLER_10_88 vgnd vpwr scs8hd_fill_1
XFILLER_19_53 vgnd vpwr scs8hd_decap_4
XFILLER_35_63 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vgnd vpwr scs8hd_fill_1
XFILLER_19_75 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_right_track_0.LATCH_4_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_145_ _145_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_32_7 vgnd vpwr scs8hd_decap_3
XANTENNA__122__B _119_/B vgnd vpwr scs8hd_diode_2
X_076_ _069_/A _077_/B _076_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_24_143 vgnd vpwr scs8hd_decap_8
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_3
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_146 vgnd vpwr scs8hd_decap_6
XFILLER_30_102 vgnd vpwr scs8hd_decap_3
XPHY_7 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB _061_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_198 vpwr vgnd scs8hd_fill_2
XFILLER_7_34 vgnd vpwr scs8hd_decap_3
XFILLER_7_56 vpwr vgnd scs8hd_fill_2
XFILLER_7_78 vpwr vgnd scs8hd_fill_2
X_128_ _128_/HI _128_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__117__B _112_/B vgnd vpwr scs8hd_diode_2
X_059_ _063_/A _077_/A _059_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_3 vpwr vgnd scs8hd_fill_2
XFILLER_21_135 vpwr vgnd scs8hd_fill_2
XFILLER_21_179 vgnd vpwr scs8hd_decap_4
XANTENNA__043__A _043_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_102 vgnd vpwr scs8hd_decap_8
XFILLER_16_43 vgnd vpwr scs8hd_decap_8
XFILLER_16_54 vgnd vpwr scs8hd_decap_8
XFILLER_16_76 vgnd vpwr scs8hd_decap_4
XFILLER_32_64 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A left_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_172 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.INVTX1_2_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_227 vgnd vpwr scs8hd_decap_6
XFILLER_27_97 vpwr vgnd scs8hd_fill_2
XFILLER_4_13 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__114__C _112_/C vgnd vpwr scs8hd_diode_2
XFILLER_4_79 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_219 vpwr vgnd scs8hd_fill_2
XFILLER_23_208 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_219 vgnd vpwr scs8hd_decap_12
XFILLER_13_66 vpwr vgnd scs8hd_fill_2
XFILLER_1_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__141__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__051__A address[6] vgnd vpwr scs8hd_diode_2
X_161_ _161_/A chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_24_32 vgnd vpwr scs8hd_fill_1
X_092_ _077_/A _090_/X _092_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_47 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_3_.latch data_in mem_right_track_8.LATCH_3_.latch/Q _071_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__136__A _136_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__046__A _046_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_23 vpwr vgnd scs8hd_fill_2
XFILLER_35_75 vgnd vpwr scs8hd_decap_12
X_144_ _144_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
X_075_ _068_/A _112_/B _068_/C _077_/B vgnd vpwr scs8hd_or3_4
XFILLER_18_141 vgnd vpwr scs8hd_decap_6
XFILLER_18_163 vgnd vpwr scs8hd_decap_8
XFILLER_18_174 vgnd vpwr scs8hd_decap_12
XFILLER_33_155 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _110_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_166 vpwr vgnd scs8hd_fill_2
XFILLER_2_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_2_.scs8hd_inv_1 chany_top_in[8] mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_77 vpwr vgnd scs8hd_fill_2
XFILLER_30_114 vgnd vpwr scs8hd_decap_12
XPHY_8 vgnd vpwr scs8hd_decap_3
XANTENNA__117__C _112_/C vgnd vpwr scs8hd_diode_2
XFILLER_15_111 vpwr vgnd scs8hd_fill_2
X_058_ address[1] _048_/Y address[0] _077_/A vgnd vpwr scs8hd_or3_4
X_127_ _127_/HI _127_/LO vgnd vpwr scs8hd_conb_1
XFILLER_16_3 vgnd vpwr scs8hd_decap_4
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_5_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_107 vpwr vgnd scs8hd_fill_2
XFILLER_8_118 vgnd vpwr scs8hd_decap_4
XFILLER_16_22 vgnd vpwr scs8hd_decap_8
XFILLER_32_87 vgnd vpwr scs8hd_decap_4
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XFILLER_20_180 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__144__A _144_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_162 vgnd vpwr scs8hd_fill_1
Xmux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _045_/A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB _093_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__054__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_17_217 vgnd vpwr scs8hd_decap_12
XFILLER_4_47 vgnd vpwr scs8hd_decap_4
XANTENNA__114__D _112_/D vgnd vpwr scs8hd_diode_2
XANTENNA__139__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__049__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_14_209 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_179 vpwr vgnd scs8hd_fill_2
XFILLER_1_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_3_.scs8hd_inv_1 right_bottom_grid_pin_1_ mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_160_ chanx_right_in[4] chany_top_out[2] vgnd vpwr scs8hd_buf_2
X_091_ _069_/A _090_/X _091_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_201 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XANTENNA__152__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__062__A _047_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_57 vgnd vpwr scs8hd_decap_12
XFILLER_19_88 vpwr vgnd scs8hd_fill_2
XFILLER_35_87 vgnd vpwr scs8hd_decap_6
XFILLER_35_32 vgnd vpwr scs8hd_decap_12
X_074_ _074_/A _073_/B _074_/Y vgnd vpwr scs8hd_nor2_4
X_143_ chanx_right_in[0] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_2_230 vgnd vpwr scs8hd_decap_3
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
XFILLER_18_7 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_120 vgnd vpwr scs8hd_decap_3
XFILLER_18_186 vgnd vpwr scs8hd_decap_12
XANTENNA__147__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_24_189 vgnd vpwr scs8hd_decap_12
XFILLER_24_134 vpwr vgnd scs8hd_fill_2
XFILLER_24_112 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.INVTX1_5_.scs8hd_inv_1 left_top_grid_pin_10_ mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__057__A _069_/A vgnd vpwr scs8hd_diode_2
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_45 vpwr vgnd scs8hd_fill_2
XFILLER_21_56 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_134 vgnd vpwr scs8hd_decap_3
XFILLER_30_137 vgnd vpwr scs8hd_decap_3
XFILLER_30_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__117__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_15_156 vpwr vgnd scs8hd_fill_2
X_126_ _126_/HI _126_/LO vgnd vpwr scs8hd_conb_1
X_057_ _069_/A _063_/A _057_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_21_159 vgnd vpwr scs8hd_fill_1
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_218 vgnd vpwr scs8hd_decap_12
XFILLER_7_130 vpwr vgnd scs8hd_fill_2
XANTENNA__160__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
X_109_ _079_/A _105_/X _109_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__054__B _048_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__070__A _077_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_77 vpwr vgnd scs8hd_fill_2
XFILLER_27_55 vgnd vpwr scs8hd_decap_4
XFILLER_17_229 vgnd vpwr scs8hd_decap_4
XFILLER_4_199 vgnd vpwr scs8hd_decap_12
XFILLER_4_133 vgnd vpwr scs8hd_decap_8
XFILLER_31_210 vgnd vpwr scs8hd_fill_1
XANTENNA__155__A _155_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__065__A _063_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_114 vpwr vgnd scs8hd_fill_2
XFILLER_0_191 vgnd vpwr scs8hd_fill_1
X_090_ address[4] _112_/B _083_/C _083_/D _090_/X vgnd vpwr scs8hd_or4_4
XFILLER_10_213 vgnd vpwr scs8hd_fill_1
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_3 vgnd vpwr scs8hd_decap_8
Xmux_right_track_0.INVTX1_6_.scs8hd_inv_1 chanx_left_in[0] mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__062__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_10_47 vgnd vpwr scs8hd_fill_1
XFILLER_27_154 vpwr vgnd scs8hd_fill_2
XFILLER_27_132 vgnd vpwr scs8hd_decap_4
XFILLER_19_23 vgnd vpwr scs8hd_decap_4
XFILLER_19_78 vgnd vpwr scs8hd_decap_3
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_44 vgnd vpwr scs8hd_decap_12
X_142_ chanx_right_in[1] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
X_073_ _073_/A _073_/B _073_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_146 vgnd vpwr scs8hd_decap_6
XFILLER_33_102 vpwr vgnd scs8hd_fill_2
XFILLER_18_198 vgnd vpwr scs8hd_decap_12
XFILLER_2_70 vgnd vpwr scs8hd_fill_1
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__057__B _063_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__073__A _073_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_24 vgnd vpwr scs8hd_decap_8
XFILLER_7_48 vpwr vgnd scs8hd_fill_2
X_125_ _125_/HI _125_/LO vgnd vpwr scs8hd_conb_1
XFILLER_30_7 vgnd vpwr scs8hd_decap_8
X_056_ address[4] _112_/B _068_/C _063_/A vgnd vpwr scs8hd_or3_4
XANTENNA__158__A _158_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_205 vgnd vpwr scs8hd_decap_12
XANTENNA__068__A _068_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_56 vgnd vpwr scs8hd_decap_6
Xmem_top_track_0.LATCH_2_.latch data_in mem_top_track_0.LATCH_2_.latch/Q _109_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_127 vgnd vpwr scs8hd_fill_1
X_108_ _071_/A _105_/X _108_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A right_bottom_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB _070_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__070__B _073_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__054__C _112_/D vgnd vpwr scs8hd_diode_2
XFILLER_8_91 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _158_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_45 vgnd vpwr scs8hd_decap_4
XFILLER_17_208 vgnd vpwr scs8hd_decap_6
Xmem_left_track_17.LATCH_5_.latch data_in mem_left_track_17.LATCH_5_.latch/Q _098_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_167 vpwr vgnd scs8hd_fill_2
XFILLER_4_145 vpwr vgnd scs8hd_fill_2
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XFILLER_16_230 vgnd vpwr scs8hd_decap_3
XFILLER_22_211 vgnd vpwr scs8hd_decap_3
XANTENNA__065__B _073_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_25 vpwr vgnd scs8hd_fill_2
XFILLER_13_58 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__081__A _074_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_7 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_24_46 vgnd vpwr scs8hd_decap_12
XANTENNA__076__A _069_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__062__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_35_56 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A right_bottom_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_177 vpwr vgnd scs8hd_fill_2
X_141_ chanx_right_in[2] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
X_072_ _079_/A _073_/B _072_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _043_/A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _067_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_3_.latch data_in mem_left_track_1.LATCH_3_.latch/Q _086_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_93 vpwr vgnd scs8hd_fill_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__073__B _073_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_103 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_180 vgnd vpwr scs8hd_decap_3
XFILLER_7_16 vgnd vpwr scs8hd_decap_3
X_124_ _074_/A _119_/B _124_/Y vgnd vpwr scs8hd_nor2_4
X_055_ enable address[5] _083_/C _068_/C vgnd vpwr scs8hd_nand3_4
Xmem_right_track_16.LATCH_4_.latch data_in mem_right_track_16.LATCH_4_.latch/Q _077_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_139 vgnd vpwr scs8hd_decap_3
XFILLER_29_217 vgnd vpwr scs8hd_decap_12
XANTENNA__068__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_32_68 vgnd vpwr scs8hd_fill_1
XFILLER_32_13 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_161 vpwr vgnd scs8hd_fill_2
XANTENNA__084__A _069_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB _098_/Y vgnd vpwr scs8hd_diode_2
X_107_ _077_/A _105_/X _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_110 vpwr vgnd scs8hd_fill_2
XFILLER_7_143 vpwr vgnd scs8hd_fill_2
XFILLER_7_154 vpwr vgnd scs8hd_fill_2
XFILLER_7_176 vgnd vpwr scs8hd_decap_6
XFILLER_7_187 vpwr vgnd scs8hd_fill_2
XANTENNA__079__A _079_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_102 vpwr vgnd scs8hd_fill_2
XFILLER_17_90 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _044_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__081__B _077_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_138 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_212 vgnd vpwr scs8hd_decap_3
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
XFILLER_5_82 vpwr vgnd scs8hd_fill_2
XFILLER_5_93 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_69 vpwr vgnd scs8hd_fill_2
XFILLER_24_58 vpwr vgnd scs8hd_fill_2
XANTENNA__076__B _077_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__092__A _077_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_29 vgnd vpwr scs8hd_decap_3
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_19_36 vpwr vgnd scs8hd_fill_2
XFILLER_27_123 vgnd vpwr scs8hd_decap_3
XFILLER_27_112 vpwr vgnd scs8hd_fill_2
XANTENNA__087__A _079_/A vgnd vpwr scs8hd_diode_2
X_140_ _140_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
X_071_ _071_/A _073_/B _071_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_4_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_33_159 vgnd vpwr scs8hd_decap_12
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_83 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_4_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 chanx_left_in[7] mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_115 vpwr vgnd scs8hd_fill_2
XFILLER_15_126 vpwr vgnd scs8hd_fill_2
X_123_ _073_/A _119_/B _123_/Y vgnd vpwr scs8hd_nor2_4
X_054_ address[1] _048_/Y _112_/D _069_/A vgnd vpwr scs8hd_or3_4
XFILLER_7_28 vgnd vpwr scs8hd_decap_4
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_229 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_3_.latch data_in mem_right_track_0.LATCH_3_.latch/Q _061_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__068__C _068_/C vgnd vpwr scs8hd_diode_2
XFILLER_32_25 vgnd vpwr scs8hd_decap_6
XANTENNA__084__B _089_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _096_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_140 vpwr vgnd scs8hd_fill_2
XFILLER_11_162 vpwr vgnd scs8hd_fill_2
X_106_ _069_/A _105_/X _106_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_195 vpwr vgnd scs8hd_fill_2
XFILLER_8_93 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__079__B _077_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_25 vpwr vgnd scs8hd_fill_2
XFILLER_27_14 vpwr vgnd scs8hd_fill_2
XFILLER_25_232 vgnd vpwr scs8hd_fill_1
XANTENNA__095__A _073_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_125 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_210 vgnd vpwr scs8hd_decap_4
XFILLER_33_90 vgnd vpwr scs8hd_decap_8
XFILLER_0_150 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_15 vpwr vgnd scs8hd_fill_2
XANTENNA__092__B _090_/X vgnd vpwr scs8hd_diode_2
XFILLER_10_205 vgnd vpwr scs8hd_decap_8
XFILLER_30_91 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__087__B _089_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_070_ _077_/A _073_/B _070_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_4_3 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.INVTX1_2_.scs8hd_inv_1 chany_top_in[6] mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_138 vpwr vgnd scs8hd_fill_2
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_left_track_9.LATCH_4_.latch data_in mem_left_track_9.LATCH_4_.latch/Q _092_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _046_/A mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_2_73 vgnd vpwr scs8hd_fill_1
XFILLER_24_138 vgnd vpwr scs8hd_decap_3
XFILLER_24_116 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_16 vpwr vgnd scs8hd_fill_2
XFILLER_21_49 vgnd vpwr scs8hd_decap_4
XANTENNA__098__A _069_/A vgnd vpwr scs8hd_diode_2
X_122_ _079_/A _119_/B _122_/Y vgnd vpwr scs8hd_nor2_4
X_053_ address[3] _112_/B vgnd vpwr scs8hd_inv_8
XFILLER_11_60 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_5_.latch data_in mem_top_track_16.LATCH_5_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_119 vgnd vpwr scs8hd_decap_8
Xmux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_105_ address[4] address[3] address[6] _083_/D _105_/X vgnd vpwr scs8hd_or4_4
XFILLER_19_230 vgnd vpwr scs8hd_decap_3
XFILLER_8_50 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__095__B _090_/X vgnd vpwr scs8hd_diode_2
XFILLER_31_225 vpwr vgnd scs8hd_fill_2
XFILLER_31_214 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_13_ mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
XFILLER_9_207 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_218 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_3_.scs8hd_inv_1 right_top_grid_pin_10_ mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_62 vgnd vpwr scs8hd_decap_3
Xmux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_5_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_81 vpwr vgnd scs8hd_fill_2
XFILLER_30_70 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_210 vpwr vgnd scs8hd_fill_2
XFILLER_5_221 vpwr vgnd scs8hd_fill_2
XFILLER_14_93 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_158 vpwr vgnd scs8hd_fill_2
XFILLER_27_136 vgnd vpwr scs8hd_fill_1
XFILLER_35_180 vgnd vpwr scs8hd_decap_6
XFILLER_2_213 vgnd vpwr scs8hd_fill_1
XFILLER_2_202 vgnd vpwr scs8hd_fill_1
XFILLER_33_106 vpwr vgnd scs8hd_fill_2
XFILLER_26_191 vgnd vpwr scs8hd_decap_12
XFILLER_18_125 vpwr vgnd scs8hd_fill_2
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__098__B _102_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_150 vgnd vpwr scs8hd_fill_1
X_121_ _071_/A _119_/B _121_/Y vgnd vpwr scs8hd_nor2_4
X_052_ address[4] _068_/A vgnd vpwr scs8hd_inv_8
XFILLER_11_83 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A left_bottom_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_161 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_8.LATCH_4_.latch data_in mem_right_track_8.LATCH_4_.latch/Q _070_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_197 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _073_/Y vgnd vpwr scs8hd_diode_2
X_104_ address[6] _083_/D _112_/C vgnd vpwr scs8hd_or2_4
XFILLER_11_175 vpwr vgnd scs8hd_fill_2
Xmem_top_track_2.LATCH_0_.latch data_in _042_/A _113_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_left_track_17.LATCH_0_.latch data_in mem_left_track_17.LATCH_0_.latch/Q _103_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_190 vgnd vpwr scs8hd_fill_1
XFILLER_8_84 vgnd vpwr scs8hd_decap_4
XFILLER_25_212 vgnd vpwr scs8hd_decap_12
XFILLER_4_149 vpwr vgnd scs8hd_fill_2
XFILLER_3_171 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _127_/HI mem_left_track_9.LATCH_2_.latch/Q
+ mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_12_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_215 vgnd vpwr scs8hd_decap_12
XFILLER_13_29 vpwr vgnd scs8hd_fill_2
XFILLER_13_204 vgnd vpwr scs8hd_decap_8
XFILLER_0_163 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ _042_/A mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_5_96 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB _077_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_93 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_5_.scs8hd_inv_1 left_bottom_grid_pin_3_ mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_4_.scs8hd_inv_1 right_bottom_grid_pin_9_ mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_19 vpwr vgnd scs8hd_fill_2
XFILLER_35_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _132_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_25_71 vpwr vgnd scs8hd_fill_2
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _154_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_97 vgnd vpwr scs8hd_fill_1
XFILLER_17_181 vpwr vgnd scs8hd_fill_2
XFILLER_15_107 vpwr vgnd scs8hd_fill_2
XFILLER_23_184 vgnd vpwr scs8hd_decap_12
X_120_ _077_/A _119_/B _120_/Y vgnd vpwr scs8hd_nor2_4
X_051_ address[6] _083_/C vgnd vpwr scs8hd_inv_8
XFILLER_11_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _043_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _132_/HI _045_/Y mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_18 vpwr vgnd scs8hd_fill_2
XFILLER_20_121 vpwr vgnd scs8hd_fill_2
XFILLER_20_165 vpwr vgnd scs8hd_fill_2
XFILLER_11_110 vpwr vgnd scs8hd_fill_2
X_103_ _074_/A _102_/B _103_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_103 vpwr vgnd scs8hd_fill_2
XFILLER_7_114 vgnd vpwr scs8hd_decap_6
XFILLER_7_147 vgnd vpwr scs8hd_decap_4
XFILLER_7_158 vpwr vgnd scs8hd_fill_2
XFILLER_22_50 vgnd vpwr scs8hd_decap_6
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_14_7 vpwr vgnd scs8hd_fill_2
XFILLER_25_224 vgnd vpwr scs8hd_decap_8
XFILLER_4_106 vgnd vpwr scs8hd_decap_4
XFILLER_22_227 vgnd vpwr scs8hd_decap_6
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _044_/A mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_93 vgnd vpwr scs8hd_decap_8
XFILLER_28_60 vpwr vgnd scs8hd_fill_2
XFILLER_8_231 vpwr vgnd scs8hd_fill_2
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_5_31 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _149_/A vgnd vpwr scs8hd_inv_1
XANTENNA__101__A _079_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_19_29 vpwr vgnd scs8hd_fill_2
XFILLER_27_116 vgnd vpwr scs8hd_decap_6
XFILLER_18_149 vgnd vpwr scs8hd_decap_4
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_25_94 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_2_43 vpwr vgnd scs8hd_fill_2
XFILLER_2_32 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_108 vpwr vgnd scs8hd_fill_2
XFILLER_2_87 vgnd vpwr scs8hd_fill_1
XFILLER_17_160 vpwr vgnd scs8hd_fill_2
XFILLER_32_174 vgnd vpwr scs8hd_decap_12
XFILLER_32_163 vgnd vpwr scs8hd_decap_8
XFILLER_32_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_130 vgnd vpwr scs8hd_decap_3
XFILLER_15_119 vgnd vpwr scs8hd_decap_3
XFILLER_23_196 vgnd vpwr scs8hd_decap_12
X_050_ enable _082_/A vgnd vpwr scs8hd_inv_8
XFILLER_11_41 vpwr vgnd scs8hd_fill_2
XFILLER_11_52 vpwr vgnd scs8hd_fill_2
XFILLER_14_141 vpwr vgnd scs8hd_fill_2
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_20_111 vgnd vpwr scs8hd_decap_8
XFILLER_20_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_144 vgnd vpwr scs8hd_decap_3
X_102_ _073_/A _102_/B _102_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_126 vpwr vgnd scs8hd_fill_2
XFILLER_11_199 vpwr vgnd scs8hd_fill_2
XFILLER_22_40 vgnd vpwr scs8hd_fill_1
XFILLER_22_84 vpwr vgnd scs8hd_fill_2
XFILLER_19_222 vgnd vpwr scs8hd_decap_8
XFILLER_27_29 vgnd vpwr scs8hd_decap_3
XFILLER_27_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_51 vgnd vpwr scs8hd_decap_8
XFILLER_17_62 vpwr vgnd scs8hd_fill_2
XFILLER_17_73 vpwr vgnd scs8hd_fill_2
XFILLER_3_195 vpwr vgnd scs8hd_fill_2
XFILLER_3_140 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB _057_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__104__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_217 vgnd vpwr scs8hd_decap_12
XFILLER_28_72 vgnd vpwr scs8hd_decap_3
XFILLER_0_187 vgnd vpwr scs8hd_decap_4
Xmem_top_track_0.LATCH_3_.latch data_in mem_top_track_0.LATCH_3_.latch/Q _108_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_24_19 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_30 vgnd vpwr scs8hd_fill_1
XANTENNA__101__B _102_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_19 vpwr vgnd scs8hd_fill_2
XFILLER_27_128 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_4_7 vgnd vpwr scs8hd_decap_6
XFILLER_2_205 vgnd vpwr scs8hd_decap_8
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 chanx_left_in[6] mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_161 vgnd vpwr scs8hd_fill_1
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_51 vpwr vgnd scs8hd_fill_2
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_2_66 vgnd vpwr scs8hd_decap_4
XFILLER_2_55 vpwr vgnd scs8hd_fill_2
XANTENNA__112__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_32_186 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_153 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_0_.latch data_in mem_top_track_16.LATCH_0_.latch/Q _124_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_86 vpwr vgnd scs8hd_fill_2
XANTENNA__107__A _077_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_197 vgnd vpwr scs8hd_decap_12
XFILLER_28_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A right_bottom_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_101 vgnd vpwr scs8hd_fill_1
XFILLER_9_190 vpwr vgnd scs8hd_fill_2
Xmux_top_track_14.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_101_ _079_/A _102_/B _101_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_123 vpwr vgnd scs8hd_fill_2
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_43 vgnd vpwr scs8hd_decap_4
XFILLER_6_182 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_119 vgnd vpwr scs8hd_decap_4
Xmux_left_track_9.INVTX1_4_.scs8hd_inv_1 chanx_right_in[5] mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_left_track_1.LATCH_4_.latch data_in mem_left_track_1.LATCH_4_.latch/Q _085_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_31_229 vgnd vpwr scs8hd_decap_4
XFILLER_31_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_73 vpwr vgnd scs8hd_fill_2
XFILLER_33_62 vgnd vpwr scs8hd_decap_8
XANTENNA__104__B _083_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _077_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_3_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_229 vgnd vpwr scs8hd_decap_4
Xmem_right_track_16.LATCH_5_.latch data_in mem_right_track_16.LATCH_5_.latch/Q _076_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_28_84 vpwr vgnd scs8hd_fill_2
XANTENNA__115__A _068_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A right_bottom_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB _091_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_30 vgnd vpwr scs8hd_fill_1
XFILLER_5_203 vpwr vgnd scs8hd_fill_2
XFILLER_5_214 vpwr vgnd scs8hd_fill_2
XFILLER_5_225 vgnd vpwr scs8hd_decap_8
XFILLER_14_75 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _135_/HI _043_/Y mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_85 vgnd vpwr scs8hd_decap_6
XFILLER_29_170 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _044_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[3] mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_18_129 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_2_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__112__B _112_/B vgnd vpwr scs8hd_diode_2
XFILLER_17_140 vgnd vpwr scs8hd_decap_4
XFILLER_17_173 vgnd vpwr scs8hd_decap_8
XFILLER_17_184 vgnd vpwr scs8hd_decap_12
XFILLER_32_198 vgnd vpwr scs8hd_decap_12
XFILLER_23_176 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_5_.scs8hd_inv_1 right_bottom_grid_pin_13_ mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__107__B _105_/X vgnd vpwr scs8hd_diode_2
XANTENNA__123__A _073_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_157 vpwr vgnd scs8hd_fill_2
XFILLER_9_180 vgnd vpwr scs8hd_fill_1
XFILLER_28_213 vgnd vpwr scs8hd_fill_1
XFILLER_11_179 vpwr vgnd scs8hd_fill_2
X_100_ _071_/A _102_/B _100_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_227 vgnd vpwr scs8hd_decap_6
XANTENNA__118__A address[4] vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_88 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _046_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_1.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_11_ mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_31 vgnd vpwr scs8hd_fill_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_175 vpwr vgnd scs8hd_fill_2
XANTENNA__120__B _119_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _080_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_178 vpwr vgnd scs8hd_fill_2
XFILLER_0_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_41 vgnd vpwr scs8hd_decap_8
Xmem_right_track_0.LATCH_4_.latch data_in mem_right_track_0.LATCH_4_.latch/Q _059_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_201 vgnd vpwr scs8hd_decap_12
XFILLER_12_230 vgnd vpwr scs8hd_decap_3
XFILLER_5_78 vpwr vgnd scs8hd_fill_2
XFILLER_5_12 vpwr vgnd scs8hd_fill_2
XFILLER_5_89 vgnd vpwr scs8hd_decap_4
XANTENNA__115__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__041__A _041_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_2_.scs8hd_inv_1 chany_top_in[7] mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_32 vpwr vgnd scs8hd_fill_2
XFILLER_14_87 vgnd vpwr scs8hd_decap_3
XFILLER_30_97 vgnd vpwr scs8hd_decap_3
XFILLER_30_53 vgnd vpwr scs8hd_decap_8
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _133_/HI mem_top_track_16.LATCH_5_.latch/Q
+ mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_193 vgnd vpwr scs8hd_decap_12
XFILLER_2_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
Xmux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_5_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_141 vgnd vpwr scs8hd_decap_12
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_18_108 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_25_75 vgnd vpwr scs8hd_decap_8
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__112__C _112_/C vgnd vpwr scs8hd_diode_2
XFILLER_2_13 vgnd vpwr scs8hd_fill_1
XFILLER_32_144 vgnd vpwr scs8hd_decap_8
XFILLER_17_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_166 vgnd vpwr scs8hd_decap_8
XFILLER_11_33 vpwr vgnd scs8hd_fill_2
XFILLER_11_66 vpwr vgnd scs8hd_fill_2
XFILLER_11_99 vpwr vgnd scs8hd_fill_2
XANTENNA__123__B _119_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_136 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_103 vpwr vgnd scs8hd_fill_2
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XFILLER_11_136 vpwr vgnd scs8hd_fill_2
XFILLER_11_158 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vpwr vgnd scs8hd_fill_2
XFILLER_19_203 vpwr vgnd scs8hd_fill_2
XFILLER_19_214 vpwr vgnd scs8hd_fill_2
XANTENNA__118__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
X_159_ chanx_right_in[5] chany_top_out[3] vgnd vpwr scs8hd_buf_2
Xmux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_left_track_9.LATCH_5_.latch data_in mem_left_track_9.LATCH_5_.latch/Q _091_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__044__A _044_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _126_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_10 vpwr vgnd scs8hd_fill_2
XFILLER_17_43 vpwr vgnd scs8hd_fill_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_31 vpwr vgnd scs8hd_fill_2
XFILLER_3_154 vpwr vgnd scs8hd_fill_2
XFILLER_3_143 vpwr vgnd scs8hd_fill_2
XFILLER_3_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_220 vgnd vpwr scs8hd_decap_12
XFILLER_0_146 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_64 vpwr vgnd scs8hd_fill_2
XFILLER_8_213 vgnd vpwr scs8hd_fill_1
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XFILLER_5_35 vpwr vgnd scs8hd_fill_2
XANTENNA__115__C _112_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_11 vpwr vgnd scs8hd_fill_2
XFILLER_14_22 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _046_/Y mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__142__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__052__A address[4] vgnd vpwr scs8hd_diode_2
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_164 vgnd vpwr scs8hd_fill_1
XFILLER_26_131 vgnd vpwr scs8hd_fill_1
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_32 vpwr vgnd scs8hd_fill_2
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XANTENNA__112__D _112_/D vgnd vpwr scs8hd_diode_2
XFILLER_2_47 vgnd vpwr scs8hd_decap_8
XANTENNA__137__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_32_123 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _130_/HI mem_right_track_8.LATCH_2_.latch/Q
+ mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__047__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_2_7 vgnd vpwr scs8hd_decap_6
XFILLER_11_56 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_101 vpwr vgnd scs8hd_fill_2
XFILLER_14_145 vgnd vpwr scs8hd_decap_8
XFILLER_14_178 vgnd vpwr scs8hd_decap_8
XFILLER_20_148 vgnd vpwr scs8hd_decap_4
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XFILLER_3_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_88 vgnd vpwr scs8hd_decap_4
XANTENNA__118__C _068_/C vgnd vpwr scs8hd_diode_2
XFILLER_8_13 vgnd vpwr scs8hd_fill_1
X_089_ _074_/A _089_/B _089_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_141 vgnd vpwr scs8hd_fill_1
XFILLER_6_152 vgnd vpwr scs8hd_fill_1
XFILLER_6_163 vpwr vgnd scs8hd_fill_2
X_158_ _158_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_26_3 vpwr vgnd scs8hd_fill_2
XANTENNA__150__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB _063_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__060__A _047_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_218 vgnd vpwr scs8hd_decap_12
XFILLER_17_77 vpwr vgnd scs8hd_fill_2
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_10 vgnd vpwr scs8hd_decap_4
XFILLER_3_199 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_210 vgnd vpwr scs8hd_decap_4
XANTENNA__145__A _145_/A vgnd vpwr scs8hd_diode_2
XANTENNA__055__A enable vgnd vpwr scs8hd_diode_2
XFILLER_21_232 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_8.LATCH_5_.latch data_in mem_right_track_8.LATCH_5_.latch/Q _069_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__115__D address[0] vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _041_/A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmem_top_track_2.LATCH_1_.latch data_in _041_/A _112_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_left_track_17.LATCH_1_.latch data_in mem_left_track_17.LATCH_1_.latch/Q _102_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_56 vgnd vpwr scs8hd_decap_8
XFILLER_29_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _129_/HI mem_right_track_16.LATCH_2_.latch/Q
+ mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_35_187 vgnd vpwr scs8hd_decap_12
XFILLER_26_110 vgnd vpwr scs8hd_decap_4
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_187 vpwr vgnd scs8hd_fill_2
XFILLER_25_99 vgnd vpwr scs8hd_decap_3
XFILLER_25_55 vgnd vpwr scs8hd_decap_4
XFILLER_25_22 vgnd vpwr scs8hd_decap_4
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_231 vpwr vgnd scs8hd_fill_2
XFILLER_17_132 vpwr vgnd scs8hd_fill_2
XANTENNA__153__A _153_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_146 vgnd vpwr scs8hd_decap_4
XFILLER_23_113 vpwr vgnd scs8hd_fill_2
XFILLER_31_190 vgnd vpwr scs8hd_fill_1
XANTENNA__063__A _063_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_79 vgnd vpwr scs8hd_decap_4
XFILLER_14_157 vpwr vgnd scs8hd_fill_2
XANTENNA__148__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_9_172 vpwr vgnd scs8hd_fill_2
XFILLER_9_194 vpwr vgnd scs8hd_fill_2
XFILLER_28_227 vgnd vpwr scs8hd_decap_6
XANTENNA__058__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_67 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
X_157_ chanx_left_in[5] chany_top_out[5] vgnd vpwr scs8hd_buf_2
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_120 vgnd vpwr scs8hd_decap_8
XFILLER_8_47 vgnd vpwr scs8hd_fill_1
XFILLER_8_69 vgnd vpwr scs8hd_decap_8
XFILLER_10_182 vpwr vgnd scs8hd_fill_2
X_088_ _073_/A _089_/B _088_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_208 vpwr vgnd scs8hd_fill_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_4
XFILLER_33_230 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__060__B address[2] vgnd vpwr scs8hd_diode_2
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_23 vpwr vgnd scs8hd_fill_2
XFILLER_33_77 vpwr vgnd scs8hd_fill_2
XFILLER_33_22 vgnd vpwr scs8hd_decap_4
Xmem_right_track_16.LATCH_0_.latch data_in mem_right_track_16.LATCH_0_.latch/Q _081_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _134_/HI _042_/Y mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__055__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _043_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__071__A _071_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_88 vgnd vpwr scs8hd_decap_4
XFILLER_0_159 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB _094_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_7 vgnd vpwr scs8hd_fill_1
XANTENNA__156__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__066__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_14_79 vgnd vpwr scs8hd_decap_8
XFILLER_29_174 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_199 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_2_16 vgnd vpwr scs8hd_decap_4
XFILLER_17_144 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.INVTX1_2_.scs8hd_inv_1 chany_top_in[6] mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _045_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_25 vpwr vgnd scs8hd_fill_2
XANTENNA__063__B _079_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_125 vgnd vpwr scs8hd_decap_3
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_184 vgnd vpwr scs8hd_decap_3
XFILLER_3_70 vpwr vgnd scs8hd_fill_2
XANTENNA__058__B _048_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__074__A _074_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_156_ chanx_left_in[4] chany_top_out[6] vgnd vpwr scs8hd_buf_2
X_087_ _079_/A _089_/B _087_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_6 vpwr vgnd scs8hd_fill_2
XANTENNA__159__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__069__A _069_/A vgnd vpwr scs8hd_diode_2
XANTENNA__060__C _112_/D vgnd vpwr scs8hd_diode_2
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_231 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _044_/Y mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_139_ chanx_right_in[4] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA__055__C _083_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _125_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_105 vpwr vgnd scs8hd_fill_2
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_0_138 vpwr vgnd scs8hd_fill_2
XANTENNA__071__B _073_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _134_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__066__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_14_36 vgnd vpwr scs8hd_decap_3
XANTENNA__082__A _082_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_153 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_4_230 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_156 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__077__A _077_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_123 vgnd vpwr scs8hd_decap_8
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_101 vpwr vgnd scs8hd_fill_2
XFILLER_32_115 vgnd vpwr scs8hd_decap_8
XFILLER_32_104 vgnd vpwr scs8hd_decap_8
XFILLER_17_156 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.INVTX1_5_.scs8hd_inv_1 right_bottom_grid_pin_11_ mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_181 vpwr vgnd scs8hd_fill_2
XFILLER_23_126 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_4_.latch data_in mem_top_track_0.LATCH_4_.latch/Q _107_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_37 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_3_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_115 vgnd vpwr scs8hd_decap_8
XFILLER_14_137 vpwr vgnd scs8hd_fill_2
XFILLER_13_192 vgnd vpwr scs8hd_fill_1
XFILLER_28_207 vgnd vpwr scs8hd_decap_6
XANTENNA__058__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__074__B _073_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_118 vgnd vpwr scs8hd_decap_4
XFILLER_22_36 vpwr vgnd scs8hd_fill_2
XFILLER_0_7 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_0_.latch data_in mem_left_track_9.LATCH_0_.latch/Q _096_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__090__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_19_207 vgnd vpwr scs8hd_decap_4
XFILLER_19_218 vpwr vgnd scs8hd_fill_2
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
X_155_ _155_/A chany_top_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_6_144 vgnd vpwr scs8hd_decap_8
XFILLER_12_80 vgnd vpwr scs8hd_decap_6
X_086_ _071_/A _089_/B _086_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_17_47 vpwr vgnd scs8hd_fill_2
XANTENNA__069__B _073_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_35 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__085__A _077_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_3_103 vpwr vgnd scs8hd_fill_2
XFILLER_3_158 vpwr vgnd scs8hd_fill_2
XFILLER_3_136 vgnd vpwr scs8hd_decap_4
Xmem_top_track_16.LATCH_1_.latch data_in mem_top_track_16.LATCH_1_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_069_ _069_/A _073_/B _069_/Y vgnd vpwr scs8hd_nor2_4
X_138_ chanx_right_in[5] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_24_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_68 vpwr vgnd scs8hd_fill_2
XFILLER_12_213 vgnd vpwr scs8hd_fill_1
XFILLER_5_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB _071_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__066__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_14_26 vpwr vgnd scs8hd_fill_2
XANTENNA__082__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_29_132 vpwr vgnd scs8hd_fill_2
XFILLER_20_91 vgnd vpwr scs8hd_fill_1
Xmem_left_track_1.LATCH_5_.latch data_in mem_left_track_1.LATCH_5_.latch/Q _084_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_3_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_168 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_60 vgnd vpwr scs8hd_decap_6
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_6_93 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _162_/A vgnd vpwr scs8hd_inv_1
XPHY_69 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_168 vgnd vpwr scs8hd_decap_8
XFILLER_26_157 vgnd vpwr scs8hd_decap_4
XANTENNA__077__B _077_/B vgnd vpwr scs8hd_diode_2
XFILLER_25_47 vpwr vgnd scs8hd_fill_2
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__093__A _071_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_127 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_31_160 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A _073_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_105 vgnd vpwr scs8hd_fill_1
XFILLER_9_142 vpwr vgnd scs8hd_fill_2
XFILLER_13_171 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_15_ mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[2] mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__090__B _112_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_154_ _154_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_6_167 vpwr vgnd scs8hd_fill_2
XFILLER_10_163 vgnd vpwr scs8hd_decap_3
XFILLER_10_174 vgnd vpwr scs8hd_decap_8
X_085_ _077_/A _089_/B _085_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_26_7 vpwr vgnd scs8hd_fill_2
XFILLER_33_222 vgnd vpwr scs8hd_decap_8
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_4_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_47 vgnd vpwr scs8hd_decap_12
XFILLER_33_14 vgnd vpwr scs8hd_fill_1
XANTENNA__085__B _089_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A right_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_8.LATCH_0_.latch data_in mem_right_track_8.LATCH_0_.latch/Q _074_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_137_ chanx_right_in[6] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
Xmux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_91 vpwr vgnd scs8hd_fill_2
XFILLER_2_181 vgnd vpwr scs8hd_decap_3
X_068_ _068_/A address[3] _068_/C _073_/B vgnd vpwr scs8hd_or3_4
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB _099_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _136_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A right_bottom_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__096__A _074_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_91 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_125 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _046_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _140_/A vgnd vpwr scs8hd_inv_1
XFILLER_6_50 vgnd vpwr scs8hd_fill_1
XPHY_59 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA__093__B _090_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_202 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_117 vgnd vpwr scs8hd_decap_3
Xmem_right_track_0.LATCH_5_.latch data_in mem_right_track_0.LATCH_5_.latch/Q _057_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_180 vgnd vpwr scs8hd_decap_8
XFILLER_31_194 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__088__B _089_/B vgnd vpwr scs8hd_diode_2
XFILLER_26_91 vgnd vpwr scs8hd_fill_1
Xmux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_176 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__090__C _083_/C vgnd vpwr scs8hd_diode_2
XANTENNA__099__A _077_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_231 vpwr vgnd scs8hd_fill_2
X_153_ _153_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_10_186 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _042_/A mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_10_197 vpwr vgnd scs8hd_fill_2
X_084_ _069_/A _089_/B _084_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_231 vpwr vgnd scs8hd_fill_2
XFILLER_19_7 vgnd vpwr scs8hd_fill_1
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 chanx_left_in[1] mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_201 vgnd vpwr scs8hd_decap_12
XFILLER_17_27 vgnd vpwr scs8hd_decap_4
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XFILLER_33_26 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _129_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_136_ _136_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_6 vgnd vpwr scs8hd_decap_4
X_067_ _063_/A _074_/A _067_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_63 vgnd vpwr scs8hd_fill_1
XFILLER_9_83 vgnd vpwr scs8hd_decap_4
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XANTENNA__096__B _090_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_219 vgnd vpwr scs8hd_decap_12
XFILLER_18_81 vpwr vgnd scs8hd_fill_2
XFILLER_34_91 vgnd vpwr scs8hd_fill_1
XFILLER_34_80 vgnd vpwr scs8hd_fill_1
X_119_ _069_/A _119_/B _119_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_29_178 vgnd vpwr scs8hd_decap_3
XFILLER_29_101 vpwr vgnd scs8hd_fill_2
XFILLER_4_211 vgnd vpwr scs8hd_decap_3
XFILLER_29_80 vpwr vgnd scs8hd_fill_2
XFILLER_20_93 vpwr vgnd scs8hd_fill_2
XFILLER_35_137 vgnd vpwr scs8hd_decap_12
XFILLER_29_91 vgnd vpwr scs8hd_decap_4
XFILLER_6_73 vpwr vgnd scs8hd_fill_2
XFILLER_6_84 vgnd vpwr scs8hd_decap_8
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_17_115 vgnd vpwr scs8hd_fill_1
XFILLER_15_82 vgnd vpwr scs8hd_decap_6
XFILLER_31_92 vpwr vgnd scs8hd_fill_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_6
XFILLER_31_173 vgnd vpwr scs8hd_decap_8
XFILLER_11_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _128_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _042_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_151 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_155 vpwr vgnd scs8hd_fill_2
XFILLER_13_184 vpwr vgnd scs8hd_fill_2
XFILLER_3_74 vgnd vpwr scs8hd_decap_3
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_17 vgnd vpwr scs8hd_decap_12
XANTENNA__090__D _083_/D vgnd vpwr scs8hd_diode_2
XANTENNA__099__B _102_/B vgnd vpwr scs8hd_diode_2
X_152_ chanx_left_in[0] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_6_103 vpwr vgnd scs8hd_fill_2
XFILLER_12_61 vgnd vpwr scs8hd_decap_8
X_083_ address[4] address[3] _083_/C _083_/D _089_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_18_210 vgnd vpwr scs8hd_decap_4
XFILLER_24_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_202 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_227 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_066_ address[1] address[2] address[0] _074_/A vgnd vpwr scs8hd_or3_4
X_135_ _135_/HI _135_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_0_53 vgnd vpwr scs8hd_decap_3
XFILLER_0_75 vpwr vgnd scs8hd_fill_2
XFILLER_9_62 vpwr vgnd scs8hd_fill_2
XFILLER_0_109 vpwr vgnd scs8hd_fill_2
XFILLER_28_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_93 vpwr vgnd scs8hd_fill_2
XFILLER_7_231 vpwr vgnd scs8hd_fill_2
X_049_ address[0] _112_/D vgnd vpwr scs8hd_inv_8
X_118_ address[4] address[3] _068_/C _119_/B vgnd vpwr scs8hd_or3_4
XFILLER_22_3 vgnd vpwr scs8hd_decap_3
XFILLER_14_18 vpwr vgnd scs8hd_fill_2
XFILLER_29_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_6_.scs8hd_inv_1 left_bottom_grid_pin_7_ mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_50 vgnd vpwr scs8hd_decap_6
XFILLER_20_72 vgnd vpwr scs8hd_decap_4
XFILLER_35_149 vgnd vpwr scs8hd_decap_6
XFILLER_6_41 vgnd vpwr scs8hd_decap_3
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_25_28 vpwr vgnd scs8hd_fill_2
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_1_215 vpwr vgnd scs8hd_fill_2
XFILLER_9_7 vgnd vpwr scs8hd_decap_3
Xmux_right_track_0.INVTX1_2_.scs8hd_inv_1 chany_top_in[8] mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_25_193 vpwr vgnd scs8hd_fill_2
XFILLER_25_182 vgnd vpwr scs8hd_fill_1
XFILLER_17_105 vpwr vgnd scs8hd_fill_2
XFILLER_31_71 vpwr vgnd scs8hd_fill_2
XFILLER_31_82 vgnd vpwr scs8hd_fill_1
Xmem_left_track_17.LATCH_2_.latch data_in mem_left_track_17.LATCH_2_.latch/Q _101_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_163 vgnd vpwr scs8hd_fill_1
XFILLER_26_93 vgnd vpwr scs8hd_decap_4
XFILLER_9_134 vpwr vgnd scs8hd_fill_2
XFILLER_3_86 vpwr vgnd scs8hd_fill_2
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
XFILLER_3_20 vgnd vpwr scs8hd_fill_1
XFILLER_22_29 vpwr vgnd scs8hd_fill_2
XFILLER_6_137 vgnd vpwr scs8hd_decap_4
X_082_ _082_/A address[5] _083_/D vgnd vpwr scs8hd_or2_4
XFILLER_10_133 vgnd vpwr scs8hd_fill_1
X_151_ chanx_left_in[1] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_33_214 vgnd vpwr scs8hd_fill_1
XFILLER_3_107 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _125_/HI mem_left_track_1.LATCH_2_.latch/Q
+ mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_214 vgnd vpwr scs8hd_fill_1
Xmux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _041_/Y mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[5] mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_065_ _063_/A _073_/A _065_/Y vgnd vpwr scs8hd_nor2_4
X_134_ _134_/HI _134_/LO vgnd vpwr scs8hd_conb_1
XFILLER_17_6 vpwr vgnd scs8hd_fill_2
XFILLER_0_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _074_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_93 vgnd vpwr scs8hd_decap_6
X_117_ _068_/A _112_/B _112_/C address[0] _117_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_048_ address[2] _048_/Y vgnd vpwr scs8hd_inv_8
Xmem_left_track_1.LATCH_0_.latch data_in mem_left_track_1.LATCH_0_.latch/Q _089_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_18 vgnd vpwr scs8hd_decap_12
XFILLER_29_136 vpwr vgnd scs8hd_fill_2
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB _086_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_106 vgnd vpwr scs8hd_decap_12
XFILLER_29_71 vgnd vpwr scs8hd_decap_3
Xmem_right_track_16.LATCH_1_.latch data_in mem_right_track_16.LATCH_1_.latch/Q _080_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_106 vpwr vgnd scs8hd_fill_2
XFILLER_25_18 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_19_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_25_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB _078_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__102__A _073_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_109 vpwr vgnd scs8hd_fill_2
XFILLER_31_164 vpwr vgnd scs8hd_fill_2
XFILLER_31_153 vgnd vpwr scs8hd_fill_1
XFILLER_31_131 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[6] mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_175 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.INVTX1_3_.scs8hd_inv_1 right_bottom_grid_pin_3_ mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_83 vpwr vgnd scs8hd_fill_2
XFILLER_13_175 vgnd vpwr scs8hd_decap_6
XFILLER_3_32 vpwr vgnd scs8hd_fill_2
XFILLER_27_223 vgnd vpwr scs8hd_decap_8
XFILLER_10_112 vpwr vgnd scs8hd_fill_2
X_150_ chanx_left_in[2] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_081_ _074_/A _077_/B _081_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_145 vgnd vpwr scs8hd_decap_6
XFILLER_12_41 vgnd vpwr scs8hd_decap_3
XFILLER_33_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _102_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_95 vpwr vgnd scs8hd_fill_2
XFILLER_23_62 vgnd vpwr scs8hd_decap_3
X_133_ _133_/HI _133_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _045_/Y vgnd vpwr
+ scs8hd_diode_2
X_064_ address[1] address[2] _112_/D _073_/A vgnd vpwr scs8hd_or3_4
XFILLER_2_141 vgnd vpwr scs8hd_decap_4
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_11 vgnd vpwr scs8hd_decap_8
XANTENNA__110__A _073_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_42 vpwr vgnd scs8hd_fill_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XFILLER_12_218 vgnd vpwr scs8hd_decap_12
XFILLER_34_83 vgnd vpwr scs8hd_decap_8
XANTENNA__105__A address[4] vgnd vpwr scs8hd_diode_2
X_116_ _068_/A _112_/B _112_/C _112_/D _116_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mem_right_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_047_ address[1] _047_/Y vgnd vpwr scs8hd_inv_8
XFILLER_20_30 vgnd vpwr scs8hd_fill_1
XFILLER_35_118 vgnd vpwr scs8hd_decap_6
XFILLER_29_50 vgnd vpwr scs8hd_decap_4
XFILLER_34_140 vgnd vpwr scs8hd_decap_12
XPHY_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_0_.latch data_in mem_right_track_0.LATCH_0_.latch/Q _067_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_top_track_8.LATCH_0_.latch data_in _044_/A _115_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_30 vpwr vgnd scs8hd_fill_2
XANTENNA__102__B _102_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_198 vgnd vpwr scs8hd_decap_12
XFILLER_31_121 vgnd vpwr scs8hd_fill_1
XFILLER_22_121 vpwr vgnd scs8hd_fill_2
XFILLER_22_154 vgnd vpwr scs8hd_decap_3
XFILLER_22_187 vgnd vpwr scs8hd_decap_12
XFILLER_7_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_103 vpwr vgnd scs8hd_fill_2
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_132 vpwr vgnd scs8hd_fill_2
XFILLER_13_154 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_3_66 vpwr vgnd scs8hd_fill_2
X_080_ _073_/A _077_/B _080_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_168 vgnd vpwr scs8hd_decap_3
XFILLER_5_3 vgnd vpwr scs8hd_decap_6
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _153_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__108__A _071_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_161 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_132_ _132_/HI _132_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_74 vgnd vpwr scs8hd_decap_3
Xmem_top_track_0.LATCH_5_.latch data_in mem_top_track_0.LATCH_5_.latch/Q _106_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_063_ _063_/A _079_/A _063_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_186 vgnd vpwr scs8hd_decap_3
XFILLER_2_120 vgnd vpwr scs8hd_decap_3
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_45 vpwr vgnd scs8hd_fill_2
XANTENNA__110__B _105_/X vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _145_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XFILLER_21_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_18_30 vgnd vpwr scs8hd_fill_1
XFILLER_18_85 vgnd vpwr scs8hd_decap_6
X_046_ _046_/A _046_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_223 vgnd vpwr scs8hd_decap_8
XANTENNA__105__B address[3] vgnd vpwr scs8hd_diode_2
X_115_ _068_/A address[3] _112_/C address[0] _115_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__121__A _071_/A vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_1_.latch data_in mem_left_track_9.LATCH_1_.latch/Q _095_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A left_bottom_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB _059_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _041_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_42 vpwr vgnd scs8hd_fill_2
XFILLER_29_40 vgnd vpwr scs8hd_decap_4
XFILLER_20_97 vgnd vpwr scs8hd_decap_4
XANTENNA__116__A _068_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_11 vgnd vpwr scs8hd_decap_3
XFILLER_6_66 vgnd vpwr scs8hd_fill_1
Xmem_top_track_16.LATCH_2_.latch data_in mem_top_track_16.LATCH_2_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_34_152 vgnd vpwr scs8hd_fill_1
XFILLER_19_182 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_4_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_174 vpwr vgnd scs8hd_fill_2
XFILLER_25_152 vpwr vgnd scs8hd_fill_2
XFILLER_31_96 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_141 vgnd vpwr scs8hd_decap_6
XFILLER_16_163 vgnd vpwr scs8hd_decap_3
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
.ends

