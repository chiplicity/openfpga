magic
tech sky130A
magscale 1 2
timestamp 1607686528
<< obsli1 >>
rect 354 2159 10106 11441
<< obsm1 >>
rect 0 2128 10460 11472
<< metal2 >>
rect 4 0 60 800
rect 1476 0 1532 800
rect 2948 0 3004 800
rect 4420 0 4476 800
rect 5984 0 6040 800
rect 7456 0 7512 800
rect 8928 0 8984 800
rect 10400 0 10456 800
<< obsm2 >>
rect 6 856 10454 11472
rect 116 800 1420 856
rect 1588 800 2892 856
rect 3060 800 4364 856
rect 4532 800 5928 856
rect 6096 800 7400 856
rect 7568 800 8872 856
rect 9040 800 10344 856
<< obsm3 >>
rect 1826 2143 8674 11457
<< metal4 >>
rect 1826 2128 2146 11472
rect 3458 2128 3778 11472
<< obsm4 >>
rect 5090 2128 8674 11472
<< labels >>
rlabel metal2 s 4 0 60 800 6 x[0]
port 1 nsew default output
rlabel metal2 s 1476 0 1532 800 6 x[1]
port 2 nsew default output
rlabel metal2 s 2948 0 3004 800 6 x[2]
port 3 nsew default output
rlabel metal2 s 4420 0 4476 800 6 x[3]
port 4 nsew default output
rlabel metal2 s 5984 0 6040 800 6 x[4]
port 5 nsew default output
rlabel metal2 s 7456 0 7512 800 6 x[5]
port 6 nsew default output
rlabel metal2 s 8928 0 8984 800 6 x[6]
port 7 nsew default output
rlabel metal2 s 10400 0 10456 800 6 x[7]
port 8 nsew default output
rlabel metal4 s 1826 2128 2146 11472 6 VPWR
port 9 nsew power input
rlabel metal4 s 3458 2128 3778 11472 6 VGND
port 10 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 10460 11472
string LEFview TRUE
<< end >>
