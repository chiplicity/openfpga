magic
tech sky130A
magscale 1 2
timestamp 1608156304
<< obsli1 >>
rect 1104 2159 21620 20145
<< obsm1 >>
rect 198 1368 22526 20176
<< metal2 >>
rect 5722 22000 5778 22800
rect 17130 22000 17186 22800
rect 202 0 258 800
rect 662 0 718 800
rect 1214 0 1270 800
rect 1766 0 1822 800
rect 2318 0 2374 800
rect 2870 0 2926 800
rect 3422 0 3478 800
rect 3974 0 4030 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5630 0 5686 800
rect 6090 0 6146 800
rect 6642 0 6698 800
rect 7194 0 7250 800
rect 7746 0 7802 800
rect 8298 0 8354 800
rect 8850 0 8906 800
rect 9402 0 9458 800
rect 9954 0 10010 800
rect 10506 0 10562 800
rect 11058 0 11114 800
rect 11610 0 11666 800
rect 12070 0 12126 800
rect 12622 0 12678 800
rect 13174 0 13230 800
rect 13726 0 13782 800
rect 14278 0 14334 800
rect 14830 0 14886 800
rect 15382 0 15438 800
rect 15934 0 15990 800
rect 16486 0 16542 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 18050 0 18106 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21914 0 21970 800
rect 22466 0 22522 800
<< obsm2 >>
rect 204 21944 5666 22545
rect 5834 21944 17074 22545
rect 17242 21944 22520 22545
rect 204 856 22520 21944
rect 314 167 606 856
rect 774 167 1158 856
rect 1326 167 1710 856
rect 1878 167 2262 856
rect 2430 167 2814 856
rect 2982 167 3366 856
rect 3534 167 3918 856
rect 4086 167 4470 856
rect 4638 167 5022 856
rect 5190 167 5574 856
rect 5742 167 6034 856
rect 6202 167 6586 856
rect 6754 167 7138 856
rect 7306 167 7690 856
rect 7858 167 8242 856
rect 8410 167 8794 856
rect 8962 167 9346 856
rect 9514 167 9898 856
rect 10066 167 10450 856
rect 10618 167 11002 856
rect 11170 167 11554 856
rect 11722 167 12014 856
rect 12182 167 12566 856
rect 12734 167 13118 856
rect 13286 167 13670 856
rect 13838 167 14222 856
rect 14390 167 14774 856
rect 14942 167 15326 856
rect 15494 167 15878 856
rect 16046 167 16430 856
rect 16598 167 16982 856
rect 17150 167 17442 856
rect 17610 167 17994 856
rect 18162 167 18546 856
rect 18714 167 19098 856
rect 19266 167 19650 856
rect 19818 167 20202 856
rect 20370 167 20754 856
rect 20922 167 21306 856
rect 21474 167 21858 856
rect 22026 167 22410 856
<< metal3 >>
rect 22000 22448 22800 22568
rect 22000 22040 22800 22160
rect 22000 21496 22800 21616
rect 22000 21088 22800 21208
rect 22000 20680 22800 20800
rect 22000 20136 22800 20256
rect 22000 19728 22800 19848
rect 22000 19320 22800 19440
rect 22000 18776 22800 18896
rect 22000 18368 22800 18488
rect 22000 17960 22800 18080
rect 22000 17416 22800 17536
rect 22000 17008 22800 17128
rect 22000 16464 22800 16584
rect 22000 16056 22800 16176
rect 22000 15648 22800 15768
rect 22000 15104 22800 15224
rect 22000 14696 22800 14816
rect 22000 14288 22800 14408
rect 22000 13744 22800 13864
rect 22000 13336 22800 13456
rect 22000 12928 22800 13048
rect 22000 12384 22800 12504
rect 22000 11976 22800 12096
rect 0 11432 800 11552
rect 22000 11568 22800 11688
rect 22000 11024 22800 11144
rect 22000 10616 22800 10736
rect 22000 10072 22800 10192
rect 22000 9664 22800 9784
rect 22000 9256 22800 9376
rect 22000 8712 22800 8832
rect 22000 8304 22800 8424
rect 22000 7896 22800 8016
rect 22000 7352 22800 7472
rect 22000 6944 22800 7064
rect 22000 6536 22800 6656
rect 22000 5992 22800 6112
rect 22000 5584 22800 5704
rect 22000 5040 22800 5160
rect 22000 4632 22800 4752
rect 22000 4224 22800 4344
rect 22000 3680 22800 3800
rect 22000 3272 22800 3392
rect 22000 2864 22800 2984
rect 22000 2320 22800 2440
rect 22000 1912 22800 2032
rect 22000 1504 22800 1624
rect 22000 960 22800 1080
rect 22000 552 22800 672
rect 22000 144 22800 264
<< obsm3 >>
rect 800 22368 21920 22541
rect 800 22240 22000 22368
rect 800 21960 21920 22240
rect 800 21696 22000 21960
rect 800 21416 21920 21696
rect 800 21288 22000 21416
rect 800 21008 21920 21288
rect 800 20880 22000 21008
rect 800 20600 21920 20880
rect 800 20336 22000 20600
rect 800 20056 21920 20336
rect 800 19928 22000 20056
rect 800 19648 21920 19928
rect 800 19520 22000 19648
rect 800 19240 21920 19520
rect 800 18976 22000 19240
rect 800 18696 21920 18976
rect 800 18568 22000 18696
rect 800 18288 21920 18568
rect 800 18160 22000 18288
rect 800 17880 21920 18160
rect 800 17616 22000 17880
rect 800 17336 21920 17616
rect 800 17208 22000 17336
rect 800 16928 21920 17208
rect 800 16664 22000 16928
rect 800 16384 21920 16664
rect 800 16256 22000 16384
rect 800 15976 21920 16256
rect 800 15848 22000 15976
rect 800 15568 21920 15848
rect 800 15304 22000 15568
rect 800 15024 21920 15304
rect 800 14896 22000 15024
rect 800 14616 21920 14896
rect 800 14488 22000 14616
rect 800 14208 21920 14488
rect 800 13944 22000 14208
rect 800 13664 21920 13944
rect 800 13536 22000 13664
rect 800 13256 21920 13536
rect 800 13128 22000 13256
rect 800 12848 21920 13128
rect 800 12584 22000 12848
rect 800 12304 21920 12584
rect 800 12176 22000 12304
rect 800 11896 21920 12176
rect 800 11768 22000 11896
rect 800 11632 21920 11768
rect 880 11488 21920 11632
rect 880 11352 22000 11488
rect 800 11224 22000 11352
rect 800 10944 21920 11224
rect 800 10816 22000 10944
rect 800 10536 21920 10816
rect 800 10272 22000 10536
rect 800 9992 21920 10272
rect 800 9864 22000 9992
rect 800 9584 21920 9864
rect 800 9456 22000 9584
rect 800 9176 21920 9456
rect 800 8912 22000 9176
rect 800 8632 21920 8912
rect 800 8504 22000 8632
rect 800 8224 21920 8504
rect 800 8096 22000 8224
rect 800 7816 21920 8096
rect 800 7552 22000 7816
rect 800 7272 21920 7552
rect 800 7144 22000 7272
rect 800 6864 21920 7144
rect 800 6736 22000 6864
rect 800 6456 21920 6736
rect 800 6192 22000 6456
rect 800 5912 21920 6192
rect 800 5784 22000 5912
rect 800 5504 21920 5784
rect 800 5240 22000 5504
rect 800 4960 21920 5240
rect 800 4832 22000 4960
rect 800 4552 21920 4832
rect 800 4424 22000 4552
rect 800 4144 21920 4424
rect 800 3880 22000 4144
rect 800 3600 21920 3880
rect 800 3472 22000 3600
rect 800 3192 21920 3472
rect 800 3064 22000 3192
rect 800 2784 21920 3064
rect 800 2520 22000 2784
rect 800 2240 21920 2520
rect 800 2112 22000 2240
rect 800 1832 21920 2112
rect 800 1704 22000 1832
rect 800 1424 21920 1704
rect 800 1160 22000 1424
rect 800 880 21920 1160
rect 800 752 22000 880
rect 800 472 21920 752
rect 800 344 22000 472
rect 800 171 21920 344
<< metal4 >>
rect 4376 2128 4696 20176
rect 7808 2128 8128 20176
<< obsm4 >>
rect 11240 2128 18424 20176
<< labels >>
rlabel metal2 s 5722 22000 5778 22800 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 22466 0 22522 800 6 SC_OUT_BOT
port 2 nsew default output
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_1_
port 3 nsew default input
rlabel metal2 s 17130 22000 17186 22800 6 ccff_head
port 4 nsew default input
rlabel metal3 s 0 11432 800 11552 6 ccff_tail
port 5 nsew default output
rlabel metal3 s 22000 3680 22800 3800 6 chanx_right_in[0]
port 6 nsew default input
rlabel metal3 s 22000 8304 22800 8424 6 chanx_right_in[10]
port 7 nsew default input
rlabel metal3 s 22000 8712 22800 8832 6 chanx_right_in[11]
port 8 nsew default input
rlabel metal3 s 22000 9256 22800 9376 6 chanx_right_in[12]
port 9 nsew default input
rlabel metal3 s 22000 9664 22800 9784 6 chanx_right_in[13]
port 10 nsew default input
rlabel metal3 s 22000 10072 22800 10192 6 chanx_right_in[14]
port 11 nsew default input
rlabel metal3 s 22000 10616 22800 10736 6 chanx_right_in[15]
port 12 nsew default input
rlabel metal3 s 22000 11024 22800 11144 6 chanx_right_in[16]
port 13 nsew default input
rlabel metal3 s 22000 11568 22800 11688 6 chanx_right_in[17]
port 14 nsew default input
rlabel metal3 s 22000 11976 22800 12096 6 chanx_right_in[18]
port 15 nsew default input
rlabel metal3 s 22000 12384 22800 12504 6 chanx_right_in[19]
port 16 nsew default input
rlabel metal3 s 22000 4224 22800 4344 6 chanx_right_in[1]
port 17 nsew default input
rlabel metal3 s 22000 4632 22800 4752 6 chanx_right_in[2]
port 18 nsew default input
rlabel metal3 s 22000 5040 22800 5160 6 chanx_right_in[3]
port 19 nsew default input
rlabel metal3 s 22000 5584 22800 5704 6 chanx_right_in[4]
port 20 nsew default input
rlabel metal3 s 22000 5992 22800 6112 6 chanx_right_in[5]
port 21 nsew default input
rlabel metal3 s 22000 6536 22800 6656 6 chanx_right_in[6]
port 22 nsew default input
rlabel metal3 s 22000 6944 22800 7064 6 chanx_right_in[7]
port 23 nsew default input
rlabel metal3 s 22000 7352 22800 7472 6 chanx_right_in[8]
port 24 nsew default input
rlabel metal3 s 22000 7896 22800 8016 6 chanx_right_in[9]
port 25 nsew default input
rlabel metal3 s 22000 12928 22800 13048 6 chanx_right_out[0]
port 26 nsew default output
rlabel metal3 s 22000 17416 22800 17536 6 chanx_right_out[10]
port 27 nsew default output
rlabel metal3 s 22000 17960 22800 18080 6 chanx_right_out[11]
port 28 nsew default output
rlabel metal3 s 22000 18368 22800 18488 6 chanx_right_out[12]
port 29 nsew default output
rlabel metal3 s 22000 18776 22800 18896 6 chanx_right_out[13]
port 30 nsew default output
rlabel metal3 s 22000 19320 22800 19440 6 chanx_right_out[14]
port 31 nsew default output
rlabel metal3 s 22000 19728 22800 19848 6 chanx_right_out[15]
port 32 nsew default output
rlabel metal3 s 22000 20136 22800 20256 6 chanx_right_out[16]
port 33 nsew default output
rlabel metal3 s 22000 20680 22800 20800 6 chanx_right_out[17]
port 34 nsew default output
rlabel metal3 s 22000 21088 22800 21208 6 chanx_right_out[18]
port 35 nsew default output
rlabel metal3 s 22000 21496 22800 21616 6 chanx_right_out[19]
port 36 nsew default output
rlabel metal3 s 22000 13336 22800 13456 6 chanx_right_out[1]
port 37 nsew default output
rlabel metal3 s 22000 13744 22800 13864 6 chanx_right_out[2]
port 38 nsew default output
rlabel metal3 s 22000 14288 22800 14408 6 chanx_right_out[3]
port 39 nsew default output
rlabel metal3 s 22000 14696 22800 14816 6 chanx_right_out[4]
port 40 nsew default output
rlabel metal3 s 22000 15104 22800 15224 6 chanx_right_out[5]
port 41 nsew default output
rlabel metal3 s 22000 15648 22800 15768 6 chanx_right_out[6]
port 42 nsew default output
rlabel metal3 s 22000 16056 22800 16176 6 chanx_right_out[7]
port 43 nsew default output
rlabel metal3 s 22000 16464 22800 16584 6 chanx_right_out[8]
port 44 nsew default output
rlabel metal3 s 22000 17008 22800 17128 6 chanx_right_out[9]
port 45 nsew default output
rlabel metal2 s 662 0 718 800 6 chany_bottom_in[0]
port 46 nsew default input
rlabel metal2 s 6090 0 6146 800 6 chany_bottom_in[10]
port 47 nsew default input
rlabel metal2 s 6642 0 6698 800 6 chany_bottom_in[11]
port 48 nsew default input
rlabel metal2 s 7194 0 7250 800 6 chany_bottom_in[12]
port 49 nsew default input
rlabel metal2 s 7746 0 7802 800 6 chany_bottom_in[13]
port 50 nsew default input
rlabel metal2 s 8298 0 8354 800 6 chany_bottom_in[14]
port 51 nsew default input
rlabel metal2 s 8850 0 8906 800 6 chany_bottom_in[15]
port 52 nsew default input
rlabel metal2 s 9402 0 9458 800 6 chany_bottom_in[16]
port 53 nsew default input
rlabel metal2 s 9954 0 10010 800 6 chany_bottom_in[17]
port 54 nsew default input
rlabel metal2 s 10506 0 10562 800 6 chany_bottom_in[18]
port 55 nsew default input
rlabel metal2 s 11058 0 11114 800 6 chany_bottom_in[19]
port 56 nsew default input
rlabel metal2 s 1214 0 1270 800 6 chany_bottom_in[1]
port 57 nsew default input
rlabel metal2 s 1766 0 1822 800 6 chany_bottom_in[2]
port 58 nsew default input
rlabel metal2 s 2318 0 2374 800 6 chany_bottom_in[3]
port 59 nsew default input
rlabel metal2 s 2870 0 2926 800 6 chany_bottom_in[4]
port 60 nsew default input
rlabel metal2 s 3422 0 3478 800 6 chany_bottom_in[5]
port 61 nsew default input
rlabel metal2 s 3974 0 4030 800 6 chany_bottom_in[6]
port 62 nsew default input
rlabel metal2 s 4526 0 4582 800 6 chany_bottom_in[7]
port 63 nsew default input
rlabel metal2 s 5078 0 5134 800 6 chany_bottom_in[8]
port 64 nsew default input
rlabel metal2 s 5630 0 5686 800 6 chany_bottom_in[9]
port 65 nsew default input
rlabel metal2 s 11610 0 11666 800 6 chany_bottom_out[0]
port 66 nsew default output
rlabel metal2 s 17038 0 17094 800 6 chany_bottom_out[10]
port 67 nsew default output
rlabel metal2 s 17498 0 17554 800 6 chany_bottom_out[11]
port 68 nsew default output
rlabel metal2 s 18050 0 18106 800 6 chany_bottom_out[12]
port 69 nsew default output
rlabel metal2 s 18602 0 18658 800 6 chany_bottom_out[13]
port 70 nsew default output
rlabel metal2 s 19154 0 19210 800 6 chany_bottom_out[14]
port 71 nsew default output
rlabel metal2 s 19706 0 19762 800 6 chany_bottom_out[15]
port 72 nsew default output
rlabel metal2 s 20258 0 20314 800 6 chany_bottom_out[16]
port 73 nsew default output
rlabel metal2 s 20810 0 20866 800 6 chany_bottom_out[17]
port 74 nsew default output
rlabel metal2 s 21362 0 21418 800 6 chany_bottom_out[18]
port 75 nsew default output
rlabel metal2 s 21914 0 21970 800 6 chany_bottom_out[19]
port 76 nsew default output
rlabel metal2 s 12070 0 12126 800 6 chany_bottom_out[1]
port 77 nsew default output
rlabel metal2 s 12622 0 12678 800 6 chany_bottom_out[2]
port 78 nsew default output
rlabel metal2 s 13174 0 13230 800 6 chany_bottom_out[3]
port 79 nsew default output
rlabel metal2 s 13726 0 13782 800 6 chany_bottom_out[4]
port 80 nsew default output
rlabel metal2 s 14278 0 14334 800 6 chany_bottom_out[5]
port 81 nsew default output
rlabel metal2 s 14830 0 14886 800 6 chany_bottom_out[6]
port 82 nsew default output
rlabel metal2 s 15382 0 15438 800 6 chany_bottom_out[7]
port 83 nsew default output
rlabel metal2 s 15934 0 15990 800 6 chany_bottom_out[8]
port 84 nsew default output
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_out[9]
port 85 nsew default output
rlabel metal3 s 22000 22040 22800 22160 6 prog_clk_0_E_in
port 86 nsew default input
rlabel metal3 s 22000 144 22800 264 6 right_bottom_grid_pin_34_
port 87 nsew default input
rlabel metal3 s 22000 552 22800 672 6 right_bottom_grid_pin_35_
port 88 nsew default input
rlabel metal3 s 22000 960 22800 1080 6 right_bottom_grid_pin_36_
port 89 nsew default input
rlabel metal3 s 22000 1504 22800 1624 6 right_bottom_grid_pin_37_
port 90 nsew default input
rlabel metal3 s 22000 1912 22800 2032 6 right_bottom_grid_pin_38_
port 91 nsew default input
rlabel metal3 s 22000 2320 22800 2440 6 right_bottom_grid_pin_39_
port 92 nsew default input
rlabel metal3 s 22000 2864 22800 2984 6 right_bottom_grid_pin_40_
port 93 nsew default input
rlabel metal3 s 22000 3272 22800 3392 6 right_bottom_grid_pin_41_
port 94 nsew default input
rlabel metal3 s 22000 22448 22800 22568 6 right_top_grid_pin_1_
port 95 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 96 nsew power input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 97 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 22800 22800
string LEFview TRUE
<< end >>
