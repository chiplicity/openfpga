* NGSPICE file created from sb_1__3_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

.subckt sb_1__3_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_left_grid_pin_13_ bottom_right_grid_pin_11_ chanx_left_in[0] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chanx_right_in[0] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chany_bottom_in[0]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_out[0] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] data_in enable left_bottom_grid_pin_12_
+ left_top_grid_pin_11_ left_top_grid_pin_13_ left_top_grid_pin_15_ left_top_grid_pin_1_
+ left_top_grid_pin_3_ left_top_grid_pin_5_ left_top_grid_pin_7_ left_top_grid_pin_9_
+ right_bottom_grid_pin_12_ right_top_grid_pin_11_ right_top_grid_pin_13_ right_top_grid_pin_15_
+ right_top_grid_pin_1_ right_top_grid_pin_3_ right_top_grid_pin_5_ right_top_grid_pin_7_
+ right_top_grid_pin_9_ vpwr vgnd
XFILLER_7_7 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_63 vgnd vpwr scs8hd_decap_6
XFILLER_26_52 vgnd vpwr scs8hd_decap_8
XFILLER_26_30 vgnd vpwr scs8hd_fill_1
XFILLER_13_100 vgnd vpwr scs8hd_decap_3
XFILLER_13_144 vpwr vgnd scs8hd_fill_2
XFILLER_13_188 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_34 vpwr vgnd scs8hd_fill_2
XFILLER_27_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_118 vgnd vpwr scs8hd_decap_4
XFILLER_10_136 vgnd vpwr scs8hd_decap_6
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XANTENNA__108__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__124__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_5_173 vgnd vpwr scs8hd_decap_4
XFILLER_5_184 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_3_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_200_ _200_/A _200_/Y vgnd vpwr scs8hd_inv_8
X_131_ _120_/A _129_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__119__A _130_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _242_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ _188_/Y mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__105__C _105_/C vgnd vpwr scs8hd_diode_2
X_114_ _114_/A address[4] _125_/C _114_/X vgnd vpwr scs8hd_or3_4
XFILLER_38_117 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[3] mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__121__B _120_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_right_track_16.LATCH_4_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_117 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_65 vgnd vpwr scs8hd_decap_8
XFILLER_20_32 vgnd vpwr scs8hd_decap_8
XANTENNA__222__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_28_172 vgnd vpwr scs8hd_decap_12
XFILLER_28_150 vgnd vpwr scs8hd_decap_3
XANTENNA__116__B _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_23 vpwr vgnd scs8hd_fill_2
XANTENNA__132__A _121_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_56 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
Xmem_right_track_8.LATCH_1_.latch data_in mem_right_track_8.LATCH_1_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_25_175 vpwr vgnd scs8hd_fill_2
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XFILLER_15_54 vpwr vgnd scs8hd_fill_2
XFILLER_15_65 vpwr vgnd scs8hd_fill_2
XFILLER_15_87 vpwr vgnd scs8hd_fill_2
XFILLER_31_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _202_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XANTENNA__127__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_167 vpwr vgnd scs8hd_fill_2
XFILLER_22_123 vpwr vgnd scs8hd_fill_2
XFILLER_13_123 vgnd vpwr scs8hd_fill_1
XFILLER_13_156 vpwr vgnd scs8hd_fill_2
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_5_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_8_182 vgnd vpwr scs8hd_decap_4
XFILLER_8_193 vpwr vgnd scs8hd_fill_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_12_22 vpwr vgnd scs8hd_fill_2
XANTENNA__230__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_215 vgnd vpwr scs8hd_decap_3
XFILLER_26_270 vgnd vpwr scs8hd_decap_4
XANTENNA__108__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _130_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB _184_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _188_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_24_229 vgnd vpwr scs8hd_decap_12
XFILLER_24_218 vgnd vpwr scs8hd_decap_8
XFILLER_17_270 vgnd vpwr scs8hd_decap_6
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[3] mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_130_ _130_/A _129_/B _130_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__225__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__119__B _120_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_58 vgnd vpwr scs8hd_decap_4
XANTENNA__135__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_9_23 vpwr vgnd scs8hd_fill_2
XFILLER_20_232 vgnd vpwr scs8hd_fill_1
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _204_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_21 vgnd vpwr scs8hd_decap_6
X_113_ address[3] _114_/A vgnd vpwr scs8hd_inv_8
XFILLER_7_236 vgnd vpwr scs8hd_decap_6
XFILLER_11_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_129 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.INVTX1_6_.scs8hd_inv_1 left_top_grid_pin_7_ mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XFILLER_4_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_184 vgnd vpwr scs8hd_decap_12
XANTENNA__116__C _116_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_13 vgnd vpwr scs8hd_fill_1
XANTENNA__132__B _129_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_68 vgnd vpwr scs8hd_decap_4
XFILLER_19_184 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB _181_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_187 vpwr vgnd scs8hd_fill_2
XFILLER_25_143 vgnd vpwr scs8hd_decap_4
XFILLER_25_132 vpwr vgnd scs8hd_fill_2
XFILLER_15_33 vpwr vgnd scs8hd_fill_2
XFILLER_31_21 vgnd vpwr scs8hd_decap_12
XFILLER_31_10 vpwr vgnd scs8hd_fill_2
XANTENNA__233__A _233_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_98 vgnd vpwr scs8hd_decap_12
XFILLER_0_231 vgnd vpwr scs8hd_decap_3
XFILLER_16_110 vgnd vpwr scs8hd_decap_8
XFILLER_31_135 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 chanx_right_in[6] mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__127__B address[5] vgnd vpwr scs8hd_diode_2
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _190_/A vgnd
+ vpwr scs8hd_diode_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_154 vpwr vgnd scs8hd_fill_2
XFILLER_16_165 vgnd vpwr scs8hd_decap_8
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_5_ mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_102 vpwr vgnd scs8hd_fill_2
XFILLER_30_190 vgnd vpwr scs8hd_decap_12
XFILLER_22_179 vgnd vpwr scs8hd_decap_4
XFILLER_22_146 vgnd vpwr scs8hd_fill_1
XANTENNA__228__A _228_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _238_/A vgnd vpwr scs8hd_inv_1
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A _137_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_161 vpwr vgnd scs8hd_fill_2
XFILLER_27_249 vgnd vpwr scs8hd_decap_6
XFILLER_12_56 vgnd vpwr scs8hd_decap_6
XFILLER_12_67 vgnd vpwr scs8hd_decap_6
XFILLER_12_89 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XFILLER_18_227 vgnd vpwr scs8hd_decap_12
XFILLER_5_153 vgnd vpwr scs8hd_fill_1
XANTENNA__140__B _138_/X vgnd vpwr scs8hd_diode_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[4] mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_263 vgnd vpwr scs8hd_decap_12
XFILLER_23_66 vgnd vpwr scs8hd_fill_1
XFILLER_23_22 vpwr vgnd scs8hd_fill_2
XFILLER_23_99 vpwr vgnd scs8hd_fill_2
XANTENNA__241__A _241_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _188_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_230 vgnd vpwr scs8hd_decap_3
XFILLER_14_252 vpwr vgnd scs8hd_fill_2
XFILLER_14_263 vgnd vpwr scs8hd_decap_12
XFILLER_9_46 vpwr vgnd scs8hd_fill_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XFILLER_9_79 vgnd vpwr scs8hd_decap_6
X_189_ _189_/A _189_/Y vgnd vpwr scs8hd_inv_8
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA__151__A _122_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A right_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_11 vgnd vpwr scs8hd_fill_1
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XFILLER_18_88 vgnd vpwr scs8hd_decap_4
X_112_ address[5] _162_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_259 vpwr vgnd scs8hd_fill_2
XFILLER_11_233 vpwr vgnd scs8hd_fill_2
XANTENNA__236__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_22_9 vgnd vpwr scs8hd_decap_3
XANTENNA__146__A _146_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
XFILLER_29_10 vpwr vgnd scs8hd_fill_2
XFILLER_20_23 vpwr vgnd scs8hd_fill_2
XFILLER_29_65 vpwr vgnd scs8hd_fill_2
XFILLER_29_32 vpwr vgnd scs8hd_fill_2
XFILLER_29_21 vgnd vpwr scs8hd_decap_8
XFILLER_28_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_273 vgnd vpwr scs8hd_decap_4
XFILLER_3_262 vgnd vpwr scs8hd_decap_4
XFILLER_3_240 vpwr vgnd scs8hd_fill_2
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_19_152 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_33 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _217_/HI mem_right_track_0.LATCH_2_.latch/Q
+ mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_16_122 vpwr vgnd scs8hd_fill_2
XFILLER_31_147 vgnd vpwr scs8hd_decap_12
XANTENNA__127__C _127_/C vgnd vpwr scs8hd_diode_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB _118_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_199 vgnd vpwr scs8hd_decap_4
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _138_/X vgnd vpwr scs8hd_diode_2
XFILLER_22_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_169 vgnd vpwr scs8hd_decap_4
XFILLER_21_191 vpwr vgnd scs8hd_fill_2
XANTENNA__244__A _244_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A right_top_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_26 vpwr vgnd scs8hd_fill_2
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
XANTENNA__154__A _153_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_7 vpwr vgnd scs8hd_fill_2
XFILLER_18_206 vgnd vpwr scs8hd_decap_6
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XFILLER_18_239 vgnd vpwr scs8hd_decap_4
XANTENNA__239__A _239_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A left_top_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__149__A _120_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _203_/A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_275 vpwr vgnd scs8hd_fill_2
XFILLER_23_78 vpwr vgnd scs8hd_fill_2
XFILLER_2_146 vpwr vgnd scs8hd_fill_2
XFILLER_2_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_27 vpwr vgnd scs8hd_fill_2
XFILLER_0_49 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_3_.latch data_in mem_left_track_17.LATCH_3_.latch/Q _157_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_188_ _188_/A _188_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__151__B _146_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XFILLER_11_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
X_111_ address[6] _161_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_216 vpwr vgnd scs8hd_fill_2
XFILLER_11_245 vpwr vgnd scs8hd_fill_2
XFILLER_11_256 vpwr vgnd scs8hd_fill_2
XANTENNA__162__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_271 vgnd vpwr scs8hd_decap_4
XFILLER_28_142 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB _175_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_13.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_37 vpwr vgnd scs8hd_fill_2
XFILLER_19_131 vpwr vgnd scs8hd_fill_2
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XANTENNA__157__A _120_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_25_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_167 vpwr vgnd scs8hd_fill_2
XFILLER_31_45 vgnd vpwr scs8hd_decap_12
XFILLER_0_244 vpwr vgnd scs8hd_fill_2
XFILLER_16_145 vgnd vpwr scs8hd_decap_6
XFILLER_31_159 vgnd vpwr scs8hd_decap_12
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_259 vpwr vgnd scs8hd_fill_2
XFILLER_11_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_1_.latch data_in mem_left_track_1.LATCH_1_.latch/Q _143_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_148 vpwr vgnd scs8hd_fill_2
XFILLER_3_38 vgnd vpwr scs8hd_decap_4
XFILLER_8_141 vgnd vpwr scs8hd_fill_1
XFILLER_12_181 vpwr vgnd scs8hd_fill_2
XANTENNA__170__A _161_/X vgnd vpwr scs8hd_diode_2
Xmem_right_track_16.LATCH_2_.latch data_in mem_right_track_16.LATCH_2_.latch/Q _132_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_36 vgnd vpwr scs8hd_decap_6
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_5_111 vpwr vgnd scs8hd_fill_2
XFILLER_5_166 vgnd vpwr scs8hd_decap_4
XFILLER_5_188 vgnd vpwr scs8hd_decap_4
XANTENNA__149__B _146_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB _172_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_240 vpwr vgnd scs8hd_fill_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_232 vgnd vpwr scs8hd_decap_12
XFILLER_23_221 vpwr vgnd scs8hd_fill_2
XFILLER_23_35 vpwr vgnd scs8hd_fill_2
XFILLER_2_169 vpwr vgnd scs8hd_fill_2
XFILLER_2_136 vpwr vgnd scs8hd_fill_2
XFILLER_2_125 vpwr vgnd scs8hd_fill_2
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _187_/A _187_/Y vgnd vpwr scs8hd_inv_8
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chanx_right_in[1] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_224 vgnd vpwr scs8hd_decap_8
XFILLER_20_213 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_46 vpwr vgnd scs8hd_fill_2
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _201_/Y vgnd
+ vpwr scs8hd_diode_2
X_110_ _097_/A _123_/A _110_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_268 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_239_ _239_/A chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_110 vgnd vpwr scs8hd_decap_12
XFILLER_1_93 vpwr vgnd scs8hd_fill_2
XFILLER_28_154 vgnd vpwr scs8hd_decap_3
XFILLER_28_121 vgnd vpwr scs8hd_fill_1
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_8 vpwr vgnd scs8hd_fill_2
XANTENNA__157__B _154_/X vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _161_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_14 vpwr vgnd scs8hd_fill_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XFILLER_25_179 vpwr vgnd scs8hd_fill_2
XANTENNA__083__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_15_58 vgnd vpwr scs8hd_decap_3
XFILLER_15_69 vgnd vpwr scs8hd_decap_4
XFILLER_31_57 vgnd vpwr scs8hd_decap_4
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _187_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__168__A _161_/X vgnd vpwr scs8hd_diode_2
XFILLER_22_149 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_26_35 vgnd vpwr scs8hd_decap_12
XFILLER_13_127 vpwr vgnd scs8hd_fill_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_182 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_160 vpwr vgnd scs8hd_fill_2
XFILLER_8_131 vpwr vgnd scs8hd_fill_2
XFILLER_8_186 vgnd vpwr scs8hd_fill_1
XANTENNA__170__B _169_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_119 vgnd vpwr scs8hd_decap_6
XFILLER_12_26 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _203_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_230 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 right_top_grid_pin_9_ mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_274 vgnd vpwr scs8hd_fill_1
Xmem_right_track_0.LATCH_1_.latch data_in mem_right_track_0.LATCH_1_.latch/Q _107_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_156 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__181__A _178_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_71 vpwr vgnd scs8hd_fill_2
XFILLER_23_58 vgnd vpwr scs8hd_decap_3
XANTENNA__091__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_3_6 vpwr vgnd scs8hd_fill_2
XFILLER_9_38 vpwr vgnd scs8hd_fill_2
X_186_ _135_/Y _162_/A _164_/X _095_/C _186_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__176__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_247 vgnd vpwr scs8hd_decap_8
XFILLER_20_236 vgnd vpwr scs8hd_decap_8
Xmux_left_track_1.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[5] mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_36 vgnd vpwr scs8hd_decap_8
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XANTENNA__086__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_7_229 vgnd vpwr scs8hd_decap_4
XFILLER_1_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _189_/A vgnd
+ vpwr scs8hd_diode_2
X_169_ _169_/A _169_/X vgnd vpwr scs8hd_buf_1
XFILLER_24_90 vpwr vgnd scs8hd_fill_2
X_238_ _238_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_6_240 vgnd vpwr scs8hd_decap_6
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_7.LATCH_0_.latch data_in _194_/A _175_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_221 vpwr vgnd scs8hd_fill_2
XFILLER_10_81 vgnd vpwr scs8hd_decap_3
Xmux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_199 vpwr vgnd scs8hd_fill_2
XFILLER_19_166 vpwr vgnd scs8hd_fill_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XANTENNA__173__B _169_/X vgnd vpwr scs8hd_diode_2
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_147 vgnd vpwr scs8hd_fill_1
XFILLER_25_136 vpwr vgnd scs8hd_fill_2
XFILLER_25_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_37 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_213 vpwr vgnd scs8hd_fill_2
XFILLER_0_202 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_191 vgnd vpwr scs8hd_decap_8
XFILLER_24_180 vgnd vpwr scs8hd_decap_8
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_track_0.LATCH_3_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_106 vpwr vgnd scs8hd_fill_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _162_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__184__A _178_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_71 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_2_.latch data_in mem_left_track_9.LATCH_2_.latch/Q _150_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_47 vpwr vgnd scs8hd_fill_2
XANTENNA__094__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_21_172 vgnd vpwr scs8hd_decap_4
XFILLER_8_121 vgnd vpwr scs8hd_fill_1
XANTENNA__170__C _137_/C vgnd vpwr scs8hd_diode_2
XANTENNA__179__A _178_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_275 vpwr vgnd scs8hd_fill_2
XFILLER_35_253 vpwr vgnd scs8hd_fill_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XFILLER_26_242 vpwr vgnd scs8hd_fill_2
XANTENNA__089__A address[3] vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[4] mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
XFILLER_27_90 vgnd vpwr scs8hd_decap_4
XFILLER_17_231 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__181__B _162_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_61 vpwr vgnd scs8hd_fill_2
XFILLER_23_245 vpwr vgnd scs8hd_fill_2
XANTENNA__091__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_256 vgnd vpwr scs8hd_decap_4
X_185_ _135_/Y _162_/A _164_/X _165_/A _185_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_13_81 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A left_top_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_6 vpwr vgnd scs8hd_fill_2
XANTENNA__176__B _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA__192__A _192_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_259 vgnd vpwr scs8hd_decap_12
XANTENNA__086__B _083_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_59 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _201_/A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_11_237 vgnd vpwr scs8hd_decap_4
X_237_ _237_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
X_168_ _161_/X _162_/X _164_/X _167_/X _168_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_10_270 vgnd vpwr scs8hd_decap_4
X_099_ _098_/Y address[2] _165_/A _099_/X vgnd vpwr scs8hd_or3_4
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
XFILLER_1_40 vpwr vgnd scs8hd_fill_2
XANTENNA__187__A _187_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_right_track_8.LATCH_5_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_27 vpwr vgnd scs8hd_fill_2
XFILLER_29_69 vgnd vpwr scs8hd_decap_12
XFILLER_29_36 vgnd vpwr scs8hd_decap_12
XFILLER_29_14 vpwr vgnd scs8hd_fill_2
XANTENNA__097__A _097_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_211 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_15.LATCH_0_.latch data_in _202_/A _184_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_156 vgnd vpwr scs8hd_fill_1
XFILLER_19_123 vgnd vpwr scs8hd_fill_1
XFILLER_19_112 vpwr vgnd scs8hd_fill_2
XANTENNA__173__C _116_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XFILLER_0_269 vpwr vgnd scs8hd_fill_2
XFILLER_0_258 vgnd vpwr scs8hd_decap_8
XFILLER_16_126 vpwr vgnd scs8hd_fill_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA__168__C _164_/X vgnd vpwr scs8hd_diode_2
XANTENNA__184__B _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_251 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_140 vpwr vgnd scs8hd_fill_2
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XFILLER_21_195 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_70 vgnd vpwr scs8hd_fill_1
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_12_140 vpwr vgnd scs8hd_fill_2
XANTENNA__170__D _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA__179__B _162_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XANTENNA__195__A _195_/A vgnd vpwr scs8hd_diode_2
XANTENNA__089__B address[4] vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_track_1.LATCH_4_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_210 vgnd vpwr scs8hd_decap_4
Xmem_right_track_8.LATCH_2_.latch data_in mem_right_track_8.LATCH_2_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _244_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XFILLER_17_254 vgnd vpwr scs8hd_decap_6
XFILLER_17_276 vgnd vpwr scs8hd_fill_1
XANTENNA__181__C _116_/C vgnd vpwr scs8hd_diode_2
XFILLER_4_84 vpwr vgnd scs8hd_fill_2
XANTENNA__091__C _137_/C vgnd vpwr scs8hd_diode_2
XFILLER_2_106 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.INVTX1_6_.scs8hd_inv_1 left_top_grid_pin_11_ mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[8] mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_213 vgnd vpwr scs8hd_fill_1
XFILLER_14_235 vgnd vpwr scs8hd_decap_8
Xmux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_right_track_16.LATCH_5_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_184_ _178_/X _162_/A _127_/C _095_/C _184_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_13_71 vgnd vpwr scs8hd_decap_4
XFILLER_1_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__176__C _164_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_261 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_15.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XANTENNA__086__C _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_216 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
X_167_ _095_/C _167_/X vgnd vpwr scs8hd_buf_1
X_098_ address[1] _098_/Y vgnd vpwr scs8hd_inv_8
X_236_ chanx_left_in[0] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_37_135 vgnd vpwr scs8hd_decap_12
XFILLER_1_74 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_48 vgnd vpwr scs8hd_decap_12
XANTENNA__097__B _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_50 vgnd vpwr scs8hd_decap_3
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
XFILLER_19_146 vgnd vpwr scs8hd_decap_4
XFILLER_19_92 vgnd vpwr scs8hd_decap_4
XANTENNA__173__D _167_/X vgnd vpwr scs8hd_diode_2
X_219_ _219_/HI _219_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_3.LATCH_0_.latch data_in _190_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_71 vpwr vgnd scs8hd_fill_2
XFILLER_39_208 vgnd vpwr scs8hd_decap_12
XFILLER_22_119 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ _204_/A mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XANTENNA__184__C _127_/C vgnd vpwr scs8hd_diode_2
XANTENNA__168__D _167_/X vgnd vpwr scs8hd_diode_2
XFILLER_15_193 vgnd vpwr scs8hd_decap_4
XFILLER_30_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _204_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_95 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _215_/HI mem_left_track_17.LATCH_2_.latch/Q
+ mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_16_93 vpwr vgnd scs8hd_fill_2
XFILLER_8_145 vgnd vpwr scs8hd_decap_6
XFILLER_8_189 vpwr vgnd scs8hd_fill_2
XFILLER_12_152 vgnd vpwr scs8hd_fill_1
XFILLER_12_185 vpwr vgnd scs8hd_fill_2
XANTENNA__179__C _137_/C vgnd vpwr scs8hd_diode_2
XFILLER_12_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XANTENNA__089__C _125_/C vgnd vpwr scs8hd_diode_2
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_115 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_15.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_81 vpwr vgnd scs8hd_fill_2
XFILLER_17_266 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _228_/A vgnd vpwr scs8hd_inv_1
XANTENNA__181__D _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_41 vgnd vpwr scs8hd_decap_3
XFILLER_4_181 vpwr vgnd scs8hd_fill_2
XFILLER_23_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _190_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_19 vpwr vgnd scs8hd_fill_2
X_183_ _178_/X _162_/A _127_/C _165_/A _183_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_1_184 vgnd vpwr scs8hd_fill_1
XFILLER_1_140 vpwr vgnd scs8hd_fill_2
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__176__D _165_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_240 vpwr vgnd scs8hd_fill_2
XFILLER_9_273 vgnd vpwr scs8hd_decap_4
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _216_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_93 vpwr vgnd scs8hd_fill_2
XFILLER_24_82 vgnd vpwr scs8hd_decap_6
XFILLER_24_71 vpwr vgnd scs8hd_fill_2
X_235_ chanx_left_in[1] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
X_097_ _097_/A _130_/A _097_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_221 vgnd vpwr scs8hd_decap_4
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_166_ _161_/X _162_/X _164_/X _165_/X _166_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mem_left_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_37_147 vgnd vpwr scs8hd_decap_12
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_125 vgnd vpwr scs8hd_decap_8
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
XFILLER_27_180 vgnd vpwr scs8hd_decap_3
X_218_ _218_/HI _218_/LO vgnd vpwr scs8hd_conb_1
X_149_ _120_/A _146_/X _149_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_31_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _188_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _240_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_227 vpwr vgnd scs8hd_fill_2
XFILLER_24_150 vgnd vpwr scs8hd_fill_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_track_11.LATCH_0_.latch data_in _198_/A _180_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XANTENNA__184__D _095_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _192_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_220 vgnd vpwr scs8hd_decap_12
XFILLER_8_102 vpwr vgnd scs8hd_fill_2
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XFILLER_8_113 vpwr vgnd scs8hd_fill_2
XFILLER_8_135 vgnd vpwr scs8hd_decap_6
XFILLER_8_157 vpwr vgnd scs8hd_fill_2
XFILLER_35_245 vgnd vpwr scs8hd_decap_8
XANTENNA__179__D _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XFILLER_5_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_201 vpwr vgnd scs8hd_fill_2
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_160 vpwr vgnd scs8hd_fill_2
XFILLER_23_259 vpwr vgnd scs8hd_fill_2
XFILLER_23_204 vpwr vgnd scs8hd_fill_2
XFILLER_23_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_119 vgnd vpwr scs8hd_decap_4
XFILLER_22_270 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_182_ _178_/X _162_/X _116_/C _095_/C _182_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_14_226 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.INVTX1_1_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__100__A _099_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _190_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_29 vpwr vgnd scs8hd_fill_2
XFILLER_11_229 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_7 vgnd vpwr scs8hd_decap_3
X_165_ _165_/A _165_/X vgnd vpwr scs8hd_buf_1
XFILLER_24_50 vgnd vpwr scs8hd_decap_6
XFILLER_6_211 vgnd vpwr scs8hd_decap_3
X_234_ chanx_left_in[2] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
X_096_ _095_/X _130_/A vgnd vpwr scs8hd_buf_1
XFILLER_37_159 vgnd vpwr scs8hd_decap_12
XFILLER_27_6 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_7.INVTX1_0_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_21 vpwr vgnd scs8hd_fill_2
XFILLER_1_65 vpwr vgnd scs8hd_fill_2
XFILLER_3_269 vpwr vgnd scs8hd_fill_2
XFILLER_3_258 vpwr vgnd scs8hd_fill_2
XFILLER_3_236 vpwr vgnd scs8hd_fill_2
XFILLER_10_30 vgnd vpwr scs8hd_fill_1
XFILLER_10_41 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _199_/A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_148_ _130_/A _146_/X _148_/Y vgnd vpwr scs8hd_nor2_4
X_217_ _217_/HI _217_/LO vgnd vpwr scs8hd_conb_1
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XFILLER_18_192 vpwr vgnd scs8hd_fill_2
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.LATCH_4_.latch data_in mem_left_track_17.LATCH_4_.latch/Q _156_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_24_140 vpwr vgnd scs8hd_fill_2
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_118 vgnd vpwr scs8hd_fill_1
XFILLER_21_51 vpwr vgnd scs8hd_fill_2
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A right_top_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_9 vgnd vpwr scs8hd_decap_3
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.INVTX1_5_.scs8hd_inv_1 left_top_grid_pin_3_ mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_151 vpwr vgnd scs8hd_fill_2
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_7_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_18 vgnd vpwr scs8hd_decap_12
XFILLER_21_187 vpwr vgnd scs8hd_fill_2
XFILLER_21_132 vpwr vgnd scs8hd_fill_2
XFILLER_29_232 vgnd vpwr scs8hd_decap_12
XFILLER_12_154 vgnd vpwr scs8hd_decap_4
XFILLER_16_40 vgnd vpwr scs8hd_fill_1
XFILLER_16_84 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _185_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A left_top_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 right_top_grid_pin_7_ mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__103__A _102_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _209_/HI _203_/Y mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_191 vpwr vgnd scs8hd_fill_2
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_27_50 vpwr vgnd scs8hd_fill_2
XFILLER_4_65 vgnd vpwr scs8hd_decap_4
XFILLER_4_10 vpwr vgnd scs8hd_fill_2
XFILLER_23_249 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_205 vpwr vgnd scs8hd_fill_2
X_181_ _178_/X _162_/X _116_/C _165_/A _181_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_13_96 vpwr vgnd scs8hd_fill_2
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
Xmem_left_track_1.LATCH_2_.latch data_in mem_left_track_1.LATCH_2_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_175 vpwr vgnd scs8hd_fill_2
XFILLER_13_260 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_231 vpwr vgnd scs8hd_fill_2
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
Xmem_right_track_16.LATCH_3_.latch data_in mem_right_track_16.LATCH_3_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_233_ _233_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
X_164_ _163_/X _164_/X vgnd vpwr scs8hd_buf_1
X_095_ address[1] _083_/Y _095_/C _095_/X vgnd vpwr scs8hd_or3_4
XANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_44 vgnd vpwr scs8hd_decap_4
XANTENNA__111__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_28_105 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_11.INVTX1_1_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_8.INVTX1_6_.scs8hd_inv_1 chanx_left_in[1] mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_11.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_64 vpwr vgnd scs8hd_fill_2
XFILLER_10_86 vgnd vpwr scs8hd_decap_4
XFILLER_19_127 vpwr vgnd scs8hd_fill_2
XFILLER_19_116 vgnd vpwr scs8hd_decap_4
XFILLER_19_73 vpwr vgnd scs8hd_fill_2
XFILLER_19_62 vpwr vgnd scs8hd_fill_2
XFILLER_19_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__106__A _105_/X vgnd vpwr scs8hd_diode_2
X_216_ _216_/HI _216_/LO vgnd vpwr scs8hd_conb_1
X_147_ _129_/A _146_/X _147_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_track_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vpwr vgnd scs8hd_fill_2
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.INVTX1_0_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_163 vpwr vgnd scs8hd_fill_2
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_15_141 vpwr vgnd scs8hd_fill_2
XFILLER_30_166 vgnd vpwr scs8hd_decap_12
XFILLER_7_43 vgnd vpwr scs8hd_decap_4
XFILLER_21_155 vpwr vgnd scs8hd_fill_2
XFILLER_16_30 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_left_track_17.LATCH_3_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_100 vgnd vpwr scs8hd_decap_3
XFILLER_12_144 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_258 vgnd vpwr scs8hd_decap_12
XFILLER_26_247 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ _202_/A mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_107 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_73 vgnd vpwr scs8hd_decap_8
XFILLER_17_214 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[4] mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_2_.scs8hd_inv_1 right_bottom_grid_pin_12_ mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_88 vpwr vgnd scs8hd_fill_2
XANTENNA__114__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_228 vpwr vgnd scs8hd_fill_2
XFILLER_23_217 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_180_ _178_/X _162_/X _137_/C _167_/X _180_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XFILLER_1_165 vgnd vpwr scs8hd_fill_1
XFILLER_1_132 vpwr vgnd scs8hd_fill_2
XFILLER_20_209 vgnd vpwr scs8hd_decap_4
XANTENNA__109__A _108_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_232_ chanx_left_in[4] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_163_ _114_/A _124_/Y _125_/C _163_/X vgnd vpwr scs8hd_or3_4
X_094_ address[0] _095_/C vgnd vpwr scs8hd_buf_1
XFILLER_10_220 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _203_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_89 vpwr vgnd scs8hd_fill_2
Xmem_right_track_0.LATCH_2_.latch data_in mem_right_track_0.LATCH_2_.latch/Q _104_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _160_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_117 vgnd vpwr scs8hd_decap_4
XFILLER_19_96 vgnd vpwr scs8hd_fill_1
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
X_215_ _215_/HI _215_/LO vgnd vpwr scs8hd_conb_1
X_146_ _146_/A _146_/X vgnd vpwr scs8hd_buf_1
XANTENNA__122__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_6 vgnd vpwr scs8hd_decap_12
XFILLER_18_150 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_75 vpwr vgnd scs8hd_fill_2
XFILLER_21_31 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_164 vpwr vgnd scs8hd_fill_2
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XFILLER_30_178 vgnd vpwr scs8hd_decap_12
XFILLER_7_11 vpwr vgnd scs8hd_fill_2
XFILLER_7_22 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _116_/X vgnd vpwr scs8hd_diode_2
X_129_ _129_/A _129_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_99 vpwr vgnd scs8hd_fill_2
XFILLER_21_178 vgnd vpwr scs8hd_decap_4
XFILLER_21_112 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _195_/A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _189_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_7.LATCH_1_.latch data_in _193_/A _174_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_64 vgnd vpwr scs8hd_decap_6
XFILLER_32_30 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_3.INVTX1_0_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_16_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _219_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_119 vgnd vpwr scs8hd_fill_1
XANTENNA__220__A _220_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_237 vgnd vpwr scs8hd_fill_1
XFILLER_40_251 vgnd vpwr scs8hd_decap_12
XANTENNA__114__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA__130__A _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_144 vpwr vgnd scs8hd_fill_2
XFILLER_8_3 vgnd vpwr scs8hd_decap_4
Xmem_left_track_9.LATCH_3_.latch data_in mem_left_track_9.LATCH_3_.latch/Q _149_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_240 vpwr vgnd scs8hd_fill_2
XANTENNA__125__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _176_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_162_ _162_/A _162_/X vgnd vpwr scs8hd_buf_1
XFILLER_24_97 vgnd vpwr scs8hd_decap_6
XFILLER_24_20 vgnd vpwr scs8hd_decap_8
X_231_ chanx_left_in[5] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_10_210 vpwr vgnd scs8hd_fill_2
X_093_ _129_/A _097_/A _093_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_203 vpwr vgnd scs8hd_fill_2
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _191_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_217 vpwr vgnd scs8hd_fill_2
XFILLER_10_22 vgnd vpwr scs8hd_decap_8
XFILLER_19_53 vpwr vgnd scs8hd_fill_2
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vgnd vpwr scs8hd_decap_12
XFILLER_27_140 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_214_ _214_/HI _214_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_right_track_0.LATCH_4_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_145_ _135_/Y _169_/A _116_/C _146_/A vgnd vpwr scs8hd_or3_4
XANTENNA__122__B _120_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_140 vpwr vgnd scs8hd_fill_2
XFILLER_33_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_209 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _205_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__223__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_121 vgnd vpwr scs8hd_fill_1
XANTENNA__133__A _122_/A vgnd vpwr scs8hd_diode_2
X_128_ _127_/X _129_/B vgnd vpwr scs8hd_buf_1
XFILLER_38_202 vgnd vpwr scs8hd_decap_12
XFILLER_23_3 vgnd vpwr scs8hd_decap_4
Xmux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _197_/A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
XFILLER_16_10 vpwr vgnd scs8hd_fill_2
XFILLER_16_43 vgnd vpwr scs8hd_decap_4
XFILLER_8_106 vgnd vpwr scs8hd_decap_4
XFILLER_8_117 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A left_top_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_15.LATCH_1_.latch data_in _201_/A _183_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__128__A _127_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_161 vpwr vgnd scs8hd_fill_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_86 vpwr vgnd scs8hd_fill_2
XFILLER_40_263 vgnd vpwr scs8hd_decap_12
XFILLER_27_97 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A left_top_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__114__C _125_/C vgnd vpwr scs8hd_diode_2
XFILLER_4_142 vgnd vpwr scs8hd_decap_4
XFILLER_4_164 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__130__B _129_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_46 vpwr vgnd scs8hd_fill_2
XFILLER_23_208 vgnd vpwr scs8hd_decap_6
XFILLER_22_274 vgnd vpwr scs8hd_fill_1
XFILLER_22_241 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _208_/HI _201_/Y mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_77 vpwr vgnd scs8hd_fill_2
XANTENNA__231__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_1_112 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__125__B _124_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_212 vpwr vgnd scs8hd_fill_2
XFILLER_9_245 vgnd vpwr scs8hd_decap_3
XANTENNA__141__A _120_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_171 vgnd vpwr scs8hd_decap_12
X_161_ _161_/A _161_/X vgnd vpwr scs8hd_buf_1
XFILLER_24_65 vgnd vpwr scs8hd_decap_4
X_230_ chanx_left_in[6] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_6_215 vpwr vgnd scs8hd_fill_2
XANTENNA__226__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_248 vpwr vgnd scs8hd_fill_2
XFILLER_6_259 vgnd vpwr scs8hd_decap_12
X_092_ _091_/X _097_/A vgnd vpwr scs8hd_buf_1
Xmem_right_track_8.LATCH_3_.latch data_in mem_right_track_8.LATCH_3_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_25 vpwr vgnd scs8hd_fill_2
XFILLER_1_69 vgnd vpwr scs8hd_decap_3
XANTENNA__136__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_36_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_27_196 vgnd vpwr scs8hd_decap_12
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_213_ _213_/HI _213_/LO vgnd vpwr scs8hd_conb_1
X_144_ _123_/A _138_/X _144_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_163 vpwr vgnd scs8hd_fill_2
XFILLER_18_196 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[0] mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_144 vgnd vpwr scs8hd_decap_6
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_55 vgnd vpwr scs8hd_decap_4
XFILLER_21_11 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_199 vpwr vgnd scs8hd_fill_2
XANTENNA__133__B _129_/B vgnd vpwr scs8hd_diode_2
X_127_ address[6] address[5] _127_/C _127_/X vgnd vpwr scs8hd_or3_4
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
XFILLER_7_79 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _246_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_136 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_5_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_125 vpwr vgnd scs8hd_fill_2
XFILLER_12_136 vpwr vgnd scs8hd_fill_2
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XANTENNA__234__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__144__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_180 vgnd vpwr scs8hd_fill_1
XFILLER_11_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__229__A _229_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_65 vpwr vgnd scs8hd_fill_2
XFILLER_27_54 vgnd vpwr scs8hd_decap_4
XFILLER_27_43 vpwr vgnd scs8hd_fill_2
XFILLER_27_32 vpwr vgnd scs8hd_fill_2
XFILLER_27_21 vpwr vgnd scs8hd_fill_2
XFILLER_27_10 vpwr vgnd scs8hd_fill_2
XFILLER_4_154 vgnd vpwr scs8hd_decap_3
Xmem_bottom_track_3.LATCH_1_.latch data_in _189_/A _170_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XANTENNA__139__A _129_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_209 vgnd vpwr scs8hd_decap_4
XFILLER_13_12 vpwr vgnd scs8hd_fill_2
XFILLER_13_34 vpwr vgnd scs8hd_fill_2
XFILLER_1_179 vpwr vgnd scs8hd_fill_2
XFILLER_1_157 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ _200_/A mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__125__C _125_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_235 vgnd vpwr scs8hd_decap_3
XFILLER_9_257 vpwr vgnd scs8hd_fill_2
XFILLER_13_264 vgnd vpwr scs8hd_decap_12
XANTENNA__141__B _138_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_13.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_90 vgnd vpwr scs8hd_decap_3
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
X_160_ _123_/A _154_/X _160_/Y vgnd vpwr scs8hd_nor2_4
X_091_ address[6] address[5] _137_/C _091_/X vgnd vpwr scs8hd_or3_4
XFILLER_6_227 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[0] mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__242__A _242_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_260 vpwr vgnd scs8hd_fill_2
XANTENNA__152__A _123_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_46 vpwr vgnd scs8hd_fill_2
XFILLER_10_68 vgnd vpwr scs8hd_decap_4
XFILLER_27_153 vgnd vpwr scs8hd_decap_4
XFILLER_19_99 vpwr vgnd scs8hd_fill_2
XFILLER_19_88 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
XANTENNA__237__A _237_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_164 vpwr vgnd scs8hd_fill_2
X_212_ _212_/HI _212_/LO vgnd vpwr scs8hd_conb_1
X_143_ _122_/A _138_/X _143_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ _204_/Y mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_18_7 vpwr vgnd scs8hd_fill_2
XANTENNA__147__A _129_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_24_167 vgnd vpwr scs8hd_decap_4
XFILLER_24_112 vgnd vpwr scs8hd_decap_8
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.INVTX1_5_.scs8hd_inv_1 left_top_grid_pin_1_ mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_89 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_112 vgnd vpwr scs8hd_decap_6
XFILLER_15_123 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_145 vgnd vpwr scs8hd_decap_4
XFILLER_7_47 vgnd vpwr scs8hd_fill_1
X_126_ _125_/X _127_/C vgnd vpwr scs8hd_buf_1
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_30_6 vgnd vpwr scs8hd_decap_8
XFILLER_21_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_21_159 vpwr vgnd scs8hd_fill_2
XFILLER_16_23 vgnd vpwr scs8hd_decap_4
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB _182_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__144__B _138_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_174 vpwr vgnd scs8hd_fill_2
XANTENNA__160__A _123_/A vgnd vpwr scs8hd_diode_2
X_109_ _108_/X _123_/A vgnd vpwr scs8hd_buf_1
XFILLER_26_218 vgnd vpwr scs8hd_decap_12
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chanx_right_in[2] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_25_240 vgnd vpwr scs8hd_decap_4
XFILLER_17_218 vpwr vgnd scs8hd_fill_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XANTENNA__245__A _245_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _193_/A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_177 vpwr vgnd scs8hd_fill_2
XFILLER_31_232 vgnd vpwr scs8hd_decap_12
XANTENNA__155__A _129_/A vgnd vpwr scs8hd_diode_2
XANTENNA__139__B _138_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_11.LATCH_1_.latch data_in _197_/A _179_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_1_136 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_232 vpwr vgnd scs8hd_fill_2
XFILLER_13_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _192_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_269 vpwr vgnd scs8hd_fill_2
XFILLER_39_184 vgnd vpwr scs8hd_decap_12
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
X_090_ _089_/X _137_/C vgnd vpwr scs8hd_buf_1
XFILLER_10_224 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.INVTX1_6_.scs8hd_inv_1 chanx_left_in[0] mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__152__B _146_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB _179_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ _190_/A mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_35_11 vgnd vpwr scs8hd_decap_12
XFILLER_27_132 vpwr vgnd scs8hd_fill_2
XFILLER_19_23 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
X_211_ _211_/HI _211_/LO vgnd vpwr scs8hd_conb_1
X_142_ _121_/A _138_/X _142_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_135 vgnd vpwr scs8hd_decap_12
XANTENNA__147__B _146_/X vgnd vpwr scs8hd_diode_2
XFILLER_18_110 vgnd vpwr scs8hd_decap_6
XFILLER_18_121 vpwr vgnd scs8hd_fill_2
XANTENNA__163__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_190 vgnd vpwr scs8hd_decap_12
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_79 vgnd vpwr scs8hd_decap_3
XFILLER_21_35 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _190_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_168 vpwr vgnd scs8hd_fill_2
XFILLER_30_105 vgnd vpwr scs8hd_decap_12
X_125_ address[3] _124_/Y _125_/C _125_/X vgnd vpwr scs8hd_or3_4
XFILLER_7_26 vpwr vgnd scs8hd_fill_2
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XANTENNA__158__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_116 vgnd vpwr scs8hd_decap_4
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XFILLER_20_182 vgnd vpwr scs8hd_decap_8
XFILLER_12_105 vgnd vpwr scs8hd_decap_3
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _194_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_271 vgnd vpwr scs8hd_decap_4
XFILLER_7_142 vpwr vgnd scs8hd_fill_2
X_108_ address[1] address[2] address[0] _108_/X vgnd vpwr scs8hd_or3_4
XANTENNA__160__B _154_/X vgnd vpwr scs8hd_diode_2
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _198_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_263 vgnd vpwr scs8hd_decap_12
XFILLER_25_252 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_5_.latch data_in mem_left_track_17.LATCH_5_.latch/Q _155_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__155__B _154_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_274 vgnd vpwr scs8hd_fill_1
XANTENNA__171__A _161_/X vgnd vpwr scs8hd_diode_2
XFILLER_22_200 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _206_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__166__A _161_/X vgnd vpwr scs8hd_diode_2
XFILLER_39_196 vgnd vpwr scs8hd_decap_12
XFILLER_24_46 vpwr vgnd scs8hd_fill_2
XFILLER_24_35 vgnd vpwr scs8hd_decap_8
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_6_207 vpwr vgnd scs8hd_fill_2
XFILLER_10_258 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A right_top_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _207_/HI _199_/Y mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_240 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ _196_/A mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_36_166 vgnd vpwr scs8hd_decap_12
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_35_23 vgnd vpwr scs8hd_decap_12
XFILLER_19_57 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
X_210_ _210_/HI _210_/LO vgnd vpwr scs8hd_conb_1
X_141_ _120_/A _138_/X _141_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_232 vgnd vpwr scs8hd_decap_12
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_147 vgnd vpwr scs8hd_decap_12
XFILLER_18_144 vgnd vpwr scs8hd_decap_6
XANTENNA__163__B _124_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _110_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_3_.latch data_in mem_left_track_1.LATCH_3_.latch/Q _141_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_71 vpwr vgnd scs8hd_fill_2
XFILLER_2_60 vgnd vpwr scs8hd_decap_8
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _210_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
X_124_ address[4] _124_/Y vgnd vpwr scs8hd_inv_8
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
XANTENNA__158__B _154_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_6 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.LATCH_4_.latch data_in mem_right_track_16.LATCH_4_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__174__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_36 vgnd vpwr scs8hd_decap_4
XFILLER_16_58 vgnd vpwr scs8hd_decap_4
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XFILLER_20_150 vgnd vpwr scs8hd_fill_1
XANTENNA__084__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB _155_/Y vgnd vpwr scs8hd_diode_2
X_107_ _097_/A _122_/A _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_187 vpwr vgnd scs8hd_fill_2
XFILLER_11_172 vpwr vgnd scs8hd_fill_2
XANTENNA__169__A _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_275 vpwr vgnd scs8hd_fill_2
XFILLER_25_220 vgnd vpwr scs8hd_decap_12
XFILLER_4_102 vgnd vpwr scs8hd_decap_8
XFILLER_4_146 vgnd vpwr scs8hd_fill_1
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__171__B _169_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_212 vpwr vgnd scs8hd_fill_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_216 vpwr vgnd scs8hd_fill_2
XFILLER_13_212 vgnd vpwr scs8hd_decap_3
XFILLER_13_245 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
XANTENNA__166__B _162_/X vgnd vpwr scs8hd_diode_2
XANTENNA__182__A _178_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_260 vgnd vpwr scs8hd_decap_12
XFILLER_5_71 vpwr vgnd scs8hd_fill_2
XFILLER_10_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB _173_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XANTENNA__092__A _091_/X vgnd vpwr scs8hd_diode_2
XFILLER_36_178 vgnd vpwr scs8hd_decap_12
XANTENNA__177__A _161_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ _198_/A mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_19_69 vpwr vgnd scs8hd_fill_2
XFILLER_19_36 vpwr vgnd scs8hd_fill_2
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_35_35 vgnd vpwr scs8hd_decap_12
XFILLER_27_112 vgnd vpwr scs8hd_decap_4
XANTENNA__087__A _086_/X vgnd vpwr scs8hd_diode_2
X_140_ _130_/A _138_/X _140_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_244 vgnd vpwr scs8hd_fill_1
XFILLER_18_167 vgnd vpwr scs8hd_decap_12
XFILLER_33_159 vgnd vpwr scs8hd_decap_12
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__163__C _125_/C vgnd vpwr scs8hd_diode_2
XFILLER_21_15 vgnd vpwr scs8hd_decap_3
XFILLER_30_129 vgnd vpwr scs8hd_decap_12
XFILLER_23_170 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_track_17.LATCH_4_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_104 vpwr vgnd scs8hd_fill_2
X_123_ _123_/A _120_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__174__B _169_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__190__A _190_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ _202_/Y mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_0.LATCH_3_.latch data_in mem_right_track_0.LATCH_3_.latch/Q _101_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_28_251 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_151 vpwr vgnd scs8hd_fill_2
X_106_ _105_/X _122_/A vgnd vpwr scs8hd_buf_1
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A _135_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_69 vpwr vgnd scs8hd_fill_2
XFILLER_27_58 vgnd vpwr scs8hd_fill_1
XFILLER_25_232 vgnd vpwr scs8hd_fill_1
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XANTENNA__095__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_125 vpwr vgnd scs8hd_fill_2
XFILLER_4_136 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_210 vgnd vpwr scs8hd_decap_4
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XANTENNA__171__C _137_/C vgnd vpwr scs8hd_diode_2
XFILLER_13_16 vpwr vgnd scs8hd_fill_2
XFILLER_13_38 vgnd vpwr scs8hd_decap_4
XFILLER_1_106 vgnd vpwr scs8hd_decap_4
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_0_161 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _191_/A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__166__C _164_/X vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_3_ mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__182__B _162_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_250 vgnd vpwr scs8hd_fill_1
XFILLER_8_272 vgnd vpwr scs8hd_decap_3
XFILLER_39_110 vgnd vpwr scs8hd_decap_12
XFILLER_6_6 vgnd vpwr scs8hd_decap_4
XFILLER_5_264 vpwr vgnd scs8hd_fill_2
XFILLER_14_70 vgnd vpwr scs8hd_decap_3
XFILLER_30_80 vgnd vpwr scs8hd_decap_12
XANTENNA__177__B _169_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__193__A _193_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_35_47 vgnd vpwr scs8hd_decap_12
XFILLER_27_168 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_212 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[2] mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_179 vpwr vgnd scs8hd_fill_2
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_25_80 vpwr vgnd scs8hd_fill_2
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_199_ _199_/A _199_/Y vgnd vpwr scs8hd_inv_8
Xmem_left_track_9.LATCH_4_.latch data_in mem_left_track_9.LATCH_4_.latch/Q _148_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_84 vpwr vgnd scs8hd_fill_2
XANTENNA__188__A _188_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _213_/HI _195_/Y mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__098__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_23_193 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ _188_/A mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_15_127 vgnd vpwr scs8hd_fill_1
X_122_ _122_/A _120_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_108 vpwr vgnd scs8hd_fill_2
XANTENNA__174__C _127_/C vgnd vpwr scs8hd_diode_2
XFILLER_29_208 vgnd vpwr scs8hd_decap_12
XFILLER_20_141 vgnd vpwr scs8hd_decap_3
XFILLER_12_119 vgnd vpwr scs8hd_decap_4
XFILLER_16_27 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _191_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_70 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_105_ address[1] address[2] _105_/C _105_/X vgnd vpwr scs8hd_or3_4
XFILLER_7_112 vgnd vpwr scs8hd_decap_4
XFILLER_7_123 vpwr vgnd scs8hd_fill_2
XFILLER_7_178 vgnd vpwr scs8hd_decap_3
XFILLER_19_263 vgnd vpwr scs8hd_decap_12
XANTENNA__185__B _162_/A vgnd vpwr scs8hd_diode_2
XANTENNA__095__B _083_/Y vgnd vpwr scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_244 vpwr vgnd scs8hd_fill_2
XFILLER_16_255 vgnd vpwr scs8hd_decap_8
XFILLER_16_266 vgnd vpwr scs8hd_decap_8
XFILLER_17_81 vgnd vpwr scs8hd_fill_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
XANTENNA__171__D _167_/X vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_7_.scs8hd_inv_1 left_top_grid_pin_15_ mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__196__A _196_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_258 vgnd vpwr scs8hd_decap_12
XFILLER_22_247 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_236 vpwr vgnd scs8hd_fill_2
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _211_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_0.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[1] mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__166__D _165_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_40 vpwr vgnd scs8hd_fill_2
XANTENNA__182__C _116_/C vgnd vpwr scs8hd_diode_2
XFILLER_5_95 vgnd vpwr scs8hd_decap_3
XFILLER_24_16 vpwr vgnd scs8hd_fill_2
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_206 vpwr vgnd scs8hd_fill_2
XFILLER_10_239 vgnd vpwr scs8hd_decap_6
Xmux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_right_track_0.LATCH_5_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_7 vpwr vgnd scs8hd_fill_2
XANTENNA__177__C _164_/X vgnd vpwr scs8hd_diode_2
XFILLER_10_18 vpwr vgnd scs8hd_fill_2
XFILLER_27_136 vpwr vgnd scs8hd_fill_2
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_2_202 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _193_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_257 vgnd vpwr scs8hd_decap_12
XFILLER_18_125 vpwr vgnd scs8hd_fill_2
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_198_ _198_/A _198_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_41 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _206_/HI _197_/Y mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _197_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_39 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ _194_/A mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_121_ _121_/A _120_/B _121_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A left_top_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XFILLER_14_150 vgnd vpwr scs8hd_fill_1
XFILLER_14_172 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__174__D _165_/X vgnd vpwr scs8hd_diode_2
XFILLER_14_194 vpwr vgnd scs8hd_fill_2
XANTENNA__199__A _199_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_220 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_4_.latch data_in mem_right_track_8.LATCH_4_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_120 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
X_104_ _097_/A _121_/A _104_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_82 vgnd vpwr scs8hd_decap_4
XFILLER_7_157 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_0_.latch data_in mem_left_track_17.LATCH_0_.latch/Q _160_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_7 vpwr vgnd scs8hd_fill_2
XFILLER_19_275 vpwr vgnd scs8hd_fill_2
XFILLER_19_220 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_6 vpwr vgnd scs8hd_fill_2
XANTENNA__185__C _164_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_62 vpwr vgnd scs8hd_fill_2
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XANTENNA__095__C _095_/C vgnd vpwr scs8hd_diode_2
XFILLER_4_149 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_71 vgnd vpwr scs8hd_decap_4
XFILLER_17_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _216_/HI mem_left_track_9.LATCH_2_.latch/Q
+ mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_12_3 vpwr vgnd scs8hd_fill_2
XFILLER_13_29 vgnd vpwr scs8hd_decap_3
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _207_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA__182__D _095_/C vgnd vpwr scs8hd_diode_2
XFILLER_8_230 vpwr vgnd scs8hd_fill_2
XFILLER_5_30 vgnd vpwr scs8hd_fill_1
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XFILLER_24_28 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_93 vgnd vpwr scs8hd_decap_12
XFILLER_5_211 vpwr vgnd scs8hd_fill_2
XANTENNA__177__D _167_/X vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_5_.scs8hd_inv_1 left_top_grid_pin_5_ mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[5] mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_27_159 vpwr vgnd scs8hd_fill_2
XFILLER_2_247 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_269 vgnd vpwr scs8hd_decap_6
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_197_ _197_/A _197_/Y vgnd vpwr scs8hd_inv_8
XFILLER_24_129 vgnd vpwr scs8hd_decap_6
XFILLER_15_118 vgnd vpwr scs8hd_fill_1
X_120_ _120_/A _120_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_173 vgnd vpwr scs8hd_decap_8
XFILLER_11_40 vpwr vgnd scs8hd_fill_2
XFILLER_11_95 vpwr vgnd scs8hd_fill_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_165 vpwr vgnd scs8hd_fill_2
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_11_132 vpwr vgnd scs8hd_fill_2
X_103_ _102_/X _121_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_136 vgnd vpwr scs8hd_decap_4
XFILLER_11_176 vgnd vpwr scs8hd_decap_4
XFILLER_11_187 vpwr vgnd scs8hd_fill_2
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_19_243 vgnd vpwr scs8hd_fill_1
XANTENNA__185__D _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_41 vgnd vpwr scs8hd_decap_8
XFILLER_27_39 vpwr vgnd scs8hd_fill_2
XFILLER_27_28 vpwr vgnd scs8hd_fill_2
XFILLER_27_17 vpwr vgnd scs8hd_fill_2
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ _200_/Y mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_3.INVTX1_2_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_11.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_5_75 vpwr vgnd scs8hd_fill_2
XFILLER_39_135 vgnd vpwr scs8hd_decap_12
XFILLER_38_190 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _233_/A vgnd vpwr scs8hd_inv_1
XFILLER_14_84 vgnd vpwr scs8hd_decap_8
XFILLER_5_245 vgnd vpwr scs8hd_decap_4
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
XANTENNA__101__A _097_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_35_171 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _189_/A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_6 vpwr vgnd scs8hd_fill_2
XFILLER_2_215 vpwr vgnd scs8hd_fill_2
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
X_196_ _196_/A _196_/Y vgnd vpwr scs8hd_inv_8
Xmux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _243_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_10 vpwr vgnd scs8hd_fill_2
XFILLER_1_270 vgnd vpwr scs8hd_decap_6
XFILLER_32_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_108 vpwr vgnd scs8hd_fill_2
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_163 vpwr vgnd scs8hd_fill_2
X_179_ _178_/X _162_/X _137_/C _165_/X _179_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_32_18 vgnd vpwr scs8hd_decap_12
XFILLER_20_199 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _212_/HI _193_/Y mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_155 vpwr vgnd scs8hd_fill_2
X_102_ _098_/Y address[2] _095_/C _102_/X vgnd vpwr scs8hd_or3_4
XFILLER_19_233 vpwr vgnd scs8hd_fill_2
XFILLER_25_203 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_25_236 vpwr vgnd scs8hd_fill_2
XFILLER_16_225 vpwr vgnd scs8hd_fill_2
XFILLER_16_236 vgnd vpwr scs8hd_decap_8
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__104__A _097_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_184 vpwr vgnd scs8hd_fill_2
XFILLER_3_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB _093_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_217 vgnd vpwr scs8hd_decap_4
XFILLER_0_198 vpwr vgnd scs8hd_fill_2
XFILLER_0_165 vpwr vgnd scs8hd_fill_2
XFILLER_8_210 vpwr vgnd scs8hd_fill_2
XFILLER_8_243 vgnd vpwr scs8hd_decap_4
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_9.LATCH_0_.latch data_in _196_/A _177_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_147 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _210_/HI _190_/Y mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _194_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_41 vgnd vpwr scs8hd_decap_3
XFILLER_14_96 vpwr vgnd scs8hd_fill_2
XFILLER_5_268 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _198_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_117 vgnd vpwr scs8hd_decap_12
XANTENNA__101__B _120_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_2_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_19 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.INVTX1_0_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_84 vpwr vgnd scs8hd_fill_2
XFILLER_25_62 vpwr vgnd scs8hd_fill_2
XFILLER_25_40 vpwr vgnd scs8hd_fill_2
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_195_ _195_/A _195_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__112__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_2_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_197 vgnd vpwr scs8hd_decap_4
XFILLER_23_153 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XFILLER_11_75 vpwr vgnd scs8hd_fill_2
XANTENNA__107__A _097_/A vgnd vpwr scs8hd_diode_2
X_178_ _135_/Y _178_/X vgnd vpwr scs8hd_buf_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_245 vgnd vpwr scs8hd_decap_12
XFILLER_20_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr
+ scs8hd_diode_2
X_101_ _097_/A _120_/A _101_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_41 vpwr vgnd scs8hd_fill_2
XFILLER_11_112 vpwr vgnd scs8hd_fill_2
XFILLER_19_245 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ _192_/A mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _196_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_182 vpwr vgnd scs8hd_fill_2
XFILLER_25_248 vpwr vgnd scs8hd_fill_2
XFILLER_25_215 vpwr vgnd scs8hd_fill_2
XFILLER_25_259 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_left_track_1.LATCH_4_.latch data_in mem_left_track_1.LATCH_4_.latch/Q _140_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_119 vgnd vpwr scs8hd_decap_4
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _200_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_215 vgnd vpwr scs8hd_fill_1
XFILLER_17_41 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XANTENNA__104__B _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_163 vgnd vpwr scs8hd_fill_1
XANTENNA__120__A _120_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
XFILLER_22_229 vgnd vpwr scs8hd_decap_12
XFILLER_22_218 vgnd vpwr scs8hd_decap_8
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_3_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _186_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_16.LATCH_5_.latch data_in mem_right_track_16.LATCH_5_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_1_ mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_240 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A right_top_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _239_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _212_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_22 vpwr vgnd scs8hd_fill_2
XANTENNA__115__A _114_/X vgnd vpwr scs8hd_diode_2
XFILLER_39_159 vgnd vpwr scs8hd_decap_12
XFILLER_10_3 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ _196_/Y mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_0_.latch data_in _204_/A _186_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_129 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XFILLER_2_206 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ _194_/A _194_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XFILLER_17_140 vgnd vpwr scs8hd_fill_1
XFILLER_17_184 vpwr vgnd scs8hd_fill_2
XFILLER_23_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB _183_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_21 vpwr vgnd scs8hd_fill_2
XFILLER_11_32 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_11.INVTX1_0_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_8.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[6] mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_132 vgnd vpwr scs8hd_decap_3
XANTENNA__107__B _122_/A vgnd vpwr scs8hd_diode_2
X_246_ _246_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
X_177_ _161_/A _169_/A _164_/X _167_/X _177_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_14_176 vgnd vpwr scs8hd_fill_1
XFILLER_14_198 vpwr vgnd scs8hd_fill_2
XANTENNA__123__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XFILLER_20_146 vgnd vpwr scs8hd_decap_4
XFILLER_9_191 vpwr vgnd scs8hd_fill_2
XFILLER_22_64 vgnd vpwr scs8hd_decap_6
X_100_ _099_/X _120_/A vgnd vpwr scs8hd_buf_1
XFILLER_11_168 vpwr vgnd scs8hd_fill_2
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _129_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_22 vgnd vpwr scs8hd_decap_4
X_229_ _229_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_8_66 vgnd vpwr scs8hd_decap_4
Xmux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_7_.scs8hd_inv_1 left_top_grid_pin_13_ mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_20 vpwr vgnd scs8hd_fill_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_271 vgnd vpwr scs8hd_decap_4
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XFILLER_17_97 vpwr vgnd scs8hd_fill_2
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XFILLER_3_175 vpwr vgnd scs8hd_fill_2
XFILLER_3_153 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _120_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
XFILLER_13_208 vpwr vgnd scs8hd_fill_2
XFILLER_21_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__221__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_0_178 vpwr vgnd scs8hd_fill_2
XFILLER_0_156 vgnd vpwr scs8hd_fill_1
XFILLER_0_112 vgnd vpwr scs8hd_decap_8
XFILLER_0_134 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_30 vgnd vpwr scs8hd_fill_1
Xmem_right_track_0.LATCH_4_.latch data_in mem_right_track_0.LATCH_4_.latch/Q _097_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _208_/HI vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ _198_/Y mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__131__A _120_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[1] mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 right_top_grid_pin_11_ mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_10 vpwr vgnd scs8hd_fill_2
XFILLER_5_215 vpwr vgnd scs8hd_fill_2
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_171 vgnd vpwr scs8hd_decap_12
XANTENNA__126__A _125_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_108 vpwr vgnd scs8hd_fill_2
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_5.LATCH_0_.latch data_in _192_/A _173_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_174 vgnd vpwr scs8hd_decap_12
XFILLER_26_163 vgnd vpwr scs8hd_decap_8
XFILLER_26_152 vgnd vpwr scs8hd_fill_1
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_5_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XFILLER_25_97 vpwr vgnd scs8hd_fill_2
X_193_ _193_/A _193_/Y vgnd vpwr scs8hd_inv_8
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_2_68 vgnd vpwr scs8hd_fill_1
XFILLER_2_46 vgnd vpwr scs8hd_decap_3
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XFILLER_17_152 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_166 vgnd vpwr scs8hd_decap_4
XFILLER_2_6 vpwr vgnd scs8hd_fill_2
XFILLER_11_99 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _187_/A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_14_100 vgnd vpwr scs8hd_decap_4
XFILLER_14_144 vgnd vpwr scs8hd_decap_6
X_245_ _245_/A chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
X_176_ _161_/A _169_/A _164_/X _165_/X _176_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__123__B _120_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XFILLER_20_169 vgnd vpwr scs8hd_decap_4
XFILLER_20_125 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__224__A _224_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_32 vgnd vpwr scs8hd_fill_1
XFILLER_22_21 vgnd vpwr scs8hd_decap_4
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XFILLER_11_136 vgnd vpwr scs8hd_decap_4
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_19_203 vpwr vgnd scs8hd_fill_2
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XANTENNA__118__B _120_/B vgnd vpwr scs8hd_diode_2
X_228_ _228_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA__134__A _123_/A vgnd vpwr scs8hd_diode_2
X_159_ _122_/A _154_/X _159_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_89 vgnd vpwr scs8hd_decap_3
Xmem_left_track_9.LATCH_5_.latch data_in mem_left_track_9.LATCH_5_.latch/Q _147_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _215_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_206 vpwr vgnd scs8hd_fill_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_132 vpwr vgnd scs8hd_fill_2
XANTENNA__129__A _129_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_261 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _211_/HI _191_/Y mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_272 vgnd vpwr scs8hd_decap_4
XFILLER_21_220 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_275 vpwr vgnd scs8hd_fill_2
XFILLER_28_64 vgnd vpwr scs8hd_decap_12
XANTENNA__131__B _129_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XANTENNA__232__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _121_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_260 vgnd vpwr scs8hd_decap_12
XFILLER_2_219 vpwr vgnd scs8hd_fill_2
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_186 vgnd vpwr scs8hd_decap_12
XFILLER_26_131 vgnd vpwr scs8hd_decap_4
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _205_/HI _188_/Y mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_21 vgnd vpwr scs8hd_decap_3
XANTENNA__227__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XPHY_32 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_192_ _192_/A _192_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_241 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_13.LATCH_0_.latch data_in _200_/A _182_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _177_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_178 vgnd vpwr scs8hd_decap_12
XANTENNA__137__A _135_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_175 vpwr vgnd scs8hd_fill_2
XFILLER_17_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_112 vgnd vpwr scs8hd_decap_4
Xmux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _219_/HI mem_right_track_8.LATCH_2_.latch/Q
+ mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_244_ _244_/A chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_14_167 vgnd vpwr scs8hd_decap_3
X_175_ _161_/A _169_/X _127_/C _167_/X _175_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_35_7 vpwr vgnd scs8hd_fill_2
XFILLER_20_137 vpwr vgnd scs8hd_fill_2
XFILLER_28_259 vgnd vpwr scs8hd_decap_12
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_88 vgnd vpwr scs8hd_decap_4
XFILLER_22_55 vpwr vgnd scs8hd_fill_2
XANTENNA__240__A _240_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_259 vpwr vgnd scs8hd_fill_2
XFILLER_19_237 vgnd vpwr scs8hd_decap_6
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XFILLER_8_79 vgnd vpwr scs8hd_decap_8
X_227_ chanx_right_in[0] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA__134__B _129_/B vgnd vpwr scs8hd_diode_2
X_158_ _121_/A _154_/X _158_/Y vgnd vpwr scs8hd_nor2_4
X_089_ address[3] address[4] _125_/C _089_/X vgnd vpwr scs8hd_or3_4
XFILLER_6_152 vgnd vpwr scs8hd_fill_1
XFILLER_6_163 vpwr vgnd scs8hd_fill_2
XFILLER_6_174 vpwr vgnd scs8hd_fill_2
XFILLER_10_181 vpwr vgnd scs8hd_fill_2
XANTENNA__150__A _121_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _193_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB _104_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_229 vgnd vpwr scs8hd_decap_4
XFILLER_17_77 vgnd vpwr scs8hd_decap_4
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vgnd vpwr scs8hd_decap_12
XFILLER_33_10 vgnd vpwr scs8hd_decap_12
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__235__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _197_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_188 vgnd vpwr scs8hd_decap_4
XANTENNA__129__B _129_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_240 vpwr vgnd scs8hd_fill_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A _135_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ _190_/A mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB _174_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_232 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_8.LATCH_5_.latch data_in mem_right_track_8.LATCH_5_.latch/Q _118_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XFILLER_28_76 vgnd vpwr scs8hd_decap_12
XFILLER_12_210 vpwr vgnd scs8hd_fill_2
XFILLER_8_247 vgnd vpwr scs8hd_fill_1
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_36 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_1_.latch data_in mem_left_track_17.LATCH_1_.latch/Q _159_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_23 vpwr vgnd scs8hd_fill_2
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XANTENNA__142__B _138_/X vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _218_/HI mem_right_track_16.LATCH_2_.latch/Q
+ mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_272 vgnd vpwr scs8hd_decap_3
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ _194_/Y mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_198 vgnd vpwr scs8hd_decap_12
XFILLER_25_66 vgnd vpwr scs8hd_decap_3
XFILLER_25_44 vgnd vpwr scs8hd_decap_6
XFILLER_25_33 vpwr vgnd scs8hd_fill_2
XFILLER_25_22 vpwr vgnd scs8hd_fill_2
XFILLER_25_11 vgnd vpwr scs8hd_decap_4
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
X_191_ _191_/A _191_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__243__A _243_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A left_top_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_110 vpwr vgnd scs8hd_fill_2
XFILLER_17_132 vpwr vgnd scs8hd_fill_2
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XANTENNA__137__B _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _195_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__153__A _135_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _199_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_79 vgnd vpwr scs8hd_decap_3
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XANTENNA__238__A _238_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_0_.latch data_in _188_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_243_ _243_/A chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
X_174_ _161_/A _169_/X _127_/C _165_/X _174_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_28_7 vgnd vpwr scs8hd_decap_8
XFILLER_20_105 vgnd vpwr scs8hd_decap_4
XANTENNA__148__A _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_227 vgnd vpwr scs8hd_decap_12
XFILLER_3_91 vpwr vgnd scs8hd_fill_2
XFILLER_11_116 vgnd vpwr scs8hd_decap_4
XFILLER_22_45 vgnd vpwr scs8hd_fill_1
XFILLER_19_216 vpwr vgnd scs8hd_fill_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
XFILLER_19_249 vgnd vpwr scs8hd_decap_4
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 chanx_right_in[5] mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_157_ _120_/A _154_/X _157_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_160 vpwr vgnd scs8hd_fill_2
X_226_ chanx_right_in[1] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
X_088_ enable _125_/C vgnd vpwr scs8hd_inv_8
XANTENNA__150__B _146_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_241 vgnd vpwr scs8hd_decap_4
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_22 vgnd vpwr scs8hd_decap_12
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_right_track_16.LATCH_0_.latch data_in mem_right_track_16.LATCH_0_.latch/Q _134_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_112 vpwr vgnd scs8hd_fill_2
X_209_ _209_/HI _209_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA__145__B _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_70 vpwr vgnd scs8hd_fill_2
XFILLER_28_88 vgnd vpwr scs8hd_decap_4
XANTENNA__246__A _246_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_244 vgnd vpwr scs8hd_fill_1
XFILLER_5_26 vgnd vpwr scs8hd_decap_4
XFILLER_8_215 vpwr vgnd scs8hd_fill_2
XFILLER_8_226 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _213_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__156__A _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_141 vgnd vpwr scs8hd_decap_12
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XFILLER_14_46 vgnd vpwr scs8hd_decap_3
XFILLER_39_98 vgnd vpwr scs8hd_decap_12
XFILLER_29_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_144 vgnd vpwr scs8hd_decap_8
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
X_190_ _190_/A _190_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_27 vpwr vgnd scs8hd_fill_2
XFILLER_1_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_254 vpwr vgnd scs8hd_fill_2
XFILLER_1_221 vpwr vgnd scs8hd_fill_2
XANTENNA__137__C _137_/C vgnd vpwr scs8hd_diode_2
XANTENNA__153__B _169_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_2_.scs8hd_inv_1 right_top_grid_pin_15_ mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_136 vpwr vgnd scs8hd_fill_2
XFILLER_11_25 vpwr vgnd scs8hd_fill_2
XFILLER_11_36 vpwr vgnd scs8hd_fill_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
X_242_ _242_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
X_173_ _161_/X _169_/X _116_/C _167_/X _173_/Y vgnd vpwr scs8hd_nor4_4
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__148__B _146_/X vgnd vpwr scs8hd_diode_2
XANTENNA__164__A _163_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_140 vpwr vgnd scs8hd_fill_2
XFILLER_9_151 vgnd vpwr scs8hd_decap_4
XFILLER_3_70 vpwr vgnd scs8hd_fill_2
XFILLER_28_239 vgnd vpwr scs8hd_decap_12
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
Xmux_left_track_1.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_156_ _130_/A _154_/X _156_/Y vgnd vpwr scs8hd_nor2_4
X_087_ _086_/X _129_/A vgnd vpwr scs8hd_buf_1
XFILLER_8_26 vgnd vpwr scs8hd_fill_1
XFILLER_10_150 vgnd vpwr scs8hd_fill_1
X_225_ chanx_right_in[2] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_33_6 vpwr vgnd scs8hd_fill_2
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
XANTENNA__159__A _122_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_34 vgnd vpwr scs8hd_decap_12
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_24 vpwr vgnd scs8hd_fill_2
XFILLER_17_46 vpwr vgnd scs8hd_fill_2
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__145__C _116_/C vgnd vpwr scs8hd_diode_2
XFILLER_15_231 vpwr vgnd scs8hd_fill_2
X_208_ _208_/HI _208_/LO vgnd vpwr scs8hd_conb_1
X_139_ _129_/A _138_/X _139_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_190 vpwr vgnd scs8hd_fill_2
XFILLER_21_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _214_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_256 vgnd vpwr scs8hd_decap_8
XFILLER_12_267 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _209_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA__156__B _154_/X vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _161_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_7_271 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _189_/Y mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _245_/A vgnd vpwr scs8hd_inv_1
XFILLER_14_58 vgnd vpwr scs8hd_decap_12
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XFILLER_5_219 vgnd vpwr scs8hd_decap_4
XFILLER_39_11 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__167__A _095_/C vgnd vpwr scs8hd_diode_2
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XFILLER_1_233 vpwr vgnd scs8hd_fill_2
XFILLER_9_3 vgnd vpwr scs8hd_decap_3
XFILLER_1_266 vpwr vgnd scs8hd_fill_2
XFILLER_17_156 vpwr vgnd scs8hd_fill_2
XANTENNA__153__C _127_/C vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[7] mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_track_9.LATCH_1_.latch data_in _195_/A _176_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_track_8.LATCH_3_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB _180_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_104 vgnd vpwr scs8hd_fill_1
X_241_ _241_/A chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
X_172_ _161_/X _169_/X _116_/C _165_/X _172_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__180__A _178_/X vgnd vpwr scs8hd_diode_2
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
XFILLER_22_36 vgnd vpwr scs8hd_decap_3
XFILLER_22_25 vgnd vpwr scs8hd_fill_1
Xmem_left_track_9.LATCH_0_.latch data_in mem_left_track_9.LATCH_0_.latch/Q _152_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__090__A _089_/X vgnd vpwr scs8hd_diode_2
X_224_ _224_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_8_49 vpwr vgnd scs8hd_fill_2
X_086_ address[1] _083_/Y _165_/A _086_/X vgnd vpwr scs8hd_or3_4
X_155_ _129_/A _154_/X _155_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_100 vpwr vgnd scs8hd_fill_2
XFILLER_33_232 vgnd vpwr scs8hd_decap_12
XANTENNA__159__B _154_/X vgnd vpwr scs8hd_diode_2
XANTENNA__175__A _161_/A vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_46 vgnd vpwr scs8hd_decap_12
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XANTENNA__085__A _105_/C vgnd vpwr scs8hd_diode_2
XFILLER_3_136 vpwr vgnd scs8hd_fill_2
XFILLER_30_202 vgnd vpwr scs8hd_decap_12
X_207_ _207_/HI _207_/LO vgnd vpwr scs8hd_conb_1
XFILLER_15_276 vgnd vpwr scs8hd_fill_1
X_138_ _137_/X _138_/X vgnd vpwr scs8hd_buf_1
XFILLER_24_3 vpwr vgnd scs8hd_fill_2
XFILLER_21_224 vpwr vgnd scs8hd_fill_2
XFILLER_0_94 vgnd vpwr scs8hd_decap_3
XFILLER_0_139 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_46 vgnd vpwr scs8hd_decap_12
XFILLER_28_35 vgnd vpwr scs8hd_decap_8
XFILLER_8_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__172__B _169_/X vgnd vpwr scs8hd_diode_2
XFILLER_38_154 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ _188_/A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_23 vgnd vpwr scs8hd_decap_12
XFILLER_29_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _196_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_231 vgnd vpwr scs8hd_decap_3
Xmem_left_track_1.LATCH_5_.latch data_in mem_left_track_1.LATCH_5_.latch/Q _139_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_135 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_3_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__183__A _178_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _200_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_102 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_36 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XANTENNA__093__A _129_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
XFILLER_15_91 vpwr vgnd scs8hd_fill_2
XFILLER_17_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__178__A _135_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_171 vgnd vpwr scs8hd_decap_12
XFILLER_23_149 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A enable vgnd vpwr scs8hd_diode_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
X_240_ _240_/A chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_22_171 vgnd vpwr scs8hd_decap_4
X_171_ _161_/X _169_/X _137_/C _167_/X _171_/Y vgnd vpwr scs8hd_nor4_4
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ _192_/Y mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_1_.latch data_in _203_/A _185_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XANTENNA__180__B _162_/X vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_12_ mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_208 vgnd vpwr scs8hd_decap_6
Xmux_right_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[2] mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XFILLER_22_59 vgnd vpwr scs8hd_decap_3
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_223_ chanx_right_in[4] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
X_154_ _153_/X _154_/X vgnd vpwr scs8hd_buf_1
X_085_ _105_/C _165_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_145 vgnd vpwr scs8hd_fill_1
XFILLER_6_167 vpwr vgnd scs8hd_fill_2
XFILLER_6_178 vpwr vgnd scs8hd_fill_2
XFILLER_10_185 vpwr vgnd scs8hd_fill_2
XFILLER_26_7 vgnd vpwr scs8hd_decap_8
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
XFILLER_18_252 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_track_9.LATCH_4_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA__175__B _169_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _241_/A vgnd vpwr scs8hd_inv_1
XANTENNA__191__A _191_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_37 vpwr vgnd scs8hd_fill_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_58 vgnd vpwr scs8hd_decap_3
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_3_159 vgnd vpwr scs8hd_decap_4
Xmem_right_track_8.LATCH_0_.latch data_in mem_right_track_8.LATCH_0_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_206_ _206_/HI _206_/LO vgnd vpwr scs8hd_conb_1
X_137_ _135_/Y _169_/A _137_/C _137_/X vgnd vpwr scs8hd_or3_4
Xmux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_3 vgnd vpwr scs8hd_decap_4
XFILLER_21_236 vpwr vgnd scs8hd_fill_2
XANTENNA__186__A _135_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _202_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_71 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _220_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_28_58 vgnd vpwr scs8hd_decap_3
XANTENNA__096__A _095_/X vgnd vpwr scs8hd_diode_2
XFILLER_12_225 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__172__C _116_/C vgnd vpwr scs8hd_diode_2
XFILLER_38_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XFILLER_39_35 vgnd vpwr scs8hd_decap_12
XFILLER_4_210 vpwr vgnd scs8hd_fill_2
XFILLER_4_243 vgnd vpwr scs8hd_decap_6
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_147 vgnd vpwr scs8hd_decap_12
XANTENNA__183__B _162_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _224_/A vgnd vpwr scs8hd_inv_1
XFILLER_6_72 vgnd vpwr scs8hd_fill_1
XPHY_59 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XANTENNA__093__B _097_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _188_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_202 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_136 vgnd vpwr scs8hd_decap_4
XFILLER_17_169 vgnd vpwr scs8hd_decap_4
XFILLER_32_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_191 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__194__A _194_/A vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_5_.latch data_in mem_right_track_0.LATCH_5_.latch/Q _093_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_22_183 vgnd vpwr scs8hd_fill_1
X_170_ _161_/X _169_/X _137_/C _165_/X _170_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_14_128 vpwr vgnd scs8hd_fill_2
XFILLER_26_80 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_187 vpwr vgnd scs8hd_fill_2
XANTENNA__180__C _137_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_95 vpwr vgnd scs8hd_fill_2
XFILLER_3_62 vgnd vpwr scs8hd_decap_3
XANTENNA__189__A _189_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__099__A _098_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_220 vgnd vpwr scs8hd_decap_12
X_222_ chanx_right_in[5] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_6_124 vpwr vgnd scs8hd_fill_2
XFILLER_6_135 vpwr vgnd scs8hd_fill_2
X_153_ _135_/Y _169_/A _127_/C _153_/X vgnd vpwr scs8hd_or3_4
XFILLER_8_18 vpwr vgnd scs8hd_fill_2
XFILLER_8_29 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_5.LATCH_1_.latch data_in _191_/A _172_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_084_ address[0] _105_/C vgnd vpwr scs8hd_inv_8
XFILLER_12_93 vgnd vpwr scs8hd_decap_4
XFILLER_19_7 vgnd vpwr scs8hd_fill_1
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
XANTENNA__175__C _127_/C vgnd vpwr scs8hd_diode_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _218_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_116 vgnd vpwr scs8hd_decap_4
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XFILLER_15_245 vgnd vpwr scs8hd_decap_3
X_205_ _205_/HI _205_/LO vgnd vpwr scs8hd_conb_1
X_136_ address[5] _169_/A vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_6 vpwr vgnd scs8hd_fill_2
XANTENNA__186__B _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_41 vpwr vgnd scs8hd_fill_2
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XFILLER_21_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_108 vpwr vgnd scs8hd_fill_2
XFILLER_12_215 vgnd vpwr scs8hd_fill_1
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
X_119_ _130_/A _120_/B _119_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__172__D _165_/X vgnd vpwr scs8hd_diode_2
XFILLER_38_178 vgnd vpwr scs8hd_decap_12
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_47 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A right_top_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_20_93 vpwr vgnd scs8hd_fill_2
XFILLER_35_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__183__C _127_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_84 vpwr vgnd scs8hd_fill_2
XFILLER_26_115 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_258 vgnd vpwr scs8hd_decap_4
XFILLER_1_225 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _187_/Y mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_32_129 vgnd vpwr scs8hd_decap_12
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_107 vpwr vgnd scs8hd_fill_2
XFILLER_14_118 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_140 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _217_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_100 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_155 vgnd vpwr scs8hd_fill_1
XFILLER_13_184 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_74 vpwr vgnd scs8hd_fill_2
XFILLER_3_30 vpwr vgnd scs8hd_fill_2
XANTENNA__180__D _167_/X vgnd vpwr scs8hd_diode_2
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[4] mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_28 vgnd vpwr scs8hd_decap_3
XANTENNA__099__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_27_232 vgnd vpwr scs8hd_decap_12
X_083_ address[2] _083_/Y vgnd vpwr scs8hd_inv_8
X_221_ chanx_right_in[6] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
X_152_ _123_/A _146_/X _152_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_154 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XANTENNA__175__D _167_/X vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_13.LATCH_1_.latch data_in _199_/A _181_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_202 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.INVTX1_1_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
X_204_ _204_/A _204_/Y vgnd vpwr scs8hd_inv_8
XFILLER_15_235 vgnd vpwr scs8hd_decap_3
XFILLER_15_257 vpwr vgnd scs8hd_fill_2
XFILLER_15_268 vpwr vgnd scs8hd_fill_2
X_135_ address[6] _135_/Y vgnd vpwr scs8hd_inv_8
XFILLER_23_82 vpwr vgnd scs8hd_fill_2
XFILLER_2_194 vpwr vgnd scs8hd_fill_2
XFILLER_2_150 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__186__C _164_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_249 vgnd vpwr scs8hd_decap_4
XFILLER_21_216 vpwr vgnd scs8hd_fill_2
XFILLER_21_205 vgnd vpwr scs8hd_decap_8
XFILLER_12_238 vgnd vpwr scs8hd_decap_6
XFILLER_20_271 vgnd vpwr scs8hd_decap_4
XFILLER_18_71 vpwr vgnd scs8hd_fill_2
XFILLER_18_93 vgnd vpwr scs8hd_decap_8
XFILLER_11_260 vpwr vgnd scs8hd_fill_2
X_118_ _129_/A _120_/B _118_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_3 vgnd vpwr scs8hd_decap_4
XFILLER_30_17 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XFILLER_29_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_6_.scs8hd_inv_1 left_top_grid_pin_9_ mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_20_61 vgnd vpwr scs8hd_fill_1
XFILLER_29_81 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_15.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__183__D _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_41 vgnd vpwr scs8hd_decap_4
XFILLER_6_96 vpwr vgnd scs8hd_fill_2
XFILLER_26_127 vpwr vgnd scs8hd_fill_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
Xmux_right_track_0.INVTX1_2_.scs8hd_inv_1 right_top_grid_pin_13_ mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_237 vgnd vpwr scs8hd_decap_4
XFILLER_25_171 vgnd vpwr scs8hd_fill_1
XFILLER_15_50 vpwr vgnd scs8hd_fill_2
XFILLER_40_141 vgnd vpwr scs8hd_decap_12
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
XFILLER_39_263 vgnd vpwr scs8hd_decap_12
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XFILLER_22_196 vpwr vgnd scs8hd_fill_2
XFILLER_22_163 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_2_.latch data_in mem_left_track_17.LATCH_2_.latch/Q _158_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_123 vpwr vgnd scs8hd_fill_2
XFILLER_13_152 vpwr vgnd scs8hd_fill_2
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
XANTENNA__099__C _165_/A vgnd vpwr scs8hd_diode_2
X_220_ _220_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_6_104 vgnd vpwr scs8hd_decap_3
XFILLER_6_148 vgnd vpwr scs8hd_decap_4
X_151_ _122_/A _146_/X _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_144 vgnd vpwr scs8hd_decap_6
XFILLER_12_84 vgnd vpwr scs8hd_decap_3
XFILLER_18_200 vgnd vpwr scs8hd_decap_3
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_170 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ _190_/Y mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _214_/HI mem_left_track_1.LATCH_2_.latch/Q
+ mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _195_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_214 vpwr vgnd scs8hd_fill_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
X_203_ _203_/A _203_/Y vgnd vpwr scs8hd_inv_8
X_134_ _123_/A _129_/B _134_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_140 vgnd vpwr scs8hd_decap_4
Xmux_right_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[5] mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_10 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_1_.latch data_in _187_/A _166_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_228 vgnd vpwr scs8hd_decap_4
XANTENNA__186__D _095_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _199_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_206 vpwr vgnd scs8hd_fill_2
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.INVTX1_1_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_272 vgnd vpwr scs8hd_decap_4
X_117_ _116_/X _120_/B vgnd vpwr scs8hd_buf_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_0_.latch data_in mem_left_track_1.LATCH_0_.latch/Q _144_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_3 vpwr vgnd scs8hd_fill_2
XFILLER_30_29 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_84 vgnd vpwr scs8hd_decap_6
XFILLER_4_202 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_93 vgnd vpwr scs8hd_decap_12
XFILLER_29_60 vgnd vpwr scs8hd_fill_1
Xmem_right_track_16.LATCH_1_.latch data_in mem_right_track_16.LATCH_1_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_29 vpwr vgnd scs8hd_fill_2
XFILLER_25_18 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_25_150 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__102__A _098_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_275 vpwr vgnd scs8hd_fill_2
XFILLER_39_253 vpwr vgnd scs8hd_fill_2
XFILLER_39_220 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[7] mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_186 vgnd vpwr scs8hd_fill_1
XFILLER_22_175 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[2] mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_131 vpwr vgnd scs8hd_fill_2
XFILLER_13_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _201_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_87 vpwr vgnd scs8hd_fill_2
XFILLER_3_10 vgnd vpwr scs8hd_decap_3
XFILLER_27_245 vgnd vpwr scs8hd_fill_1
X_150_ _121_/A _146_/X _150_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_259 vgnd vpwr scs8hd_decap_12
XFILLER_24_248 vgnd vpwr scs8hd_decap_8
XFILLER_3_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__200__A _200_/A vgnd vpwr scs8hd_diode_2
X_133_ _122_/A _129_/B _133_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_95 vpwr vgnd scs8hd_fill_2
XFILLER_23_62 vgnd vpwr scs8hd_decap_4
X_202_ _202_/A _202_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_163 vgnd vpwr scs8hd_decap_4
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__110__A _097_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_66 vpwr vgnd scs8hd_fill_2
XFILLER_9_42 vpwr vgnd scs8hd_fill_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XFILLER_9_75 vpwr vgnd scs8hd_fill_2
XFILLER_28_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _187_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_84 vpwr vgnd scs8hd_fill_2
X_116_ _161_/A _162_/A _116_/C _116_/X vgnd vpwr scs8hd_or3_4
XANTENNA__105__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_7_233 vgnd vpwr scs8hd_fill_1
XFILLER_7_255 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_159 vgnd vpwr scs8hd_decap_12
XFILLER_6_10 vgnd vpwr scs8hd_fill_1
XFILLER_6_32 vpwr vgnd scs8hd_fill_2
XFILLER_26_107 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_3.INVTX1_1_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_170 vgnd vpwr scs8hd_decap_3
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_right_track_0.LATCH_0_.latch data_in mem_right_track_0.LATCH_0_.latch/Q _110_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XANTENNA__102__B address[2] vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_31_110 vgnd vpwr scs8hd_decap_12
XFILLER_16_173 vgnd vpwr scs8hd_fill_1
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_195 vpwr vgnd scs8hd_fill_2
XFILLER_39_232 vgnd vpwr scs8hd_decap_12
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_9_136 vpwr vgnd scs8hd_fill_2
XFILLER_9_147 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_257 vgnd vpwr scs8hd_decap_12
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_10_102 vgnd vpwr scs8hd_decap_6
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _237_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_3 vpwr vgnd scs8hd_fill_2
XFILLER_6_139 vgnd vpwr scs8hd_decap_6
XFILLER_12_42 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__108__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
X_132_ _121_/A _129_/B _132_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_52 vgnd vpwr scs8hd_decap_4
X_201_ _201_/A _201_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _229_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_45 vpwr vgnd scs8hd_fill_2
XANTENNA__110__B _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_12_219 vgnd vpwr scs8hd_decap_4
XFILLER_11_241 vgnd vpwr scs8hd_fill_1
XANTENNA__105__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_7_212 vpwr vgnd scs8hd_fill_2
XFILLER_7_245 vgnd vpwr scs8hd_fill_1
XFILLER_7_267 vpwr vgnd scs8hd_fill_2
X_115_ _114_/X _116_/C vgnd vpwr scs8hd_buf_1
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A left_top_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__121__A _121_/A vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_1_.latch data_in mem_left_track_9.LATCH_1_.latch/Q _151_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB _097_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_171 vgnd vpwr scs8hd_decap_12
XFILLER_4_226 vgnd vpwr scs8hd_decap_3
XFILLER_20_97 vgnd vpwr scs8hd_fill_1
XFILLER_20_53 vgnd vpwr scs8hd_decap_8
XFILLER_28_160 vgnd vpwr scs8hd_decap_12
XANTENNA__116__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_3 vgnd vpwr scs8hd_decap_3
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_right_track_8.LATCH_4_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_25_163 vpwr vgnd scs8hd_fill_2
XFILLER_15_75 vgnd vpwr scs8hd_fill_1
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
XANTENNA__102__C _095_/C vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_273 vgnd vpwr scs8hd_decap_4
XFILLER_0_240 vpwr vgnd scs8hd_fill_2
XFILLER_16_141 vpwr vgnd scs8hd_fill_2
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
.ends

