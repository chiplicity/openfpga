magic
tech EFS8A
magscale 1 2
timestamp 1602530114
<< locali >>
rect 6009 23647 6043 23749
rect 6745 23137 6906 23171
rect 22511 23137 22546 23171
rect 6745 22967 6779 23137
rect 9631 22049 9758 22083
rect 7843 21097 7849 21131
rect 19067 21097 19073 21131
rect 7843 21029 7877 21097
rect 19067 21029 19101 21097
rect 10885 20383 10919 20553
rect 20855 19873 20982 19907
rect 6469 19159 6503 19261
rect 11707 18921 11713 18955
rect 11707 18853 11741 18921
rect 6009 18071 6043 18173
rect 18515 17833 18521 17867
rect 7791 17765 7836 17799
rect 18515 17765 18549 17833
rect 9321 17119 9355 17289
rect 11707 15657 11713 15691
rect 3341 15419 3375 15657
rect 11707 15589 11741 15657
rect 3709 15351 3743 15521
rect 12075 14569 12081 14603
rect 12075 14501 12109 14569
rect 22971 14433 23006 14467
rect 3893 13719 3927 13889
rect 4813 13175 4847 13277
rect 18699 12631 18733 12699
rect 18699 12597 18705 12631
rect 17233 11611 17267 11781
rect 13087 11543 13121 11611
rect 13087 11509 13093 11543
rect 13455 11305 13461 11339
rect 6135 11237 6180 11271
rect 13455 11237 13489 11305
rect 20855 11169 20982 11203
rect 5457 10999 5491 11101
rect 15439 10217 15577 10251
rect 1547 10149 1685 10183
rect 14231 10081 14266 10115
rect 15243 10081 15370 10115
rect 8079 2601 8217 2635
rect 21327 2601 21465 2635
<< viali >>
rect 11596 25313 11630 25347
rect 12700 25313 12734 25347
rect 11667 25109 11701 25143
rect 12771 25109 12805 25143
rect 12725 24905 12759 24939
rect 13093 24905 13127 24939
rect 1460 24701 1494 24735
rect 1869 24701 1903 24735
rect 11412 24701 11446 24735
rect 12909 24701 12943 24735
rect 13461 24701 13495 24735
rect 14800 24701 14834 24735
rect 15209 24701 15243 24735
rect 1547 24633 1581 24667
rect 11897 24633 11931 24667
rect 14887 24633 14921 24667
rect 11483 24565 11517 24599
rect 12173 24565 12207 24599
rect 11621 24361 11655 24395
rect 13461 24361 13495 24395
rect 1476 24225 1510 24259
rect 5917 24225 5951 24259
rect 6929 24225 6963 24259
rect 11437 24225 11471 24259
rect 13277 24225 13311 24259
rect 15368 24225 15402 24259
rect 16380 24225 16414 24259
rect 17392 24225 17426 24259
rect 18404 24225 18438 24259
rect 20980 24225 21014 24259
rect 2421 24157 2455 24191
rect 6101 24089 6135 24123
rect 15945 24089 15979 24123
rect 17463 24089 17497 24123
rect 1547 24021 1581 24055
rect 7113 24021 7147 24055
rect 10609 24021 10643 24055
rect 14197 24021 14231 24055
rect 15439 24021 15473 24055
rect 16451 24021 16485 24055
rect 18475 24021 18509 24055
rect 21051 24021 21085 24055
rect 2329 23817 2363 23851
rect 5825 23817 5859 23851
rect 11529 23817 11563 23851
rect 13461 23817 13495 23851
rect 15393 23817 15427 23851
rect 18245 23817 18279 23851
rect 19901 23817 19935 23851
rect 21465 23817 21499 23851
rect 21833 23817 21867 23851
rect 25145 23817 25179 23851
rect 6009 23749 6043 23783
rect 6285 23749 6319 23783
rect 17417 23749 17451 23783
rect 18613 23749 18647 23783
rect 6561 23681 6595 23715
rect 12541 23681 12575 23715
rect 12817 23681 12851 23715
rect 14657 23681 14691 23715
rect 15945 23681 15979 23715
rect 16221 23681 16255 23715
rect 1409 23613 1443 23647
rect 1961 23613 1995 23647
rect 2548 23613 2582 23647
rect 2973 23613 3007 23647
rect 3560 23613 3594 23647
rect 3985 23613 4019 23647
rect 5641 23613 5675 23647
rect 6009 23613 6043 23647
rect 7424 23613 7458 23647
rect 7849 23613 7883 23647
rect 8468 23613 8502 23647
rect 8861 23613 8895 23647
rect 10609 23613 10643 23647
rect 10977 23613 11011 23647
rect 14013 23613 14047 23647
rect 14105 23613 14139 23647
rect 14565 23613 14599 23647
rect 17877 23613 17911 23647
rect 18061 23613 18095 23647
rect 19717 23613 19751 23647
rect 20269 23613 20303 23647
rect 20980 23613 21014 23647
rect 24660 23613 24694 23647
rect 2651 23545 2685 23579
rect 7021 23545 7055 23579
rect 11253 23545 11287 23579
rect 12633 23545 12667 23579
rect 16037 23545 16071 23579
rect 16957 23545 16991 23579
rect 1593 23477 1627 23511
rect 3663 23477 3697 23511
rect 7527 23477 7561 23511
rect 8539 23477 8573 23511
rect 10425 23477 10459 23511
rect 12265 23477 12299 23511
rect 15761 23477 15795 23511
rect 21051 23477 21085 23511
rect 24731 23477 24765 23511
rect 8677 23273 8711 23307
rect 12541 23273 12575 23307
rect 16313 23273 16347 23307
rect 18889 23273 18923 23307
rect 6975 23205 7009 23239
rect 11621 23205 11655 23239
rect 15485 23205 15519 23239
rect 16957 23205 16991 23239
rect 17049 23205 17083 23239
rect 21097 23205 21131 23239
rect 1409 23137 1443 23171
rect 2580 23137 2614 23171
rect 4788 23137 4822 23171
rect 7916 23137 7950 23171
rect 13737 23137 13771 23171
rect 14197 23137 14231 23171
rect 18464 23137 18498 23171
rect 22477 23137 22511 23171
rect 5733 23069 5767 23103
rect 10425 23069 10459 23103
rect 11529 23069 11563 23103
rect 14381 23069 14415 23103
rect 15393 23069 15427 23103
rect 15669 23069 15703 23103
rect 17233 23069 17267 23103
rect 21005 23069 21039 23103
rect 21281 23069 21315 23103
rect 7987 23001 8021 23035
rect 12081 23001 12115 23035
rect 1593 22933 1627 22967
rect 2053 22933 2087 22967
rect 2651 22933 2685 22967
rect 4859 22933 4893 22967
rect 5273 22933 5307 22967
rect 6745 22933 6779 22967
rect 8401 22933 8435 22967
rect 12817 22933 12851 22967
rect 18567 22933 18601 22967
rect 22615 22933 22649 22967
rect 2789 22729 2823 22763
rect 11713 22729 11747 22763
rect 13737 22729 13771 22763
rect 17233 22729 17267 22763
rect 18245 22729 18279 22763
rect 21649 22729 21683 22763
rect 22569 22729 22603 22763
rect 4813 22661 4847 22695
rect 13093 22661 13127 22695
rect 19073 22661 19107 22695
rect 21373 22661 21407 22695
rect 8309 22593 8343 22627
rect 14381 22593 14415 22627
rect 15025 22593 15059 22627
rect 15945 22593 15979 22627
rect 16221 22593 16255 22627
rect 16957 22593 16991 22627
rect 18521 22593 18555 22627
rect 20361 22593 20395 22627
rect 21005 22593 21039 22627
rect 1961 22525 1995 22559
rect 3341 22525 3375 22559
rect 3801 22525 3835 22559
rect 5273 22525 5307 22559
rect 7272 22525 7306 22559
rect 10609 22525 10643 22559
rect 10977 22525 11011 22559
rect 11253 22525 11287 22559
rect 1777 22457 1811 22491
rect 5917 22457 5951 22491
rect 8401 22457 8435 22491
rect 8953 22457 8987 22491
rect 12541 22457 12575 22491
rect 12633 22457 12667 22491
rect 14473 22457 14507 22491
rect 15393 22457 15427 22491
rect 15761 22457 15795 22491
rect 16037 22457 16071 22491
rect 17877 22457 17911 22491
rect 18613 22457 18647 22491
rect 20085 22457 20119 22491
rect 20453 22457 20487 22491
rect 1685 22389 1719 22423
rect 3525 22389 3559 22423
rect 7021 22389 7055 22423
rect 7343 22389 7377 22423
rect 7757 22389 7791 22423
rect 8033 22389 8067 22423
rect 10977 22389 11011 22423
rect 12173 22389 12207 22423
rect 14105 22389 14139 22423
rect 7849 22185 7883 22219
rect 12081 22185 12115 22219
rect 12541 22185 12575 22219
rect 14657 22185 14691 22219
rect 15117 22185 15151 22219
rect 20361 22185 20395 22219
rect 1869 22117 1903 22151
rect 6101 22117 6135 22151
rect 6193 22117 6227 22151
rect 8125 22117 8159 22151
rect 8217 22117 8251 22151
rect 11482 22117 11516 22151
rect 13093 22117 13127 22151
rect 14289 22117 14323 22151
rect 15577 22117 15611 22151
rect 16129 22117 16163 22151
rect 18337 22117 18371 22151
rect 18429 22117 18463 22151
rect 21097 22117 21131 22151
rect 4629 22049 4663 22083
rect 9597 22049 9631 22083
rect 1777 21981 1811 22015
rect 2421 21981 2455 22015
rect 3065 21981 3099 22015
rect 6377 21981 6411 22015
rect 8769 21981 8803 22015
rect 11161 21981 11195 22015
rect 13001 21981 13035 22015
rect 13277 21981 13311 22015
rect 15485 21981 15519 22015
rect 16957 21981 16991 22015
rect 18981 21981 19015 22015
rect 21005 21981 21039 22015
rect 21281 21981 21315 22015
rect 2697 21913 2731 21947
rect 13921 21913 13955 21947
rect 19901 21913 19935 21947
rect 3617 21845 3651 21879
rect 4721 21845 4755 21879
rect 5549 21845 5583 21879
rect 9827 21845 9861 21879
rect 10149 21845 10183 21879
rect 10793 21845 10827 21879
rect 16405 21845 16439 21879
rect 18061 21845 18095 21879
rect 1777 21641 1811 21675
rect 4629 21641 4663 21675
rect 5089 21641 5123 21675
rect 6193 21641 6227 21675
rect 11529 21641 11563 21675
rect 15577 21641 15611 21675
rect 15945 21641 15979 21675
rect 17509 21641 17543 21675
rect 18981 21641 19015 21675
rect 20913 21641 20947 21675
rect 21925 21641 21959 21675
rect 25145 21641 25179 21675
rect 2973 21573 3007 21607
rect 21511 21573 21545 21607
rect 2053 21505 2087 21539
rect 2513 21505 2547 21539
rect 3893 21505 3927 21539
rect 5273 21505 5307 21539
rect 5917 21505 5951 21539
rect 8493 21505 8527 21539
rect 8769 21505 8803 21539
rect 10333 21505 10367 21539
rect 12541 21505 12575 21539
rect 13185 21505 13219 21539
rect 14657 21505 14691 21539
rect 17141 21505 17175 21539
rect 18061 21505 18095 21539
rect 19901 21505 19935 21539
rect 6653 21437 6687 21471
rect 6837 21437 6871 21471
rect 7297 21437 7331 21471
rect 16497 21437 16531 21471
rect 16865 21437 16899 21471
rect 21440 21437 21474 21471
rect 24660 21437 24694 21471
rect 2145 21369 2179 21403
rect 3341 21369 3375 21403
rect 3617 21369 3651 21403
rect 3709 21369 3743 21403
rect 5365 21369 5399 21403
rect 7573 21369 7607 21403
rect 8585 21369 8619 21403
rect 10057 21369 10091 21403
rect 10149 21369 10183 21403
rect 12633 21369 12667 21403
rect 13829 21369 13863 21403
rect 15019 21369 15053 21403
rect 16313 21369 16347 21403
rect 18382 21369 18416 21403
rect 19993 21369 20027 21403
rect 20545 21369 20579 21403
rect 8033 21301 8067 21335
rect 9689 21301 9723 21335
rect 11253 21301 11287 21335
rect 12173 21301 12207 21335
rect 13461 21301 13495 21335
rect 14565 21301 14599 21335
rect 17785 21301 17819 21335
rect 19717 21301 19751 21335
rect 24731 21301 24765 21335
rect 3709 21097 3743 21131
rect 5825 21097 5859 21131
rect 6101 21097 6135 21131
rect 6837 21097 6871 21131
rect 7849 21097 7883 21131
rect 9045 21097 9079 21131
rect 11989 21097 12023 21131
rect 14657 21097 14691 21131
rect 15117 21097 15151 21131
rect 16221 21097 16255 21131
rect 16589 21097 16623 21131
rect 18337 21097 18371 21131
rect 19073 21097 19107 21131
rect 19625 21097 19659 21131
rect 19993 21097 20027 21131
rect 21373 21097 21407 21131
rect 1777 21029 1811 21063
rect 2053 21029 2087 21063
rect 2605 21029 2639 21063
rect 3249 21029 3283 21063
rect 5226 21029 5260 21063
rect 10149 21029 10183 21063
rect 11431 21029 11465 21063
rect 13179 21029 13213 21063
rect 15622 21029 15656 21063
rect 9724 20961 9758 20995
rect 11069 20961 11103 20995
rect 15301 20961 15335 20995
rect 17141 20961 17175 20995
rect 17601 20961 17635 20995
rect 1961 20893 1995 20927
rect 4905 20893 4939 20927
rect 7481 20893 7515 20927
rect 12817 20893 12851 20927
rect 17877 20893 17911 20927
rect 18705 20893 18739 20927
rect 20913 20893 20947 20927
rect 2973 20757 3007 20791
rect 8401 20757 8435 20791
rect 8769 20757 8803 20791
rect 9827 20757 9861 20791
rect 12541 20757 12575 20791
rect 13737 20757 13771 20791
rect 14105 20757 14139 20791
rect 1593 20553 1627 20587
rect 4629 20553 4663 20587
rect 10885 20553 10919 20587
rect 11069 20553 11103 20587
rect 13829 20553 13863 20587
rect 16773 20553 16807 20587
rect 17141 20553 17175 20587
rect 18981 20553 19015 20587
rect 21281 20553 21315 20587
rect 3801 20485 3835 20519
rect 6101 20485 6135 20519
rect 10241 20485 10275 20519
rect 2881 20417 2915 20451
rect 3341 20417 3375 20451
rect 5181 20417 5215 20451
rect 5549 20417 5583 20451
rect 7389 20417 7423 20451
rect 16405 20485 16439 20519
rect 11299 20417 11333 20451
rect 12541 20417 12575 20451
rect 12817 20417 12851 20451
rect 15853 20417 15887 20451
rect 18061 20417 18095 20451
rect 19809 20417 19843 20451
rect 19993 20417 20027 20451
rect 20637 20417 20671 20451
rect 21833 20417 21867 20451
rect 1409 20349 1443 20383
rect 6904 20349 6938 20383
rect 7849 20349 7883 20383
rect 10885 20349 10919 20383
rect 11196 20349 11230 20383
rect 11621 20349 11655 20383
rect 14105 20349 14139 20383
rect 14473 20349 14507 20383
rect 2973 20281 3007 20315
rect 4905 20281 4939 20315
rect 5273 20281 5307 20315
rect 7665 20281 7699 20315
rect 8170 20281 8204 20315
rect 9689 20281 9723 20315
rect 9781 20281 9815 20315
rect 12265 20281 12299 20315
rect 12633 20281 12667 20315
rect 15945 20281 15979 20315
rect 18382 20281 18416 20315
rect 19257 20281 19291 20315
rect 20085 20281 20119 20315
rect 21557 20281 21591 20315
rect 21649 20281 21683 20315
rect 1961 20213 1995 20247
rect 2421 20213 2455 20247
rect 4261 20213 4295 20247
rect 6975 20213 7009 20247
rect 8769 20213 8803 20247
rect 9137 20213 9171 20247
rect 9413 20213 9447 20247
rect 10609 20213 10643 20247
rect 13553 20213 13587 20247
rect 14105 20213 14139 20247
rect 15393 20213 15427 20247
rect 17785 20213 17819 20247
rect 1547 20009 1581 20043
rect 5641 20009 5675 20043
rect 5917 20009 5951 20043
rect 7481 20009 7515 20043
rect 7849 20009 7883 20043
rect 9781 20009 9815 20043
rect 11069 20009 11103 20043
rect 12817 20009 12851 20043
rect 15025 20009 15059 20043
rect 18613 20009 18647 20043
rect 19257 20009 19291 20043
rect 20269 20009 20303 20043
rect 21051 20009 21085 20043
rect 21557 20009 21591 20043
rect 2513 19941 2547 19975
rect 2605 19941 2639 19975
rect 5042 19941 5076 19975
rect 8125 19941 8159 19975
rect 8217 19941 8251 19975
rect 8769 19941 8803 19975
rect 9505 19941 9539 19975
rect 11983 19941 12017 19975
rect 15663 19941 15697 19975
rect 18337 19941 18371 19975
rect 18981 19941 19015 19975
rect 1476 19873 1510 19907
rect 6561 19873 6595 19907
rect 9689 19873 9723 19907
rect 10241 19873 10275 19907
rect 12541 19873 12575 19907
rect 13645 19873 13679 19907
rect 14197 19873 14231 19907
rect 17601 19873 17635 19907
rect 18061 19873 18095 19907
rect 19165 19873 19199 19907
rect 19625 19873 19659 19907
rect 20821 19873 20855 19907
rect 24660 19873 24694 19907
rect 3157 19805 3191 19839
rect 4721 19805 4755 19839
rect 6469 19805 6503 19839
rect 11621 19805 11655 19839
rect 14381 19805 14415 19839
rect 15301 19805 15335 19839
rect 16497 19737 16531 19771
rect 2145 19669 2179 19703
rect 3433 19669 3467 19703
rect 3801 19669 3835 19703
rect 4537 19669 4571 19703
rect 14749 19669 14783 19703
rect 16221 19669 16255 19703
rect 24731 19669 24765 19703
rect 2973 19465 3007 19499
rect 3249 19465 3283 19499
rect 3709 19465 3743 19499
rect 6285 19465 6319 19499
rect 9413 19465 9447 19499
rect 15393 19465 15427 19499
rect 16589 19465 16623 19499
rect 17417 19465 17451 19499
rect 19625 19465 19659 19499
rect 25145 19465 25179 19499
rect 25513 19465 25547 19499
rect 13093 19397 13127 19431
rect 17049 19397 17083 19431
rect 18981 19397 19015 19431
rect 1685 19329 1719 19363
rect 2053 19329 2087 19363
rect 4353 19329 4387 19363
rect 5549 19329 5583 19363
rect 8401 19329 8435 19363
rect 9965 19329 9999 19363
rect 11345 19329 11379 19363
rect 13553 19329 13587 19363
rect 15669 19329 15703 19363
rect 19901 19329 19935 19363
rect 20545 19329 20579 19363
rect 21511 19329 21545 19363
rect 3985 19261 4019 19295
rect 4721 19261 4755 19295
rect 4997 19261 5031 19295
rect 6469 19261 6503 19295
rect 7021 19261 7055 19295
rect 7389 19261 7423 19295
rect 14013 19261 14047 19295
rect 14473 19261 14507 19295
rect 17785 19261 17819 19295
rect 18061 19261 18095 19295
rect 21424 19261 21458 19295
rect 21925 19261 21959 19295
rect 24660 19261 24694 19295
rect 2415 19193 2449 19227
rect 3801 19193 3835 19227
rect 5273 19193 5307 19227
rect 5365 19193 5399 19227
rect 6837 19193 6871 19227
rect 7665 19193 7699 19227
rect 8493 19193 8527 19227
rect 9045 19193 9079 19227
rect 10057 19193 10091 19227
rect 10609 19193 10643 19227
rect 12541 19193 12575 19227
rect 12633 19193 12667 19227
rect 15761 19193 15795 19227
rect 16313 19193 16347 19227
rect 18382 19193 18416 19227
rect 19993 19193 20027 19227
rect 6469 19125 6503 19159
rect 6561 19125 6595 19159
rect 8217 19125 8251 19159
rect 9689 19125 9723 19159
rect 10885 19125 10919 19159
rect 11713 19125 11747 19159
rect 12265 19125 12299 19159
rect 13829 19125 13863 19159
rect 14105 19125 14139 19159
rect 19257 19125 19291 19159
rect 20913 19125 20947 19159
rect 24731 19125 24765 19159
rect 2605 18921 2639 18955
rect 4445 18921 4479 18955
rect 6193 18921 6227 18955
rect 7205 18921 7239 18955
rect 9137 18921 9171 18955
rect 11713 18921 11747 18955
rect 15025 18921 15059 18955
rect 18521 18921 18555 18955
rect 2047 18853 2081 18887
rect 8217 18853 8251 18887
rect 9781 18853 9815 18887
rect 9873 18853 9907 18887
rect 12633 18853 12667 18887
rect 13277 18853 13311 18887
rect 15761 18853 15795 18887
rect 19165 18853 19199 18887
rect 19717 18853 19751 18887
rect 1685 18785 1719 18819
rect 4629 18785 4663 18819
rect 5181 18785 5215 18819
rect 5365 18785 5399 18819
rect 6285 18785 6319 18819
rect 6469 18785 6503 18819
rect 7573 18785 7607 18819
rect 10793 18785 10827 18819
rect 12265 18785 12299 18819
rect 17693 18785 17727 18819
rect 17877 18785 17911 18819
rect 2973 18717 3007 18751
rect 5733 18717 5767 18751
rect 6837 18717 6871 18751
rect 8125 18717 8159 18751
rect 8769 18717 8803 18751
rect 11345 18717 11379 18751
rect 13185 18717 13219 18751
rect 15669 18717 15703 18751
rect 16037 18717 16071 18751
rect 18153 18717 18187 18751
rect 18797 18717 18831 18751
rect 19073 18717 19107 18751
rect 20913 18717 20947 18751
rect 10333 18649 10367 18683
rect 13737 18649 13771 18683
rect 14565 18649 14599 18683
rect 3341 18581 3375 18615
rect 3617 18581 3651 18615
rect 7849 18581 7883 18615
rect 13001 18581 13035 18615
rect 14197 18581 14231 18615
rect 19993 18581 20027 18615
rect 2697 18377 2731 18411
rect 2973 18377 3007 18411
rect 3985 18377 4019 18411
rect 4353 18377 4387 18411
rect 6561 18377 6595 18411
rect 7757 18377 7791 18411
rect 10609 18377 10643 18411
rect 11989 18377 12023 18411
rect 13829 18377 13863 18411
rect 17509 18377 17543 18411
rect 18521 18377 18555 18411
rect 19625 18377 19659 18411
rect 10241 18309 10275 18343
rect 13093 18309 13127 18343
rect 19901 18309 19935 18343
rect 2513 18241 2547 18275
rect 3525 18241 3559 18275
rect 9689 18241 9723 18275
rect 11299 18241 11333 18275
rect 12541 18241 12575 18275
rect 16497 18241 16531 18275
rect 16773 18241 16807 18275
rect 18705 18241 18739 18275
rect 20821 18241 20855 18275
rect 1869 18173 1903 18207
rect 2421 18173 2455 18207
rect 4629 18173 4663 18207
rect 5273 18173 5307 18207
rect 5457 18173 5491 18207
rect 5825 18173 5859 18207
rect 6009 18173 6043 18207
rect 6872 18173 6906 18207
rect 7297 18173 7331 18207
rect 7849 18173 7883 18207
rect 8769 18173 8803 18207
rect 11212 18173 11246 18207
rect 11621 18173 11655 18207
rect 14657 18173 14691 18207
rect 8170 18105 8204 18139
rect 9137 18105 9171 18139
rect 9505 18105 9539 18139
rect 9781 18105 9815 18139
rect 12633 18105 12667 18139
rect 14565 18105 14599 18139
rect 14978 18105 15012 18139
rect 16589 18105 16623 18139
rect 19026 18105 19060 18139
rect 20545 18105 20579 18139
rect 20637 18105 20671 18139
rect 4537 18037 4571 18071
rect 6009 18037 6043 18071
rect 6193 18037 6227 18071
rect 6975 18037 7009 18071
rect 10977 18037 11011 18071
rect 13553 18037 13587 18071
rect 15577 18037 15611 18071
rect 15853 18037 15887 18071
rect 16221 18037 16255 18071
rect 17877 18037 17911 18071
rect 20361 18037 20395 18071
rect 2605 17833 2639 17867
rect 2973 17833 3007 17867
rect 3893 17833 3927 17867
rect 4813 17833 4847 17867
rect 7389 17833 7423 17867
rect 8401 17833 8435 17867
rect 8677 17833 8711 17867
rect 9965 17833 9999 17867
rect 11345 17833 11379 17867
rect 11621 17833 11655 17867
rect 16221 17833 16255 17867
rect 16497 17833 16531 17867
rect 17233 17833 17267 17867
rect 18521 17833 18555 17867
rect 19073 17833 19107 17867
rect 19349 17833 19383 17867
rect 20545 17833 20579 17867
rect 5733 17765 5767 17799
rect 6929 17765 6963 17799
rect 7757 17765 7791 17799
rect 10977 17765 11011 17799
rect 11989 17765 12023 17799
rect 15663 17765 15697 17799
rect 1777 17697 1811 17731
rect 2329 17697 2363 17731
rect 2513 17697 2547 17731
rect 4353 17697 4387 17731
rect 4629 17697 4663 17731
rect 6101 17697 6135 17731
rect 6469 17697 6503 17731
rect 10241 17697 10275 17731
rect 10701 17697 10735 17731
rect 13645 17697 13679 17731
rect 14105 17697 14139 17731
rect 15117 17697 15151 17731
rect 17049 17697 17083 17731
rect 20980 17697 21014 17731
rect 4445 17629 4479 17663
rect 6653 17629 6687 17663
rect 7481 17629 7515 17663
rect 11897 17629 11931 17663
rect 12173 17629 12207 17663
rect 14381 17629 14415 17663
rect 15301 17629 15335 17663
rect 18153 17629 18187 17663
rect 14749 17561 14783 17595
rect 3433 17493 3467 17527
rect 5457 17493 5491 17527
rect 12909 17493 12943 17527
rect 21051 17493 21085 17527
rect 1685 17289 1719 17323
rect 5641 17289 5675 17323
rect 6193 17289 6227 17323
rect 7941 17289 7975 17323
rect 8309 17289 8343 17323
rect 9321 17289 9355 17323
rect 9505 17289 9539 17323
rect 16313 17289 16347 17323
rect 17049 17289 17083 17323
rect 17509 17289 17543 17323
rect 19441 17289 19475 17323
rect 20039 17289 20073 17323
rect 21051 17289 21085 17323
rect 25145 17289 25179 17323
rect 4077 17221 4111 17255
rect 4813 17221 4847 17255
rect 9137 17221 9171 17255
rect 2053 17153 2087 17187
rect 3617 17153 3651 17187
rect 3948 17153 3982 17187
rect 4169 17153 4203 17187
rect 4537 17153 4571 17187
rect 7665 17153 7699 17187
rect 8585 17153 8619 17187
rect 17877 17221 17911 17255
rect 18981 17221 19015 17255
rect 10885 17153 10919 17187
rect 11529 17153 11563 17187
rect 12817 17153 12851 17187
rect 18429 17153 18463 17187
rect 2881 17085 2915 17119
rect 2973 17085 3007 17119
rect 5181 17085 5215 17119
rect 5549 17085 5583 17119
rect 6653 17085 6687 17119
rect 7205 17085 7239 17119
rect 7389 17085 7423 17119
rect 9321 17085 9355 17119
rect 10609 17085 10643 17119
rect 14749 17085 14783 17119
rect 16564 17085 16598 17119
rect 19968 17085 20002 17119
rect 20980 17085 21014 17119
rect 21373 17085 21407 17119
rect 21741 17085 21775 17119
rect 24660 17085 24694 17119
rect 3341 17017 3375 17051
rect 3801 17017 3835 17051
rect 5365 17017 5399 17051
rect 8677 17017 8711 17051
rect 9965 17017 9999 17051
rect 10977 17017 11011 17051
rect 12541 17017 12575 17051
rect 12633 17017 12667 17051
rect 14657 17017 14691 17051
rect 15111 17017 15145 17051
rect 16037 17017 16071 17051
rect 18521 17017 18555 17051
rect 10241 16949 10275 16983
rect 11897 16949 11931 16983
rect 12265 16949 12299 16983
rect 13645 16949 13679 16983
rect 14105 16949 14139 16983
rect 15669 16949 15703 16983
rect 16635 16949 16669 16983
rect 20361 16949 20395 16983
rect 24731 16949 24765 16983
rect 1547 16745 1581 16779
rect 3433 16745 3467 16779
rect 6469 16745 6503 16779
rect 6929 16745 6963 16779
rect 7481 16745 7515 16779
rect 11069 16745 11103 16779
rect 12817 16745 12851 16779
rect 16773 16745 16807 16779
rect 18705 16745 18739 16779
rect 18981 16745 19015 16779
rect 24777 16745 24811 16779
rect 2329 16677 2363 16711
rect 2421 16677 2455 16711
rect 3801 16677 3835 16711
rect 4537 16677 4571 16711
rect 10511 16677 10545 16711
rect 12219 16677 12253 16711
rect 13093 16677 13127 16711
rect 14381 16677 14415 16711
rect 14749 16677 14783 16711
rect 15577 16677 15611 16711
rect 16129 16677 16163 16711
rect 18061 16677 18095 16711
rect 1476 16609 1510 16643
rect 2568 16609 2602 16643
rect 4629 16609 4663 16643
rect 5181 16609 5215 16643
rect 5457 16609 5491 16643
rect 6009 16609 6043 16643
rect 7941 16609 7975 16643
rect 13645 16609 13679 16643
rect 14197 16609 14231 16643
rect 17325 16609 17359 16643
rect 17877 16609 17911 16643
rect 18889 16609 18923 16643
rect 19441 16609 19475 16643
rect 20913 16609 20947 16643
rect 21960 16609 21994 16643
rect 24593 16609 24627 16643
rect 2789 16541 2823 16575
rect 6101 16541 6135 16575
rect 10149 16541 10183 16575
rect 11897 16541 11931 16575
rect 15485 16541 15519 16575
rect 16405 16541 16439 16575
rect 2697 16473 2731 16507
rect 1961 16405 1995 16439
rect 3065 16405 3099 16439
rect 8309 16405 8343 16439
rect 8861 16405 8895 16439
rect 11805 16405 11839 16439
rect 18337 16405 18371 16439
rect 21097 16405 21131 16439
rect 22063 16405 22097 16439
rect 3157 16201 3191 16235
rect 3525 16201 3559 16235
rect 3985 16201 4019 16235
rect 4353 16201 4387 16235
rect 7757 16201 7791 16235
rect 8401 16201 8435 16235
rect 10241 16201 10275 16235
rect 11897 16201 11931 16235
rect 14105 16201 14139 16235
rect 15853 16201 15887 16235
rect 17509 16201 17543 16235
rect 17877 16201 17911 16235
rect 19257 16201 19291 16235
rect 19717 16201 19751 16235
rect 22293 16201 22327 16235
rect 23811 16201 23845 16235
rect 24685 16201 24719 16235
rect 15485 16133 15519 16167
rect 21971 16133 22005 16167
rect 6837 16065 6871 16099
rect 11345 16065 11379 16099
rect 14749 16065 14783 16099
rect 20361 16065 20395 16099
rect 20637 16065 20671 16099
rect 1961 15997 1995 16031
rect 2329 15997 2363 16031
rect 2421 15997 2455 16031
rect 2881 15997 2915 16031
rect 4445 15997 4479 16031
rect 5181 15997 5215 16031
rect 5457 15997 5491 16031
rect 5825 15997 5859 16031
rect 8033 15997 8067 16031
rect 10701 15997 10735 16031
rect 10793 15997 10827 16031
rect 11253 15997 11287 16031
rect 12633 15997 12667 16031
rect 12909 15997 12943 16031
rect 16313 15997 16347 16031
rect 16405 15997 16439 16031
rect 16865 15997 16899 16031
rect 18061 15997 18095 16031
rect 21868 15997 21902 16031
rect 22661 15997 22695 16031
rect 23740 15997 23774 16031
rect 24133 15997 24167 16031
rect 5917 15929 5951 15963
rect 6653 15929 6687 15963
rect 7199 15929 7233 15963
rect 8677 15929 8711 15963
rect 8769 15929 8803 15963
rect 9321 15929 9355 15963
rect 13645 15929 13679 15963
rect 14933 15929 14967 15963
rect 15025 15929 15059 15963
rect 17141 15929 17175 15963
rect 18382 15929 18416 15963
rect 20085 15929 20119 15963
rect 20453 15929 20487 15963
rect 6193 15861 6227 15895
rect 9781 15861 9815 15895
rect 12541 15861 12575 15895
rect 18981 15861 19015 15895
rect 21281 15861 21315 15895
rect 3065 15657 3099 15691
rect 3341 15657 3375 15691
rect 3525 15657 3559 15691
rect 5457 15657 5491 15691
rect 7297 15657 7331 15691
rect 7941 15657 7975 15691
rect 9781 15657 9815 15691
rect 10793 15657 10827 15691
rect 11713 15657 11747 15691
rect 12265 15657 12299 15691
rect 13001 15657 13035 15691
rect 17417 15657 17451 15691
rect 18981 15657 19015 15691
rect 20361 15657 20395 15691
rect 21925 15657 21959 15691
rect 24777 15657 24811 15691
rect 1777 15589 1811 15623
rect 2053 15521 2087 15555
rect 2329 15521 2363 15555
rect 2789 15453 2823 15487
rect 5825 15589 5859 15623
rect 6463 15589 6497 15623
rect 8217 15589 8251 15623
rect 8769 15589 8803 15623
rect 13829 15589 13863 15623
rect 15485 15589 15519 15623
rect 18382 15589 18416 15623
rect 21097 15589 21131 15623
rect 22477 15589 22511 15623
rect 2145 15385 2179 15419
rect 3341 15385 3375 15419
rect 3709 15521 3743 15555
rect 4065 15521 4099 15555
rect 4353 15521 4387 15555
rect 9965 15521 9999 15555
rect 10241 15521 10275 15555
rect 16865 15521 16899 15555
rect 18061 15521 18095 15555
rect 19876 15521 19910 15555
rect 24593 15521 24627 15555
rect 4169 15453 4203 15487
rect 4813 15453 4847 15487
rect 6101 15453 6135 15487
rect 8125 15453 8159 15487
rect 11345 15453 11379 15487
rect 13737 15453 13771 15487
rect 15393 15453 15427 15487
rect 15669 15453 15703 15487
rect 21005 15453 21039 15487
rect 21649 15453 21683 15487
rect 14289 15385 14323 15419
rect 17049 15385 17083 15419
rect 19947 15385 19981 15419
rect 3709 15317 3743 15351
rect 3801 15317 3835 15351
rect 5089 15317 5123 15351
rect 7021 15317 7055 15351
rect 11161 15317 11195 15351
rect 12633 15317 12667 15351
rect 14841 15317 14875 15351
rect 16497 15317 16531 15351
rect 19349 15317 19383 15351
rect 2513 15113 2547 15147
rect 3341 15113 3375 15147
rect 4537 15113 4571 15147
rect 5227 15113 5261 15147
rect 5365 15113 5399 15147
rect 6469 15113 6503 15147
rect 8401 15113 8435 15147
rect 10057 15113 10091 15147
rect 10425 15113 10459 15147
rect 12173 15113 12207 15147
rect 14519 15113 14553 15147
rect 16773 15113 16807 15147
rect 17417 15113 17451 15147
rect 17785 15113 17819 15147
rect 18245 15113 18279 15147
rect 21097 15113 21131 15147
rect 21373 15113 21407 15147
rect 22661 15113 22695 15147
rect 24685 15113 24719 15147
rect 24961 15113 24995 15147
rect 3617 15045 3651 15079
rect 6193 15045 6227 15079
rect 14197 15045 14231 15079
rect 16037 15045 16071 15079
rect 20637 15045 20671 15079
rect 2881 14977 2915 15011
rect 5457 14977 5491 15011
rect 7481 14977 7515 15011
rect 8125 14977 8159 15011
rect 10885 14977 10919 15011
rect 12909 14977 12943 15011
rect 13185 14977 13219 15011
rect 15485 14977 15519 15011
rect 17095 14977 17129 15011
rect 18521 14977 18555 15011
rect 19901 14977 19935 15011
rect 20085 14977 20119 15011
rect 21649 14977 21683 15011
rect 22017 14977 22051 15011
rect 1501 14909 1535 14943
rect 3525 14909 3559 14943
rect 3801 14909 3835 14943
rect 4905 14909 4939 14943
rect 5089 14909 5123 14943
rect 8861 14909 8895 14943
rect 9045 14909 9079 14943
rect 14448 14909 14482 14943
rect 16992 14909 17026 14943
rect 24184 14909 24218 14943
rect 2145 14841 2179 14875
rect 5825 14841 5859 14875
rect 7573 14841 7607 14875
rect 8953 14841 8987 14875
rect 10977 14841 11011 14875
rect 11529 14841 11563 14875
rect 12725 14841 12759 14875
rect 13001 14841 13035 14875
rect 15586 14841 15620 14875
rect 16405 14841 16439 14875
rect 18613 14841 18647 14875
rect 19165 14841 19199 14875
rect 20177 14841 20211 14875
rect 21741 14841 21775 14875
rect 24271 14841 24305 14875
rect 3985 14773 4019 14807
rect 7297 14773 7331 14807
rect 11897 14773 11931 14807
rect 13921 14773 13955 14807
rect 14933 14773 14967 14807
rect 15301 14773 15335 14807
rect 19533 14773 19567 14807
rect 1593 14569 1627 14603
rect 3065 14569 3099 14603
rect 4353 14569 4387 14603
rect 5457 14569 5491 14603
rect 6653 14569 6687 14603
rect 7389 14569 7423 14603
rect 12081 14569 12115 14603
rect 12633 14569 12667 14603
rect 14749 14569 14783 14603
rect 18613 14569 18647 14603
rect 21051 14569 21085 14603
rect 24777 14569 24811 14603
rect 7941 14501 7975 14535
rect 12909 14501 12943 14535
rect 13645 14501 13679 14535
rect 15117 14501 15151 14535
rect 15669 14501 15703 14535
rect 17877 14501 17911 14535
rect 18797 14501 18831 14535
rect 18889 14501 18923 14535
rect 20085 14501 20119 14535
rect 23075 14501 23109 14535
rect 2053 14433 2087 14467
rect 2329 14433 2363 14467
rect 4261 14433 4295 14467
rect 5089 14433 5123 14467
rect 5733 14433 5767 14467
rect 10425 14433 10459 14467
rect 10701 14433 10735 14467
rect 17141 14433 17175 14467
rect 17693 14433 17727 14467
rect 20361 14433 20395 14467
rect 20980 14433 21014 14467
rect 21992 14433 22026 14467
rect 22937 14433 22971 14467
rect 24593 14433 24627 14467
rect 2513 14365 2547 14399
rect 5641 14365 5675 14399
rect 7113 14365 7147 14399
rect 7849 14365 7883 14399
rect 8125 14365 8159 14399
rect 8769 14365 8803 14399
rect 10885 14365 10919 14399
rect 11713 14365 11747 14399
rect 13553 14365 13587 14399
rect 15577 14365 15611 14399
rect 15853 14365 15887 14399
rect 19165 14365 19199 14399
rect 2145 14297 2179 14331
rect 14105 14297 14139 14331
rect 22063 14297 22097 14331
rect 3617 14229 3651 14263
rect 11253 14229 11287 14263
rect 18245 14229 18279 14263
rect 21465 14229 21499 14263
rect 21741 14229 21775 14263
rect 1593 14025 1627 14059
rect 2053 14025 2087 14059
rect 2421 14025 2455 14059
rect 5181 14025 5215 14059
rect 6193 14025 6227 14059
rect 8585 14025 8619 14059
rect 10149 14025 10183 14059
rect 11529 14025 11563 14059
rect 13461 14025 13495 14059
rect 13829 14025 13863 14059
rect 17141 14025 17175 14059
rect 17877 14025 17911 14059
rect 19073 14025 19107 14059
rect 21005 14025 21039 14059
rect 2697 13957 2731 13991
rect 5917 13957 5951 13991
rect 11897 13957 11931 13991
rect 14933 13957 14967 13991
rect 15761 13957 15795 13991
rect 3065 13889 3099 13923
rect 3893 13889 3927 13923
rect 4261 13889 4295 13923
rect 5549 13889 5583 13923
rect 6561 13889 6595 13923
rect 9781 13889 9815 13923
rect 10609 13889 10643 13923
rect 12541 13889 12575 13923
rect 13185 13889 13219 13923
rect 16681 13889 16715 13923
rect 22937 13889 22971 13923
rect 1409 13821 1443 13855
rect 2605 13821 2639 13855
rect 2881 13821 2915 13855
rect 4169 13821 4203 13855
rect 4445 13821 4479 13855
rect 5733 13821 5767 13855
rect 7757 13821 7791 13855
rect 7941 13821 7975 13855
rect 9045 13821 9079 13855
rect 9505 13821 9539 13855
rect 14013 13821 14047 13855
rect 14473 13821 14507 13855
rect 18061 13821 18095 13855
rect 18613 13821 18647 13855
rect 21373 13821 21407 13855
rect 21649 13821 21683 13855
rect 8217 13753 8251 13787
rect 10517 13753 10551 13787
rect 10971 13753 11005 13787
rect 12633 13753 12667 13787
rect 15209 13753 15243 13787
rect 15301 13753 15335 13787
rect 19717 13753 19751 13787
rect 19809 13753 19843 13787
rect 20361 13753 20395 13787
rect 3617 13685 3651 13719
rect 3893 13685 3927 13719
rect 3985 13685 4019 13719
rect 4629 13685 4663 13719
rect 7389 13685 7423 13719
rect 8953 13685 8987 13719
rect 12173 13685 12207 13719
rect 14197 13685 14231 13719
rect 16129 13685 16163 13719
rect 16497 13685 16531 13719
rect 18153 13685 18187 13719
rect 19441 13685 19475 13719
rect 21281 13685 21315 13719
rect 22201 13685 22235 13719
rect 24593 13685 24627 13719
rect 3801 13481 3835 13515
rect 10149 13481 10183 13515
rect 10793 13481 10827 13515
rect 11897 13481 11931 13515
rect 12265 13481 12299 13515
rect 12541 13481 12575 13515
rect 13645 13481 13679 13515
rect 17141 13481 17175 13515
rect 18337 13481 18371 13515
rect 19717 13481 19751 13515
rect 2421 13413 2455 13447
rect 3525 13413 3559 13447
rect 4077 13413 4111 13447
rect 5911 13413 5945 13447
rect 8211 13413 8245 13447
rect 11339 13413 11373 13447
rect 13087 13413 13121 13447
rect 15669 13413 15703 13447
rect 19118 13413 19152 13447
rect 21005 13413 21039 13447
rect 21097 13413 21131 13447
rect 2329 13345 2363 13379
rect 4261 13345 4295 13379
rect 4997 13345 5031 13379
rect 8769 13345 8803 13379
rect 9965 13345 9999 13379
rect 14657 13345 14691 13379
rect 17325 13345 17359 13379
rect 17509 13345 17543 13379
rect 18797 13345 18831 13379
rect 4813 13277 4847 13311
rect 5549 13277 5583 13311
rect 7849 13277 7883 13311
rect 9137 13277 9171 13311
rect 10977 13277 11011 13311
rect 12725 13277 12759 13311
rect 15117 13277 15151 13311
rect 15577 13277 15611 13311
rect 15853 13277 15887 13311
rect 21281 13277 21315 13311
rect 2697 13141 2731 13175
rect 3065 13141 3099 13175
rect 4353 13141 4387 13175
rect 4813 13141 4847 13175
rect 5273 13141 5307 13175
rect 6469 13141 6503 13175
rect 6837 13141 6871 13175
rect 7481 13141 7515 13175
rect 10425 13141 10459 13175
rect 13921 13141 13955 13175
rect 19993 13141 20027 13175
rect 1593 12937 1627 12971
rect 2053 12937 2087 12971
rect 2697 12937 2731 12971
rect 7849 12937 7883 12971
rect 8401 12937 8435 12971
rect 9505 12937 9539 12971
rect 13645 12937 13679 12971
rect 15301 12937 15335 12971
rect 17141 12937 17175 12971
rect 19257 12937 19291 12971
rect 21281 12937 21315 12971
rect 9781 12869 9815 12903
rect 11437 12869 11471 12903
rect 16129 12869 16163 12903
rect 22477 12869 22511 12903
rect 2421 12801 2455 12835
rect 2973 12801 3007 12835
rect 7205 12801 7239 12835
rect 8585 12801 8619 12835
rect 11069 12801 11103 12835
rect 11713 12801 11747 12835
rect 14197 12801 14231 12835
rect 15577 12801 15611 12835
rect 16589 12801 16623 12835
rect 24731 12801 24765 12835
rect 1409 12733 1443 12767
rect 2881 12733 2915 12767
rect 3157 12733 3191 12767
rect 5089 12733 5123 12767
rect 5549 12733 5583 12767
rect 10149 12733 10183 12767
rect 10333 12733 10367 12767
rect 10793 12733 10827 12767
rect 12449 12733 12483 12767
rect 13277 12733 13311 12767
rect 17877 12733 17911 12767
rect 18337 12733 18371 12767
rect 20085 12733 20119 12767
rect 21005 12733 21039 12767
rect 21649 12733 21683 12767
rect 24644 12733 24678 12767
rect 5825 12665 5859 12699
rect 6929 12665 6963 12699
rect 7021 12665 7055 12699
rect 8906 12665 8940 12699
rect 13921 12665 13955 12699
rect 14013 12665 14047 12699
rect 14933 12665 14967 12699
rect 15669 12665 15703 12699
rect 20406 12665 20440 12699
rect 21925 12665 21959 12699
rect 22017 12665 22051 12699
rect 3341 12597 3375 12631
rect 4077 12597 4111 12631
rect 4537 12597 4571 12631
rect 4997 12597 5031 12631
rect 6101 12597 6135 12631
rect 6653 12597 6687 12631
rect 12633 12597 12667 12631
rect 13001 12597 13035 12631
rect 17509 12597 17543 12631
rect 18705 12597 18739 12631
rect 19533 12597 19567 12631
rect 19901 12597 19935 12631
rect 25145 12597 25179 12631
rect 3801 12393 3835 12427
rect 4261 12393 4295 12427
rect 4721 12393 4755 12427
rect 5089 12393 5123 12427
rect 6193 12393 6227 12427
rect 7205 12393 7239 12427
rect 7849 12393 7883 12427
rect 9045 12393 9079 12427
rect 10793 12393 10827 12427
rect 11437 12393 11471 12427
rect 15485 12393 15519 12427
rect 19533 12393 19567 12427
rect 20637 12393 20671 12427
rect 10517 12325 10551 12359
rect 12725 12325 12759 12359
rect 13829 12325 13863 12359
rect 16497 12325 16531 12359
rect 18607 12325 18641 12359
rect 21097 12325 21131 12359
rect 21649 12325 21683 12359
rect 1501 12257 1535 12291
rect 2973 12257 3007 12291
rect 4077 12257 4111 12291
rect 5365 12257 5399 12291
rect 5641 12257 5675 12291
rect 7021 12257 7055 12291
rect 8033 12257 8067 12291
rect 8493 12257 8527 12291
rect 9781 12257 9815 12291
rect 10241 12257 10275 12291
rect 11345 12257 11379 12291
rect 11805 12257 11839 12291
rect 15301 12257 15335 12291
rect 18245 12257 18279 12291
rect 2145 12189 2179 12223
rect 5917 12189 5951 12223
rect 8769 12189 8803 12223
rect 13737 12189 13771 12223
rect 14105 12189 14139 12223
rect 16405 12189 16439 12223
rect 21005 12189 21039 12223
rect 3433 12121 3467 12155
rect 16957 12121 16991 12155
rect 2605 12053 2639 12087
rect 3157 12053 3191 12087
rect 6929 12053 6963 12087
rect 13093 12053 13127 12087
rect 15853 12053 15887 12087
rect 19165 12053 19199 12087
rect 20085 12053 20119 12087
rect 21925 12053 21959 12087
rect 3065 11849 3099 11883
rect 4629 11849 4663 11883
rect 6285 11849 6319 11883
rect 11805 11849 11839 11883
rect 13921 11849 13955 11883
rect 14657 11849 14691 11883
rect 16129 11849 16163 11883
rect 16497 11849 16531 11883
rect 16865 11849 16899 11883
rect 17877 11849 17911 11883
rect 18337 11849 18371 11883
rect 19901 11849 19935 11883
rect 21097 11849 21131 11883
rect 22017 11849 22051 11883
rect 5089 11781 5123 11815
rect 8585 11781 8619 11815
rect 14381 11781 14415 11815
rect 17233 11781 17267 11815
rect 2789 11713 2823 11747
rect 8769 11713 8803 11747
rect 11529 11713 11563 11747
rect 12725 11713 12759 11747
rect 17095 11713 17129 11747
rect 2053 11645 2087 11679
rect 2145 11645 2179 11679
rect 2329 11645 2363 11679
rect 3709 11645 3743 11679
rect 4077 11645 4111 11679
rect 5365 11645 5399 11679
rect 5733 11645 5767 11679
rect 6837 11645 6871 11679
rect 7297 11645 7331 11679
rect 10701 11645 10735 11679
rect 10793 11645 10827 11679
rect 11253 11645 11287 11679
rect 12173 11645 12207 11679
rect 15209 11645 15243 11679
rect 16992 11645 17026 11679
rect 19165 11713 19199 11747
rect 20729 11713 20763 11747
rect 17417 11645 17451 11679
rect 21624 11645 21658 11679
rect 3433 11577 3467 11611
rect 5917 11577 5951 11611
rect 6653 11577 6687 11611
rect 9090 11577 9124 11611
rect 9965 11577 9999 11611
rect 15117 11577 15151 11611
rect 15571 11577 15605 11611
rect 17233 11577 17267 11611
rect 18521 11577 18555 11611
rect 18613 11577 18647 11611
rect 19533 11577 19567 11611
rect 20085 11577 20119 11611
rect 20177 11577 20211 11611
rect 1593 11509 1627 11543
rect 3893 11509 3927 11543
rect 6929 11509 6963 11543
rect 8033 11509 8067 11543
rect 9689 11509 9723 11543
rect 13093 11509 13127 11543
rect 13645 11509 13679 11543
rect 21373 11509 21407 11543
rect 21695 11509 21729 11543
rect 1593 11305 1627 11339
rect 3893 11305 3927 11339
rect 5273 11305 5307 11339
rect 7389 11305 7423 11339
rect 7849 11305 7883 11339
rect 8953 11305 8987 11339
rect 12817 11305 12851 11339
rect 13461 11305 13495 11339
rect 14013 11305 14047 11339
rect 15485 11305 15519 11339
rect 17601 11305 17635 11339
rect 18889 11305 18923 11339
rect 21051 11305 21085 11339
rect 4261 11237 4295 11271
rect 6101 11237 6135 11271
rect 9413 11237 9447 11271
rect 9873 11237 9907 11271
rect 11707 11237 11741 11271
rect 16123 11237 16157 11271
rect 18613 11237 18647 11271
rect 19809 11237 19843 11271
rect 1409 11169 1443 11203
rect 2421 11169 2455 11203
rect 2881 11169 2915 11203
rect 5825 11169 5859 11203
rect 7849 11169 7883 11203
rect 8033 11169 8067 11203
rect 11345 11169 11379 11203
rect 15761 11169 15795 11203
rect 17509 11169 17543 11203
rect 17969 11169 18003 11203
rect 19073 11169 19107 11203
rect 19533 11169 19567 11203
rect 20821 11169 20855 11203
rect 24593 11169 24627 11203
rect 3157 11101 3191 11135
rect 4169 11101 4203 11135
rect 4813 11101 4847 11135
rect 5457 11101 5491 11135
rect 7021 11101 7055 11135
rect 9781 11101 9815 11135
rect 13093 11101 13127 11135
rect 6745 11033 6779 11067
rect 10333 11033 10367 11067
rect 2053 10965 2087 10999
rect 3433 10965 3467 10999
rect 5457 10965 5491 10999
rect 5549 10965 5583 10999
rect 8585 10965 8619 10999
rect 10793 10965 10827 10999
rect 12265 10965 12299 10999
rect 16681 10965 16715 10999
rect 24777 10965 24811 10999
rect 4261 10761 4295 10795
rect 4537 10761 4571 10795
rect 8401 10761 8435 10795
rect 9413 10761 9447 10795
rect 10057 10761 10091 10795
rect 12173 10761 12207 10795
rect 13369 10761 13403 10795
rect 17095 10761 17129 10795
rect 17785 10761 17819 10795
rect 19073 10761 19107 10795
rect 19441 10761 19475 10795
rect 19763 10761 19797 10795
rect 20177 10761 20211 10795
rect 24409 10761 24443 10795
rect 8999 10693 9033 10727
rect 11897 10693 11931 10727
rect 14105 10693 14139 10727
rect 16773 10693 16807 10727
rect 24777 10693 24811 10727
rect 2513 10625 2547 10659
rect 3341 10625 3375 10659
rect 5917 10625 5951 10659
rect 6837 10625 6871 10659
rect 13553 10625 13587 10659
rect 15761 10625 15795 10659
rect 16405 10625 16439 10659
rect 1685 10557 1719 10591
rect 2053 10557 2087 10591
rect 8928 10557 8962 10591
rect 10701 10557 10735 10591
rect 11069 10557 11103 10591
rect 11253 10557 11287 10591
rect 12516 10557 12550 10591
rect 17024 10557 17058 10591
rect 18061 10557 18095 10591
rect 18613 10557 18647 10591
rect 19692 10557 19726 10591
rect 24593 10557 24627 10591
rect 25145 10557 25179 10591
rect 3249 10489 3283 10523
rect 3662 10489 3696 10523
rect 5273 10489 5307 10523
rect 5365 10489 5399 10523
rect 7158 10489 7192 10523
rect 8033 10489 8067 10523
rect 11529 10489 11563 10523
rect 13645 10489 13679 10523
rect 14933 10489 14967 10523
rect 15485 10489 15519 10523
rect 15577 10489 15611 10523
rect 17509 10489 17543 10523
rect 2881 10421 2915 10455
rect 5089 10421 5123 10455
rect 6193 10421 6227 10455
rect 6561 10421 6595 10455
rect 7757 10421 7791 10455
rect 9689 10421 9723 10455
rect 12587 10421 12621 10455
rect 13001 10421 13035 10455
rect 14473 10421 14507 10455
rect 15301 10421 15335 10455
rect 18337 10421 18371 10455
rect 20913 10421 20947 10455
rect 2237 10217 2271 10251
rect 3801 10217 3835 10251
rect 4261 10217 4295 10251
rect 6101 10217 6135 10251
rect 8769 10217 8803 10251
rect 10517 10217 10551 10251
rect 14013 10217 14047 10251
rect 14335 10217 14369 10251
rect 15577 10217 15611 10251
rect 15761 10217 15795 10251
rect 17601 10217 17635 10251
rect 18153 10217 18187 10251
rect 1685 10149 1719 10183
rect 5267 10149 5301 10183
rect 6837 10149 6871 10183
rect 12817 10149 12851 10183
rect 13369 10149 13403 10183
rect 13645 10149 13679 10183
rect 16773 10149 16807 10183
rect 1476 10081 1510 10115
rect 1869 10081 1903 10115
rect 2421 10081 2455 10115
rect 2513 10081 2547 10115
rect 2697 10081 2731 10115
rect 3433 10081 3467 10115
rect 8585 10081 8619 10115
rect 10333 10081 10367 10115
rect 14197 10081 14231 10115
rect 15209 10081 15243 10115
rect 3157 10013 3191 10047
rect 4905 10013 4939 10047
rect 6745 10013 6779 10047
rect 12725 10013 12759 10047
rect 16681 10013 16715 10047
rect 16957 10013 16991 10047
rect 7297 9945 7331 9979
rect 10793 9945 10827 9979
rect 4813 9877 4847 9911
rect 5825 9877 5859 9911
rect 1593 9673 1627 9707
rect 2789 9673 2823 9707
rect 6285 9673 6319 9707
rect 6561 9673 6595 9707
rect 8861 9673 8895 9707
rect 10333 9673 10367 9707
rect 12725 9673 12759 9707
rect 13093 9673 13127 9707
rect 14289 9673 14323 9707
rect 16083 9673 16117 9707
rect 16773 9673 16807 9707
rect 5917 9605 5951 9639
rect 16497 9605 16531 9639
rect 2513 9537 2547 9571
rect 4261 9537 4295 9571
rect 6929 9537 6963 9571
rect 7205 9537 7239 9571
rect 8401 9537 8435 9571
rect 9413 9537 9447 9571
rect 13369 9537 13403 9571
rect 13829 9537 13863 9571
rect 1409 9469 1443 9503
rect 1869 9469 1903 9503
rect 3316 9469 3350 9503
rect 3709 9469 3743 9503
rect 16012 9469 16046 9503
rect 24660 9469 24694 9503
rect 4169 9401 4203 9435
rect 4582 9401 4616 9435
rect 5457 9401 5491 9435
rect 7021 9401 7055 9435
rect 13461 9401 13495 9435
rect 15393 9401 15427 9435
rect 3387 9333 3421 9367
rect 5181 9333 5215 9367
rect 7849 9333 7883 9367
rect 12173 9333 12207 9367
rect 17233 9333 17267 9367
rect 24731 9333 24765 9367
rect 25145 9333 25179 9367
rect 1593 9129 1627 9163
rect 2421 9129 2455 9163
rect 4261 9129 4295 9163
rect 6561 9129 6595 9163
rect 7757 9129 7791 9163
rect 13369 9129 13403 9163
rect 24777 9129 24811 9163
rect 5181 9061 5215 9095
rect 5733 9061 5767 9095
rect 1409 8993 1443 9027
rect 2973 8993 3007 9027
rect 7573 8993 7607 9027
rect 24593 8993 24627 9027
rect 5089 8925 5123 8959
rect 3157 8857 3191 8891
rect 7021 8789 7055 8823
rect 1547 8585 1581 8619
rect 3341 8585 3375 8619
rect 5089 8585 5123 8619
rect 5319 8585 5353 8619
rect 7573 8585 7607 8619
rect 24685 8585 24719 8619
rect 2973 8517 3007 8551
rect 4353 8517 4387 8551
rect 6009 8517 6043 8551
rect 2329 8449 2363 8483
rect 5733 8449 5767 8483
rect 1476 8381 1510 8415
rect 1869 8381 1903 8415
rect 3157 8381 3191 8415
rect 3617 8381 3651 8415
rect 4178 8381 4212 8415
rect 4629 8381 4663 8415
rect 5248 8381 5282 8415
rect 1593 8041 1627 8075
rect 4261 8041 4295 8075
rect 5273 8041 5307 8075
rect 1409 7905 1443 7939
rect 4077 7905 4111 7939
rect 5089 7905 5123 7939
rect 1593 7497 1627 7531
rect 4077 7497 4111 7531
rect 5089 7497 5123 7531
rect 24777 7429 24811 7463
rect 24593 7293 24627 7327
rect 25145 7293 25179 7327
rect 1593 6953 1627 6987
rect 1409 6817 1443 6851
rect 1593 6409 1627 6443
rect 24777 5865 24811 5899
rect 24593 5729 24627 5763
rect 24685 5321 24719 5355
rect 3928 2941 3962 2975
rect 4353 2941 4387 2975
rect 4031 2805 4065 2839
rect 7067 2601 7101 2635
rect 8217 2601 8251 2635
rect 11667 2601 11701 2635
rect 21465 2601 21499 2635
rect 24777 2601 24811 2635
rect 6996 2465 7030 2499
rect 8008 2465 8042 2499
rect 11596 2465 11630 2499
rect 11989 2465 12023 2499
rect 14105 2465 14139 2499
rect 14657 2465 14691 2499
rect 18337 2465 18371 2499
rect 21256 2465 21290 2499
rect 22820 2465 22854 2499
rect 23213 2465 23247 2499
rect 24593 2465 24627 2499
rect 25145 2465 25179 2499
rect 18889 2397 18923 2431
rect 14289 2329 14323 2363
rect 18521 2329 18555 2363
rect 7389 2261 7423 2295
rect 8493 2261 8527 2295
rect 21741 2261 21775 2295
rect 22891 2261 22925 2295
<< metal1 >>
rect 24946 27480 24952 27532
rect 25004 27520 25010 27532
rect 25958 27520 25964 27532
rect 25004 27492 25964 27520
rect 25004 27480 25010 27492
rect 25958 27480 25964 27492
rect 26016 27480 26022 27532
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 11584 25347 11642 25353
rect 11584 25313 11596 25347
rect 11630 25344 11642 25347
rect 12158 25344 12164 25356
rect 11630 25316 12164 25344
rect 11630 25313 11642 25316
rect 11584 25307 11642 25313
rect 12158 25304 12164 25316
rect 12216 25304 12222 25356
rect 12710 25353 12716 25356
rect 12688 25347 12716 25353
rect 12688 25344 12700 25347
rect 12623 25316 12700 25344
rect 12688 25313 12700 25316
rect 12768 25344 12774 25356
rect 27614 25344 27620 25356
rect 12768 25316 27620 25344
rect 12688 25307 12716 25313
rect 12710 25304 12716 25307
rect 12768 25304 12774 25316
rect 27614 25304 27620 25316
rect 27672 25304 27678 25356
rect 5626 25168 5632 25220
rect 5684 25208 5690 25220
rect 6546 25208 6552 25220
rect 5684 25180 6552 25208
rect 5684 25168 5690 25180
rect 6546 25168 6552 25180
rect 6604 25168 6610 25220
rect 9398 25168 9404 25220
rect 9456 25208 9462 25220
rect 13538 25208 13544 25220
rect 9456 25180 13544 25208
rect 9456 25168 9462 25180
rect 13538 25168 13544 25180
rect 13596 25168 13602 25220
rect 11655 25143 11713 25149
rect 11655 25109 11667 25143
rect 11701 25140 11713 25143
rect 12434 25140 12440 25152
rect 11701 25112 12440 25140
rect 11701 25109 11713 25112
rect 11655 25103 11713 25109
rect 12434 25100 12440 25112
rect 12492 25100 12498 25152
rect 12526 25100 12532 25152
rect 12584 25140 12590 25152
rect 12759 25143 12817 25149
rect 12759 25140 12771 25143
rect 12584 25112 12771 25140
rect 12584 25100 12590 25112
rect 12759 25109 12771 25112
rect 12805 25109 12817 25143
rect 12759 25103 12817 25109
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 12710 24936 12716 24948
rect 12671 24908 12716 24936
rect 12710 24896 12716 24908
rect 12768 24896 12774 24948
rect 13081 24939 13139 24945
rect 13081 24905 13093 24939
rect 13127 24936 13139 24939
rect 13262 24936 13268 24948
rect 13127 24908 13268 24936
rect 13127 24905 13139 24908
rect 13081 24899 13139 24905
rect 13262 24896 13268 24908
rect 13320 24896 13326 24948
rect 1448 24735 1506 24741
rect 1448 24701 1460 24735
rect 1494 24732 1506 24735
rect 1854 24732 1860 24744
rect 1494 24704 1860 24732
rect 1494 24701 1506 24704
rect 1448 24695 1506 24701
rect 1854 24692 1860 24704
rect 1912 24692 1918 24744
rect 11400 24735 11458 24741
rect 11400 24701 11412 24735
rect 11446 24732 11458 24735
rect 12897 24735 12955 24741
rect 11446 24704 11928 24732
rect 11446 24701 11458 24704
rect 11400 24695 11458 24701
rect 1535 24667 1593 24673
rect 1535 24633 1547 24667
rect 1581 24664 1593 24667
rect 8662 24664 8668 24676
rect 1581 24636 8668 24664
rect 1581 24633 1593 24636
rect 1535 24627 1593 24633
rect 8662 24624 8668 24636
rect 8720 24624 8726 24676
rect 11900 24673 11928 24704
rect 12897 24701 12909 24735
rect 12943 24732 12955 24735
rect 13449 24735 13507 24741
rect 13449 24732 13461 24735
rect 12943 24704 13461 24732
rect 12943 24701 12955 24704
rect 12897 24695 12955 24701
rect 13449 24701 13461 24704
rect 13495 24732 13507 24735
rect 14090 24732 14096 24744
rect 13495 24704 14096 24732
rect 13495 24701 13507 24704
rect 13449 24695 13507 24701
rect 14090 24692 14096 24704
rect 14148 24692 14154 24744
rect 14788 24735 14846 24741
rect 14788 24701 14800 24735
rect 14834 24732 14846 24735
rect 15194 24732 15200 24744
rect 14834 24704 15200 24732
rect 14834 24701 14846 24704
rect 14788 24695 14846 24701
rect 15194 24692 15200 24704
rect 15252 24692 15258 24744
rect 11885 24667 11943 24673
rect 11885 24633 11897 24667
rect 11931 24664 11943 24667
rect 12250 24664 12256 24676
rect 11931 24636 12256 24664
rect 11931 24633 11943 24636
rect 11885 24627 11943 24633
rect 12250 24624 12256 24636
rect 12308 24624 12314 24676
rect 14875 24667 14933 24673
rect 14875 24633 14887 24667
rect 14921 24664 14933 24667
rect 15378 24664 15384 24676
rect 14921 24636 15384 24664
rect 14921 24633 14933 24636
rect 14875 24627 14933 24633
rect 15378 24624 15384 24636
rect 15436 24624 15442 24676
rect 11330 24556 11336 24608
rect 11388 24596 11394 24608
rect 11471 24599 11529 24605
rect 11471 24596 11483 24599
rect 11388 24568 11483 24596
rect 11388 24556 11394 24568
rect 11471 24565 11483 24568
rect 11517 24565 11529 24599
rect 12158 24596 12164 24608
rect 12119 24568 12164 24596
rect 11471 24559 11529 24565
rect 12158 24556 12164 24568
rect 12216 24556 12222 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 11606 24392 11612 24404
rect 11567 24364 11612 24392
rect 11606 24352 11612 24364
rect 11664 24352 11670 24404
rect 13449 24395 13507 24401
rect 13449 24361 13461 24395
rect 13495 24392 13507 24395
rect 14550 24392 14556 24404
rect 13495 24364 14556 24392
rect 13495 24361 13507 24364
rect 13449 24355 13507 24361
rect 14550 24352 14556 24364
rect 14608 24352 14614 24404
rect 1464 24259 1522 24265
rect 1464 24225 1476 24259
rect 1510 24225 1522 24259
rect 1464 24219 1522 24225
rect 5905 24259 5963 24265
rect 5905 24225 5917 24259
rect 5951 24256 5963 24259
rect 6086 24256 6092 24268
rect 5951 24228 6092 24256
rect 5951 24225 5963 24228
rect 5905 24219 5963 24225
rect 106 24148 112 24200
rect 164 24188 170 24200
rect 1479 24188 1507 24219
rect 6086 24216 6092 24228
rect 6144 24216 6150 24268
rect 6914 24256 6920 24268
rect 6875 24228 6920 24256
rect 6914 24216 6920 24228
rect 6972 24216 6978 24268
rect 11330 24216 11336 24268
rect 11388 24256 11394 24268
rect 11425 24259 11483 24265
rect 11425 24256 11437 24259
rect 11388 24228 11437 24256
rect 11388 24216 11394 24228
rect 11425 24225 11437 24228
rect 11471 24225 11483 24259
rect 11425 24219 11483 24225
rect 12434 24216 12440 24268
rect 12492 24256 12498 24268
rect 13265 24259 13323 24265
rect 13265 24256 13277 24259
rect 12492 24228 13277 24256
rect 12492 24216 12498 24228
rect 13265 24225 13277 24228
rect 13311 24256 13323 24259
rect 13446 24256 13452 24268
rect 13311 24228 13452 24256
rect 13311 24225 13323 24228
rect 13265 24219 13323 24225
rect 13446 24216 13452 24228
rect 13504 24216 13510 24268
rect 15356 24259 15414 24265
rect 15356 24225 15368 24259
rect 15402 24256 15414 24259
rect 15746 24256 15752 24268
rect 15402 24228 15752 24256
rect 15402 24225 15414 24228
rect 15356 24219 15414 24225
rect 15746 24216 15752 24228
rect 15804 24216 15810 24268
rect 16368 24259 16426 24265
rect 16368 24225 16380 24259
rect 16414 24256 16426 24259
rect 16942 24256 16948 24268
rect 16414 24228 16948 24256
rect 16414 24225 16426 24228
rect 16368 24219 16426 24225
rect 16942 24216 16948 24228
rect 17000 24216 17006 24268
rect 17380 24259 17438 24265
rect 17380 24225 17392 24259
rect 17426 24256 17438 24259
rect 18392 24259 18450 24265
rect 18392 24256 18404 24259
rect 17426 24228 18404 24256
rect 17426 24225 17438 24228
rect 17380 24219 17438 24225
rect 18392 24225 18404 24228
rect 18438 24256 18450 24259
rect 18598 24256 18604 24268
rect 18438 24228 18604 24256
rect 18438 24225 18450 24228
rect 18392 24219 18450 24225
rect 18598 24216 18604 24228
rect 18656 24216 18662 24268
rect 20968 24259 21026 24265
rect 20968 24225 20980 24259
rect 21014 24256 21026 24259
rect 21450 24256 21456 24268
rect 21014 24228 21456 24256
rect 21014 24225 21026 24228
rect 20968 24219 21026 24225
rect 21450 24216 21456 24228
rect 21508 24216 21514 24268
rect 1946 24188 1952 24200
rect 164 24160 1952 24188
rect 164 24148 170 24160
rect 1946 24148 1952 24160
rect 2004 24148 2010 24200
rect 2038 24148 2044 24200
rect 2096 24188 2102 24200
rect 2409 24191 2467 24197
rect 2409 24188 2421 24191
rect 2096 24160 2421 24188
rect 2096 24148 2102 24160
rect 2409 24157 2421 24160
rect 2455 24157 2467 24191
rect 2409 24151 2467 24157
rect 6089 24123 6147 24129
rect 6089 24089 6101 24123
rect 6135 24120 6147 24123
rect 6822 24120 6828 24132
rect 6135 24092 6828 24120
rect 6135 24089 6147 24092
rect 6089 24083 6147 24089
rect 6822 24080 6828 24092
rect 6880 24080 6886 24132
rect 15930 24120 15936 24132
rect 15843 24092 15936 24120
rect 15930 24080 15936 24092
rect 15988 24120 15994 24132
rect 17451 24123 17509 24129
rect 17451 24120 17463 24123
rect 15988 24092 17463 24120
rect 15988 24080 15994 24092
rect 17451 24089 17463 24092
rect 17497 24089 17509 24123
rect 17451 24083 17509 24089
rect 1535 24055 1593 24061
rect 1535 24021 1547 24055
rect 1581 24052 1593 24055
rect 5994 24052 6000 24064
rect 1581 24024 6000 24052
rect 1581 24021 1593 24024
rect 1535 24015 1593 24021
rect 5994 24012 6000 24024
rect 6052 24012 6058 24064
rect 6454 24012 6460 24064
rect 6512 24052 6518 24064
rect 7101 24055 7159 24061
rect 7101 24052 7113 24055
rect 6512 24024 7113 24052
rect 6512 24012 6518 24024
rect 7101 24021 7113 24024
rect 7147 24021 7159 24055
rect 10594 24052 10600 24064
rect 10555 24024 10600 24052
rect 7101 24015 7159 24021
rect 10594 24012 10600 24024
rect 10652 24012 10658 24064
rect 14182 24052 14188 24064
rect 14143 24024 14188 24052
rect 14182 24012 14188 24024
rect 14240 24012 14246 24064
rect 15427 24055 15485 24061
rect 15427 24021 15439 24055
rect 15473 24052 15485 24055
rect 16206 24052 16212 24064
rect 15473 24024 16212 24052
rect 15473 24021 15485 24024
rect 15427 24015 15485 24021
rect 16206 24012 16212 24024
rect 16264 24012 16270 24064
rect 16298 24012 16304 24064
rect 16356 24052 16362 24064
rect 16439 24055 16497 24061
rect 16439 24052 16451 24055
rect 16356 24024 16451 24052
rect 16356 24012 16362 24024
rect 16439 24021 16451 24024
rect 16485 24021 16497 24055
rect 16439 24015 16497 24021
rect 18463 24055 18521 24061
rect 18463 24021 18475 24055
rect 18509 24052 18521 24055
rect 18874 24052 18880 24064
rect 18509 24024 18880 24052
rect 18509 24021 18521 24024
rect 18463 24015 18521 24021
rect 18874 24012 18880 24024
rect 18932 24012 18938 24064
rect 20346 24012 20352 24064
rect 20404 24052 20410 24064
rect 21039 24055 21097 24061
rect 21039 24052 21051 24055
rect 20404 24024 21051 24052
rect 20404 24012 20410 24024
rect 21039 24021 21051 24024
rect 21085 24021 21097 24055
rect 21039 24015 21097 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1946 23808 1952 23860
rect 2004 23848 2010 23860
rect 2317 23851 2375 23857
rect 2317 23848 2329 23851
rect 2004 23820 2329 23848
rect 2004 23808 2010 23820
rect 2317 23817 2329 23820
rect 2363 23817 2375 23851
rect 2317 23811 2375 23817
rect 5813 23851 5871 23857
rect 5813 23817 5825 23851
rect 5859 23848 5871 23851
rect 6638 23848 6644 23860
rect 5859 23820 6644 23848
rect 5859 23817 5871 23820
rect 5813 23811 5871 23817
rect 6638 23808 6644 23820
rect 6696 23808 6702 23860
rect 11330 23808 11336 23860
rect 11388 23848 11394 23860
rect 11517 23851 11575 23857
rect 11517 23848 11529 23851
rect 11388 23820 11529 23848
rect 11388 23808 11394 23820
rect 11517 23817 11529 23820
rect 11563 23817 11575 23851
rect 13446 23848 13452 23860
rect 13407 23820 13452 23848
rect 11517 23811 11575 23817
rect 13446 23808 13452 23820
rect 13504 23808 13510 23860
rect 15381 23851 15439 23857
rect 15381 23817 15393 23851
rect 15427 23848 15439 23851
rect 15746 23848 15752 23860
rect 15427 23820 15752 23848
rect 15427 23817 15439 23820
rect 15381 23811 15439 23817
rect 15746 23808 15752 23820
rect 15804 23848 15810 23860
rect 17310 23848 17316 23860
rect 15804 23820 17316 23848
rect 15804 23808 15810 23820
rect 17310 23808 17316 23820
rect 17368 23808 17374 23860
rect 18233 23851 18291 23857
rect 18233 23817 18245 23851
rect 18279 23848 18291 23851
rect 19334 23848 19340 23860
rect 18279 23820 19340 23848
rect 18279 23817 18291 23820
rect 18233 23811 18291 23817
rect 19334 23808 19340 23820
rect 19392 23808 19398 23860
rect 19889 23851 19947 23857
rect 19889 23817 19901 23851
rect 19935 23848 19947 23851
rect 20898 23848 20904 23860
rect 19935 23820 20904 23848
rect 19935 23817 19947 23820
rect 19889 23811 19947 23817
rect 20898 23808 20904 23820
rect 20956 23808 20962 23860
rect 21450 23848 21456 23860
rect 21411 23820 21456 23848
rect 21450 23808 21456 23820
rect 21508 23808 21514 23860
rect 21821 23851 21879 23857
rect 21821 23817 21833 23851
rect 21867 23848 21879 23851
rect 24670 23848 24676 23860
rect 21867 23820 24676 23848
rect 21867 23817 21879 23820
rect 21821 23811 21879 23817
rect 5997 23783 6055 23789
rect 5997 23749 6009 23783
rect 6043 23780 6055 23783
rect 6273 23783 6331 23789
rect 6273 23780 6285 23783
rect 6043 23752 6285 23780
rect 6043 23749 6055 23752
rect 5997 23743 6055 23749
rect 6273 23749 6285 23752
rect 6319 23780 6331 23783
rect 8202 23780 8208 23792
rect 6319 23752 8208 23780
rect 6319 23749 6331 23752
rect 6273 23743 6331 23749
rect 8202 23740 8208 23752
rect 8260 23740 8266 23792
rect 17405 23783 17463 23789
rect 17405 23749 17417 23783
rect 17451 23780 17463 23783
rect 18598 23780 18604 23792
rect 17451 23752 18604 23780
rect 17451 23749 17463 23752
rect 17405 23743 17463 23749
rect 18598 23740 18604 23752
rect 18656 23740 18662 23792
rect 4798 23672 4804 23724
rect 4856 23712 4862 23724
rect 6086 23712 6092 23724
rect 4856 23684 6092 23712
rect 4856 23672 4862 23684
rect 6086 23672 6092 23684
rect 6144 23712 6150 23724
rect 6549 23715 6607 23721
rect 6549 23712 6561 23715
rect 6144 23684 6561 23712
rect 6144 23672 6150 23684
rect 6549 23681 6561 23684
rect 6595 23681 6607 23715
rect 12526 23712 12532 23724
rect 12487 23684 12532 23712
rect 6549 23675 6607 23681
rect 12526 23672 12532 23684
rect 12584 23672 12590 23724
rect 12802 23712 12808 23724
rect 12763 23684 12808 23712
rect 12802 23672 12808 23684
rect 12860 23672 12866 23724
rect 14642 23712 14648 23724
rect 14603 23684 14648 23712
rect 14642 23672 14648 23684
rect 14700 23672 14706 23724
rect 15930 23712 15936 23724
rect 15891 23684 15936 23712
rect 15930 23672 15936 23684
rect 15988 23672 15994 23724
rect 16114 23672 16120 23724
rect 16172 23712 16178 23724
rect 16209 23715 16267 23721
rect 16209 23712 16221 23715
rect 16172 23684 16221 23712
rect 16172 23672 16178 23684
rect 16209 23681 16221 23684
rect 16255 23681 16267 23715
rect 16209 23675 16267 23681
rect 1397 23647 1455 23653
rect 1397 23613 1409 23647
rect 1443 23644 1455 23647
rect 1486 23644 1492 23656
rect 1443 23616 1492 23644
rect 1443 23613 1455 23616
rect 1397 23607 1455 23613
rect 1486 23604 1492 23616
rect 1544 23644 1550 23656
rect 1949 23647 2007 23653
rect 1949 23644 1961 23647
rect 1544 23616 1961 23644
rect 1544 23604 1550 23616
rect 1949 23613 1961 23616
rect 1995 23613 2007 23647
rect 1949 23607 2007 23613
rect 2222 23604 2228 23656
rect 2280 23644 2286 23656
rect 2536 23647 2594 23653
rect 2536 23644 2548 23647
rect 2280 23616 2548 23644
rect 2280 23604 2286 23616
rect 2536 23613 2548 23616
rect 2582 23644 2594 23647
rect 2961 23647 3019 23653
rect 2961 23644 2973 23647
rect 2582 23616 2973 23644
rect 2582 23613 2594 23616
rect 2536 23607 2594 23613
rect 2961 23613 2973 23616
rect 3007 23613 3019 23647
rect 2961 23607 3019 23613
rect 3142 23604 3148 23656
rect 3200 23644 3206 23656
rect 3548 23647 3606 23653
rect 3548 23644 3560 23647
rect 3200 23616 3560 23644
rect 3200 23604 3206 23616
rect 3548 23613 3560 23616
rect 3594 23644 3606 23647
rect 3973 23647 4031 23653
rect 3973 23644 3985 23647
rect 3594 23616 3985 23644
rect 3594 23613 3606 23616
rect 3548 23607 3606 23613
rect 3973 23613 3985 23616
rect 4019 23613 4031 23647
rect 3973 23607 4031 23613
rect 5629 23647 5687 23653
rect 5629 23613 5641 23647
rect 5675 23644 5687 23647
rect 5997 23647 6055 23653
rect 5997 23644 6009 23647
rect 5675 23616 6009 23644
rect 5675 23613 5687 23616
rect 5629 23607 5687 23613
rect 5997 23613 6009 23616
rect 6043 23613 6055 23647
rect 5997 23607 6055 23613
rect 6638 23604 6644 23656
rect 6696 23644 6702 23656
rect 8478 23653 8484 23656
rect 7412 23647 7470 23653
rect 7412 23644 7424 23647
rect 6696 23616 7424 23644
rect 6696 23604 6702 23616
rect 7412 23613 7424 23616
rect 7458 23644 7470 23647
rect 7837 23647 7895 23653
rect 7837 23644 7849 23647
rect 7458 23616 7849 23644
rect 7458 23613 7470 23616
rect 7412 23607 7470 23613
rect 7837 23613 7849 23616
rect 7883 23613 7895 23647
rect 8456 23647 8484 23653
rect 8456 23644 8468 23647
rect 8391 23616 8468 23644
rect 7837 23607 7895 23613
rect 8456 23613 8468 23616
rect 8536 23644 8542 23656
rect 8849 23647 8907 23653
rect 8849 23644 8861 23647
rect 8536 23616 8861 23644
rect 8456 23607 8484 23613
rect 8478 23604 8484 23607
rect 8536 23604 8542 23616
rect 8849 23613 8861 23616
rect 8895 23613 8907 23647
rect 10594 23644 10600 23656
rect 10555 23616 10600 23644
rect 8849 23607 8907 23613
rect 10594 23604 10600 23616
rect 10652 23604 10658 23656
rect 10962 23644 10968 23656
rect 10923 23616 10968 23644
rect 10962 23604 10968 23616
rect 11020 23604 11026 23656
rect 13814 23604 13820 23656
rect 13872 23644 13878 23656
rect 14001 23647 14059 23653
rect 14001 23644 14013 23647
rect 13872 23616 14013 23644
rect 13872 23604 13878 23616
rect 14001 23613 14013 23616
rect 14047 23644 14059 23647
rect 14093 23647 14151 23653
rect 14093 23644 14105 23647
rect 14047 23616 14105 23644
rect 14047 23613 14059 23616
rect 14001 23607 14059 23613
rect 14093 23613 14105 23616
rect 14139 23613 14151 23647
rect 14093 23607 14151 23613
rect 14182 23604 14188 23656
rect 14240 23644 14246 23656
rect 14553 23647 14611 23653
rect 14553 23644 14565 23647
rect 14240 23616 14565 23644
rect 14240 23604 14246 23616
rect 14553 23613 14565 23616
rect 14599 23613 14611 23647
rect 14553 23607 14611 23613
rect 17770 23604 17776 23656
rect 17828 23644 17834 23656
rect 17865 23647 17923 23653
rect 17865 23644 17877 23647
rect 17828 23616 17877 23644
rect 17828 23604 17834 23616
rect 17865 23613 17877 23616
rect 17911 23644 17923 23647
rect 18049 23647 18107 23653
rect 18049 23644 18061 23647
rect 17911 23616 18061 23644
rect 17911 23613 17923 23616
rect 17865 23607 17923 23613
rect 18049 23613 18061 23616
rect 18095 23613 18107 23647
rect 18049 23607 18107 23613
rect 19334 23604 19340 23656
rect 19392 23644 19398 23656
rect 19705 23647 19763 23653
rect 19705 23644 19717 23647
rect 19392 23616 19717 23644
rect 19392 23604 19398 23616
rect 19705 23613 19717 23616
rect 19751 23644 19763 23647
rect 20257 23647 20315 23653
rect 20257 23644 20269 23647
rect 19751 23616 20269 23644
rect 19751 23613 19763 23616
rect 19705 23607 19763 23613
rect 20257 23613 20269 23616
rect 20303 23613 20315 23647
rect 20257 23607 20315 23613
rect 20968 23647 21026 23653
rect 20968 23613 20980 23647
rect 21014 23644 21026 23647
rect 21836 23644 21864 23811
rect 24670 23808 24676 23820
rect 24728 23808 24734 23860
rect 25133 23851 25191 23857
rect 25133 23817 25145 23851
rect 25179 23848 25191 23851
rect 27246 23848 27252 23860
rect 25179 23820 27252 23848
rect 25179 23817 25191 23820
rect 25133 23811 25191 23817
rect 21014 23616 21864 23644
rect 24648 23647 24706 23653
rect 21014 23613 21026 23616
rect 20968 23607 21026 23613
rect 24648 23613 24660 23647
rect 24694 23644 24706 23647
rect 25148 23644 25176 23811
rect 27246 23808 27252 23820
rect 27304 23808 27310 23860
rect 24694 23616 25176 23644
rect 24694 23613 24706 23616
rect 24648 23607 24706 23613
rect 2639 23579 2697 23585
rect 2639 23545 2651 23579
rect 2685 23576 2697 23579
rect 2685 23548 3556 23576
rect 2685 23545 2697 23548
rect 2639 23539 2697 23545
rect 3528 23520 3556 23548
rect 6270 23536 6276 23588
rect 6328 23576 6334 23588
rect 6914 23576 6920 23588
rect 6328 23548 6920 23576
rect 6328 23536 6334 23548
rect 6914 23536 6920 23548
rect 6972 23576 6978 23588
rect 7009 23579 7067 23585
rect 7009 23576 7021 23579
rect 6972 23548 7021 23576
rect 6972 23536 6978 23548
rect 7009 23545 7021 23548
rect 7055 23545 7067 23579
rect 7009 23539 7067 23545
rect 11054 23536 11060 23588
rect 11112 23576 11118 23588
rect 11241 23579 11299 23585
rect 11241 23576 11253 23579
rect 11112 23548 11253 23576
rect 11112 23536 11118 23548
rect 11241 23545 11253 23548
rect 11287 23545 11299 23579
rect 11241 23539 11299 23545
rect 12621 23579 12679 23585
rect 12621 23545 12633 23579
rect 12667 23545 12679 23579
rect 12621 23539 12679 23545
rect 16025 23579 16083 23585
rect 16025 23545 16037 23579
rect 16071 23545 16083 23579
rect 16942 23576 16948 23588
rect 16855 23548 16948 23576
rect 16025 23539 16083 23545
rect 106 23468 112 23520
rect 164 23508 170 23520
rect 1581 23511 1639 23517
rect 1581 23508 1593 23511
rect 164 23480 1593 23508
rect 164 23468 170 23480
rect 1581 23477 1593 23480
rect 1627 23477 1639 23511
rect 1581 23471 1639 23477
rect 3510 23468 3516 23520
rect 3568 23468 3574 23520
rect 3651 23511 3709 23517
rect 3651 23477 3663 23511
rect 3697 23508 3709 23511
rect 3786 23508 3792 23520
rect 3697 23480 3792 23508
rect 3697 23477 3709 23480
rect 3651 23471 3709 23477
rect 3786 23468 3792 23480
rect 3844 23468 3850 23520
rect 7515 23511 7573 23517
rect 7515 23477 7527 23511
rect 7561 23508 7573 23511
rect 7742 23508 7748 23520
rect 7561 23480 7748 23508
rect 7561 23477 7573 23480
rect 7515 23471 7573 23477
rect 7742 23468 7748 23480
rect 7800 23468 7806 23520
rect 8386 23468 8392 23520
rect 8444 23508 8450 23520
rect 8527 23511 8585 23517
rect 8527 23508 8539 23511
rect 8444 23480 8539 23508
rect 8444 23468 8450 23480
rect 8527 23477 8539 23480
rect 8573 23477 8585 23511
rect 8527 23471 8585 23477
rect 10413 23511 10471 23517
rect 10413 23477 10425 23511
rect 10459 23508 10471 23511
rect 10962 23508 10968 23520
rect 10459 23480 10968 23508
rect 10459 23477 10471 23480
rect 10413 23471 10471 23477
rect 10962 23468 10968 23480
rect 11020 23508 11026 23520
rect 11330 23508 11336 23520
rect 11020 23480 11336 23508
rect 11020 23468 11026 23480
rect 11330 23468 11336 23480
rect 11388 23468 11394 23520
rect 12253 23511 12311 23517
rect 12253 23477 12265 23511
rect 12299 23508 12311 23511
rect 12636 23508 12664 23539
rect 12710 23508 12716 23520
rect 12299 23480 12716 23508
rect 12299 23477 12311 23480
rect 12253 23471 12311 23477
rect 12710 23468 12716 23480
rect 12768 23468 12774 23520
rect 15746 23508 15752 23520
rect 15659 23480 15752 23508
rect 15746 23468 15752 23480
rect 15804 23508 15810 23520
rect 16040 23508 16068 23539
rect 16942 23536 16948 23548
rect 17000 23576 17006 23588
rect 23382 23576 23388 23588
rect 17000 23548 23388 23576
rect 17000 23536 17006 23548
rect 23382 23536 23388 23548
rect 23440 23536 23446 23588
rect 15804 23480 16068 23508
rect 15804 23468 15810 23480
rect 20898 23468 20904 23520
rect 20956 23508 20962 23520
rect 21039 23511 21097 23517
rect 21039 23508 21051 23511
rect 20956 23480 21051 23508
rect 20956 23468 20962 23480
rect 21039 23477 21051 23480
rect 21085 23477 21097 23511
rect 21039 23471 21097 23477
rect 22738 23468 22744 23520
rect 22796 23508 22802 23520
rect 24719 23511 24777 23517
rect 24719 23508 24731 23511
rect 22796 23480 24731 23508
rect 22796 23468 22802 23480
rect 24719 23477 24731 23480
rect 24765 23477 24777 23511
rect 24719 23471 24777 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 8662 23304 8668 23316
rect 8623 23276 8668 23304
rect 8662 23264 8668 23276
rect 8720 23264 8726 23316
rect 12526 23304 12532 23316
rect 12487 23276 12532 23304
rect 12526 23264 12532 23276
rect 12584 23264 12590 23316
rect 16298 23304 16304 23316
rect 16259 23276 16304 23304
rect 16298 23264 16304 23276
rect 16356 23264 16362 23316
rect 18874 23304 18880 23316
rect 18835 23276 18880 23304
rect 18874 23264 18880 23276
rect 18932 23264 18938 23316
rect 6963 23239 7021 23245
rect 6963 23205 6975 23239
rect 7009 23236 7021 23239
rect 10410 23236 10416 23248
rect 7009 23208 10416 23236
rect 7009 23205 7021 23208
rect 6963 23199 7021 23205
rect 10410 23196 10416 23208
rect 10468 23196 10474 23248
rect 11609 23239 11667 23245
rect 11609 23205 11621 23239
rect 11655 23236 11667 23239
rect 12710 23236 12716 23248
rect 11655 23208 12716 23236
rect 11655 23205 11667 23208
rect 11609 23199 11667 23205
rect 12710 23196 12716 23208
rect 12768 23196 12774 23248
rect 15470 23236 15476 23248
rect 15431 23208 15476 23236
rect 15470 23196 15476 23208
rect 15528 23196 15534 23248
rect 16206 23196 16212 23248
rect 16264 23236 16270 23248
rect 16942 23236 16948 23248
rect 16264 23208 16948 23236
rect 16264 23196 16270 23208
rect 16942 23196 16948 23208
rect 17000 23196 17006 23248
rect 17034 23196 17040 23248
rect 17092 23236 17098 23248
rect 17092 23208 17137 23236
rect 17092 23196 17098 23208
rect 17310 23196 17316 23248
rect 17368 23236 17374 23248
rect 18230 23236 18236 23248
rect 17368 23208 18236 23236
rect 17368 23196 17374 23208
rect 18230 23196 18236 23208
rect 18288 23236 18294 23248
rect 21085 23239 21143 23245
rect 18288 23208 18495 23236
rect 18288 23196 18294 23208
rect 1397 23171 1455 23177
rect 1397 23137 1409 23171
rect 1443 23168 1455 23171
rect 1443 23140 2084 23168
rect 1443 23137 1455 23140
rect 1397 23131 1455 23137
rect 14 22924 20 22976
rect 72 22964 78 22976
rect 2056 22973 2084 23140
rect 2314 23128 2320 23180
rect 2372 23168 2378 23180
rect 2568 23171 2626 23177
rect 2568 23168 2580 23171
rect 2372 23140 2580 23168
rect 2372 23128 2378 23140
rect 2568 23137 2580 23140
rect 2614 23168 2626 23171
rect 2774 23168 2780 23180
rect 2614 23140 2780 23168
rect 2614 23137 2626 23140
rect 2568 23131 2626 23137
rect 2774 23128 2780 23140
rect 2832 23128 2838 23180
rect 4776 23171 4834 23177
rect 4776 23137 4788 23171
rect 4822 23168 4834 23171
rect 4890 23168 4896 23180
rect 4822 23140 4896 23168
rect 4822 23137 4834 23140
rect 4776 23131 4834 23137
rect 4890 23128 4896 23140
rect 4948 23128 4954 23180
rect 7904 23171 7962 23177
rect 7904 23137 7916 23171
rect 7950 23168 7962 23171
rect 8018 23168 8024 23180
rect 7950 23140 8024 23168
rect 7950 23137 7962 23140
rect 7904 23131 7962 23137
rect 8018 23128 8024 23140
rect 8076 23128 8082 23180
rect 13722 23168 13728 23180
rect 13683 23140 13728 23168
rect 13722 23128 13728 23140
rect 13780 23128 13786 23180
rect 14182 23168 14188 23180
rect 14143 23140 14188 23168
rect 14182 23128 14188 23140
rect 14240 23128 14246 23180
rect 18467 23177 18495 23208
rect 21085 23205 21097 23239
rect 21131 23236 21143 23239
rect 21358 23236 21364 23248
rect 21131 23208 21364 23236
rect 21131 23205 21143 23208
rect 21085 23199 21143 23205
rect 21358 23196 21364 23208
rect 21416 23196 21422 23248
rect 18452 23171 18510 23177
rect 18452 23137 18464 23171
rect 18498 23137 18510 23171
rect 18452 23131 18510 23137
rect 22465 23171 22523 23177
rect 22465 23137 22477 23171
rect 22511 23168 22523 23171
rect 22554 23168 22560 23180
rect 22511 23140 22560 23168
rect 22511 23137 22523 23140
rect 22465 23131 22523 23137
rect 22554 23128 22560 23140
rect 22612 23128 22618 23180
rect 5721 23103 5779 23109
rect 5721 23069 5733 23103
rect 5767 23100 5779 23103
rect 6086 23100 6092 23112
rect 5767 23072 6092 23100
rect 5767 23069 5779 23072
rect 5721 23063 5779 23069
rect 6086 23060 6092 23072
rect 6144 23060 6150 23112
rect 10413 23103 10471 23109
rect 10413 23069 10425 23103
rect 10459 23100 10471 23103
rect 11517 23103 11575 23109
rect 11517 23100 11529 23103
rect 10459 23072 11529 23100
rect 10459 23069 10471 23072
rect 10413 23063 10471 23069
rect 11517 23069 11529 23072
rect 11563 23100 11575 23103
rect 11698 23100 11704 23112
rect 11563 23072 11704 23100
rect 11563 23069 11575 23072
rect 11517 23063 11575 23069
rect 11698 23060 11704 23072
rect 11756 23060 11762 23112
rect 14369 23103 14427 23109
rect 14369 23069 14381 23103
rect 14415 23100 14427 23103
rect 14826 23100 14832 23112
rect 14415 23072 14832 23100
rect 14415 23069 14427 23072
rect 14369 23063 14427 23069
rect 14826 23060 14832 23072
rect 14884 23060 14890 23112
rect 15378 23100 15384 23112
rect 15339 23072 15384 23100
rect 15378 23060 15384 23072
rect 15436 23060 15442 23112
rect 15654 23100 15660 23112
rect 15615 23072 15660 23100
rect 15654 23060 15660 23072
rect 15712 23060 15718 23112
rect 16114 23060 16120 23112
rect 16172 23100 16178 23112
rect 17221 23103 17279 23109
rect 17221 23100 17233 23103
rect 16172 23072 17233 23100
rect 16172 23060 16178 23072
rect 17221 23069 17233 23072
rect 17267 23069 17279 23103
rect 20990 23100 20996 23112
rect 20951 23072 20996 23100
rect 17221 23063 17279 23069
rect 20990 23060 20996 23072
rect 21048 23060 21054 23112
rect 21266 23100 21272 23112
rect 21227 23072 21272 23100
rect 21266 23060 21272 23072
rect 21324 23060 21330 23112
rect 7975 23035 8033 23041
rect 7975 23001 7987 23035
rect 8021 23032 8033 23035
rect 9490 23032 9496 23044
rect 8021 23004 9496 23032
rect 8021 23001 8033 23004
rect 7975 22995 8033 23001
rect 9490 22992 9496 23004
rect 9548 22992 9554 23044
rect 12066 23032 12072 23044
rect 12027 23004 12072 23032
rect 12066 22992 12072 23004
rect 12124 22992 12130 23044
rect 1581 22967 1639 22973
rect 1581 22964 1593 22967
rect 72 22936 1593 22964
rect 72 22924 78 22936
rect 1581 22933 1593 22936
rect 1627 22933 1639 22967
rect 1581 22927 1639 22933
rect 2041 22967 2099 22973
rect 2041 22933 2053 22967
rect 2087 22964 2099 22967
rect 2314 22964 2320 22976
rect 2087 22936 2320 22964
rect 2087 22933 2099 22936
rect 2041 22927 2099 22933
rect 2314 22924 2320 22936
rect 2372 22924 2378 22976
rect 2639 22967 2697 22973
rect 2639 22933 2651 22967
rect 2685 22964 2697 22967
rect 3234 22964 3240 22976
rect 2685 22936 3240 22964
rect 2685 22933 2697 22936
rect 2639 22927 2697 22933
rect 3234 22924 3240 22936
rect 3292 22924 3298 22976
rect 4847 22967 4905 22973
rect 4847 22933 4859 22967
rect 4893 22964 4905 22967
rect 4982 22964 4988 22976
rect 4893 22936 4988 22964
rect 4893 22933 4905 22936
rect 4847 22927 4905 22933
rect 4982 22924 4988 22936
rect 5040 22924 5046 22976
rect 5258 22964 5264 22976
rect 5219 22936 5264 22964
rect 5258 22924 5264 22936
rect 5316 22924 5322 22976
rect 6730 22964 6736 22976
rect 6691 22936 6736 22964
rect 6730 22924 6736 22936
rect 6788 22924 6794 22976
rect 8389 22967 8447 22973
rect 8389 22933 8401 22967
rect 8435 22964 8447 22967
rect 8570 22964 8576 22976
rect 8435 22936 8576 22964
rect 8435 22933 8447 22936
rect 8389 22927 8447 22933
rect 8570 22924 8576 22936
rect 8628 22924 8634 22976
rect 12526 22924 12532 22976
rect 12584 22964 12590 22976
rect 12802 22964 12808 22976
rect 12584 22936 12808 22964
rect 12584 22924 12590 22936
rect 12802 22924 12808 22936
rect 12860 22924 12866 22976
rect 18322 22924 18328 22976
rect 18380 22964 18386 22976
rect 18555 22967 18613 22973
rect 18555 22964 18567 22967
rect 18380 22936 18567 22964
rect 18380 22924 18386 22936
rect 18555 22933 18567 22936
rect 18601 22933 18613 22967
rect 18555 22927 18613 22933
rect 21082 22924 21088 22976
rect 21140 22964 21146 22976
rect 22603 22967 22661 22973
rect 22603 22964 22615 22967
rect 21140 22936 22615 22964
rect 21140 22924 21146 22936
rect 22603 22933 22615 22936
rect 22649 22933 22661 22967
rect 22603 22927 22661 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 2774 22760 2780 22772
rect 2735 22732 2780 22760
rect 2774 22720 2780 22732
rect 2832 22720 2838 22772
rect 11698 22760 11704 22772
rect 11659 22732 11704 22760
rect 11698 22720 11704 22732
rect 11756 22720 11762 22772
rect 13722 22760 13728 22772
rect 13683 22732 13728 22760
rect 13722 22720 13728 22732
rect 13780 22720 13786 22772
rect 16942 22720 16948 22772
rect 17000 22760 17006 22772
rect 17221 22763 17279 22769
rect 17221 22760 17233 22763
rect 17000 22732 17233 22760
rect 17000 22720 17006 22732
rect 17221 22729 17233 22732
rect 17267 22729 17279 22763
rect 18230 22760 18236 22772
rect 18191 22732 18236 22760
rect 17221 22723 17279 22729
rect 18230 22720 18236 22732
rect 18288 22720 18294 22772
rect 20990 22720 20996 22772
rect 21048 22760 21054 22772
rect 21637 22763 21695 22769
rect 21637 22760 21649 22763
rect 21048 22732 21649 22760
rect 21048 22720 21054 22732
rect 21637 22729 21649 22732
rect 21683 22729 21695 22763
rect 22554 22760 22560 22772
rect 22515 22732 22560 22760
rect 21637 22723 21695 22729
rect 22554 22720 22560 22732
rect 22612 22720 22618 22772
rect 4801 22695 4859 22701
rect 4801 22661 4813 22695
rect 4847 22692 4859 22695
rect 4890 22692 4896 22704
rect 4847 22664 4896 22692
rect 4847 22661 4859 22664
rect 4801 22655 4859 22661
rect 4890 22652 4896 22664
rect 4948 22692 4954 22704
rect 8478 22692 8484 22704
rect 4948 22664 8484 22692
rect 4948 22652 4954 22664
rect 8478 22652 8484 22664
rect 8536 22652 8542 22704
rect 12158 22652 12164 22704
rect 12216 22692 12222 22704
rect 13081 22695 13139 22701
rect 13081 22692 13093 22695
rect 12216 22664 13093 22692
rect 12216 22652 12222 22664
rect 13081 22661 13093 22664
rect 13127 22692 13139 22695
rect 13262 22692 13268 22704
rect 13127 22664 13268 22692
rect 13127 22661 13139 22664
rect 13081 22655 13139 22661
rect 13262 22652 13268 22664
rect 13320 22652 13326 22704
rect 16298 22692 16304 22704
rect 15948 22664 16304 22692
rect 8297 22627 8355 22633
rect 8297 22593 8309 22627
rect 8343 22624 8355 22627
rect 8662 22624 8668 22636
rect 8343 22596 8668 22624
rect 8343 22593 8355 22596
rect 8297 22587 8355 22593
rect 8662 22584 8668 22596
rect 8720 22584 8726 22636
rect 13906 22624 13912 22636
rect 10980 22596 13912 22624
rect 1949 22559 2007 22565
rect 1949 22525 1961 22559
rect 1995 22525 2007 22559
rect 1949 22519 2007 22525
rect 1762 22488 1768 22500
rect 1723 22460 1768 22488
rect 1762 22448 1768 22460
rect 1820 22448 1826 22500
rect 1964 22432 1992 22519
rect 3142 22516 3148 22568
rect 3200 22556 3206 22568
rect 3329 22559 3387 22565
rect 3329 22556 3341 22559
rect 3200 22528 3341 22556
rect 3200 22516 3206 22528
rect 3329 22525 3341 22528
rect 3375 22556 3387 22559
rect 3789 22559 3847 22565
rect 3789 22556 3801 22559
rect 3375 22528 3801 22556
rect 3375 22525 3387 22528
rect 3329 22519 3387 22525
rect 3789 22525 3801 22528
rect 3835 22525 3847 22559
rect 5258 22556 5264 22568
rect 5219 22528 5264 22556
rect 3789 22519 3847 22525
rect 5258 22516 5264 22528
rect 5316 22516 5322 22568
rect 10980 22565 11008 22596
rect 13906 22584 13912 22596
rect 13964 22584 13970 22636
rect 14366 22624 14372 22636
rect 14327 22596 14372 22624
rect 14366 22584 14372 22596
rect 14424 22584 14430 22636
rect 15013 22627 15071 22633
rect 15013 22593 15025 22627
rect 15059 22624 15071 22627
rect 15654 22624 15660 22636
rect 15059 22596 15660 22624
rect 15059 22593 15071 22596
rect 15013 22587 15071 22593
rect 15654 22584 15660 22596
rect 15712 22584 15718 22636
rect 15948 22633 15976 22664
rect 16298 22652 16304 22664
rect 16356 22652 16362 22704
rect 18874 22692 18880 22704
rect 18524 22664 18880 22692
rect 15933 22627 15991 22633
rect 15933 22593 15945 22627
rect 15979 22593 15991 22627
rect 16206 22624 16212 22636
rect 16167 22596 16212 22624
rect 15933 22587 15991 22593
rect 16206 22584 16212 22596
rect 16264 22584 16270 22636
rect 16945 22627 17003 22633
rect 16945 22593 16957 22627
rect 16991 22624 17003 22627
rect 17034 22624 17040 22636
rect 16991 22596 17040 22624
rect 16991 22593 17003 22596
rect 16945 22587 17003 22593
rect 7260 22559 7318 22565
rect 7260 22525 7272 22559
rect 7306 22556 7318 22559
rect 10597 22559 10655 22565
rect 7306 22528 7788 22556
rect 7306 22525 7318 22528
rect 7260 22519 7318 22525
rect 5905 22491 5963 22497
rect 5905 22457 5917 22491
rect 5951 22488 5963 22491
rect 6178 22488 6184 22500
rect 5951 22460 6184 22488
rect 5951 22457 5963 22460
rect 5905 22451 5963 22457
rect 6178 22448 6184 22460
rect 6236 22448 6242 22500
rect 1673 22423 1731 22429
rect 1673 22389 1685 22423
rect 1719 22420 1731 22423
rect 1946 22420 1952 22432
rect 1719 22392 1952 22420
rect 1719 22389 1731 22392
rect 1673 22383 1731 22389
rect 1946 22380 1952 22392
rect 2004 22380 2010 22432
rect 3050 22380 3056 22432
rect 3108 22420 3114 22432
rect 3513 22423 3571 22429
rect 3513 22420 3525 22423
rect 3108 22392 3525 22420
rect 3108 22380 3114 22392
rect 3513 22389 3525 22392
rect 3559 22389 3571 22423
rect 3513 22383 3571 22389
rect 6362 22380 6368 22432
rect 6420 22420 6426 22432
rect 6730 22420 6736 22432
rect 6420 22392 6736 22420
rect 6420 22380 6426 22392
rect 6730 22380 6736 22392
rect 6788 22420 6794 22432
rect 7009 22423 7067 22429
rect 7009 22420 7021 22423
rect 6788 22392 7021 22420
rect 6788 22380 6794 22392
rect 7009 22389 7021 22392
rect 7055 22389 7067 22423
rect 7009 22383 7067 22389
rect 7331 22423 7389 22429
rect 7331 22389 7343 22423
rect 7377 22420 7389 22423
rect 7558 22420 7564 22432
rect 7377 22392 7564 22420
rect 7377 22389 7389 22392
rect 7331 22383 7389 22389
rect 7558 22380 7564 22392
rect 7616 22380 7622 22432
rect 7760 22429 7788 22528
rect 10597 22525 10609 22559
rect 10643 22556 10655 22559
rect 10965 22559 11023 22565
rect 10965 22556 10977 22559
rect 10643 22528 10977 22556
rect 10643 22525 10655 22528
rect 10597 22519 10655 22525
rect 10965 22525 10977 22528
rect 11011 22525 11023 22559
rect 10965 22519 11023 22525
rect 11241 22559 11299 22565
rect 11241 22525 11253 22559
rect 11287 22556 11299 22559
rect 11330 22556 11336 22568
rect 11287 22528 11336 22556
rect 11287 22525 11299 22528
rect 11241 22519 11299 22525
rect 11330 22516 11336 22528
rect 11388 22516 11394 22568
rect 8389 22491 8447 22497
rect 8389 22457 8401 22491
rect 8435 22488 8447 22491
rect 8570 22488 8576 22500
rect 8435 22460 8576 22488
rect 8435 22457 8447 22460
rect 8389 22451 8447 22457
rect 8570 22448 8576 22460
rect 8628 22448 8634 22500
rect 8938 22488 8944 22500
rect 8899 22460 8944 22488
rect 8938 22448 8944 22460
rect 8996 22488 9002 22500
rect 12526 22488 12532 22500
rect 8996 22460 12532 22488
rect 8996 22448 9002 22460
rect 12526 22448 12532 22460
rect 12584 22448 12590 22500
rect 12618 22448 12624 22500
rect 12676 22488 12682 22500
rect 14458 22488 14464 22500
rect 12676 22460 12721 22488
rect 14419 22460 14464 22488
rect 12676 22448 12682 22460
rect 14458 22448 14464 22460
rect 14516 22448 14522 22500
rect 15381 22491 15439 22497
rect 15381 22457 15393 22491
rect 15427 22488 15439 22491
rect 15470 22488 15476 22500
rect 15427 22460 15476 22488
rect 15427 22457 15439 22460
rect 15381 22451 15439 22457
rect 15470 22448 15476 22460
rect 15528 22488 15534 22500
rect 15749 22491 15807 22497
rect 15749 22488 15761 22491
rect 15528 22460 15761 22488
rect 15528 22448 15534 22460
rect 15749 22457 15761 22460
rect 15795 22488 15807 22491
rect 16025 22491 16083 22497
rect 16025 22488 16037 22491
rect 15795 22460 16037 22488
rect 15795 22457 15807 22460
rect 15749 22451 15807 22457
rect 16025 22457 16037 22460
rect 16071 22457 16083 22491
rect 16025 22451 16083 22457
rect 7745 22423 7803 22429
rect 7745 22389 7757 22423
rect 7791 22420 7803 22423
rect 7834 22420 7840 22432
rect 7791 22392 7840 22420
rect 7791 22389 7803 22392
rect 7745 22383 7803 22389
rect 7834 22380 7840 22392
rect 7892 22380 7898 22432
rect 8018 22420 8024 22432
rect 7979 22392 8024 22420
rect 8018 22380 8024 22392
rect 8076 22380 8082 22432
rect 10965 22423 11023 22429
rect 10965 22389 10977 22423
rect 11011 22420 11023 22423
rect 11146 22420 11152 22432
rect 11011 22392 11152 22420
rect 11011 22389 11023 22392
rect 10965 22383 11023 22389
rect 11146 22380 11152 22392
rect 11204 22380 11210 22432
rect 12161 22423 12219 22429
rect 12161 22389 12173 22423
rect 12207 22420 12219 22423
rect 12710 22420 12716 22432
rect 12207 22392 12716 22420
rect 12207 22389 12219 22392
rect 12161 22383 12219 22389
rect 12710 22380 12716 22392
rect 12768 22380 12774 22432
rect 14093 22423 14151 22429
rect 14093 22389 14105 22423
rect 14139 22420 14151 22423
rect 14182 22420 14188 22432
rect 14139 22392 14188 22420
rect 14139 22389 14151 22392
rect 14093 22383 14151 22389
rect 14182 22380 14188 22392
rect 14240 22380 14246 22432
rect 16040 22420 16068 22451
rect 16960 22420 16988 22587
rect 17034 22584 17040 22596
rect 17092 22584 17098 22636
rect 18524 22633 18552 22664
rect 18874 22652 18880 22664
rect 18932 22652 18938 22704
rect 18966 22652 18972 22704
rect 19024 22692 19030 22704
rect 19061 22695 19119 22701
rect 19061 22692 19073 22695
rect 19024 22664 19073 22692
rect 19024 22652 19030 22664
rect 19061 22661 19073 22664
rect 19107 22661 19119 22695
rect 21358 22692 21364 22704
rect 21319 22664 21364 22692
rect 19061 22655 19119 22661
rect 21358 22652 21364 22664
rect 21416 22652 21422 22704
rect 18509 22627 18567 22633
rect 18509 22593 18521 22627
rect 18555 22593 18567 22627
rect 20346 22624 20352 22636
rect 20307 22596 20352 22624
rect 18509 22587 18567 22593
rect 20346 22584 20352 22596
rect 20404 22584 20410 22636
rect 20993 22627 21051 22633
rect 20993 22593 21005 22627
rect 21039 22624 21051 22627
rect 21266 22624 21272 22636
rect 21039 22596 21272 22624
rect 21039 22593 21051 22596
rect 20993 22587 21051 22593
rect 21266 22584 21272 22596
rect 21324 22584 21330 22636
rect 17865 22491 17923 22497
rect 17865 22457 17877 22491
rect 17911 22488 17923 22491
rect 18601 22491 18659 22497
rect 18601 22488 18613 22491
rect 17911 22460 18613 22488
rect 17911 22457 17923 22460
rect 17865 22451 17923 22457
rect 18601 22457 18613 22460
rect 18647 22488 18659 22491
rect 19978 22488 19984 22500
rect 18647 22460 19984 22488
rect 18647 22457 18659 22460
rect 18601 22451 18659 22457
rect 19978 22448 19984 22460
rect 20036 22488 20042 22500
rect 20073 22491 20131 22497
rect 20073 22488 20085 22491
rect 20036 22460 20085 22488
rect 20036 22448 20042 22460
rect 20073 22457 20085 22460
rect 20119 22488 20131 22491
rect 20441 22491 20499 22497
rect 20441 22488 20453 22491
rect 20119 22460 20453 22488
rect 20119 22457 20131 22460
rect 20073 22451 20131 22457
rect 20441 22457 20453 22460
rect 20487 22457 20499 22491
rect 20441 22451 20499 22457
rect 16040 22392 16988 22420
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 7742 22176 7748 22228
rect 7800 22216 7806 22228
rect 7837 22219 7895 22225
rect 7837 22216 7849 22219
rect 7800 22188 7849 22216
rect 7800 22176 7806 22188
rect 7837 22185 7849 22188
rect 7883 22185 7895 22219
rect 7837 22179 7895 22185
rect 1857 22151 1915 22157
rect 1857 22117 1869 22151
rect 1903 22148 1915 22151
rect 1946 22148 1952 22160
rect 1903 22120 1952 22148
rect 1903 22117 1915 22120
rect 1857 22111 1915 22117
rect 1946 22108 1952 22120
rect 2004 22108 2010 22160
rect 6086 22148 6092 22160
rect 6047 22120 6092 22148
rect 6086 22108 6092 22120
rect 6144 22108 6150 22160
rect 6178 22108 6184 22160
rect 6236 22148 6242 22160
rect 7852 22148 7880 22179
rect 7926 22176 7932 22228
rect 7984 22216 7990 22228
rect 12069 22219 12127 22225
rect 7984 22188 8248 22216
rect 7984 22176 7990 22188
rect 8220 22157 8248 22188
rect 12069 22185 12081 22219
rect 12115 22216 12127 22219
rect 12529 22219 12587 22225
rect 12529 22216 12541 22219
rect 12115 22188 12541 22216
rect 12115 22185 12127 22188
rect 12069 22179 12127 22185
rect 12529 22185 12541 22188
rect 12575 22216 12587 22219
rect 12618 22216 12624 22228
rect 12575 22188 12624 22216
rect 12575 22185 12587 22188
rect 12529 22179 12587 22185
rect 12618 22176 12624 22188
rect 12676 22176 12682 22228
rect 14366 22176 14372 22228
rect 14424 22216 14430 22228
rect 14645 22219 14703 22225
rect 14645 22216 14657 22219
rect 14424 22188 14657 22216
rect 14424 22176 14430 22188
rect 14645 22185 14657 22188
rect 14691 22185 14703 22219
rect 14645 22179 14703 22185
rect 15105 22219 15163 22225
rect 15105 22185 15117 22219
rect 15151 22216 15163 22219
rect 15378 22216 15384 22228
rect 15151 22188 15384 22216
rect 15151 22185 15163 22188
rect 15105 22179 15163 22185
rect 15378 22176 15384 22188
rect 15436 22176 15442 22228
rect 20346 22216 20352 22228
rect 20307 22188 20352 22216
rect 20346 22176 20352 22188
rect 20404 22176 20410 22228
rect 8113 22151 8171 22157
rect 8113 22148 8125 22151
rect 6236 22120 6281 22148
rect 7852 22120 8125 22148
rect 6236 22108 6242 22120
rect 8113 22117 8125 22120
rect 8159 22117 8171 22151
rect 8113 22111 8171 22117
rect 8205 22151 8263 22157
rect 8205 22117 8217 22151
rect 8251 22117 8263 22151
rect 8205 22111 8263 22117
rect 11238 22108 11244 22160
rect 11296 22148 11302 22160
rect 11470 22151 11528 22157
rect 11470 22148 11482 22151
rect 11296 22120 11482 22148
rect 11296 22108 11302 22120
rect 11470 22117 11482 22120
rect 11516 22117 11528 22151
rect 11470 22111 11528 22117
rect 13081 22151 13139 22157
rect 13081 22117 13093 22151
rect 13127 22148 13139 22151
rect 13446 22148 13452 22160
rect 13127 22120 13452 22148
rect 13127 22117 13139 22120
rect 13081 22111 13139 22117
rect 13446 22108 13452 22120
rect 13504 22108 13510 22160
rect 14277 22151 14335 22157
rect 14277 22117 14289 22151
rect 14323 22148 14335 22151
rect 14458 22148 14464 22160
rect 14323 22120 14464 22148
rect 14323 22117 14335 22120
rect 14277 22111 14335 22117
rect 14458 22108 14464 22120
rect 14516 22148 14522 22160
rect 15286 22148 15292 22160
rect 14516 22120 15292 22148
rect 14516 22108 14522 22120
rect 15286 22108 15292 22120
rect 15344 22148 15350 22160
rect 15565 22151 15623 22157
rect 15565 22148 15577 22151
rect 15344 22120 15577 22148
rect 15344 22108 15350 22120
rect 15565 22117 15577 22120
rect 15611 22148 15623 22151
rect 15746 22148 15752 22160
rect 15611 22120 15752 22148
rect 15611 22117 15623 22120
rect 15565 22111 15623 22117
rect 15746 22108 15752 22120
rect 15804 22108 15810 22160
rect 16117 22151 16175 22157
rect 16117 22117 16129 22151
rect 16163 22148 16175 22151
rect 16206 22148 16212 22160
rect 16163 22120 16212 22148
rect 16163 22117 16175 22120
rect 16117 22111 16175 22117
rect 16206 22108 16212 22120
rect 16264 22108 16270 22160
rect 18322 22148 18328 22160
rect 18283 22120 18328 22148
rect 18322 22108 18328 22120
rect 18380 22108 18386 22160
rect 18414 22108 18420 22160
rect 18472 22148 18478 22160
rect 18472 22120 18517 22148
rect 18472 22108 18478 22120
rect 20990 22108 20996 22160
rect 21048 22148 21054 22160
rect 21085 22151 21143 22157
rect 21085 22148 21097 22151
rect 21048 22120 21097 22148
rect 21048 22108 21054 22120
rect 21085 22117 21097 22120
rect 21131 22117 21143 22151
rect 21085 22111 21143 22117
rect 4614 22080 4620 22092
rect 4575 22052 4620 22080
rect 4614 22040 4620 22052
rect 4672 22040 4678 22092
rect 9582 22080 9588 22092
rect 9543 22052 9588 22080
rect 9582 22040 9588 22052
rect 9640 22040 9646 22092
rect 1765 22015 1823 22021
rect 1765 21981 1777 22015
rect 1811 22012 1823 22015
rect 1854 22012 1860 22024
rect 1811 21984 1860 22012
rect 1811 21981 1823 21984
rect 1765 21975 1823 21981
rect 1854 21972 1860 21984
rect 1912 21972 1918 22024
rect 2409 22015 2467 22021
rect 2409 21981 2421 22015
rect 2455 22012 2467 22015
rect 2498 22012 2504 22024
rect 2455 21984 2504 22012
rect 2455 21981 2467 21984
rect 2409 21975 2467 21981
rect 2498 21972 2504 21984
rect 2556 22012 2562 22024
rect 3053 22015 3111 22021
rect 3053 22012 3065 22015
rect 2556 21984 3065 22012
rect 2556 21972 2562 21984
rect 3053 21981 3065 21984
rect 3099 21981 3111 22015
rect 6362 22012 6368 22024
rect 6323 21984 6368 22012
rect 3053 21975 3111 21981
rect 6362 21972 6368 21984
rect 6420 21972 6426 22024
rect 8754 22012 8760 22024
rect 8715 21984 8760 22012
rect 8754 21972 8760 21984
rect 8812 21972 8818 22024
rect 11146 22012 11152 22024
rect 11107 21984 11152 22012
rect 11146 21972 11152 21984
rect 11204 21972 11210 22024
rect 12986 22012 12992 22024
rect 12947 21984 12992 22012
rect 12986 21972 12992 21984
rect 13044 21972 13050 22024
rect 13262 22012 13268 22024
rect 13223 21984 13268 22012
rect 13262 21972 13268 21984
rect 13320 21972 13326 22024
rect 15473 22015 15531 22021
rect 15473 21981 15485 22015
rect 15519 22012 15531 22015
rect 15930 22012 15936 22024
rect 15519 21984 15936 22012
rect 15519 21981 15531 21984
rect 15473 21975 15531 21981
rect 15930 21972 15936 21984
rect 15988 22012 15994 22024
rect 16945 22015 17003 22021
rect 16945 22012 16957 22015
rect 15988 21984 16957 22012
rect 15988 21972 15994 21984
rect 16945 21981 16957 21984
rect 16991 21981 17003 22015
rect 18966 22012 18972 22024
rect 18927 21984 18972 22012
rect 16945 21975 17003 21981
rect 18966 21972 18972 21984
rect 19024 21972 19030 22024
rect 20993 22015 21051 22021
rect 20993 21981 21005 22015
rect 21039 22012 21051 22015
rect 21082 22012 21088 22024
rect 21039 21984 21088 22012
rect 21039 21981 21051 21984
rect 20993 21975 21051 21981
rect 21082 21972 21088 21984
rect 21140 21972 21146 22024
rect 21266 22012 21272 22024
rect 21227 21984 21272 22012
rect 21266 21972 21272 21984
rect 21324 21972 21330 22024
rect 1872 21944 1900 21972
rect 2685 21947 2743 21953
rect 2685 21944 2697 21947
rect 1872 21916 2697 21944
rect 2685 21913 2697 21916
rect 2731 21913 2743 21947
rect 2685 21907 2743 21913
rect 6822 21904 6828 21956
rect 6880 21944 6886 21956
rect 11330 21944 11336 21956
rect 6880 21916 11336 21944
rect 6880 21904 6886 21916
rect 10796 21888 10824 21916
rect 11330 21904 11336 21916
rect 11388 21904 11394 21956
rect 12066 21904 12072 21956
rect 12124 21944 12130 21956
rect 13909 21947 13967 21953
rect 13909 21944 13921 21947
rect 12124 21916 13921 21944
rect 12124 21904 12130 21916
rect 13909 21913 13921 21916
rect 13955 21913 13967 21947
rect 19886 21944 19892 21956
rect 19799 21916 19892 21944
rect 13909 21907 13967 21913
rect 19886 21904 19892 21916
rect 19944 21944 19950 21956
rect 21284 21944 21312 21972
rect 19944 21916 21312 21944
rect 19944 21904 19950 21916
rect 3602 21876 3608 21888
rect 3563 21848 3608 21876
rect 3602 21836 3608 21848
rect 3660 21836 3666 21888
rect 4706 21876 4712 21888
rect 4667 21848 4712 21876
rect 4706 21836 4712 21848
rect 4764 21836 4770 21888
rect 5534 21876 5540 21888
rect 5495 21848 5540 21876
rect 5534 21836 5540 21848
rect 5592 21836 5598 21888
rect 9398 21836 9404 21888
rect 9456 21876 9462 21888
rect 9815 21879 9873 21885
rect 9815 21876 9827 21879
rect 9456 21848 9827 21876
rect 9456 21836 9462 21848
rect 9815 21845 9827 21848
rect 9861 21845 9873 21879
rect 9815 21839 9873 21845
rect 10042 21836 10048 21888
rect 10100 21876 10106 21888
rect 10137 21879 10195 21885
rect 10137 21876 10149 21879
rect 10100 21848 10149 21876
rect 10100 21836 10106 21848
rect 10137 21845 10149 21848
rect 10183 21845 10195 21879
rect 10778 21876 10784 21888
rect 10739 21848 10784 21876
rect 10137 21839 10195 21845
rect 10778 21836 10784 21848
rect 10836 21836 10842 21888
rect 13814 21836 13820 21888
rect 13872 21876 13878 21888
rect 16393 21879 16451 21885
rect 16393 21876 16405 21879
rect 13872 21848 16405 21876
rect 13872 21836 13878 21848
rect 16393 21845 16405 21848
rect 16439 21876 16451 21879
rect 16482 21876 16488 21888
rect 16439 21848 16488 21876
rect 16439 21845 16451 21848
rect 16393 21839 16451 21845
rect 16482 21836 16488 21848
rect 16540 21836 16546 21888
rect 18046 21876 18052 21888
rect 18007 21848 18052 21876
rect 18046 21836 18052 21848
rect 18104 21836 18110 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1762 21672 1768 21684
rect 1723 21644 1768 21672
rect 1762 21632 1768 21644
rect 1820 21632 1826 21684
rect 4614 21672 4620 21684
rect 4575 21644 4620 21672
rect 4614 21632 4620 21644
rect 4672 21632 4678 21684
rect 5077 21675 5135 21681
rect 5077 21641 5089 21675
rect 5123 21672 5135 21675
rect 5258 21672 5264 21684
rect 5123 21644 5264 21672
rect 5123 21641 5135 21644
rect 5077 21635 5135 21641
rect 5258 21632 5264 21644
rect 5316 21632 5322 21684
rect 6178 21672 6184 21684
rect 6139 21644 6184 21672
rect 6178 21632 6184 21644
rect 6236 21632 6242 21684
rect 11146 21632 11152 21684
rect 11204 21672 11210 21684
rect 11517 21675 11575 21681
rect 11517 21672 11529 21675
rect 11204 21644 11529 21672
rect 11204 21632 11210 21644
rect 11517 21641 11529 21644
rect 11563 21641 11575 21675
rect 11517 21635 11575 21641
rect 12434 21632 12440 21684
rect 12492 21672 12498 21684
rect 13538 21672 13544 21684
rect 12492 21644 13544 21672
rect 12492 21632 12498 21644
rect 13538 21632 13544 21644
rect 13596 21632 13602 21684
rect 15470 21632 15476 21684
rect 15528 21672 15534 21684
rect 15565 21675 15623 21681
rect 15565 21672 15577 21675
rect 15528 21644 15577 21672
rect 15528 21632 15534 21644
rect 15565 21641 15577 21644
rect 15611 21641 15623 21675
rect 15930 21672 15936 21684
rect 15891 21644 15936 21672
rect 15565 21635 15623 21641
rect 15930 21632 15936 21644
rect 15988 21632 15994 21684
rect 17497 21675 17555 21681
rect 17497 21641 17509 21675
rect 17543 21672 17555 21675
rect 18322 21672 18328 21684
rect 17543 21644 18328 21672
rect 17543 21641 17555 21644
rect 17497 21635 17555 21641
rect 18322 21632 18328 21644
rect 18380 21632 18386 21684
rect 18414 21632 18420 21684
rect 18472 21672 18478 21684
rect 18969 21675 19027 21681
rect 18969 21672 18981 21675
rect 18472 21644 18981 21672
rect 18472 21632 18478 21644
rect 18969 21641 18981 21644
rect 19015 21672 19027 21675
rect 20901 21675 20959 21681
rect 20901 21672 20913 21675
rect 19015 21644 20913 21672
rect 19015 21641 19027 21644
rect 18969 21635 19027 21641
rect 20901 21641 20913 21644
rect 20947 21672 20959 21675
rect 20990 21672 20996 21684
rect 20947 21644 20996 21672
rect 20947 21641 20959 21644
rect 20901 21635 20959 21641
rect 20990 21632 20996 21644
rect 21048 21632 21054 21684
rect 21910 21672 21916 21684
rect 21871 21644 21916 21672
rect 21910 21632 21916 21644
rect 21968 21632 21974 21684
rect 25130 21672 25136 21684
rect 25091 21644 25136 21672
rect 25130 21632 25136 21644
rect 25188 21632 25194 21684
rect 2961 21607 3019 21613
rect 2961 21604 2973 21607
rect 2056 21576 2973 21604
rect 2056 21548 2084 21576
rect 2961 21573 2973 21576
rect 3007 21573 3019 21607
rect 2961 21567 3019 21573
rect 8386 21564 8392 21616
rect 8444 21604 8450 21616
rect 12066 21604 12072 21616
rect 8444 21576 8524 21604
rect 8444 21564 8450 21576
rect 2038 21536 2044 21548
rect 1999 21508 2044 21536
rect 2038 21496 2044 21508
rect 2096 21496 2102 21548
rect 2498 21536 2504 21548
rect 2459 21508 2504 21536
rect 2498 21496 2504 21508
rect 2556 21496 2562 21548
rect 3878 21536 3884 21548
rect 3839 21508 3884 21536
rect 3878 21496 3884 21508
rect 3936 21496 3942 21548
rect 5261 21539 5319 21545
rect 5261 21505 5273 21539
rect 5307 21536 5319 21539
rect 5534 21536 5540 21548
rect 5307 21508 5540 21536
rect 5307 21505 5319 21508
rect 5261 21499 5319 21505
rect 5534 21496 5540 21508
rect 5592 21496 5598 21548
rect 5905 21539 5963 21545
rect 5905 21505 5917 21539
rect 5951 21536 5963 21539
rect 6362 21536 6368 21548
rect 5951 21508 6368 21536
rect 5951 21505 5963 21508
rect 5905 21499 5963 21505
rect 6362 21496 6368 21508
rect 6420 21496 6426 21548
rect 8496 21545 8524 21576
rect 8772 21576 12072 21604
rect 8772 21548 8800 21576
rect 12066 21564 12072 21576
rect 12124 21604 12130 21616
rect 12124 21576 12572 21604
rect 12124 21564 12130 21576
rect 8481 21539 8539 21545
rect 8481 21505 8493 21539
rect 8527 21505 8539 21539
rect 8754 21536 8760 21548
rect 8715 21508 8760 21536
rect 8481 21499 8539 21505
rect 8754 21496 8760 21508
rect 8812 21496 8818 21548
rect 8938 21496 8944 21548
rect 8996 21536 9002 21548
rect 12544 21545 12572 21576
rect 16574 21564 16580 21616
rect 16632 21604 16638 21616
rect 21499 21607 21557 21613
rect 21499 21604 21511 21607
rect 16632 21576 21511 21604
rect 16632 21564 16638 21576
rect 21499 21573 21511 21576
rect 21545 21573 21557 21607
rect 21499 21567 21557 21573
rect 10321 21539 10379 21545
rect 10321 21536 10333 21539
rect 8996 21508 10333 21536
rect 8996 21496 9002 21508
rect 10321 21505 10333 21508
rect 10367 21505 10379 21539
rect 10321 21499 10379 21505
rect 12529 21539 12587 21545
rect 12529 21505 12541 21539
rect 12575 21505 12587 21539
rect 12529 21499 12587 21505
rect 13173 21539 13231 21545
rect 13173 21505 13185 21539
rect 13219 21536 13231 21539
rect 13262 21536 13268 21548
rect 13219 21508 13268 21536
rect 13219 21505 13231 21508
rect 13173 21499 13231 21505
rect 13262 21496 13268 21508
rect 13320 21496 13326 21548
rect 14642 21536 14648 21548
rect 14603 21508 14648 21536
rect 14642 21496 14648 21508
rect 14700 21496 14706 21548
rect 17129 21539 17187 21545
rect 17129 21505 17141 21539
rect 17175 21536 17187 21539
rect 18046 21536 18052 21548
rect 17175 21508 18052 21536
rect 17175 21505 17187 21508
rect 17129 21499 17187 21505
rect 18046 21496 18052 21508
rect 18104 21496 18110 21548
rect 19886 21536 19892 21548
rect 19847 21508 19892 21536
rect 19886 21496 19892 21508
rect 19944 21496 19950 21548
rect 5994 21428 6000 21480
rect 6052 21468 6058 21480
rect 6641 21471 6699 21477
rect 6641 21468 6653 21471
rect 6052 21440 6653 21468
rect 6052 21428 6058 21440
rect 6641 21437 6653 21440
rect 6687 21468 6699 21471
rect 6825 21471 6883 21477
rect 6825 21468 6837 21471
rect 6687 21440 6837 21468
rect 6687 21437 6699 21440
rect 6641 21431 6699 21437
rect 6825 21437 6837 21440
rect 6871 21437 6883 21471
rect 6825 21431 6883 21437
rect 6914 21428 6920 21480
rect 6972 21468 6978 21480
rect 7285 21471 7343 21477
rect 7285 21468 7297 21471
rect 6972 21440 7297 21468
rect 6972 21428 6978 21440
rect 7285 21437 7297 21440
rect 7331 21437 7343 21471
rect 7285 21431 7343 21437
rect 13538 21428 13544 21480
rect 13596 21468 13602 21480
rect 16482 21468 16488 21480
rect 13596 21440 14596 21468
rect 16443 21440 16488 21468
rect 13596 21428 13602 21440
rect 1762 21360 1768 21412
rect 1820 21400 1826 21412
rect 2133 21403 2191 21409
rect 2133 21400 2145 21403
rect 1820 21372 2145 21400
rect 1820 21360 1826 21372
rect 2133 21369 2145 21372
rect 2179 21400 2191 21403
rect 3329 21403 3387 21409
rect 3329 21400 3341 21403
rect 2179 21372 3341 21400
rect 2179 21369 2191 21372
rect 2133 21363 2191 21369
rect 3329 21369 3341 21372
rect 3375 21369 3387 21403
rect 3602 21400 3608 21412
rect 3563 21372 3608 21400
rect 3329 21363 3387 21369
rect 3344 21332 3372 21363
rect 3602 21360 3608 21372
rect 3660 21360 3666 21412
rect 3697 21403 3755 21409
rect 3697 21369 3709 21403
rect 3743 21369 3755 21403
rect 3697 21363 3755 21369
rect 3712 21332 3740 21363
rect 5350 21360 5356 21412
rect 5408 21400 5414 21412
rect 5408 21372 5453 21400
rect 5408 21360 5414 21372
rect 7466 21360 7472 21412
rect 7524 21400 7530 21412
rect 7561 21403 7619 21409
rect 7561 21400 7573 21403
rect 7524 21372 7573 21400
rect 7524 21360 7530 21372
rect 7561 21369 7573 21372
rect 7607 21369 7619 21403
rect 8570 21400 8576 21412
rect 8531 21372 8576 21400
rect 7561 21363 7619 21369
rect 8570 21360 8576 21372
rect 8628 21360 8634 21412
rect 9766 21360 9772 21412
rect 9824 21400 9830 21412
rect 10042 21400 10048 21412
rect 9824 21372 10048 21400
rect 9824 21360 9830 21372
rect 10042 21360 10048 21372
rect 10100 21360 10106 21412
rect 10134 21360 10140 21412
rect 10192 21400 10198 21412
rect 12621 21403 12679 21409
rect 10192 21372 10237 21400
rect 10192 21360 10198 21372
rect 12621 21369 12633 21403
rect 12667 21369 12679 21403
rect 12621 21363 12679 21369
rect 3344 21304 3740 21332
rect 7926 21292 7932 21344
rect 7984 21332 7990 21344
rect 8021 21335 8079 21341
rect 8021 21332 8033 21335
rect 7984 21304 8033 21332
rect 7984 21292 7990 21304
rect 8021 21301 8033 21304
rect 8067 21301 8079 21335
rect 8021 21295 8079 21301
rect 8662 21292 8668 21344
rect 8720 21332 8726 21344
rect 9582 21332 9588 21344
rect 8720 21304 9588 21332
rect 8720 21292 8726 21304
rect 9582 21292 9588 21304
rect 9640 21332 9646 21344
rect 9677 21335 9735 21341
rect 9677 21332 9689 21335
rect 9640 21304 9689 21332
rect 9640 21292 9646 21304
rect 9677 21301 9689 21304
rect 9723 21301 9735 21335
rect 11238 21332 11244 21344
rect 11199 21304 11244 21332
rect 9677 21295 9735 21301
rect 11238 21292 11244 21304
rect 11296 21292 11302 21344
rect 12158 21332 12164 21344
rect 12119 21304 12164 21332
rect 12158 21292 12164 21304
rect 12216 21332 12222 21344
rect 12636 21332 12664 21363
rect 12986 21360 12992 21412
rect 13044 21400 13050 21412
rect 13817 21403 13875 21409
rect 13817 21400 13829 21403
rect 13044 21372 13829 21400
rect 13044 21360 13050 21372
rect 13817 21369 13829 21372
rect 13863 21369 13875 21403
rect 13817 21363 13875 21369
rect 13446 21332 13452 21344
rect 12216 21304 12664 21332
rect 13407 21304 13452 21332
rect 12216 21292 12222 21304
rect 13446 21292 13452 21304
rect 13504 21292 13510 21344
rect 14568 21341 14596 21440
rect 16482 21428 16488 21440
rect 16540 21428 16546 21480
rect 16853 21471 16911 21477
rect 16853 21437 16865 21471
rect 16899 21437 16911 21471
rect 16853 21431 16911 21437
rect 21428 21471 21486 21477
rect 21428 21437 21440 21471
rect 21474 21468 21486 21471
rect 21910 21468 21916 21480
rect 21474 21440 21916 21468
rect 21474 21437 21486 21440
rect 21428 21431 21486 21437
rect 15007 21403 15065 21409
rect 15007 21369 15019 21403
rect 15053 21369 15065 21403
rect 15007 21363 15065 21369
rect 16301 21403 16359 21409
rect 16301 21369 16313 21403
rect 16347 21400 16359 21403
rect 16868 21400 16896 21431
rect 21910 21428 21916 21440
rect 21968 21428 21974 21480
rect 24648 21471 24706 21477
rect 24648 21437 24660 21471
rect 24694 21468 24706 21471
rect 25130 21468 25136 21480
rect 24694 21440 25136 21468
rect 24694 21437 24706 21440
rect 24648 21431 24706 21437
rect 25130 21428 25136 21440
rect 25188 21428 25194 21480
rect 17126 21400 17132 21412
rect 16347 21372 17132 21400
rect 16347 21369 16359 21372
rect 16301 21363 16359 21369
rect 14553 21335 14611 21341
rect 14553 21301 14565 21335
rect 14599 21332 14611 21335
rect 15022 21332 15050 21363
rect 17126 21360 17132 21372
rect 17184 21360 17190 21412
rect 18370 21403 18428 21409
rect 18370 21369 18382 21403
rect 18416 21369 18428 21403
rect 18370 21363 18428 21369
rect 19981 21403 20039 21409
rect 19981 21369 19993 21403
rect 20027 21369 20039 21403
rect 20530 21400 20536 21412
rect 20491 21372 20536 21400
rect 19981 21363 20039 21369
rect 15378 21332 15384 21344
rect 14599 21304 15384 21332
rect 14599 21301 14611 21304
rect 14553 21295 14611 21301
rect 15378 21292 15384 21304
rect 15436 21292 15442 21344
rect 17770 21332 17776 21344
rect 17731 21304 17776 21332
rect 17770 21292 17776 21304
rect 17828 21332 17834 21344
rect 18385 21332 18413 21363
rect 17828 21304 18413 21332
rect 17828 21292 17834 21304
rect 19518 21292 19524 21344
rect 19576 21332 19582 21344
rect 19705 21335 19763 21341
rect 19705 21332 19717 21335
rect 19576 21304 19717 21332
rect 19576 21292 19582 21304
rect 19705 21301 19717 21304
rect 19751 21332 19763 21335
rect 19996 21332 20024 21363
rect 20530 21360 20536 21372
rect 20588 21360 20594 21412
rect 19751 21304 20024 21332
rect 19751 21301 19763 21304
rect 19705 21295 19763 21301
rect 20438 21292 20444 21344
rect 20496 21332 20502 21344
rect 24719 21335 24777 21341
rect 24719 21332 24731 21335
rect 20496 21304 24731 21332
rect 20496 21292 20502 21304
rect 24719 21301 24731 21304
rect 24765 21301 24777 21335
rect 24719 21295 24777 21301
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 2866 21128 2872 21140
rect 2608 21100 2872 21128
rect 1765 21063 1823 21069
rect 1765 21029 1777 21063
rect 1811 21060 1823 21063
rect 2038 21060 2044 21072
rect 1811 21032 2044 21060
rect 1811 21029 1823 21032
rect 1765 21023 1823 21029
rect 2038 21020 2044 21032
rect 2096 21020 2102 21072
rect 2608 21069 2636 21100
rect 2866 21088 2872 21100
rect 2924 21128 2930 21140
rect 3697 21131 3755 21137
rect 3697 21128 3709 21131
rect 2924 21100 3709 21128
rect 2924 21088 2930 21100
rect 3697 21097 3709 21100
rect 3743 21128 3755 21131
rect 3878 21128 3884 21140
rect 3743 21100 3884 21128
rect 3743 21097 3755 21100
rect 3697 21091 3755 21097
rect 3878 21088 3884 21100
rect 3936 21088 3942 21140
rect 5350 21088 5356 21140
rect 5408 21128 5414 21140
rect 5813 21131 5871 21137
rect 5813 21128 5825 21131
rect 5408 21100 5825 21128
rect 5408 21088 5414 21100
rect 5813 21097 5825 21100
rect 5859 21097 5871 21131
rect 6086 21128 6092 21140
rect 6047 21100 6092 21128
rect 5813 21091 5871 21097
rect 6086 21088 6092 21100
rect 6144 21088 6150 21140
rect 6822 21128 6828 21140
rect 6783 21100 6828 21128
rect 6822 21088 6828 21100
rect 6880 21088 6886 21140
rect 7742 21088 7748 21140
rect 7800 21128 7806 21140
rect 7837 21131 7895 21137
rect 7837 21128 7849 21131
rect 7800 21100 7849 21128
rect 7800 21088 7806 21100
rect 7837 21097 7849 21100
rect 7883 21097 7895 21131
rect 7837 21091 7895 21097
rect 8386 21088 8392 21140
rect 8444 21128 8450 21140
rect 9033 21131 9091 21137
rect 9033 21128 9045 21131
rect 8444 21100 9045 21128
rect 8444 21088 8450 21100
rect 9033 21097 9045 21100
rect 9079 21097 9091 21131
rect 9033 21091 9091 21097
rect 11977 21131 12035 21137
rect 11977 21097 11989 21131
rect 12023 21128 12035 21131
rect 12158 21128 12164 21140
rect 12023 21100 12164 21128
rect 12023 21097 12035 21100
rect 11977 21091 12035 21097
rect 12158 21088 12164 21100
rect 12216 21088 12222 21140
rect 14642 21128 14648 21140
rect 14603 21100 14648 21128
rect 14642 21088 14648 21100
rect 14700 21088 14706 21140
rect 15105 21131 15163 21137
rect 15105 21097 15117 21131
rect 15151 21128 15163 21131
rect 15286 21128 15292 21140
rect 15151 21100 15292 21128
rect 15151 21097 15163 21100
rect 15105 21091 15163 21097
rect 15286 21088 15292 21100
rect 15344 21128 15350 21140
rect 16209 21131 16267 21137
rect 16209 21128 16221 21131
rect 15344 21100 16221 21128
rect 15344 21088 15350 21100
rect 16209 21097 16221 21100
rect 16255 21097 16267 21131
rect 16574 21128 16580 21140
rect 16535 21100 16580 21128
rect 16209 21091 16267 21097
rect 16574 21088 16580 21100
rect 16632 21088 16638 21140
rect 18325 21131 18383 21137
rect 18325 21097 18337 21131
rect 18371 21128 18383 21131
rect 18414 21128 18420 21140
rect 18371 21100 18420 21128
rect 18371 21097 18383 21100
rect 18325 21091 18383 21097
rect 18414 21088 18420 21100
rect 18472 21088 18478 21140
rect 19058 21128 19064 21140
rect 19019 21100 19064 21128
rect 19058 21088 19064 21100
rect 19116 21088 19122 21140
rect 19518 21088 19524 21140
rect 19576 21128 19582 21140
rect 19613 21131 19671 21137
rect 19613 21128 19625 21131
rect 19576 21100 19625 21128
rect 19576 21088 19582 21100
rect 19613 21097 19625 21100
rect 19659 21097 19671 21131
rect 19978 21128 19984 21140
rect 19939 21100 19984 21128
rect 19613 21091 19671 21097
rect 19978 21088 19984 21100
rect 20036 21088 20042 21140
rect 21082 21088 21088 21140
rect 21140 21128 21146 21140
rect 21361 21131 21419 21137
rect 21361 21128 21373 21131
rect 21140 21100 21373 21128
rect 21140 21088 21146 21100
rect 21361 21097 21373 21100
rect 21407 21097 21419 21131
rect 21361 21091 21419 21097
rect 2593 21063 2651 21069
rect 2593 21029 2605 21063
rect 2639 21029 2651 21063
rect 3234 21060 3240 21072
rect 3195 21032 3240 21060
rect 2593 21023 2651 21029
rect 3234 21020 3240 21032
rect 3292 21020 3298 21072
rect 3510 21020 3516 21072
rect 3568 21060 3574 21072
rect 3568 21032 4154 21060
rect 3568 21020 3574 21032
rect 1949 20927 2007 20933
rect 1949 20893 1961 20927
rect 1995 20924 2007 20927
rect 3252 20924 3280 21020
rect 4126 20992 4154 21032
rect 4890 21020 4896 21072
rect 4948 21060 4954 21072
rect 5214 21063 5272 21069
rect 5214 21060 5226 21063
rect 4948 21032 5226 21060
rect 4948 21020 4954 21032
rect 5214 21029 5226 21032
rect 5260 21029 5272 21063
rect 5214 21023 5272 21029
rect 7926 21020 7932 21072
rect 7984 21060 7990 21072
rect 10134 21060 10140 21072
rect 7984 21032 10140 21060
rect 7984 21020 7990 21032
rect 10134 21020 10140 21032
rect 10192 21020 10198 21072
rect 11238 21020 11244 21072
rect 11296 21060 11302 21072
rect 11419 21063 11477 21069
rect 11419 21060 11431 21063
rect 11296 21032 11431 21060
rect 11296 21020 11302 21032
rect 11419 21029 11431 21032
rect 11465 21060 11477 21063
rect 13167 21063 13225 21069
rect 13167 21060 13179 21063
rect 11465 21032 13179 21060
rect 11465 21029 11477 21032
rect 11419 21023 11477 21029
rect 13167 21029 13179 21032
rect 13213 21060 13225 21063
rect 13538 21060 13544 21072
rect 13213 21032 13544 21060
rect 13213 21029 13225 21032
rect 13167 21023 13225 21029
rect 13538 21020 13544 21032
rect 13596 21020 13602 21072
rect 15378 21020 15384 21072
rect 15436 21060 15442 21072
rect 15610 21063 15668 21069
rect 15610 21060 15622 21063
rect 15436 21032 15622 21060
rect 15436 21020 15442 21032
rect 15610 21029 15622 21032
rect 15656 21029 15668 21063
rect 15610 21023 15668 21029
rect 8110 20992 8116 21004
rect 4126 20964 8116 20992
rect 8110 20952 8116 20964
rect 8168 20952 8174 21004
rect 8202 20952 8208 21004
rect 8260 20992 8266 21004
rect 9306 20992 9312 21004
rect 8260 20964 9312 20992
rect 8260 20952 8266 20964
rect 9306 20952 9312 20964
rect 9364 20992 9370 21004
rect 9712 20995 9770 21001
rect 9712 20992 9724 20995
rect 9364 20964 9724 20992
rect 9364 20952 9370 20964
rect 9712 20961 9724 20964
rect 9758 20961 9770 20995
rect 11054 20992 11060 21004
rect 11015 20964 11060 20992
rect 9712 20955 9770 20961
rect 11054 20952 11060 20964
rect 11112 20952 11118 21004
rect 14826 20952 14832 21004
rect 14884 20992 14890 21004
rect 15289 20995 15347 21001
rect 15289 20992 15301 20995
rect 14884 20964 15301 20992
rect 14884 20952 14890 20964
rect 15289 20961 15301 20964
rect 15335 20961 15347 20995
rect 15289 20955 15347 20961
rect 16758 20952 16764 21004
rect 16816 20992 16822 21004
rect 17129 20995 17187 21001
rect 17129 20992 17141 20995
rect 16816 20964 17141 20992
rect 16816 20952 16822 20964
rect 17129 20961 17141 20964
rect 17175 20961 17187 20995
rect 17129 20955 17187 20961
rect 17218 20952 17224 21004
rect 17276 20992 17282 21004
rect 17589 20995 17647 21001
rect 17589 20992 17601 20995
rect 17276 20964 17601 20992
rect 17276 20952 17282 20964
rect 17589 20961 17601 20964
rect 17635 20961 17647 20995
rect 17589 20955 17647 20961
rect 1995 20896 3280 20924
rect 1995 20893 2007 20896
rect 1949 20887 2007 20893
rect 4522 20884 4528 20936
rect 4580 20924 4586 20936
rect 4893 20927 4951 20933
rect 4893 20924 4905 20927
rect 4580 20896 4905 20924
rect 4580 20884 4586 20896
rect 4893 20893 4905 20896
rect 4939 20893 4951 20927
rect 7466 20924 7472 20936
rect 7427 20896 7472 20924
rect 4893 20887 4951 20893
rect 7466 20884 7472 20896
rect 7524 20884 7530 20936
rect 12802 20924 12808 20936
rect 12763 20896 12808 20924
rect 12802 20884 12808 20896
rect 12860 20884 12866 20936
rect 17862 20924 17868 20936
rect 17823 20896 17868 20924
rect 17862 20884 17868 20896
rect 17920 20884 17926 20936
rect 18690 20924 18696 20936
rect 18651 20896 18696 20924
rect 18690 20884 18696 20896
rect 18748 20884 18754 20936
rect 19978 20884 19984 20936
rect 20036 20924 20042 20936
rect 20901 20927 20959 20933
rect 20901 20924 20913 20927
rect 20036 20896 20913 20924
rect 20036 20884 20042 20896
rect 20901 20893 20913 20896
rect 20947 20893 20959 20927
rect 20901 20887 20959 20893
rect 2958 20788 2964 20800
rect 2919 20760 2964 20788
rect 2958 20748 2964 20760
rect 3016 20748 3022 20800
rect 8389 20791 8447 20797
rect 8389 20757 8401 20791
rect 8435 20788 8447 20791
rect 8570 20788 8576 20800
rect 8435 20760 8576 20788
rect 8435 20757 8447 20760
rect 8389 20751 8447 20757
rect 8570 20748 8576 20760
rect 8628 20788 8634 20800
rect 8757 20791 8815 20797
rect 8757 20788 8769 20791
rect 8628 20760 8769 20788
rect 8628 20748 8634 20760
rect 8757 20757 8769 20760
rect 8803 20788 8815 20791
rect 9582 20788 9588 20800
rect 8803 20760 9588 20788
rect 8803 20757 8815 20760
rect 8757 20751 8815 20757
rect 9582 20748 9588 20760
rect 9640 20748 9646 20800
rect 9674 20748 9680 20800
rect 9732 20788 9738 20800
rect 9815 20791 9873 20797
rect 9815 20788 9827 20791
rect 9732 20760 9827 20788
rect 9732 20748 9738 20760
rect 9815 20757 9827 20760
rect 9861 20757 9873 20791
rect 12526 20788 12532 20800
rect 12487 20760 12532 20788
rect 9815 20751 9873 20757
rect 12526 20748 12532 20760
rect 12584 20748 12590 20800
rect 12618 20748 12624 20800
rect 12676 20788 12682 20800
rect 13725 20791 13783 20797
rect 13725 20788 13737 20791
rect 12676 20760 13737 20788
rect 12676 20748 12682 20760
rect 13725 20757 13737 20760
rect 13771 20757 13783 20791
rect 13725 20751 13783 20757
rect 14093 20791 14151 20797
rect 14093 20757 14105 20791
rect 14139 20788 14151 20791
rect 14366 20788 14372 20800
rect 14139 20760 14372 20788
rect 14139 20757 14151 20760
rect 14093 20751 14151 20757
rect 14366 20748 14372 20760
rect 14424 20748 14430 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1578 20584 1584 20596
rect 1539 20556 1584 20584
rect 1578 20544 1584 20556
rect 1636 20544 1642 20596
rect 4617 20587 4675 20593
rect 4617 20553 4629 20587
rect 4663 20584 4675 20587
rect 4706 20584 4712 20596
rect 4663 20556 4712 20584
rect 4663 20553 4675 20556
rect 4617 20547 4675 20553
rect 4706 20544 4712 20556
rect 4764 20584 4770 20596
rect 5258 20584 5264 20596
rect 4764 20556 5264 20584
rect 4764 20544 4770 20556
rect 5258 20544 5264 20556
rect 5316 20544 5322 20596
rect 8018 20544 8024 20596
rect 8076 20584 8082 20596
rect 10873 20587 10931 20593
rect 10873 20584 10885 20587
rect 8076 20556 10885 20584
rect 8076 20544 8082 20556
rect 10873 20553 10885 20556
rect 10919 20553 10931 20587
rect 10873 20547 10931 20553
rect 11057 20587 11115 20593
rect 11057 20553 11069 20587
rect 11103 20584 11115 20587
rect 11238 20584 11244 20596
rect 11103 20556 11244 20584
rect 11103 20553 11115 20556
rect 11057 20547 11115 20553
rect 11238 20544 11244 20556
rect 11296 20544 11302 20596
rect 13722 20544 13728 20596
rect 13780 20584 13786 20596
rect 13817 20587 13875 20593
rect 13817 20584 13829 20587
rect 13780 20556 13829 20584
rect 13780 20544 13786 20556
rect 13817 20553 13829 20556
rect 13863 20584 13875 20587
rect 16758 20584 16764 20596
rect 13863 20556 16764 20584
rect 13863 20553 13875 20556
rect 13817 20547 13875 20553
rect 3789 20519 3847 20525
rect 3789 20516 3801 20519
rect 1412 20488 3801 20516
rect 1412 20392 1440 20488
rect 3789 20485 3801 20488
rect 3835 20485 3847 20519
rect 6089 20519 6147 20525
rect 6089 20516 6101 20519
rect 3789 20479 3847 20485
rect 5184 20488 6101 20516
rect 2866 20448 2872 20460
rect 2827 20420 2872 20448
rect 2866 20408 2872 20420
rect 2924 20408 2930 20460
rect 3326 20448 3332 20460
rect 3287 20420 3332 20448
rect 3326 20408 3332 20420
rect 3384 20408 3390 20460
rect 4982 20408 4988 20460
rect 5040 20448 5046 20460
rect 5184 20457 5212 20488
rect 6089 20485 6101 20488
rect 6135 20485 6147 20519
rect 6089 20479 6147 20485
rect 8754 20476 8760 20528
rect 8812 20516 8818 20528
rect 10229 20519 10287 20525
rect 10229 20516 10241 20519
rect 8812 20488 10241 20516
rect 8812 20476 8818 20488
rect 10229 20485 10241 20488
rect 10275 20516 10287 20519
rect 12986 20516 12992 20528
rect 10275 20488 12020 20516
rect 10275 20485 10287 20488
rect 10229 20479 10287 20485
rect 5169 20451 5227 20457
rect 5169 20448 5181 20451
rect 5040 20420 5181 20448
rect 5040 20408 5046 20420
rect 5169 20417 5181 20420
rect 5215 20417 5227 20451
rect 5534 20448 5540 20460
rect 5495 20420 5540 20448
rect 5169 20411 5227 20417
rect 5534 20408 5540 20420
rect 5592 20408 5598 20460
rect 7377 20451 7435 20457
rect 7377 20417 7389 20451
rect 7423 20448 7435 20451
rect 8662 20448 8668 20460
rect 7423 20420 8668 20448
rect 7423 20417 7435 20420
rect 7377 20411 7435 20417
rect 1394 20380 1400 20392
rect 1355 20352 1400 20380
rect 1394 20340 1400 20352
rect 1452 20340 1458 20392
rect 6892 20383 6950 20389
rect 6892 20349 6904 20383
rect 6938 20380 6950 20383
rect 7392 20380 7420 20411
rect 8662 20408 8668 20420
rect 8720 20408 8726 20460
rect 9214 20408 9220 20460
rect 9272 20448 9278 20460
rect 11287 20451 11345 20457
rect 11287 20448 11299 20451
rect 9272 20420 11299 20448
rect 9272 20408 9278 20420
rect 11287 20417 11299 20420
rect 11333 20417 11345 20451
rect 11992 20448 12020 20488
rect 12268 20488 12992 20516
rect 12268 20448 12296 20488
rect 12526 20448 12532 20460
rect 11992 20420 12296 20448
rect 12487 20420 12532 20448
rect 11287 20411 11345 20417
rect 12526 20408 12532 20420
rect 12584 20408 12590 20460
rect 12820 20457 12848 20488
rect 12986 20476 12992 20488
rect 13044 20476 13050 20528
rect 12805 20451 12863 20457
rect 12805 20417 12817 20451
rect 12851 20417 12863 20451
rect 13832 20448 13860 20547
rect 16758 20544 16764 20556
rect 16816 20544 16822 20596
rect 17126 20584 17132 20596
rect 17087 20556 17132 20584
rect 17126 20544 17132 20556
rect 17184 20544 17190 20596
rect 18969 20587 19027 20593
rect 18969 20553 18981 20587
rect 19015 20584 19027 20587
rect 19886 20584 19892 20596
rect 19015 20556 19892 20584
rect 19015 20553 19027 20556
rect 18969 20547 19027 20553
rect 19886 20544 19892 20556
rect 19944 20544 19950 20596
rect 20990 20544 20996 20596
rect 21048 20584 21054 20596
rect 21269 20587 21327 20593
rect 21269 20584 21281 20587
rect 21048 20556 21281 20584
rect 21048 20544 21054 20556
rect 21269 20553 21281 20556
rect 21315 20584 21327 20587
rect 21634 20584 21640 20596
rect 21315 20556 21640 20584
rect 21315 20553 21327 20556
rect 21269 20547 21327 20553
rect 21634 20544 21640 20556
rect 21692 20544 21698 20596
rect 16206 20476 16212 20528
rect 16264 20516 16270 20528
rect 16393 20519 16451 20525
rect 16393 20516 16405 20519
rect 16264 20488 16405 20516
rect 16264 20476 16270 20488
rect 16393 20485 16405 20488
rect 16439 20485 16451 20519
rect 16393 20479 16451 20485
rect 13998 20448 14004 20460
rect 13832 20420 14004 20448
rect 12805 20411 12863 20417
rect 13998 20408 14004 20420
rect 14056 20448 14062 20460
rect 15841 20451 15899 20457
rect 14056 20420 14136 20448
rect 14056 20408 14062 20420
rect 14108 20389 14136 20420
rect 15841 20417 15853 20451
rect 15887 20448 15899 20451
rect 16574 20448 16580 20460
rect 15887 20420 16580 20448
rect 15887 20417 15899 20420
rect 15841 20411 15899 20417
rect 16574 20408 16580 20420
rect 16632 20408 16638 20460
rect 17862 20408 17868 20460
rect 17920 20448 17926 20460
rect 18049 20451 18107 20457
rect 18049 20448 18061 20451
rect 17920 20420 18061 20448
rect 17920 20408 17926 20420
rect 18049 20417 18061 20420
rect 18095 20417 18107 20451
rect 18049 20411 18107 20417
rect 19797 20451 19855 20457
rect 19797 20417 19809 20451
rect 19843 20448 19855 20451
rect 19978 20448 19984 20460
rect 19843 20420 19984 20448
rect 19843 20417 19855 20420
rect 19797 20411 19855 20417
rect 19978 20408 19984 20420
rect 20036 20408 20042 20460
rect 20254 20408 20260 20460
rect 20312 20448 20318 20460
rect 20625 20451 20683 20457
rect 20625 20448 20637 20451
rect 20312 20420 20637 20448
rect 20312 20408 20318 20420
rect 20625 20417 20637 20420
rect 20671 20448 20683 20451
rect 21821 20451 21879 20457
rect 21821 20448 21833 20451
rect 20671 20420 21833 20448
rect 20671 20417 20683 20420
rect 20625 20411 20683 20417
rect 21821 20417 21833 20420
rect 21867 20417 21879 20451
rect 21821 20411 21879 20417
rect 6938 20352 7420 20380
rect 7837 20383 7895 20389
rect 6938 20349 6950 20352
rect 6892 20343 6950 20349
rect 7837 20349 7849 20383
rect 7883 20380 7895 20383
rect 10873 20383 10931 20389
rect 7883 20352 9168 20380
rect 7883 20349 7895 20352
rect 7837 20343 7895 20349
rect 2958 20312 2964 20324
rect 2919 20284 2964 20312
rect 2958 20272 2964 20284
rect 3016 20272 3022 20324
rect 3694 20272 3700 20324
rect 3752 20312 3758 20324
rect 4890 20312 4896 20324
rect 3752 20284 4896 20312
rect 3752 20272 3758 20284
rect 4890 20272 4896 20284
rect 4948 20272 4954 20324
rect 5258 20272 5264 20324
rect 5316 20312 5322 20324
rect 7653 20315 7711 20321
rect 7653 20312 7665 20315
rect 5316 20284 5361 20312
rect 6104 20284 7665 20312
rect 5316 20272 5322 20284
rect 1946 20244 1952 20256
rect 1907 20216 1952 20244
rect 1946 20204 1952 20216
rect 2004 20204 2010 20256
rect 2038 20204 2044 20256
rect 2096 20244 2102 20256
rect 2409 20247 2467 20253
rect 2409 20244 2421 20247
rect 2096 20216 2421 20244
rect 2096 20204 2102 20216
rect 2409 20213 2421 20216
rect 2455 20244 2467 20247
rect 2590 20244 2596 20256
rect 2455 20216 2596 20244
rect 2455 20213 2467 20216
rect 2409 20207 2467 20213
rect 2590 20204 2596 20216
rect 2648 20204 2654 20256
rect 4249 20247 4307 20253
rect 4249 20213 4261 20247
rect 4295 20244 4307 20247
rect 4522 20244 4528 20256
rect 4295 20216 4528 20244
rect 4295 20213 4307 20216
rect 4249 20207 4307 20213
rect 4522 20204 4528 20216
rect 4580 20204 4586 20256
rect 4908 20244 4936 20272
rect 6104 20244 6132 20284
rect 7653 20281 7665 20284
rect 7699 20312 7711 20315
rect 7742 20312 7748 20324
rect 7699 20284 7748 20312
rect 7699 20281 7711 20284
rect 7653 20275 7711 20281
rect 7742 20272 7748 20284
rect 7800 20312 7806 20324
rect 8158 20315 8216 20321
rect 8158 20312 8170 20315
rect 7800 20284 8170 20312
rect 7800 20272 7806 20284
rect 8158 20281 8170 20284
rect 8204 20281 8216 20315
rect 8158 20275 8216 20281
rect 9140 20256 9168 20352
rect 10873 20349 10885 20383
rect 10919 20380 10931 20383
rect 11184 20383 11242 20389
rect 11184 20380 11196 20383
rect 10919 20352 11196 20380
rect 10919 20349 10931 20352
rect 10873 20343 10931 20349
rect 11184 20349 11196 20352
rect 11230 20380 11242 20383
rect 11609 20383 11667 20389
rect 11609 20380 11621 20383
rect 11230 20352 11621 20380
rect 11230 20349 11242 20352
rect 11184 20343 11242 20349
rect 11609 20349 11621 20352
rect 11655 20349 11667 20383
rect 11609 20343 11667 20349
rect 14093 20383 14151 20389
rect 14093 20349 14105 20383
rect 14139 20349 14151 20383
rect 14093 20343 14151 20349
rect 14366 20340 14372 20392
rect 14424 20380 14430 20392
rect 14461 20383 14519 20389
rect 14461 20380 14473 20383
rect 14424 20352 14473 20380
rect 14424 20340 14430 20352
rect 14461 20349 14473 20352
rect 14507 20349 14519 20383
rect 14461 20343 14519 20349
rect 9490 20272 9496 20324
rect 9548 20312 9554 20324
rect 9677 20315 9735 20321
rect 9677 20312 9689 20315
rect 9548 20284 9689 20312
rect 9548 20272 9554 20284
rect 9677 20281 9689 20284
rect 9723 20281 9735 20315
rect 9677 20275 9735 20281
rect 9769 20315 9827 20321
rect 9769 20281 9781 20315
rect 9815 20281 9827 20315
rect 9769 20275 9827 20281
rect 12253 20315 12311 20321
rect 12253 20281 12265 20315
rect 12299 20312 12311 20315
rect 12618 20312 12624 20324
rect 12299 20284 12624 20312
rect 12299 20281 12311 20284
rect 12253 20275 12311 20281
rect 4908 20216 6132 20244
rect 6178 20204 6184 20256
rect 6236 20244 6242 20256
rect 6963 20247 7021 20253
rect 6963 20244 6975 20247
rect 6236 20216 6975 20244
rect 6236 20204 6242 20216
rect 6963 20213 6975 20216
rect 7009 20213 7021 20247
rect 6963 20207 7021 20213
rect 7926 20204 7932 20256
rect 7984 20244 7990 20256
rect 8757 20247 8815 20253
rect 8757 20244 8769 20247
rect 7984 20216 8769 20244
rect 7984 20204 7990 20216
rect 8757 20213 8769 20216
rect 8803 20213 8815 20247
rect 9122 20244 9128 20256
rect 9083 20216 9128 20244
rect 8757 20207 8815 20213
rect 9122 20204 9128 20216
rect 9180 20204 9186 20256
rect 9306 20204 9312 20256
rect 9364 20244 9370 20256
rect 9401 20247 9459 20253
rect 9401 20244 9413 20247
rect 9364 20216 9413 20244
rect 9364 20204 9370 20216
rect 9401 20213 9413 20216
rect 9447 20213 9459 20247
rect 9401 20207 9459 20213
rect 9582 20204 9588 20256
rect 9640 20244 9646 20256
rect 9784 20244 9812 20275
rect 12618 20272 12624 20284
rect 12676 20272 12682 20324
rect 15933 20315 15991 20321
rect 15933 20281 15945 20315
rect 15979 20281 15991 20315
rect 18370 20315 18428 20321
rect 18370 20312 18382 20315
rect 15933 20275 15991 20281
rect 17788 20284 18382 20312
rect 10597 20247 10655 20253
rect 10597 20244 10609 20247
rect 9640 20216 10609 20244
rect 9640 20204 9646 20216
rect 10597 20213 10609 20216
rect 10643 20213 10655 20247
rect 13538 20244 13544 20256
rect 13499 20216 13544 20244
rect 10597 20207 10655 20213
rect 13538 20204 13544 20216
rect 13596 20204 13602 20256
rect 14090 20244 14096 20256
rect 14051 20216 14096 20244
rect 14090 20204 14096 20216
rect 14148 20204 14154 20256
rect 15378 20244 15384 20256
rect 15339 20216 15384 20244
rect 15378 20204 15384 20216
rect 15436 20204 15442 20256
rect 15746 20204 15752 20256
rect 15804 20244 15810 20256
rect 15948 20244 15976 20275
rect 17788 20256 17816 20284
rect 18370 20281 18382 20284
rect 18416 20312 18428 20315
rect 19058 20312 19064 20324
rect 18416 20284 19064 20312
rect 18416 20281 18428 20284
rect 18370 20275 18428 20281
rect 19058 20272 19064 20284
rect 19116 20312 19122 20324
rect 19245 20315 19303 20321
rect 19245 20312 19257 20315
rect 19116 20284 19257 20312
rect 19116 20272 19122 20284
rect 19245 20281 19257 20284
rect 19291 20281 19303 20315
rect 19245 20275 19303 20281
rect 19978 20272 19984 20324
rect 20036 20312 20042 20324
rect 20073 20315 20131 20321
rect 20073 20312 20085 20315
rect 20036 20284 20085 20312
rect 20036 20272 20042 20284
rect 20073 20281 20085 20284
rect 20119 20281 20131 20315
rect 21542 20312 21548 20324
rect 21503 20284 21548 20312
rect 20073 20275 20131 20281
rect 21542 20272 21548 20284
rect 21600 20272 21606 20324
rect 21634 20272 21640 20324
rect 21692 20312 21698 20324
rect 21692 20284 21737 20312
rect 21692 20272 21698 20284
rect 17770 20244 17776 20256
rect 15804 20216 15976 20244
rect 17731 20216 17776 20244
rect 15804 20204 15810 20216
rect 17770 20204 17776 20216
rect 17828 20204 17834 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1535 20043 1593 20049
rect 1535 20009 1547 20043
rect 1581 20040 1593 20043
rect 3602 20040 3608 20052
rect 1581 20012 3608 20040
rect 1581 20009 1593 20012
rect 1535 20003 1593 20009
rect 3602 20000 3608 20012
rect 3660 20000 3666 20052
rect 4614 20000 4620 20052
rect 4672 20040 4678 20052
rect 5350 20040 5356 20052
rect 4672 20012 5356 20040
rect 4672 20000 4678 20012
rect 5350 20000 5356 20012
rect 5408 20040 5414 20052
rect 5629 20043 5687 20049
rect 5629 20040 5641 20043
rect 5408 20012 5641 20040
rect 5408 20000 5414 20012
rect 5629 20009 5641 20012
rect 5675 20040 5687 20043
rect 5905 20043 5963 20049
rect 5905 20040 5917 20043
rect 5675 20012 5917 20040
rect 5675 20009 5687 20012
rect 5629 20003 5687 20009
rect 5905 20009 5917 20012
rect 5951 20009 5963 20043
rect 7466 20040 7472 20052
rect 7427 20012 7472 20040
rect 5905 20003 5963 20009
rect 7466 20000 7472 20012
rect 7524 20000 7530 20052
rect 7742 20000 7748 20052
rect 7800 20040 7806 20052
rect 7837 20043 7895 20049
rect 7837 20040 7849 20043
rect 7800 20012 7849 20040
rect 7800 20000 7806 20012
rect 7837 20009 7849 20012
rect 7883 20009 7895 20043
rect 7837 20003 7895 20009
rect 7926 20000 7932 20052
rect 7984 20040 7990 20052
rect 7984 20012 8248 20040
rect 7984 20000 7990 20012
rect 2498 19972 2504 19984
rect 2459 19944 2504 19972
rect 2498 19932 2504 19944
rect 2556 19932 2562 19984
rect 2593 19975 2651 19981
rect 2593 19941 2605 19975
rect 2639 19972 2651 19975
rect 3234 19972 3240 19984
rect 2639 19944 3240 19972
rect 2639 19941 2651 19944
rect 2593 19935 2651 19941
rect 3234 19932 3240 19944
rect 3292 19932 3298 19984
rect 4890 19932 4896 19984
rect 4948 19972 4954 19984
rect 5030 19975 5088 19981
rect 5030 19972 5042 19975
rect 4948 19944 5042 19972
rect 4948 19932 4954 19944
rect 5030 19941 5042 19944
rect 5076 19941 5088 19975
rect 5030 19935 5088 19941
rect 6454 19932 6460 19984
rect 6512 19972 6518 19984
rect 6730 19972 6736 19984
rect 6512 19944 6736 19972
rect 6512 19932 6518 19944
rect 6730 19932 6736 19944
rect 6788 19932 6794 19984
rect 7558 19932 7564 19984
rect 7616 19972 7622 19984
rect 8220 19981 8248 20012
rect 9122 20000 9128 20052
rect 9180 20040 9186 20052
rect 9769 20043 9827 20049
rect 9769 20040 9781 20043
rect 9180 20012 9781 20040
rect 9180 20000 9186 20012
rect 9769 20009 9781 20012
rect 9815 20009 9827 20043
rect 11054 20040 11060 20052
rect 11015 20012 11060 20040
rect 9769 20003 9827 20009
rect 11054 20000 11060 20012
rect 11112 20000 11118 20052
rect 12802 20040 12808 20052
rect 12763 20012 12808 20040
rect 12802 20000 12808 20012
rect 12860 20040 12866 20052
rect 14090 20040 14096 20052
rect 12860 20012 14096 20040
rect 12860 20000 12866 20012
rect 14090 20000 14096 20012
rect 14148 20000 14154 20052
rect 14826 20000 14832 20052
rect 14884 20040 14890 20052
rect 15013 20043 15071 20049
rect 15013 20040 15025 20043
rect 14884 20012 15025 20040
rect 14884 20000 14890 20012
rect 15013 20009 15025 20012
rect 15059 20009 15071 20043
rect 15013 20003 15071 20009
rect 15378 20000 15384 20052
rect 15436 20040 15442 20052
rect 17770 20040 17776 20052
rect 15436 20012 17776 20040
rect 15436 20000 15442 20012
rect 8113 19975 8171 19981
rect 8113 19972 8125 19975
rect 7616 19944 8125 19972
rect 7616 19932 7622 19944
rect 8113 19941 8125 19944
rect 8159 19941 8171 19975
rect 8113 19935 8171 19941
rect 8205 19975 8263 19981
rect 8205 19941 8217 19975
rect 8251 19941 8263 19975
rect 8754 19972 8760 19984
rect 8715 19944 8760 19972
rect 8205 19935 8263 19941
rect 8754 19932 8760 19944
rect 8812 19932 8818 19984
rect 9490 19972 9496 19984
rect 9451 19944 9496 19972
rect 9490 19932 9496 19944
rect 9548 19932 9554 19984
rect 11971 19975 12029 19981
rect 11971 19941 11983 19975
rect 12017 19972 12029 19975
rect 13538 19972 13544 19984
rect 12017 19944 13544 19972
rect 12017 19941 12029 19944
rect 11971 19935 12029 19941
rect 13538 19932 13544 19944
rect 13596 19932 13602 19984
rect 15666 19981 15694 20012
rect 17770 20000 17776 20012
rect 17828 20000 17834 20052
rect 17862 20000 17868 20052
rect 17920 20040 17926 20052
rect 18601 20043 18659 20049
rect 18601 20040 18613 20043
rect 17920 20012 18613 20040
rect 17920 20000 17926 20012
rect 18601 20009 18613 20012
rect 18647 20009 18659 20043
rect 19242 20040 19248 20052
rect 19203 20012 19248 20040
rect 18601 20003 18659 20009
rect 19242 20000 19248 20012
rect 19300 20000 19306 20052
rect 20254 20040 20260 20052
rect 20215 20012 20260 20040
rect 20254 20000 20260 20012
rect 20312 20000 20318 20052
rect 21039 20043 21097 20049
rect 21039 20009 21051 20043
rect 21085 20040 21097 20043
rect 21542 20040 21548 20052
rect 21085 20012 21548 20040
rect 21085 20009 21097 20012
rect 21039 20003 21097 20009
rect 21542 20000 21548 20012
rect 21600 20000 21606 20052
rect 15651 19975 15709 19981
rect 15651 19941 15663 19975
rect 15697 19941 15709 19975
rect 18325 19975 18383 19981
rect 15651 19935 15709 19941
rect 17420 19944 18184 19972
rect 1464 19907 1522 19913
rect 1464 19873 1476 19907
rect 1510 19904 1522 19907
rect 1762 19904 1768 19916
rect 1510 19876 1768 19904
rect 1510 19873 1522 19876
rect 1464 19867 1522 19873
rect 1762 19864 1768 19876
rect 1820 19864 1826 19916
rect 6270 19904 6276 19916
rect 4356 19876 6276 19904
rect 3145 19839 3203 19845
rect 3145 19805 3157 19839
rect 3191 19836 3203 19839
rect 3326 19836 3332 19848
rect 3191 19808 3332 19836
rect 3191 19805 3203 19808
rect 3145 19799 3203 19805
rect 3326 19796 3332 19808
rect 3384 19796 3390 19848
rect 3510 19796 3516 19848
rect 3568 19836 3574 19848
rect 3786 19836 3792 19848
rect 3568 19808 3792 19836
rect 3568 19796 3574 19808
rect 3786 19796 3792 19808
rect 3844 19796 3850 19848
rect 2958 19728 2964 19780
rect 3016 19768 3022 19780
rect 4356 19768 4384 19876
rect 6270 19864 6276 19876
rect 6328 19904 6334 19916
rect 6549 19907 6607 19913
rect 6549 19904 6561 19907
rect 6328 19876 6561 19904
rect 6328 19864 6334 19876
rect 6549 19873 6561 19876
rect 6595 19873 6607 19907
rect 6549 19867 6607 19873
rect 9582 19864 9588 19916
rect 9640 19904 9646 19916
rect 9677 19907 9735 19913
rect 9677 19904 9689 19907
rect 9640 19876 9689 19904
rect 9640 19864 9646 19876
rect 9677 19873 9689 19876
rect 9723 19873 9735 19907
rect 10226 19904 10232 19916
rect 10139 19876 10232 19904
rect 9677 19867 9735 19873
rect 4709 19839 4767 19845
rect 4709 19836 4721 19839
rect 3016 19740 4384 19768
rect 4540 19808 4721 19836
rect 3016 19728 3022 19740
rect 2130 19700 2136 19712
rect 2091 19672 2136 19700
rect 2130 19660 2136 19672
rect 2188 19660 2194 19712
rect 3418 19700 3424 19712
rect 3379 19672 3424 19700
rect 3418 19660 3424 19672
rect 3476 19660 3482 19712
rect 3602 19660 3608 19712
rect 3660 19700 3666 19712
rect 3789 19703 3847 19709
rect 3789 19700 3801 19703
rect 3660 19672 3801 19700
rect 3660 19660 3666 19672
rect 3789 19669 3801 19672
rect 3835 19669 3847 19703
rect 3789 19663 3847 19669
rect 4062 19660 4068 19712
rect 4120 19700 4126 19712
rect 4540 19709 4568 19808
rect 4709 19805 4721 19808
rect 4755 19805 4767 19839
rect 6454 19836 6460 19848
rect 6415 19808 6460 19836
rect 4709 19799 4767 19805
rect 6454 19796 6460 19808
rect 6512 19796 6518 19848
rect 9692 19768 9720 19867
rect 10226 19864 10232 19876
rect 10284 19904 10290 19916
rect 10778 19904 10784 19916
rect 10284 19876 10784 19904
rect 10284 19864 10290 19876
rect 10778 19864 10784 19876
rect 10836 19904 10842 19916
rect 12529 19907 12587 19913
rect 10836 19876 11744 19904
rect 10836 19864 10842 19876
rect 11606 19836 11612 19848
rect 11567 19808 11612 19836
rect 11606 19796 11612 19808
rect 11664 19796 11670 19848
rect 11716 19836 11744 19876
rect 12529 19873 12541 19907
rect 12575 19904 12587 19907
rect 13446 19904 13452 19916
rect 12575 19876 13452 19904
rect 12575 19873 12587 19876
rect 12529 19867 12587 19873
rect 13446 19864 13452 19876
rect 13504 19864 13510 19916
rect 13630 19904 13636 19916
rect 13591 19876 13636 19904
rect 13630 19864 13636 19876
rect 13688 19864 13694 19916
rect 14182 19904 14188 19916
rect 14143 19876 14188 19904
rect 14182 19864 14188 19876
rect 14240 19864 14246 19916
rect 17420 19904 17448 19944
rect 17586 19904 17592 19916
rect 15672 19876 17448 19904
rect 17547 19876 17592 19904
rect 13354 19836 13360 19848
rect 11716 19808 13360 19836
rect 13354 19796 13360 19808
rect 13412 19796 13418 19848
rect 14369 19839 14427 19845
rect 14369 19805 14381 19839
rect 14415 19836 14427 19839
rect 14826 19836 14832 19848
rect 14415 19808 14832 19836
rect 14415 19805 14427 19808
rect 14369 19799 14427 19805
rect 14826 19796 14832 19808
rect 14884 19836 14890 19848
rect 15289 19839 15347 19845
rect 15289 19836 15301 19839
rect 14884 19808 15301 19836
rect 14884 19796 14890 19808
rect 15289 19805 15301 19808
rect 15335 19805 15347 19839
rect 15289 19799 15347 19805
rect 15672 19768 15700 19876
rect 17586 19864 17592 19876
rect 17644 19864 17650 19916
rect 18049 19907 18107 19913
rect 18049 19873 18061 19907
rect 18095 19873 18107 19907
rect 18156 19904 18184 19944
rect 18325 19941 18337 19975
rect 18371 19972 18383 19975
rect 18690 19972 18696 19984
rect 18371 19944 18696 19972
rect 18371 19941 18383 19944
rect 18325 19935 18383 19941
rect 18690 19932 18696 19944
rect 18748 19972 18754 19984
rect 18969 19975 19027 19981
rect 18969 19972 18981 19975
rect 18748 19944 18981 19972
rect 18748 19932 18754 19944
rect 18969 19941 18981 19944
rect 19015 19941 19027 19975
rect 18969 19935 19027 19941
rect 19150 19904 19156 19916
rect 18156 19876 19156 19904
rect 18049 19867 18107 19873
rect 17126 19796 17132 19848
rect 17184 19836 17190 19848
rect 17862 19836 17868 19848
rect 17184 19808 17868 19836
rect 17184 19796 17190 19808
rect 17862 19796 17868 19808
rect 17920 19836 17926 19848
rect 18064 19836 18092 19867
rect 19150 19864 19156 19876
rect 19208 19864 19214 19916
rect 19613 19907 19671 19913
rect 19613 19873 19625 19907
rect 19659 19873 19671 19907
rect 20806 19904 20812 19916
rect 20767 19876 20812 19904
rect 19613 19867 19671 19873
rect 19628 19836 19656 19867
rect 20806 19864 20812 19876
rect 20864 19864 20870 19916
rect 24648 19907 24706 19913
rect 24648 19873 24660 19907
rect 24694 19904 24706 19907
rect 25498 19904 25504 19916
rect 24694 19876 25504 19904
rect 24694 19873 24706 19876
rect 24648 19867 24706 19873
rect 25498 19864 25504 19876
rect 25556 19864 25562 19916
rect 17920 19808 19656 19836
rect 17920 19796 17926 19808
rect 9692 19740 15700 19768
rect 15746 19728 15752 19780
rect 15804 19768 15810 19780
rect 16485 19771 16543 19777
rect 16485 19768 16497 19771
rect 15804 19740 16497 19768
rect 15804 19728 15810 19740
rect 16485 19737 16497 19740
rect 16531 19737 16543 19771
rect 16485 19731 16543 19737
rect 4525 19703 4583 19709
rect 4525 19700 4537 19703
rect 4120 19672 4537 19700
rect 4120 19660 4126 19672
rect 4525 19669 4537 19672
rect 4571 19669 4583 19703
rect 14734 19700 14740 19712
rect 14695 19672 14740 19700
rect 4525 19663 4583 19669
rect 14734 19660 14740 19672
rect 14792 19660 14798 19712
rect 16206 19700 16212 19712
rect 16167 19672 16212 19700
rect 16206 19660 16212 19672
rect 16264 19660 16270 19712
rect 18598 19660 18604 19712
rect 18656 19700 18662 19712
rect 24719 19703 24777 19709
rect 24719 19700 24731 19703
rect 18656 19672 24731 19700
rect 18656 19660 18662 19672
rect 24719 19669 24731 19672
rect 24765 19669 24777 19703
rect 24719 19663 24777 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 2958 19496 2964 19508
rect 2919 19468 2964 19496
rect 2958 19456 2964 19468
rect 3016 19456 3022 19508
rect 3234 19496 3240 19508
rect 3195 19468 3240 19496
rect 3234 19456 3240 19468
rect 3292 19456 3298 19508
rect 3697 19499 3755 19505
rect 3697 19465 3709 19499
rect 3743 19496 3755 19499
rect 3970 19496 3976 19508
rect 3743 19468 3976 19496
rect 3743 19465 3755 19468
rect 3697 19459 3755 19465
rect 3970 19456 3976 19468
rect 4028 19456 4034 19508
rect 6270 19496 6276 19508
rect 6231 19468 6276 19496
rect 6270 19456 6276 19468
rect 6328 19456 6334 19508
rect 9401 19499 9459 19505
rect 9401 19465 9413 19499
rect 9447 19496 9459 19499
rect 10226 19496 10232 19508
rect 9447 19468 10232 19496
rect 9447 19465 9459 19468
rect 9401 19459 9459 19465
rect 10226 19456 10232 19468
rect 10284 19456 10290 19508
rect 10686 19456 10692 19508
rect 10744 19496 10750 19508
rect 13630 19496 13636 19508
rect 10744 19468 13636 19496
rect 10744 19456 10750 19468
rect 13630 19456 13636 19468
rect 13688 19456 13694 19508
rect 15378 19496 15384 19508
rect 15339 19468 15384 19496
rect 15378 19456 15384 19468
rect 15436 19456 15442 19508
rect 16206 19456 16212 19508
rect 16264 19496 16270 19508
rect 16577 19499 16635 19505
rect 16577 19496 16589 19499
rect 16264 19468 16589 19496
rect 16264 19456 16270 19468
rect 16577 19465 16589 19468
rect 16623 19465 16635 19499
rect 16577 19459 16635 19465
rect 17126 19456 17132 19508
rect 17184 19496 17190 19508
rect 17405 19499 17463 19505
rect 17405 19496 17417 19499
rect 17184 19468 17417 19496
rect 17184 19456 17190 19468
rect 17405 19465 17417 19468
rect 17451 19465 17463 19499
rect 17405 19459 17463 19465
rect 18874 19456 18880 19508
rect 18932 19496 18938 19508
rect 19150 19496 19156 19508
rect 18932 19468 19156 19496
rect 18932 19456 18938 19468
rect 19150 19456 19156 19468
rect 19208 19496 19214 19508
rect 19613 19499 19671 19505
rect 19613 19496 19625 19499
rect 19208 19468 19625 19496
rect 19208 19456 19214 19468
rect 19613 19465 19625 19468
rect 19659 19465 19671 19499
rect 25130 19496 25136 19508
rect 25091 19468 25136 19496
rect 19613 19459 19671 19465
rect 25130 19456 25136 19468
rect 25188 19456 25194 19508
rect 25498 19496 25504 19508
rect 25459 19468 25504 19496
rect 25498 19456 25504 19468
rect 25556 19456 25562 19508
rect 3252 19428 3280 19456
rect 6454 19428 6460 19440
rect 3252 19400 6460 19428
rect 6454 19388 6460 19400
rect 6512 19388 6518 19440
rect 12342 19388 12348 19440
rect 12400 19428 12406 19440
rect 13081 19431 13139 19437
rect 13081 19428 13093 19431
rect 12400 19400 13093 19428
rect 12400 19388 12406 19400
rect 13081 19397 13093 19400
rect 13127 19397 13139 19431
rect 13081 19391 13139 19397
rect 13906 19388 13912 19440
rect 13964 19428 13970 19440
rect 17037 19431 17095 19437
rect 17037 19428 17049 19431
rect 13964 19400 17049 19428
rect 13964 19388 13970 19400
rect 17037 19397 17049 19400
rect 17083 19428 17095 19431
rect 17586 19428 17592 19440
rect 17083 19400 17592 19428
rect 17083 19397 17095 19400
rect 17037 19391 17095 19397
rect 17586 19388 17592 19400
rect 17644 19388 17650 19440
rect 18506 19388 18512 19440
rect 18564 19428 18570 19440
rect 18969 19431 19027 19437
rect 18969 19428 18981 19431
rect 18564 19400 18981 19428
rect 18564 19388 18570 19400
rect 18969 19397 18981 19400
rect 19015 19428 19027 19431
rect 21358 19428 21364 19440
rect 19015 19400 21364 19428
rect 19015 19397 19027 19400
rect 18969 19391 19027 19397
rect 21358 19388 21364 19400
rect 21416 19388 21422 19440
rect 1673 19363 1731 19369
rect 1673 19329 1685 19363
rect 1719 19360 1731 19363
rect 1762 19360 1768 19372
rect 1719 19332 1768 19360
rect 1719 19329 1731 19332
rect 1673 19323 1731 19329
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 2041 19363 2099 19369
rect 2041 19329 2053 19363
rect 2087 19360 2099 19363
rect 2682 19360 2688 19372
rect 2087 19332 2688 19360
rect 2087 19329 2099 19332
rect 2041 19323 2099 19329
rect 2682 19320 2688 19332
rect 2740 19360 2746 19372
rect 3602 19360 3608 19372
rect 2740 19332 3608 19360
rect 2740 19320 2746 19332
rect 3602 19320 3608 19332
rect 3660 19320 3666 19372
rect 3878 19320 3884 19372
rect 3936 19360 3942 19372
rect 4341 19363 4399 19369
rect 3936 19332 4154 19360
rect 3936 19320 3942 19332
rect 3694 19252 3700 19304
rect 3752 19252 3758 19304
rect 3970 19292 3976 19304
rect 3931 19264 3976 19292
rect 3970 19252 3976 19264
rect 4028 19252 4034 19304
rect 4126 19292 4154 19332
rect 4341 19329 4353 19363
rect 4387 19360 4399 19363
rect 4614 19360 4620 19372
rect 4387 19332 4620 19360
rect 4387 19329 4399 19332
rect 4341 19323 4399 19329
rect 4614 19320 4620 19332
rect 4672 19360 4678 19372
rect 5258 19360 5264 19372
rect 4672 19332 5264 19360
rect 4672 19320 4678 19332
rect 5258 19320 5264 19332
rect 5316 19320 5322 19372
rect 5534 19360 5540 19372
rect 5495 19332 5540 19360
rect 5534 19320 5540 19332
rect 5592 19320 5598 19372
rect 8389 19363 8447 19369
rect 8389 19329 8401 19363
rect 8435 19360 8447 19363
rect 9214 19360 9220 19372
rect 8435 19332 9220 19360
rect 8435 19329 8447 19332
rect 8389 19323 8447 19329
rect 9214 19320 9220 19332
rect 9272 19320 9278 19372
rect 9953 19363 10011 19369
rect 9953 19329 9965 19363
rect 9999 19360 10011 19363
rect 10778 19360 10784 19372
rect 9999 19332 10784 19360
rect 9999 19329 10011 19332
rect 9953 19323 10011 19329
rect 10778 19320 10784 19332
rect 10836 19320 10842 19372
rect 11333 19363 11391 19369
rect 11333 19329 11345 19363
rect 11379 19360 11391 19363
rect 11606 19360 11612 19372
rect 11379 19332 11612 19360
rect 11379 19329 11391 19332
rect 11333 19323 11391 19329
rect 11606 19320 11612 19332
rect 11664 19360 11670 19372
rect 11664 19332 13308 19360
rect 11664 19320 11670 19332
rect 4709 19295 4767 19301
rect 4709 19292 4721 19295
rect 4126 19264 4721 19292
rect 4709 19261 4721 19264
rect 4755 19261 4767 19295
rect 4709 19255 4767 19261
rect 4890 19252 4896 19304
rect 4948 19292 4954 19304
rect 4985 19295 5043 19301
rect 4985 19292 4997 19295
rect 4948 19264 4997 19292
rect 4948 19252 4954 19264
rect 4985 19261 4997 19264
rect 5031 19261 5043 19295
rect 4985 19255 5043 19261
rect 6457 19295 6515 19301
rect 6457 19261 6469 19295
rect 6503 19292 6515 19295
rect 7009 19295 7067 19301
rect 7009 19292 7021 19295
rect 6503 19264 7021 19292
rect 6503 19261 6515 19264
rect 6457 19255 6515 19261
rect 7009 19261 7021 19264
rect 7055 19261 7067 19295
rect 7374 19292 7380 19304
rect 7335 19264 7380 19292
rect 7009 19255 7067 19261
rect 7374 19252 7380 19264
rect 7432 19252 7438 19304
rect 2130 19184 2136 19236
rect 2188 19224 2194 19236
rect 2403 19227 2461 19233
rect 2403 19224 2415 19227
rect 2188 19196 2415 19224
rect 2188 19184 2194 19196
rect 2403 19193 2415 19196
rect 2449 19224 2461 19227
rect 2958 19224 2964 19236
rect 2449 19196 2964 19224
rect 2449 19193 2461 19196
rect 2403 19187 2461 19193
rect 2958 19184 2964 19196
rect 3016 19224 3022 19236
rect 3712 19224 3740 19252
rect 3016 19196 3740 19224
rect 3789 19227 3847 19233
rect 3016 19184 3022 19196
rect 3789 19193 3801 19227
rect 3835 19224 3847 19227
rect 3878 19224 3884 19236
rect 3835 19196 3884 19224
rect 3835 19193 3847 19196
rect 3789 19187 3847 19193
rect 3878 19184 3884 19196
rect 3936 19184 3942 19236
rect 5261 19227 5319 19233
rect 5261 19193 5273 19227
rect 5307 19193 5319 19227
rect 5261 19187 5319 19193
rect 5276 19156 5304 19187
rect 5350 19184 5356 19236
rect 5408 19224 5414 19236
rect 5408 19196 5453 19224
rect 5408 19184 5414 19196
rect 5534 19184 5540 19236
rect 5592 19224 5598 19236
rect 6825 19227 6883 19233
rect 6825 19224 6837 19227
rect 5592 19196 6837 19224
rect 5592 19184 5598 19196
rect 6825 19193 6837 19196
rect 6871 19224 6883 19227
rect 7653 19227 7711 19233
rect 7653 19224 7665 19227
rect 6871 19196 7665 19224
rect 6871 19193 6883 19196
rect 6825 19187 6883 19193
rect 7653 19193 7665 19196
rect 7699 19193 7711 19227
rect 7653 19187 7711 19193
rect 8481 19227 8539 19233
rect 8481 19193 8493 19227
rect 8527 19193 8539 19227
rect 9030 19224 9036 19236
rect 8991 19196 9036 19224
rect 8481 19187 8539 19193
rect 6086 19156 6092 19168
rect 5276 19128 6092 19156
rect 6086 19116 6092 19128
rect 6144 19116 6150 19168
rect 6270 19116 6276 19168
rect 6328 19156 6334 19168
rect 6457 19159 6515 19165
rect 6457 19156 6469 19159
rect 6328 19128 6469 19156
rect 6328 19116 6334 19128
rect 6457 19125 6469 19128
rect 6503 19156 6515 19159
rect 6549 19159 6607 19165
rect 6549 19156 6561 19159
rect 6503 19128 6561 19156
rect 6503 19125 6515 19128
rect 6457 19119 6515 19125
rect 6549 19125 6561 19128
rect 6595 19125 6607 19159
rect 8202 19156 8208 19168
rect 8115 19128 8208 19156
rect 6549 19119 6607 19125
rect 8202 19116 8208 19128
rect 8260 19156 8266 19168
rect 8496 19156 8524 19187
rect 9030 19184 9036 19196
rect 9088 19184 9094 19236
rect 10045 19227 10103 19233
rect 10045 19193 10057 19227
rect 10091 19193 10103 19227
rect 10045 19187 10103 19193
rect 10597 19227 10655 19233
rect 10597 19193 10609 19227
rect 10643 19224 10655 19227
rect 11422 19224 11428 19236
rect 10643 19196 11428 19224
rect 10643 19193 10655 19196
rect 10597 19187 10655 19193
rect 8260 19128 8524 19156
rect 8260 19116 8266 19128
rect 8570 19116 8576 19168
rect 8628 19156 8634 19168
rect 9582 19156 9588 19168
rect 8628 19128 9588 19156
rect 8628 19116 8634 19128
rect 9582 19116 9588 19128
rect 9640 19156 9646 19168
rect 9677 19159 9735 19165
rect 9677 19156 9689 19159
rect 9640 19128 9689 19156
rect 9640 19116 9646 19128
rect 9677 19125 9689 19128
rect 9723 19125 9735 19159
rect 9677 19119 9735 19125
rect 9858 19116 9864 19168
rect 9916 19156 9922 19168
rect 10060 19156 10088 19187
rect 11422 19184 11428 19196
rect 11480 19184 11486 19236
rect 12526 19224 12532 19236
rect 12487 19196 12532 19224
rect 12526 19184 12532 19196
rect 12584 19184 12590 19236
rect 12618 19184 12624 19236
rect 12676 19224 12682 19236
rect 13280 19224 13308 19332
rect 13354 19320 13360 19372
rect 13412 19360 13418 19372
rect 13541 19363 13599 19369
rect 13541 19360 13553 19363
rect 13412 19332 13553 19360
rect 13412 19320 13418 19332
rect 13541 19329 13553 19332
rect 13587 19360 13599 19363
rect 14366 19360 14372 19372
rect 13587 19332 14372 19360
rect 13587 19329 13599 19332
rect 13541 19323 13599 19329
rect 14366 19320 14372 19332
rect 14424 19320 14430 19372
rect 14734 19320 14740 19372
rect 14792 19360 14798 19372
rect 15657 19363 15715 19369
rect 15657 19360 15669 19363
rect 14792 19332 15669 19360
rect 14792 19320 14798 19332
rect 15657 19329 15669 19332
rect 15703 19360 15715 19363
rect 16114 19360 16120 19372
rect 15703 19332 16120 19360
rect 15703 19329 15715 19332
rect 15657 19323 15715 19329
rect 16114 19320 16120 19332
rect 16172 19320 16178 19372
rect 19889 19363 19947 19369
rect 19889 19329 19901 19363
rect 19935 19360 19947 19363
rect 20254 19360 20260 19372
rect 19935 19332 20260 19360
rect 19935 19329 19947 19332
rect 19889 19323 19947 19329
rect 20254 19320 20260 19332
rect 20312 19320 20318 19372
rect 20530 19360 20536 19372
rect 20491 19332 20536 19360
rect 20530 19320 20536 19332
rect 20588 19320 20594 19372
rect 21266 19320 21272 19372
rect 21324 19360 21330 19372
rect 21499 19363 21557 19369
rect 21499 19360 21511 19363
rect 21324 19332 21511 19360
rect 21324 19320 21330 19332
rect 21499 19329 21511 19332
rect 21545 19329 21557 19363
rect 21499 19323 21557 19329
rect 13722 19252 13728 19304
rect 13780 19292 13786 19304
rect 14001 19295 14059 19301
rect 14001 19292 14013 19295
rect 13780 19264 14013 19292
rect 13780 19252 13786 19264
rect 14001 19261 14013 19264
rect 14047 19261 14059 19295
rect 14458 19292 14464 19304
rect 14419 19264 14464 19292
rect 14001 19255 14059 19261
rect 14458 19252 14464 19264
rect 14516 19252 14522 19304
rect 17770 19292 17776 19304
rect 17731 19264 17776 19292
rect 17770 19252 17776 19264
rect 17828 19252 17834 19304
rect 18046 19292 18052 19304
rect 18007 19264 18052 19292
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 21412 19295 21470 19301
rect 21412 19261 21424 19295
rect 21458 19292 21470 19295
rect 21913 19295 21971 19301
rect 21913 19292 21925 19295
rect 21458 19264 21925 19292
rect 21458 19261 21470 19264
rect 21412 19255 21470 19261
rect 21913 19261 21925 19264
rect 21959 19292 21971 19295
rect 22094 19292 22100 19304
rect 21959 19264 22100 19292
rect 21959 19261 21971 19264
rect 21913 19255 21971 19261
rect 22094 19252 22100 19264
rect 22152 19252 22158 19304
rect 24648 19295 24706 19301
rect 24648 19261 24660 19295
rect 24694 19292 24706 19295
rect 25130 19292 25136 19304
rect 24694 19264 25136 19292
rect 24694 19261 24706 19264
rect 24648 19255 24706 19261
rect 25130 19252 25136 19264
rect 25188 19252 25194 19304
rect 15749 19227 15807 19233
rect 12676 19196 12721 19224
rect 13280 19196 14044 19224
rect 12676 19184 12682 19196
rect 10873 19159 10931 19165
rect 10873 19156 10885 19159
rect 9916 19128 10885 19156
rect 9916 19116 9922 19128
rect 10873 19125 10885 19128
rect 10919 19125 10931 19159
rect 11698 19156 11704 19168
rect 11659 19128 11704 19156
rect 10873 19119 10931 19125
rect 11698 19116 11704 19128
rect 11756 19116 11762 19168
rect 12253 19159 12311 19165
rect 12253 19125 12265 19159
rect 12299 19156 12311 19159
rect 12636 19156 12664 19184
rect 12299 19128 12664 19156
rect 12299 19125 12311 19128
rect 12253 19119 12311 19125
rect 13722 19116 13728 19168
rect 13780 19156 13786 19168
rect 13817 19159 13875 19165
rect 13817 19156 13829 19159
rect 13780 19128 13829 19156
rect 13780 19116 13786 19128
rect 13817 19125 13829 19128
rect 13863 19125 13875 19159
rect 14016 19156 14044 19196
rect 15749 19193 15761 19227
rect 15795 19224 15807 19227
rect 16114 19224 16120 19236
rect 15795 19196 16120 19224
rect 15795 19193 15807 19196
rect 15749 19187 15807 19193
rect 16114 19184 16120 19196
rect 16172 19184 16178 19236
rect 16301 19227 16359 19233
rect 16301 19193 16313 19227
rect 16347 19224 16359 19227
rect 16758 19224 16764 19236
rect 16347 19196 16764 19224
rect 16347 19193 16359 19196
rect 16301 19187 16359 19193
rect 16758 19184 16764 19196
rect 16816 19184 16822 19236
rect 17788 19224 17816 19252
rect 18414 19233 18420 19236
rect 18370 19227 18420 19233
rect 18370 19224 18382 19227
rect 17788 19196 18382 19224
rect 18370 19193 18382 19196
rect 18416 19193 18420 19227
rect 18370 19187 18420 19193
rect 18414 19184 18420 19187
rect 18472 19184 18478 19236
rect 19978 19184 19984 19236
rect 20036 19224 20042 19236
rect 20036 19196 20081 19224
rect 20036 19184 20042 19196
rect 14093 19159 14151 19165
rect 14093 19156 14105 19159
rect 14016 19128 14105 19156
rect 13817 19119 13875 19125
rect 14093 19125 14105 19128
rect 14139 19125 14151 19159
rect 14093 19119 14151 19125
rect 17862 19116 17868 19168
rect 17920 19156 17926 19168
rect 19245 19159 19303 19165
rect 19245 19156 19257 19159
rect 17920 19128 19257 19156
rect 17920 19116 17926 19128
rect 19245 19125 19257 19128
rect 19291 19125 19303 19159
rect 19245 19119 19303 19125
rect 20070 19116 20076 19168
rect 20128 19156 20134 19168
rect 20806 19156 20812 19168
rect 20128 19128 20812 19156
rect 20128 19116 20134 19128
rect 20806 19116 20812 19128
rect 20864 19156 20870 19168
rect 20901 19159 20959 19165
rect 20901 19156 20913 19159
rect 20864 19128 20913 19156
rect 20864 19116 20870 19128
rect 20901 19125 20913 19128
rect 20947 19125 20959 19159
rect 20901 19119 20959 19125
rect 21910 19116 21916 19168
rect 21968 19156 21974 19168
rect 24719 19159 24777 19165
rect 24719 19156 24731 19159
rect 21968 19128 24731 19156
rect 21968 19116 21974 19128
rect 24719 19125 24731 19128
rect 24765 19125 24777 19159
rect 24719 19119 24777 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 2590 18952 2596 18964
rect 2551 18924 2596 18952
rect 2590 18912 2596 18924
rect 2648 18912 2654 18964
rect 4062 18912 4068 18964
rect 4120 18952 4126 18964
rect 4433 18955 4491 18961
rect 4433 18952 4445 18955
rect 4120 18924 4445 18952
rect 4120 18912 4126 18924
rect 4433 18921 4445 18924
rect 4479 18921 4491 18955
rect 6178 18952 6184 18964
rect 6139 18924 6184 18952
rect 4433 18915 4491 18921
rect 6178 18912 6184 18924
rect 6236 18912 6242 18964
rect 7193 18955 7251 18961
rect 7193 18921 7205 18955
rect 7239 18952 7251 18955
rect 7558 18952 7564 18964
rect 7239 18924 7564 18952
rect 7239 18921 7251 18924
rect 7193 18915 7251 18921
rect 7558 18912 7564 18924
rect 7616 18912 7622 18964
rect 9125 18955 9183 18961
rect 9125 18921 9137 18955
rect 9171 18952 9183 18955
rect 9214 18952 9220 18964
rect 9171 18924 9220 18952
rect 9171 18921 9183 18924
rect 9125 18915 9183 18921
rect 9214 18912 9220 18924
rect 9272 18912 9278 18964
rect 9674 18912 9680 18964
rect 9732 18952 9738 18964
rect 11698 18952 11704 18964
rect 9732 18924 9812 18952
rect 11659 18924 11704 18952
rect 9732 18912 9738 18924
rect 2035 18887 2093 18893
rect 2035 18853 2047 18887
rect 2081 18884 2093 18887
rect 2130 18884 2136 18896
rect 2081 18856 2136 18884
rect 2081 18853 2093 18856
rect 2035 18847 2093 18853
rect 2130 18844 2136 18856
rect 2188 18844 2194 18896
rect 3786 18844 3792 18896
rect 3844 18884 3850 18896
rect 8202 18884 8208 18896
rect 3844 18856 6500 18884
rect 8163 18856 8208 18884
rect 3844 18844 3850 18856
rect 1673 18819 1731 18825
rect 1673 18785 1685 18819
rect 1719 18816 1731 18819
rect 2590 18816 2596 18828
rect 1719 18788 2596 18816
rect 1719 18785 1731 18788
rect 1673 18779 1731 18785
rect 2590 18776 2596 18788
rect 2648 18816 2654 18828
rect 3418 18816 3424 18828
rect 2648 18788 3424 18816
rect 2648 18776 2654 18788
rect 3418 18776 3424 18788
rect 3476 18776 3482 18828
rect 4614 18816 4620 18828
rect 4575 18788 4620 18816
rect 4614 18776 4620 18788
rect 4672 18776 4678 18828
rect 4706 18776 4712 18828
rect 4764 18816 4770 18828
rect 5169 18819 5227 18825
rect 5169 18816 5181 18819
rect 4764 18788 5181 18816
rect 4764 18776 4770 18788
rect 5169 18785 5181 18788
rect 5215 18785 5227 18819
rect 5169 18779 5227 18785
rect 5353 18819 5411 18825
rect 5353 18785 5365 18819
rect 5399 18816 5411 18819
rect 5442 18816 5448 18828
rect 5399 18788 5448 18816
rect 5399 18785 5411 18788
rect 5353 18779 5411 18785
rect 2406 18708 2412 18760
rect 2464 18748 2470 18760
rect 2961 18751 3019 18757
rect 2961 18748 2973 18751
rect 2464 18720 2973 18748
rect 2464 18708 2470 18720
rect 2961 18717 2973 18720
rect 3007 18748 3019 18751
rect 5074 18748 5080 18760
rect 3007 18720 5080 18748
rect 3007 18717 3019 18720
rect 2961 18711 3019 18717
rect 5074 18708 5080 18720
rect 5132 18708 5138 18760
rect 5184 18748 5212 18779
rect 5442 18776 5448 18788
rect 5500 18776 5506 18828
rect 6270 18816 6276 18828
rect 6231 18788 6276 18816
rect 6270 18776 6276 18788
rect 6328 18776 6334 18828
rect 6472 18825 6500 18856
rect 8202 18844 8208 18856
rect 8260 18844 8266 18896
rect 9784 18893 9812 18924
rect 11698 18912 11704 18924
rect 11756 18912 11762 18964
rect 14826 18912 14832 18964
rect 14884 18952 14890 18964
rect 15013 18955 15071 18961
rect 15013 18952 15025 18955
rect 14884 18924 15025 18952
rect 14884 18912 14890 18924
rect 15013 18921 15025 18924
rect 15059 18921 15071 18955
rect 15013 18915 15071 18921
rect 18046 18912 18052 18964
rect 18104 18952 18110 18964
rect 18509 18955 18567 18961
rect 18509 18952 18521 18955
rect 18104 18924 18521 18952
rect 18104 18912 18110 18924
rect 18509 18921 18521 18924
rect 18555 18952 18567 18955
rect 19242 18952 19248 18964
rect 18555 18924 19248 18952
rect 18555 18921 18567 18924
rect 18509 18915 18567 18921
rect 19242 18912 19248 18924
rect 19300 18912 19306 18964
rect 9769 18887 9827 18893
rect 9769 18853 9781 18887
rect 9815 18853 9827 18887
rect 9769 18847 9827 18853
rect 9858 18844 9864 18896
rect 9916 18884 9922 18896
rect 12618 18884 12624 18896
rect 9916 18856 9961 18884
rect 12531 18856 12624 18884
rect 9916 18844 9922 18856
rect 12618 18844 12624 18856
rect 12676 18884 12682 18896
rect 13265 18887 13323 18893
rect 13265 18884 13277 18887
rect 12676 18856 13277 18884
rect 12676 18844 12682 18856
rect 13265 18853 13277 18856
rect 13311 18884 13323 18887
rect 13814 18884 13820 18896
rect 13311 18856 13820 18884
rect 13311 18853 13323 18856
rect 13265 18847 13323 18853
rect 13814 18844 13820 18856
rect 13872 18844 13878 18896
rect 15746 18884 15752 18896
rect 15707 18856 15752 18884
rect 15746 18844 15752 18856
rect 15804 18844 15810 18896
rect 19150 18884 19156 18896
rect 19111 18856 19156 18884
rect 19150 18844 19156 18856
rect 19208 18844 19214 18896
rect 19705 18887 19763 18893
rect 19705 18853 19717 18887
rect 19751 18884 19763 18887
rect 20162 18884 20168 18896
rect 19751 18856 20168 18884
rect 19751 18853 19763 18856
rect 19705 18847 19763 18853
rect 20162 18844 20168 18856
rect 20220 18884 20226 18896
rect 20530 18884 20536 18896
rect 20220 18856 20536 18884
rect 20220 18844 20226 18856
rect 20530 18844 20536 18856
rect 20588 18844 20594 18896
rect 6457 18819 6515 18825
rect 6457 18785 6469 18819
rect 6503 18816 6515 18819
rect 6546 18816 6552 18828
rect 6503 18788 6552 18816
rect 6503 18785 6515 18788
rect 6457 18779 6515 18785
rect 6546 18776 6552 18788
rect 6604 18776 6610 18828
rect 7561 18819 7619 18825
rect 7561 18785 7573 18819
rect 7607 18816 7619 18819
rect 7926 18816 7932 18828
rect 7607 18788 7932 18816
rect 7607 18785 7619 18788
rect 7561 18779 7619 18785
rect 7926 18776 7932 18788
rect 7984 18776 7990 18828
rect 10778 18816 10784 18828
rect 10739 18788 10784 18816
rect 10778 18776 10784 18788
rect 10836 18776 10842 18828
rect 12253 18819 12311 18825
rect 12253 18785 12265 18819
rect 12299 18816 12311 18819
rect 12636 18816 12664 18844
rect 12299 18788 12664 18816
rect 17681 18819 17739 18825
rect 12299 18785 12311 18788
rect 12253 18779 12311 18785
rect 17681 18785 17693 18819
rect 17727 18785 17739 18819
rect 17862 18816 17868 18828
rect 17823 18788 17868 18816
rect 17681 18779 17739 18785
rect 5721 18751 5779 18757
rect 5721 18748 5733 18751
rect 5184 18720 5733 18748
rect 5721 18717 5733 18720
rect 5767 18748 5779 18751
rect 5994 18748 6000 18760
rect 5767 18720 6000 18748
rect 5767 18717 5779 18720
rect 5721 18711 5779 18717
rect 5994 18708 6000 18720
rect 6052 18708 6058 18760
rect 6822 18748 6828 18760
rect 6783 18720 6828 18748
rect 6822 18708 6828 18720
rect 6880 18708 6886 18760
rect 8110 18748 8116 18760
rect 8071 18720 8116 18748
rect 8110 18708 8116 18720
rect 8168 18708 8174 18760
rect 8757 18751 8815 18757
rect 8757 18717 8769 18751
rect 8803 18748 8815 18751
rect 8803 18720 10916 18748
rect 8803 18717 8815 18720
rect 8757 18711 8815 18717
rect 1946 18640 1952 18692
rect 2004 18680 2010 18692
rect 4706 18680 4712 18692
rect 2004 18652 4712 18680
rect 2004 18640 2010 18652
rect 4706 18640 4712 18652
rect 4764 18640 4770 18692
rect 9122 18640 9128 18692
rect 9180 18680 9186 18692
rect 10321 18683 10379 18689
rect 10321 18680 10333 18683
rect 9180 18652 10333 18680
rect 9180 18640 9186 18652
rect 10321 18649 10333 18652
rect 10367 18649 10379 18683
rect 10888 18680 10916 18720
rect 10962 18708 10968 18760
rect 11020 18748 11026 18760
rect 11333 18751 11391 18757
rect 11333 18748 11345 18751
rect 11020 18720 11345 18748
rect 11020 18708 11026 18720
rect 11333 18717 11345 18720
rect 11379 18717 11391 18751
rect 11333 18711 11391 18717
rect 13173 18751 13231 18757
rect 13173 18717 13185 18751
rect 13219 18748 13231 18751
rect 13538 18748 13544 18760
rect 13219 18720 13544 18748
rect 13219 18717 13231 18720
rect 13173 18711 13231 18717
rect 13538 18708 13544 18720
rect 13596 18708 13602 18760
rect 15470 18708 15476 18760
rect 15528 18748 15534 18760
rect 15657 18751 15715 18757
rect 15657 18748 15669 18751
rect 15528 18720 15669 18748
rect 15528 18708 15534 18720
rect 15657 18717 15669 18720
rect 15703 18717 15715 18751
rect 16022 18748 16028 18760
rect 15983 18720 16028 18748
rect 15657 18711 15715 18717
rect 16022 18708 16028 18720
rect 16080 18708 16086 18760
rect 17696 18748 17724 18779
rect 17862 18776 17868 18788
rect 17920 18776 17926 18828
rect 17954 18748 17960 18760
rect 16592 18720 17960 18748
rect 11422 18680 11428 18692
rect 10888 18652 11428 18680
rect 10321 18643 10379 18649
rect 3329 18615 3387 18621
rect 3329 18581 3341 18615
rect 3375 18612 3387 18615
rect 3605 18615 3663 18621
rect 3605 18612 3617 18615
rect 3375 18584 3617 18612
rect 3375 18581 3387 18584
rect 3329 18575 3387 18581
rect 3605 18581 3617 18584
rect 3651 18612 3663 18615
rect 3786 18612 3792 18624
rect 3651 18584 3792 18612
rect 3651 18581 3663 18584
rect 3605 18575 3663 18581
rect 3786 18572 3792 18584
rect 3844 18572 3850 18624
rect 7650 18572 7656 18624
rect 7708 18612 7714 18624
rect 7837 18615 7895 18621
rect 7837 18612 7849 18615
rect 7708 18584 7849 18612
rect 7708 18572 7714 18584
rect 7837 18581 7849 18584
rect 7883 18581 7895 18615
rect 10336 18612 10364 18643
rect 11422 18640 11428 18652
rect 11480 18680 11486 18692
rect 13725 18683 13783 18689
rect 13725 18680 13737 18683
rect 11480 18652 13737 18680
rect 11480 18640 11486 18652
rect 13725 18649 13737 18652
rect 13771 18649 13783 18683
rect 14550 18680 14556 18692
rect 14463 18652 14556 18680
rect 13725 18643 13783 18649
rect 14550 18640 14556 18652
rect 14608 18680 14614 18692
rect 16592 18680 16620 18720
rect 17954 18708 17960 18720
rect 18012 18708 18018 18760
rect 18141 18751 18199 18757
rect 18141 18717 18153 18751
rect 18187 18748 18199 18751
rect 18690 18748 18696 18760
rect 18187 18720 18696 18748
rect 18187 18717 18199 18720
rect 18141 18711 18199 18717
rect 18690 18708 18696 18720
rect 18748 18748 18754 18760
rect 18785 18751 18843 18757
rect 18785 18748 18797 18751
rect 18748 18720 18797 18748
rect 18748 18708 18754 18720
rect 18785 18717 18797 18720
rect 18831 18717 18843 18751
rect 19058 18748 19064 18760
rect 19019 18720 19064 18748
rect 18785 18711 18843 18717
rect 19058 18708 19064 18720
rect 19116 18708 19122 18760
rect 19242 18708 19248 18760
rect 19300 18748 19306 18760
rect 20901 18751 20959 18757
rect 20901 18748 20913 18751
rect 19300 18720 20913 18748
rect 19300 18708 19306 18720
rect 20901 18717 20913 18720
rect 20947 18717 20959 18751
rect 20901 18711 20959 18717
rect 14608 18652 16620 18680
rect 14608 18640 14614 18652
rect 16666 18640 16672 18692
rect 16724 18680 16730 18692
rect 21726 18680 21732 18692
rect 16724 18652 21732 18680
rect 16724 18640 16730 18652
rect 21726 18640 21732 18652
rect 21784 18640 21790 18692
rect 12342 18612 12348 18624
rect 10336 18584 12348 18612
rect 7837 18575 7895 18581
rect 12342 18572 12348 18584
rect 12400 18572 12406 18624
rect 12526 18572 12532 18624
rect 12584 18612 12590 18624
rect 12986 18612 12992 18624
rect 12584 18584 12992 18612
rect 12584 18572 12590 18584
rect 12986 18572 12992 18584
rect 13044 18572 13050 18624
rect 14182 18612 14188 18624
rect 14143 18584 14188 18612
rect 14182 18572 14188 18584
rect 14240 18572 14246 18624
rect 19978 18612 19984 18624
rect 19939 18584 19984 18612
rect 19978 18572 19984 18584
rect 20036 18572 20042 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 2682 18368 2688 18420
rect 2740 18408 2746 18420
rect 2958 18408 2964 18420
rect 2740 18380 2785 18408
rect 2919 18380 2964 18408
rect 2740 18368 2746 18380
rect 2958 18368 2964 18380
rect 3016 18368 3022 18420
rect 3973 18411 4031 18417
rect 3973 18377 3985 18411
rect 4019 18408 4031 18411
rect 4341 18411 4399 18417
rect 4341 18408 4353 18411
rect 4019 18380 4353 18408
rect 4019 18377 4031 18380
rect 3973 18371 4031 18377
rect 4341 18377 4353 18380
rect 4387 18408 4399 18411
rect 4614 18408 4620 18420
rect 4387 18380 4620 18408
rect 4387 18377 4399 18380
rect 4341 18371 4399 18377
rect 4614 18368 4620 18380
rect 4672 18368 4678 18420
rect 6546 18408 6552 18420
rect 6507 18380 6552 18408
rect 6546 18368 6552 18380
rect 6604 18368 6610 18420
rect 7742 18408 7748 18420
rect 7703 18380 7748 18408
rect 7742 18368 7748 18380
rect 7800 18368 7806 18420
rect 9674 18368 9680 18420
rect 9732 18408 9738 18420
rect 10597 18411 10655 18417
rect 10597 18408 10609 18411
rect 9732 18380 10609 18408
rect 9732 18368 9738 18380
rect 10597 18377 10609 18380
rect 10643 18377 10655 18411
rect 10597 18371 10655 18377
rect 11698 18368 11704 18420
rect 11756 18408 11762 18420
rect 11977 18411 12035 18417
rect 11977 18408 11989 18411
rect 11756 18380 11989 18408
rect 11756 18368 11762 18380
rect 11977 18377 11989 18380
rect 12023 18377 12035 18411
rect 11977 18371 12035 18377
rect 13814 18368 13820 18420
rect 13872 18408 13878 18420
rect 13872 18380 13917 18408
rect 13872 18368 13878 18380
rect 17218 18368 17224 18420
rect 17276 18408 17282 18420
rect 17497 18411 17555 18417
rect 17497 18408 17509 18411
rect 17276 18380 17509 18408
rect 17276 18368 17282 18380
rect 17497 18377 17509 18380
rect 17543 18408 17555 18411
rect 17862 18408 17868 18420
rect 17543 18380 17868 18408
rect 17543 18377 17555 18380
rect 17497 18371 17555 18377
rect 17862 18368 17868 18380
rect 17920 18368 17926 18420
rect 18414 18368 18420 18420
rect 18472 18408 18478 18420
rect 18509 18411 18567 18417
rect 18509 18408 18521 18411
rect 18472 18380 18521 18408
rect 18472 18368 18478 18380
rect 18509 18377 18521 18380
rect 18555 18377 18567 18411
rect 18509 18371 18567 18377
rect 19613 18411 19671 18417
rect 19613 18377 19625 18411
rect 19659 18408 19671 18411
rect 19978 18408 19984 18420
rect 19659 18380 19984 18408
rect 19659 18377 19671 18380
rect 19613 18371 19671 18377
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 9030 18300 9036 18352
rect 9088 18340 9094 18352
rect 10229 18343 10287 18349
rect 10229 18340 10241 18343
rect 9088 18312 10241 18340
rect 9088 18300 9094 18312
rect 10229 18309 10241 18312
rect 10275 18340 10287 18343
rect 11606 18340 11612 18352
rect 10275 18312 11612 18340
rect 10275 18309 10287 18312
rect 10229 18303 10287 18309
rect 11606 18300 11612 18312
rect 11664 18340 11670 18352
rect 13081 18343 13139 18349
rect 13081 18340 13093 18343
rect 11664 18312 13093 18340
rect 11664 18300 11670 18312
rect 13081 18309 13093 18312
rect 13127 18309 13139 18343
rect 13081 18303 13139 18309
rect 13630 18300 13636 18352
rect 13688 18340 13694 18352
rect 13906 18340 13912 18352
rect 13688 18312 13912 18340
rect 13688 18300 13694 18312
rect 13906 18300 13912 18312
rect 13964 18300 13970 18352
rect 19058 18300 19064 18352
rect 19116 18340 19122 18352
rect 19889 18343 19947 18349
rect 19889 18340 19901 18343
rect 19116 18312 19901 18340
rect 19116 18300 19122 18312
rect 19889 18309 19901 18312
rect 19935 18309 19947 18343
rect 19889 18303 19947 18309
rect 2501 18275 2559 18281
rect 2501 18241 2513 18275
rect 2547 18272 2559 18275
rect 3050 18272 3056 18284
rect 2547 18244 3056 18272
rect 2547 18241 2559 18244
rect 2501 18235 2559 18241
rect 3050 18232 3056 18244
rect 3108 18272 3114 18284
rect 3513 18275 3571 18281
rect 3513 18272 3525 18275
rect 3108 18244 3525 18272
rect 3108 18232 3114 18244
rect 3513 18241 3525 18244
rect 3559 18272 3571 18275
rect 9677 18275 9735 18281
rect 3559 18244 5488 18272
rect 3559 18241 3571 18244
rect 3513 18235 3571 18241
rect 5460 18216 5488 18244
rect 9677 18241 9689 18275
rect 9723 18272 9735 18275
rect 9950 18272 9956 18284
rect 9723 18244 9956 18272
rect 9723 18241 9735 18244
rect 9677 18235 9735 18241
rect 9950 18232 9956 18244
rect 10008 18272 10014 18284
rect 11287 18275 11345 18281
rect 11287 18272 11299 18275
rect 10008 18244 11299 18272
rect 10008 18232 10014 18244
rect 11287 18241 11299 18244
rect 11333 18241 11345 18275
rect 11287 18235 11345 18241
rect 12529 18275 12587 18281
rect 12529 18241 12541 18275
rect 12575 18272 12587 18275
rect 12894 18272 12900 18284
rect 12575 18244 12900 18272
rect 12575 18241 12587 18244
rect 12529 18235 12587 18241
rect 12894 18232 12900 18244
rect 12952 18232 12958 18284
rect 16022 18232 16028 18284
rect 16080 18272 16086 18284
rect 16482 18272 16488 18284
rect 16080 18244 16488 18272
rect 16080 18232 16086 18244
rect 16482 18232 16488 18244
rect 16540 18232 16546 18284
rect 16758 18272 16764 18284
rect 16719 18244 16764 18272
rect 16758 18232 16764 18244
rect 16816 18232 16822 18284
rect 18690 18272 18696 18284
rect 18651 18244 18696 18272
rect 18690 18232 18696 18244
rect 18748 18232 18754 18284
rect 20254 18232 20260 18284
rect 20312 18272 20318 18284
rect 20809 18275 20867 18281
rect 20809 18272 20821 18275
rect 20312 18244 20821 18272
rect 20312 18232 20318 18244
rect 20809 18241 20821 18244
rect 20855 18241 20867 18275
rect 20809 18235 20867 18241
rect 1857 18207 1915 18213
rect 1857 18173 1869 18207
rect 1903 18173 1915 18207
rect 2406 18204 2412 18216
rect 2367 18176 2412 18204
rect 1857 18167 1915 18173
rect 1762 18096 1768 18148
rect 1820 18136 1826 18148
rect 1872 18136 1900 18167
rect 2406 18164 2412 18176
rect 2464 18164 2470 18216
rect 4614 18204 4620 18216
rect 4575 18176 4620 18204
rect 4614 18164 4620 18176
rect 4672 18164 4678 18216
rect 5074 18164 5080 18216
rect 5132 18204 5138 18216
rect 5261 18207 5319 18213
rect 5261 18204 5273 18207
rect 5132 18176 5273 18204
rect 5132 18164 5138 18176
rect 5261 18173 5273 18176
rect 5307 18173 5319 18207
rect 5442 18204 5448 18216
rect 5403 18176 5448 18204
rect 5261 18167 5319 18173
rect 3786 18136 3792 18148
rect 1820 18108 3792 18136
rect 1820 18096 1826 18108
rect 3786 18096 3792 18108
rect 3844 18096 3850 18148
rect 5276 18136 5304 18167
rect 5442 18164 5448 18176
rect 5500 18204 5506 18216
rect 5813 18207 5871 18213
rect 5813 18204 5825 18207
rect 5500 18176 5825 18204
rect 5500 18164 5506 18176
rect 5813 18173 5825 18176
rect 5859 18173 5871 18207
rect 5813 18167 5871 18173
rect 5997 18207 6055 18213
rect 5997 18173 6009 18207
rect 6043 18204 6055 18207
rect 6638 18204 6644 18216
rect 6043 18176 6644 18204
rect 6043 18173 6055 18176
rect 5997 18167 6055 18173
rect 6638 18164 6644 18176
rect 6696 18204 6702 18216
rect 6860 18207 6918 18213
rect 6860 18204 6872 18207
rect 6696 18176 6872 18204
rect 6696 18164 6702 18176
rect 6860 18173 6872 18176
rect 6906 18204 6918 18207
rect 7285 18207 7343 18213
rect 7285 18204 7297 18207
rect 6906 18176 7297 18204
rect 6906 18173 6918 18176
rect 6860 18167 6918 18173
rect 7285 18173 7297 18176
rect 7331 18173 7343 18207
rect 7285 18167 7343 18173
rect 7650 18164 7656 18216
rect 7708 18204 7714 18216
rect 7837 18207 7895 18213
rect 7837 18204 7849 18207
rect 7708 18176 7849 18204
rect 7708 18164 7714 18176
rect 7837 18173 7849 18176
rect 7883 18173 7895 18207
rect 7837 18167 7895 18173
rect 8757 18207 8815 18213
rect 8757 18173 8769 18207
rect 8803 18173 8815 18207
rect 8757 18167 8815 18173
rect 11200 18207 11258 18213
rect 11200 18173 11212 18207
rect 11246 18204 11258 18207
rect 11514 18204 11520 18216
rect 11246 18176 11520 18204
rect 11246 18173 11258 18176
rect 11200 18167 11258 18173
rect 5276 18108 6224 18136
rect 6196 18080 6224 18108
rect 7742 18096 7748 18148
rect 7800 18136 7806 18148
rect 8158 18139 8216 18145
rect 8158 18136 8170 18139
rect 7800 18108 8170 18136
rect 7800 18096 7806 18108
rect 8158 18105 8170 18108
rect 8204 18105 8216 18139
rect 8772 18136 8800 18167
rect 11514 18164 11520 18176
rect 11572 18204 11578 18216
rect 11609 18207 11667 18213
rect 11609 18204 11621 18207
rect 11572 18176 11621 18204
rect 11572 18164 11578 18176
rect 11609 18173 11621 18176
rect 11655 18173 11667 18207
rect 14642 18204 14648 18216
rect 14603 18176 14648 18204
rect 11609 18167 11667 18173
rect 14642 18164 14648 18176
rect 14700 18164 14706 18216
rect 9125 18139 9183 18145
rect 9125 18136 9137 18139
rect 8772 18108 9137 18136
rect 8158 18099 8216 18105
rect 9125 18105 9137 18108
rect 9171 18136 9183 18139
rect 9493 18139 9551 18145
rect 9493 18136 9505 18139
rect 9171 18108 9505 18136
rect 9171 18105 9183 18108
rect 9125 18099 9183 18105
rect 9493 18105 9505 18108
rect 9539 18136 9551 18139
rect 9769 18139 9827 18145
rect 9769 18136 9781 18139
rect 9539 18108 9781 18136
rect 9539 18105 9551 18108
rect 9493 18099 9551 18105
rect 9769 18105 9781 18108
rect 9815 18136 9827 18139
rect 9858 18136 9864 18148
rect 9815 18108 9864 18136
rect 9815 18105 9827 18108
rect 9769 18099 9827 18105
rect 9858 18096 9864 18108
rect 9916 18096 9922 18148
rect 12618 18096 12624 18148
rect 12676 18136 12682 18148
rect 14550 18136 14556 18148
rect 12676 18108 12721 18136
rect 14511 18108 14556 18136
rect 12676 18096 12682 18108
rect 14550 18096 14556 18108
rect 14608 18136 14614 18148
rect 14966 18139 15024 18145
rect 14966 18136 14978 18139
rect 14608 18108 14978 18136
rect 14608 18096 14614 18108
rect 14966 18105 14978 18108
rect 15012 18105 15024 18139
rect 14966 18099 15024 18105
rect 16577 18139 16635 18145
rect 16577 18105 16589 18139
rect 16623 18105 16635 18139
rect 16577 18099 16635 18105
rect 4522 18068 4528 18080
rect 4483 18040 4528 18068
rect 4522 18028 4528 18040
rect 4580 18028 4586 18080
rect 4614 18028 4620 18080
rect 4672 18068 4678 18080
rect 5997 18071 6055 18077
rect 5997 18068 6009 18071
rect 4672 18040 6009 18068
rect 4672 18028 4678 18040
rect 5997 18037 6009 18040
rect 6043 18037 6055 18071
rect 6178 18068 6184 18080
rect 6139 18040 6184 18068
rect 5997 18031 6055 18037
rect 6178 18028 6184 18040
rect 6236 18028 6242 18080
rect 6963 18071 7021 18077
rect 6963 18037 6975 18071
rect 7009 18068 7021 18071
rect 7190 18068 7196 18080
rect 7009 18040 7196 18068
rect 7009 18037 7021 18040
rect 6963 18031 7021 18037
rect 7190 18028 7196 18040
rect 7248 18028 7254 18080
rect 10962 18068 10968 18080
rect 10923 18040 10968 18068
rect 10962 18028 10968 18040
rect 11020 18028 11026 18080
rect 13538 18068 13544 18080
rect 13499 18040 13544 18068
rect 13538 18028 13544 18040
rect 13596 18028 13602 18080
rect 15562 18068 15568 18080
rect 15523 18040 15568 18068
rect 15562 18028 15568 18040
rect 15620 18068 15626 18080
rect 15746 18068 15752 18080
rect 15620 18040 15752 18068
rect 15620 18028 15626 18040
rect 15746 18028 15752 18040
rect 15804 18068 15810 18080
rect 15841 18071 15899 18077
rect 15841 18068 15853 18071
rect 15804 18040 15853 18068
rect 15804 18028 15810 18040
rect 15841 18037 15853 18040
rect 15887 18037 15899 18071
rect 16206 18068 16212 18080
rect 16167 18040 16212 18068
rect 15841 18031 15899 18037
rect 16206 18028 16212 18040
rect 16264 18068 16270 18080
rect 16592 18068 16620 18099
rect 18414 18096 18420 18148
rect 18472 18136 18478 18148
rect 19014 18139 19072 18145
rect 19014 18136 19026 18139
rect 18472 18108 19026 18136
rect 18472 18096 18478 18108
rect 19014 18105 19026 18108
rect 19060 18105 19072 18139
rect 20530 18136 20536 18148
rect 20491 18108 20536 18136
rect 19014 18099 19072 18105
rect 20530 18096 20536 18108
rect 20588 18096 20594 18148
rect 20625 18139 20683 18145
rect 20625 18105 20637 18139
rect 20671 18136 20683 18139
rect 21358 18136 21364 18148
rect 20671 18108 21364 18136
rect 20671 18105 20683 18108
rect 20625 18099 20683 18105
rect 16264 18040 16620 18068
rect 17865 18071 17923 18077
rect 16264 18028 16270 18040
rect 17865 18037 17877 18071
rect 17911 18068 17923 18071
rect 17954 18068 17960 18080
rect 17911 18040 17960 18068
rect 17911 18037 17923 18040
rect 17865 18031 17923 18037
rect 17954 18028 17960 18040
rect 18012 18028 18018 18080
rect 20349 18071 20407 18077
rect 20349 18037 20361 18071
rect 20395 18068 20407 18071
rect 20640 18068 20668 18099
rect 21358 18096 21364 18108
rect 21416 18096 21422 18148
rect 20395 18040 20668 18068
rect 20395 18037 20407 18040
rect 20349 18031 20407 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2590 17864 2596 17876
rect 2551 17836 2596 17864
rect 2590 17824 2596 17836
rect 2648 17824 2654 17876
rect 2961 17867 3019 17873
rect 2961 17833 2973 17867
rect 3007 17864 3019 17867
rect 3050 17864 3056 17876
rect 3007 17836 3056 17864
rect 3007 17833 3019 17836
rect 2961 17827 3019 17833
rect 2976 17796 3004 17827
rect 3050 17824 3056 17836
rect 3108 17824 3114 17876
rect 3881 17867 3939 17873
rect 3881 17833 3893 17867
rect 3927 17864 3939 17867
rect 3970 17864 3976 17876
rect 3927 17836 3976 17864
rect 3927 17833 3939 17836
rect 3881 17827 3939 17833
rect 3970 17824 3976 17836
rect 4028 17864 4034 17876
rect 4522 17864 4528 17876
rect 4028 17836 4528 17864
rect 4028 17824 4034 17836
rect 4522 17824 4528 17836
rect 4580 17824 4586 17876
rect 4798 17864 4804 17876
rect 4759 17836 4804 17864
rect 4798 17824 4804 17836
rect 4856 17824 4862 17876
rect 7377 17867 7435 17873
rect 7377 17833 7389 17867
rect 7423 17864 7435 17867
rect 8110 17864 8116 17876
rect 7423 17836 8116 17864
rect 7423 17833 7435 17836
rect 7377 17827 7435 17833
rect 8110 17824 8116 17836
rect 8168 17824 8174 17876
rect 8202 17824 8208 17876
rect 8260 17864 8266 17876
rect 8389 17867 8447 17873
rect 8389 17864 8401 17867
rect 8260 17836 8401 17864
rect 8260 17824 8266 17836
rect 8389 17833 8401 17836
rect 8435 17864 8447 17867
rect 8665 17867 8723 17873
rect 8665 17864 8677 17867
rect 8435 17836 8677 17864
rect 8435 17833 8447 17836
rect 8389 17827 8447 17833
rect 8665 17833 8677 17836
rect 8711 17833 8723 17867
rect 9950 17864 9956 17876
rect 9911 17836 9956 17864
rect 8665 17827 8723 17833
rect 9950 17824 9956 17836
rect 10008 17824 10014 17876
rect 11333 17867 11391 17873
rect 11333 17833 11345 17867
rect 11379 17864 11391 17867
rect 11422 17864 11428 17876
rect 11379 17836 11428 17864
rect 11379 17833 11391 17836
rect 11333 17827 11391 17833
rect 11422 17824 11428 17836
rect 11480 17824 11486 17876
rect 11606 17864 11612 17876
rect 11567 17836 11612 17864
rect 11606 17824 11612 17836
rect 11664 17824 11670 17876
rect 16206 17864 16212 17876
rect 16167 17836 16212 17864
rect 16206 17824 16212 17836
rect 16264 17824 16270 17876
rect 16482 17864 16488 17876
rect 16443 17836 16488 17864
rect 16482 17824 16488 17836
rect 16540 17824 16546 17876
rect 17218 17864 17224 17876
rect 17179 17836 17224 17864
rect 17218 17824 17224 17836
rect 17276 17824 17282 17876
rect 18414 17824 18420 17876
rect 18472 17864 18478 17876
rect 18509 17867 18567 17873
rect 18509 17864 18521 17867
rect 18472 17836 18521 17864
rect 18472 17824 18478 17836
rect 18509 17833 18521 17836
rect 18555 17833 18567 17867
rect 18509 17827 18567 17833
rect 19061 17867 19119 17873
rect 19061 17833 19073 17867
rect 19107 17864 19119 17867
rect 19150 17864 19156 17876
rect 19107 17836 19156 17864
rect 19107 17833 19119 17836
rect 19061 17827 19119 17833
rect 19150 17824 19156 17836
rect 19208 17864 19214 17876
rect 19337 17867 19395 17873
rect 19337 17864 19349 17867
rect 19208 17836 19349 17864
rect 19208 17824 19214 17836
rect 19337 17833 19349 17836
rect 19383 17833 19395 17867
rect 20530 17864 20536 17876
rect 20491 17836 20536 17864
rect 19337 17827 19395 17833
rect 20530 17824 20536 17836
rect 20588 17824 20594 17876
rect 5721 17799 5779 17805
rect 5721 17796 5733 17799
rect 2516 17768 3004 17796
rect 4356 17768 5733 17796
rect 2516 17740 2544 17768
rect 1762 17728 1768 17740
rect 1723 17700 1768 17728
rect 1762 17688 1768 17700
rect 1820 17688 1826 17740
rect 1946 17688 1952 17740
rect 2004 17728 2010 17740
rect 2317 17731 2375 17737
rect 2317 17728 2329 17731
rect 2004 17700 2329 17728
rect 2004 17688 2010 17700
rect 2317 17697 2329 17700
rect 2363 17697 2375 17731
rect 2317 17691 2375 17697
rect 2332 17660 2360 17691
rect 2498 17688 2504 17740
rect 2556 17728 2562 17740
rect 2556 17700 2649 17728
rect 2556 17688 2562 17700
rect 2866 17688 2872 17740
rect 2924 17728 2930 17740
rect 4356 17737 4384 17768
rect 5721 17765 5733 17768
rect 5767 17796 5779 17799
rect 6270 17796 6276 17808
rect 5767 17768 6276 17796
rect 5767 17765 5779 17768
rect 5721 17759 5779 17765
rect 6270 17756 6276 17768
rect 6328 17796 6334 17808
rect 6917 17799 6975 17805
rect 6917 17796 6929 17799
rect 6328 17768 6929 17796
rect 6328 17756 6334 17768
rect 6917 17765 6929 17768
rect 6963 17765 6975 17799
rect 7742 17796 7748 17808
rect 7703 17768 7748 17796
rect 6917 17759 6975 17765
rect 7742 17756 7748 17768
rect 7800 17756 7806 17808
rect 10962 17796 10968 17808
rect 10923 17768 10968 17796
rect 10962 17756 10968 17768
rect 11020 17756 11026 17808
rect 11882 17756 11888 17808
rect 11940 17796 11946 17808
rect 11977 17799 12035 17805
rect 11977 17796 11989 17799
rect 11940 17768 11989 17796
rect 11940 17756 11946 17768
rect 11977 17765 11989 17768
rect 12023 17765 12035 17799
rect 11977 17759 12035 17765
rect 15651 17799 15709 17805
rect 15651 17765 15663 17799
rect 15697 17796 15709 17799
rect 16022 17796 16028 17808
rect 15697 17768 16028 17796
rect 15697 17765 15709 17768
rect 15651 17759 15709 17765
rect 16022 17756 16028 17768
rect 16080 17756 16086 17808
rect 16868 17768 18092 17796
rect 4341 17731 4399 17737
rect 4341 17728 4353 17731
rect 2924 17700 4353 17728
rect 2924 17688 2930 17700
rect 4341 17697 4353 17700
rect 4387 17697 4399 17731
rect 4341 17691 4399 17697
rect 4522 17688 4528 17740
rect 4580 17728 4586 17740
rect 4617 17731 4675 17737
rect 4617 17728 4629 17731
rect 4580 17700 4629 17728
rect 4580 17688 4586 17700
rect 4617 17697 4629 17700
rect 4663 17697 4675 17731
rect 6086 17728 6092 17740
rect 6047 17700 6092 17728
rect 4617 17691 4675 17697
rect 6086 17688 6092 17700
rect 6144 17688 6150 17740
rect 6457 17731 6515 17737
rect 6457 17697 6469 17731
rect 6503 17728 6515 17731
rect 6730 17728 6736 17740
rect 6503 17700 6736 17728
rect 6503 17697 6515 17700
rect 6457 17691 6515 17697
rect 6730 17688 6736 17700
rect 6788 17688 6794 17740
rect 10134 17688 10140 17740
rect 10192 17728 10198 17740
rect 10229 17731 10287 17737
rect 10229 17728 10241 17731
rect 10192 17700 10241 17728
rect 10192 17688 10198 17700
rect 10229 17697 10241 17700
rect 10275 17697 10287 17731
rect 10229 17691 10287 17697
rect 2590 17660 2596 17672
rect 2332 17632 2596 17660
rect 2590 17620 2596 17632
rect 2648 17620 2654 17672
rect 4433 17663 4491 17669
rect 4433 17660 4445 17663
rect 3436 17632 4445 17660
rect 3436 17536 3464 17632
rect 4433 17629 4445 17632
rect 4479 17629 4491 17663
rect 4433 17623 4491 17629
rect 6641 17663 6699 17669
rect 6641 17629 6653 17663
rect 6687 17660 6699 17663
rect 7466 17660 7472 17672
rect 6687 17632 7472 17660
rect 6687 17629 6699 17632
rect 6641 17623 6699 17629
rect 7466 17620 7472 17632
rect 7524 17620 7530 17672
rect 3510 17552 3516 17604
rect 3568 17592 3574 17604
rect 6914 17592 6920 17604
rect 3568 17564 6920 17592
rect 3568 17552 3574 17564
rect 6914 17552 6920 17564
rect 6972 17552 6978 17604
rect 10244 17592 10272 17691
rect 10594 17688 10600 17740
rect 10652 17728 10658 17740
rect 10689 17731 10747 17737
rect 10689 17728 10701 17731
rect 10652 17700 10701 17728
rect 10652 17688 10658 17700
rect 10689 17697 10701 17700
rect 10735 17697 10747 17731
rect 10689 17691 10747 17697
rect 13538 17688 13544 17740
rect 13596 17728 13602 17740
rect 13633 17731 13691 17737
rect 13633 17728 13645 17731
rect 13596 17700 13645 17728
rect 13596 17688 13602 17700
rect 13633 17697 13645 17700
rect 13679 17728 13691 17731
rect 13722 17728 13728 17740
rect 13679 17700 13728 17728
rect 13679 17697 13691 17700
rect 13633 17691 13691 17697
rect 13722 17688 13728 17700
rect 13780 17688 13786 17740
rect 14090 17728 14096 17740
rect 14051 17700 14096 17728
rect 14090 17688 14096 17700
rect 14148 17688 14154 17740
rect 15105 17731 15163 17737
rect 15105 17697 15117 17731
rect 15151 17728 15163 17731
rect 15470 17728 15476 17740
rect 15151 17700 15476 17728
rect 15151 17697 15163 17700
rect 15105 17691 15163 17697
rect 15470 17688 15476 17700
rect 15528 17728 15534 17740
rect 16868 17728 16896 17768
rect 17034 17728 17040 17740
rect 15528 17700 16896 17728
rect 16995 17700 17040 17728
rect 15528 17688 15534 17700
rect 17034 17688 17040 17700
rect 17092 17688 17098 17740
rect 18064 17728 18092 17768
rect 20622 17728 20628 17740
rect 18064 17700 20628 17728
rect 20622 17688 20628 17700
rect 20680 17688 20686 17740
rect 20968 17731 21026 17737
rect 20968 17697 20980 17731
rect 21014 17728 21026 17731
rect 21358 17728 21364 17740
rect 21014 17700 21364 17728
rect 21014 17697 21026 17700
rect 20968 17691 21026 17697
rect 21358 17688 21364 17700
rect 21416 17688 21422 17740
rect 11606 17620 11612 17672
rect 11664 17660 11670 17672
rect 11885 17663 11943 17669
rect 11885 17660 11897 17663
rect 11664 17632 11897 17660
rect 11664 17620 11670 17632
rect 11885 17629 11897 17632
rect 11931 17629 11943 17663
rect 12158 17660 12164 17672
rect 12119 17632 12164 17660
rect 11885 17623 11943 17629
rect 12158 17620 12164 17632
rect 12216 17620 12222 17672
rect 14369 17663 14427 17669
rect 14369 17629 14381 17663
rect 14415 17660 14427 17663
rect 15289 17663 15347 17669
rect 15289 17660 15301 17663
rect 14415 17632 15301 17660
rect 14415 17629 14427 17632
rect 14369 17623 14427 17629
rect 15289 17629 15301 17632
rect 15335 17660 15347 17663
rect 16298 17660 16304 17672
rect 15335 17632 16304 17660
rect 15335 17629 15347 17632
rect 15289 17623 15347 17629
rect 16298 17620 16304 17632
rect 16356 17620 16362 17672
rect 18138 17660 18144 17672
rect 18099 17632 18144 17660
rect 18138 17620 18144 17632
rect 18196 17620 18202 17672
rect 10244 17564 13814 17592
rect 3418 17524 3424 17536
rect 3379 17496 3424 17524
rect 3418 17484 3424 17496
rect 3476 17484 3482 17536
rect 5445 17527 5503 17533
rect 5445 17493 5457 17527
rect 5491 17524 5503 17527
rect 5534 17524 5540 17536
rect 5491 17496 5540 17524
rect 5491 17493 5503 17496
rect 5445 17487 5503 17493
rect 5534 17484 5540 17496
rect 5592 17484 5598 17536
rect 12894 17524 12900 17536
rect 12855 17496 12900 17524
rect 12894 17484 12900 17496
rect 12952 17484 12958 17536
rect 13786 17524 13814 17564
rect 14642 17552 14648 17604
rect 14700 17592 14706 17604
rect 14737 17595 14795 17601
rect 14737 17592 14749 17595
rect 14700 17564 14749 17592
rect 14700 17552 14706 17564
rect 14737 17561 14749 17564
rect 14783 17592 14795 17595
rect 18966 17592 18972 17604
rect 14783 17564 18972 17592
rect 14783 17561 14795 17564
rect 14737 17555 14795 17561
rect 18966 17552 18972 17564
rect 19024 17552 19030 17604
rect 13998 17524 14004 17536
rect 13786 17496 14004 17524
rect 13998 17484 14004 17496
rect 14056 17524 14062 17536
rect 15930 17524 15936 17536
rect 14056 17496 15936 17524
rect 14056 17484 14062 17496
rect 15930 17484 15936 17496
rect 15988 17484 15994 17536
rect 19426 17484 19432 17536
rect 19484 17524 19490 17536
rect 21039 17527 21097 17533
rect 21039 17524 21051 17527
rect 19484 17496 21051 17524
rect 19484 17484 19490 17496
rect 21039 17493 21051 17496
rect 21085 17493 21097 17527
rect 21039 17487 21097 17493
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1673 17323 1731 17329
rect 1673 17289 1685 17323
rect 1719 17320 1731 17323
rect 2498 17320 2504 17332
rect 1719 17292 2504 17320
rect 1719 17289 1731 17292
rect 1673 17283 1731 17289
rect 2498 17280 2504 17292
rect 2556 17280 2562 17332
rect 4246 17280 4252 17332
rect 4304 17320 4310 17332
rect 4982 17320 4988 17332
rect 4304 17292 4988 17320
rect 4304 17280 4310 17292
rect 4982 17280 4988 17292
rect 5040 17320 5046 17332
rect 5629 17323 5687 17329
rect 5629 17320 5641 17323
rect 5040 17292 5641 17320
rect 5040 17280 5046 17292
rect 5629 17289 5641 17292
rect 5675 17289 5687 17323
rect 5629 17283 5687 17289
rect 6086 17280 6092 17332
rect 6144 17320 6150 17332
rect 6181 17323 6239 17329
rect 6181 17320 6193 17323
rect 6144 17292 6193 17320
rect 6144 17280 6150 17292
rect 6181 17289 6193 17292
rect 6227 17320 6239 17323
rect 7098 17320 7104 17332
rect 6227 17292 7104 17320
rect 6227 17289 6239 17292
rect 6181 17283 6239 17289
rect 7098 17280 7104 17292
rect 7156 17280 7162 17332
rect 7742 17280 7748 17332
rect 7800 17320 7806 17332
rect 7929 17323 7987 17329
rect 7929 17320 7941 17323
rect 7800 17292 7941 17320
rect 7800 17280 7806 17292
rect 7929 17289 7941 17292
rect 7975 17289 7987 17323
rect 7929 17283 7987 17289
rect 8202 17280 8208 17332
rect 8260 17320 8266 17332
rect 8297 17323 8355 17329
rect 8297 17320 8309 17323
rect 8260 17292 8309 17320
rect 8260 17280 8266 17292
rect 8297 17289 8309 17292
rect 8343 17289 8355 17323
rect 9309 17323 9367 17329
rect 9309 17320 9321 17323
rect 8297 17283 8355 17289
rect 8956 17292 9321 17320
rect 4065 17255 4123 17261
rect 4065 17252 4077 17255
rect 3620 17224 4077 17252
rect 1670 17144 1676 17196
rect 1728 17184 1734 17196
rect 2041 17187 2099 17193
rect 2041 17184 2053 17187
rect 1728 17156 2053 17184
rect 1728 17144 1734 17156
rect 2041 17153 2053 17156
rect 2087 17184 2099 17187
rect 2682 17184 2688 17196
rect 2087 17156 2688 17184
rect 2087 17153 2099 17156
rect 2041 17147 2099 17153
rect 2682 17144 2688 17156
rect 2740 17184 2746 17196
rect 3620 17193 3648 17224
rect 4065 17221 4077 17224
rect 4111 17221 4123 17255
rect 4801 17255 4859 17261
rect 4801 17252 4813 17255
rect 4065 17215 4123 17221
rect 4448 17224 4813 17252
rect 4448 17196 4476 17224
rect 4801 17221 4813 17224
rect 4847 17221 4859 17255
rect 8956 17252 8984 17292
rect 9309 17289 9321 17292
rect 9355 17289 9367 17323
rect 9309 17283 9367 17289
rect 9398 17280 9404 17332
rect 9456 17320 9462 17332
rect 9493 17323 9551 17329
rect 9493 17320 9505 17323
rect 9456 17292 9505 17320
rect 9456 17280 9462 17292
rect 9493 17289 9505 17292
rect 9539 17289 9551 17323
rect 16298 17320 16304 17332
rect 16259 17292 16304 17320
rect 9493 17283 9551 17289
rect 16298 17280 16304 17292
rect 16356 17280 16362 17332
rect 17034 17320 17040 17332
rect 16995 17292 17040 17320
rect 17034 17280 17040 17292
rect 17092 17280 17098 17332
rect 17497 17323 17555 17329
rect 17497 17289 17509 17323
rect 17543 17320 17555 17323
rect 18138 17320 18144 17332
rect 17543 17292 18144 17320
rect 17543 17289 17555 17292
rect 17497 17283 17555 17289
rect 18138 17280 18144 17292
rect 18196 17280 18202 17332
rect 18414 17320 18420 17332
rect 18248 17292 18420 17320
rect 9122 17252 9128 17264
rect 4801 17215 4859 17221
rect 7392 17224 8984 17252
rect 9083 17224 9128 17252
rect 3605 17187 3663 17193
rect 3605 17184 3617 17187
rect 2740 17156 3617 17184
rect 2740 17144 2746 17156
rect 2884 17125 2912 17156
rect 3605 17153 3617 17156
rect 3651 17153 3663 17187
rect 3605 17147 3663 17153
rect 3878 17144 3884 17196
rect 3936 17193 3942 17196
rect 3936 17187 3994 17193
rect 3936 17153 3948 17187
rect 3982 17153 3994 17187
rect 3936 17147 3994 17153
rect 4157 17187 4215 17193
rect 4157 17153 4169 17187
rect 4203 17184 4215 17187
rect 4430 17184 4436 17196
rect 4203 17156 4436 17184
rect 4203 17153 4215 17156
rect 4157 17147 4215 17153
rect 3936 17144 3942 17147
rect 4430 17144 4436 17156
rect 4488 17144 4494 17196
rect 4525 17187 4583 17193
rect 4525 17153 4537 17187
rect 4571 17184 4583 17187
rect 6362 17184 6368 17196
rect 4571 17156 6368 17184
rect 4571 17153 4583 17156
rect 4525 17147 4583 17153
rect 6362 17144 6368 17156
rect 6420 17144 6426 17196
rect 6730 17144 6736 17196
rect 6788 17184 6794 17196
rect 7392 17184 7420 17224
rect 9122 17212 9128 17224
rect 9180 17212 9186 17264
rect 7650 17184 7656 17196
rect 6788 17156 7420 17184
rect 7611 17156 7656 17184
rect 6788 17144 6794 17156
rect 2869 17119 2927 17125
rect 2869 17116 2881 17119
rect 2847 17088 2881 17116
rect 2869 17085 2881 17088
rect 2915 17085 2927 17119
rect 2869 17079 2927 17085
rect 2961 17119 3019 17125
rect 2961 17085 2973 17119
rect 3007 17116 3019 17119
rect 3418 17116 3424 17128
rect 3007 17088 3424 17116
rect 3007 17085 3019 17088
rect 2961 17079 3019 17085
rect 3418 17076 3424 17088
rect 3476 17076 3482 17128
rect 3694 17076 3700 17128
rect 3752 17116 3758 17128
rect 7392 17125 7420 17156
rect 7650 17144 7656 17156
rect 7708 17144 7714 17196
rect 8573 17187 8631 17193
rect 8573 17153 8585 17187
rect 8619 17184 8631 17187
rect 9416 17184 9444 17280
rect 10594 17212 10600 17264
rect 10652 17252 10658 17264
rect 10778 17252 10784 17264
rect 10652 17224 10784 17252
rect 10652 17212 10658 17224
rect 10778 17212 10784 17224
rect 10836 17212 10842 17264
rect 11422 17252 11428 17264
rect 10888 17224 11428 17252
rect 10888 17193 10916 17224
rect 11422 17212 11428 17224
rect 11480 17212 11486 17264
rect 16666 17252 16672 17264
rect 12820 17224 16672 17252
rect 8619 17156 9444 17184
rect 10873 17187 10931 17193
rect 8619 17153 8631 17156
rect 8573 17147 8631 17153
rect 10873 17153 10885 17187
rect 10919 17153 10931 17187
rect 10873 17147 10931 17153
rect 11517 17187 11575 17193
rect 11517 17153 11529 17187
rect 11563 17184 11575 17187
rect 12158 17184 12164 17196
rect 11563 17156 12164 17184
rect 11563 17153 11575 17156
rect 11517 17147 11575 17153
rect 12158 17144 12164 17156
rect 12216 17184 12222 17196
rect 12820 17193 12848 17224
rect 16666 17212 16672 17224
rect 16724 17212 16730 17264
rect 17865 17255 17923 17261
rect 17865 17221 17877 17255
rect 17911 17252 17923 17255
rect 18046 17252 18052 17264
rect 17911 17224 18052 17252
rect 17911 17221 17923 17224
rect 17865 17215 17923 17221
rect 18046 17212 18052 17224
rect 18104 17252 18110 17264
rect 18248 17252 18276 17292
rect 18414 17280 18420 17292
rect 18472 17280 18478 17332
rect 19426 17320 19432 17332
rect 19387 17292 19432 17320
rect 19426 17280 19432 17292
rect 19484 17280 19490 17332
rect 20027 17323 20085 17329
rect 20027 17289 20039 17323
rect 20073 17320 20085 17323
rect 20530 17320 20536 17332
rect 20073 17292 20536 17320
rect 20073 17289 20085 17292
rect 20027 17283 20085 17289
rect 20530 17280 20536 17292
rect 20588 17280 20594 17332
rect 20622 17280 20628 17332
rect 20680 17320 20686 17332
rect 21039 17323 21097 17329
rect 21039 17320 21051 17323
rect 20680 17292 21051 17320
rect 20680 17280 20686 17292
rect 21039 17289 21051 17292
rect 21085 17289 21097 17323
rect 25130 17320 25136 17332
rect 25091 17292 25136 17320
rect 21039 17283 21097 17289
rect 25130 17280 25136 17292
rect 25188 17280 25194 17332
rect 18104 17224 18276 17252
rect 18969 17255 19027 17261
rect 18104 17212 18110 17224
rect 18969 17221 18981 17255
rect 19015 17252 19027 17255
rect 19058 17252 19064 17264
rect 19015 17224 19064 17252
rect 19015 17221 19027 17224
rect 18969 17215 19027 17221
rect 19058 17212 19064 17224
rect 19116 17212 19122 17264
rect 12805 17187 12863 17193
rect 12805 17184 12817 17187
rect 12216 17156 12817 17184
rect 12216 17144 12222 17156
rect 12805 17153 12817 17156
rect 12851 17153 12863 17187
rect 17310 17184 17316 17196
rect 12805 17147 12863 17153
rect 13648 17156 17316 17184
rect 5169 17119 5227 17125
rect 5169 17116 5181 17119
rect 3752 17088 5181 17116
rect 3752 17076 3758 17088
rect 5169 17085 5181 17088
rect 5215 17116 5227 17119
rect 5537 17119 5595 17125
rect 5537 17116 5549 17119
rect 5215 17088 5549 17116
rect 5215 17085 5227 17088
rect 5169 17079 5227 17085
rect 5537 17085 5549 17088
rect 5583 17085 5595 17119
rect 5537 17079 5595 17085
rect 6641 17119 6699 17125
rect 6641 17085 6653 17119
rect 6687 17116 6699 17119
rect 7193 17119 7251 17125
rect 7193 17116 7205 17119
rect 6687 17088 7205 17116
rect 6687 17085 6699 17088
rect 6641 17079 6699 17085
rect 7193 17085 7205 17088
rect 7239 17085 7251 17119
rect 7193 17079 7251 17085
rect 7377 17119 7435 17125
rect 7377 17085 7389 17119
rect 7423 17085 7435 17119
rect 7377 17079 7435 17085
rect 9309 17119 9367 17125
rect 9309 17085 9321 17119
rect 9355 17116 9367 17119
rect 10594 17116 10600 17128
rect 9355 17088 10600 17116
rect 9355 17085 9367 17088
rect 9309 17079 9367 17085
rect 2406 17008 2412 17060
rect 2464 17048 2470 17060
rect 3329 17051 3387 17057
rect 3329 17048 3341 17051
rect 2464 17020 3341 17048
rect 2464 17008 2470 17020
rect 3329 17017 3341 17020
rect 3375 17048 3387 17051
rect 3789 17051 3847 17057
rect 3789 17048 3801 17051
rect 3375 17020 3801 17048
rect 3375 17017 3387 17020
rect 3329 17011 3387 17017
rect 3789 17017 3801 17020
rect 3835 17048 3847 17051
rect 4246 17048 4252 17060
rect 3835 17020 4252 17048
rect 3835 17017 3847 17020
rect 3789 17011 3847 17017
rect 4246 17008 4252 17020
rect 4304 17008 4310 17060
rect 5353 17051 5411 17057
rect 5353 17017 5365 17051
rect 5399 17017 5411 17051
rect 7208 17048 7236 17079
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 7650 17048 7656 17060
rect 7208 17020 7656 17048
rect 5353 17011 5411 17017
rect 5368 16980 5396 17011
rect 7650 17008 7656 17020
rect 7708 17048 7714 17060
rect 8570 17048 8576 17060
rect 7708 17020 8576 17048
rect 7708 17008 7714 17020
rect 8570 17008 8576 17020
rect 8628 17008 8634 17060
rect 8665 17051 8723 17057
rect 8665 17017 8677 17051
rect 8711 17017 8723 17051
rect 8665 17011 8723 17017
rect 9953 17051 10011 17057
rect 9953 17017 9965 17051
rect 9999 17048 10011 17051
rect 10965 17051 11023 17057
rect 9999 17020 10824 17048
rect 9999 17017 10011 17020
rect 9953 17011 10011 17017
rect 5534 16980 5540 16992
rect 5368 16952 5540 16980
rect 5534 16940 5540 16952
rect 5592 16940 5598 16992
rect 8202 16940 8208 16992
rect 8260 16980 8266 16992
rect 8680 16980 8708 17011
rect 8260 16952 8708 16980
rect 8260 16940 8266 16952
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 10229 16983 10287 16989
rect 10229 16980 10241 16983
rect 10192 16952 10241 16980
rect 10192 16940 10198 16952
rect 10229 16949 10241 16952
rect 10275 16949 10287 16983
rect 10796 16980 10824 17020
rect 10965 17017 10977 17051
rect 11011 17017 11023 17051
rect 10965 17011 11023 17017
rect 10980 16980 11008 17011
rect 12342 17008 12348 17060
rect 12400 17048 12406 17060
rect 12529 17051 12587 17057
rect 12529 17048 12541 17051
rect 12400 17020 12541 17048
rect 12400 17008 12406 17020
rect 12529 17017 12541 17020
rect 12575 17017 12587 17051
rect 12529 17011 12587 17017
rect 12621 17051 12679 17057
rect 12621 17017 12633 17051
rect 12667 17017 12679 17051
rect 12621 17011 12679 17017
rect 11054 16980 11060 16992
rect 10796 16952 11060 16980
rect 10229 16943 10287 16949
rect 11054 16940 11060 16952
rect 11112 16940 11118 16992
rect 11882 16980 11888 16992
rect 11843 16952 11888 16980
rect 11882 16940 11888 16952
rect 11940 16940 11946 16992
rect 12253 16983 12311 16989
rect 12253 16949 12265 16983
rect 12299 16980 12311 16983
rect 12636 16980 12664 17011
rect 12802 16980 12808 16992
rect 12299 16952 12808 16980
rect 12299 16949 12311 16952
rect 12253 16943 12311 16949
rect 12802 16940 12808 16952
rect 12860 16940 12866 16992
rect 13538 16940 13544 16992
rect 13596 16980 13602 16992
rect 13648 16989 13676 17156
rect 17310 17144 17316 17156
rect 17368 17144 17374 17196
rect 18417 17187 18475 17193
rect 18417 17153 18429 17187
rect 18463 17184 18475 17187
rect 19444 17184 19472 17280
rect 18463 17156 19472 17184
rect 18463 17153 18475 17156
rect 18417 17147 18475 17153
rect 14734 17116 14740 17128
rect 14695 17088 14740 17116
rect 14734 17076 14740 17088
rect 14792 17076 14798 17128
rect 16552 17119 16610 17125
rect 16552 17085 16564 17119
rect 16598 17116 16610 17119
rect 16758 17116 16764 17128
rect 16598 17088 16764 17116
rect 16598 17085 16610 17088
rect 16552 17079 16610 17085
rect 16758 17076 16764 17088
rect 16816 17076 16822 17128
rect 19956 17119 20014 17125
rect 19956 17085 19968 17119
rect 20002 17116 20014 17119
rect 20968 17119 21026 17125
rect 20002 17088 20392 17116
rect 20002 17085 20014 17088
rect 19956 17079 20014 17085
rect 14550 17008 14556 17060
rect 14608 17048 14614 17060
rect 14645 17051 14703 17057
rect 14645 17048 14657 17051
rect 14608 17020 14657 17048
rect 14608 17008 14614 17020
rect 14645 17017 14657 17020
rect 14691 17048 14703 17051
rect 15099 17051 15157 17057
rect 15099 17048 15111 17051
rect 14691 17020 15111 17048
rect 14691 17017 14703 17020
rect 14645 17011 14703 17017
rect 15099 17017 15111 17020
rect 15145 17048 15157 17051
rect 16022 17048 16028 17060
rect 15145 17020 16028 17048
rect 15145 17017 15157 17020
rect 15099 17011 15157 17017
rect 16022 17008 16028 17020
rect 16080 17048 16086 17060
rect 18046 17048 18052 17060
rect 16080 17020 18052 17048
rect 16080 17008 16086 17020
rect 18046 17008 18052 17020
rect 18104 17008 18110 17060
rect 18506 17048 18512 17060
rect 18467 17020 18512 17048
rect 18506 17008 18512 17020
rect 18564 17008 18570 17060
rect 20364 16992 20392 17088
rect 20968 17085 20980 17119
rect 21014 17116 21026 17119
rect 21358 17116 21364 17128
rect 21014 17088 21364 17116
rect 21014 17085 21026 17088
rect 20968 17079 21026 17085
rect 21358 17076 21364 17088
rect 21416 17116 21422 17128
rect 21729 17119 21787 17125
rect 21729 17116 21741 17119
rect 21416 17088 21741 17116
rect 21416 17076 21422 17088
rect 21729 17085 21741 17088
rect 21775 17085 21787 17119
rect 21729 17079 21787 17085
rect 24648 17119 24706 17125
rect 24648 17085 24660 17119
rect 24694 17116 24706 17119
rect 25130 17116 25136 17128
rect 24694 17088 25136 17116
rect 24694 17085 24706 17088
rect 24648 17079 24706 17085
rect 25130 17076 25136 17088
rect 25188 17076 25194 17128
rect 13633 16983 13691 16989
rect 13633 16980 13645 16983
rect 13596 16952 13645 16980
rect 13596 16940 13602 16952
rect 13633 16949 13645 16952
rect 13679 16949 13691 16983
rect 14090 16980 14096 16992
rect 14051 16952 14096 16980
rect 13633 16943 13691 16949
rect 14090 16940 14096 16952
rect 14148 16940 14154 16992
rect 15657 16983 15715 16989
rect 15657 16949 15669 16983
rect 15703 16980 15715 16983
rect 15838 16980 15844 16992
rect 15703 16952 15844 16980
rect 15703 16949 15715 16952
rect 15657 16943 15715 16949
rect 15838 16940 15844 16952
rect 15896 16940 15902 16992
rect 16623 16983 16681 16989
rect 16623 16949 16635 16983
rect 16669 16980 16681 16983
rect 16850 16980 16856 16992
rect 16669 16952 16856 16980
rect 16669 16949 16681 16952
rect 16623 16943 16681 16949
rect 16850 16940 16856 16952
rect 16908 16940 16914 16992
rect 20346 16980 20352 16992
rect 20307 16952 20352 16980
rect 20346 16940 20352 16952
rect 20404 16940 20410 16992
rect 22646 16940 22652 16992
rect 22704 16980 22710 16992
rect 24719 16983 24777 16989
rect 24719 16980 24731 16983
rect 22704 16952 24731 16980
rect 22704 16940 22710 16952
rect 24719 16949 24731 16952
rect 24765 16949 24777 16983
rect 24719 16943 24777 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1394 16736 1400 16788
rect 1452 16776 1458 16788
rect 1535 16779 1593 16785
rect 1535 16776 1547 16779
rect 1452 16748 1547 16776
rect 1452 16736 1458 16748
rect 1535 16745 1547 16748
rect 1581 16745 1593 16779
rect 3418 16776 3424 16788
rect 3379 16748 3424 16776
rect 1535 16739 1593 16745
rect 3418 16736 3424 16748
rect 3476 16776 3482 16788
rect 5166 16776 5172 16788
rect 3476 16748 5172 16776
rect 3476 16736 3482 16748
rect 5166 16736 5172 16748
rect 5224 16736 5230 16788
rect 6457 16779 6515 16785
rect 6457 16745 6469 16779
rect 6503 16776 6515 16779
rect 6730 16776 6736 16788
rect 6503 16748 6736 16776
rect 6503 16745 6515 16748
rect 6457 16739 6515 16745
rect 6730 16736 6736 16748
rect 6788 16776 6794 16788
rect 6917 16779 6975 16785
rect 6917 16776 6929 16779
rect 6788 16748 6929 16776
rect 6788 16736 6794 16748
rect 6917 16745 6929 16748
rect 6963 16745 6975 16779
rect 7466 16776 7472 16788
rect 7427 16748 7472 16776
rect 6917 16739 6975 16745
rect 7466 16736 7472 16748
rect 7524 16736 7530 16788
rect 11054 16776 11060 16788
rect 11015 16748 11060 16776
rect 11054 16736 11060 16748
rect 11112 16736 11118 16788
rect 12802 16776 12808 16788
rect 12763 16748 12808 16776
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 16758 16776 16764 16788
rect 16132 16748 16764 16776
rect 2317 16711 2375 16717
rect 2317 16677 2329 16711
rect 2363 16708 2375 16711
rect 2406 16708 2412 16720
rect 2363 16680 2412 16708
rect 2363 16677 2375 16680
rect 2317 16671 2375 16677
rect 2406 16668 2412 16680
rect 2464 16668 2470 16720
rect 2774 16708 2780 16720
rect 2571 16680 2780 16708
rect 1464 16643 1522 16649
rect 1464 16609 1476 16643
rect 1510 16640 1522 16643
rect 2222 16640 2228 16652
rect 1510 16612 2228 16640
rect 1510 16609 1522 16612
rect 1464 16603 1522 16609
rect 2222 16600 2228 16612
rect 2280 16600 2286 16652
rect 2571 16649 2599 16680
rect 2774 16668 2780 16680
rect 2832 16708 2838 16720
rect 3789 16711 3847 16717
rect 3789 16708 3801 16711
rect 2832 16680 3801 16708
rect 2832 16668 2838 16680
rect 3789 16677 3801 16680
rect 3835 16708 3847 16711
rect 3878 16708 3884 16720
rect 3835 16680 3884 16708
rect 3835 16677 3847 16680
rect 3789 16671 3847 16677
rect 3878 16668 3884 16680
rect 3936 16668 3942 16720
rect 4525 16711 4583 16717
rect 4525 16677 4537 16711
rect 4571 16708 4583 16711
rect 10499 16711 10557 16717
rect 4571 16680 5488 16708
rect 4571 16677 4583 16680
rect 4525 16671 4583 16677
rect 5460 16652 5488 16680
rect 10499 16677 10511 16711
rect 10545 16708 10557 16711
rect 11698 16708 11704 16720
rect 10545 16680 11704 16708
rect 10545 16677 10557 16680
rect 10499 16671 10557 16677
rect 11698 16668 11704 16680
rect 11756 16708 11762 16720
rect 12207 16711 12265 16717
rect 12207 16708 12219 16711
rect 11756 16680 12219 16708
rect 11756 16668 11762 16680
rect 12207 16677 12219 16680
rect 12253 16677 12265 16711
rect 12207 16671 12265 16677
rect 12342 16668 12348 16720
rect 12400 16708 12406 16720
rect 13081 16711 13139 16717
rect 13081 16708 13093 16711
rect 12400 16680 13093 16708
rect 12400 16668 12406 16680
rect 13081 16677 13093 16680
rect 13127 16677 13139 16711
rect 13081 16671 13139 16677
rect 14369 16711 14427 16717
rect 14369 16677 14381 16711
rect 14415 16708 14427 16711
rect 14734 16708 14740 16720
rect 14415 16680 14740 16708
rect 14415 16677 14427 16680
rect 14369 16671 14427 16677
rect 14734 16668 14740 16680
rect 14792 16668 14798 16720
rect 15565 16711 15623 16717
rect 15565 16677 15577 16711
rect 15611 16708 15623 16711
rect 15838 16708 15844 16720
rect 15611 16680 15844 16708
rect 15611 16677 15623 16680
rect 15565 16671 15623 16677
rect 15838 16668 15844 16680
rect 15896 16668 15902 16720
rect 16132 16717 16160 16748
rect 16758 16736 16764 16748
rect 16816 16736 16822 16788
rect 18506 16736 18512 16788
rect 18564 16776 18570 16788
rect 18693 16779 18751 16785
rect 18693 16776 18705 16779
rect 18564 16748 18705 16776
rect 18564 16736 18570 16748
rect 18693 16745 18705 16748
rect 18739 16745 18751 16779
rect 18966 16776 18972 16788
rect 18927 16748 18972 16776
rect 18693 16739 18751 16745
rect 18966 16736 18972 16748
rect 19024 16736 19030 16788
rect 24762 16776 24768 16788
rect 24723 16748 24768 16776
rect 24762 16736 24768 16748
rect 24820 16736 24826 16788
rect 16117 16711 16175 16717
rect 16117 16677 16129 16711
rect 16163 16677 16175 16711
rect 16117 16671 16175 16677
rect 18049 16711 18107 16717
rect 18049 16677 18061 16711
rect 18095 16708 18107 16711
rect 18138 16708 18144 16720
rect 18095 16680 18144 16708
rect 18095 16677 18107 16680
rect 18049 16671 18107 16677
rect 18138 16668 18144 16680
rect 18196 16668 18202 16720
rect 2556 16643 2614 16649
rect 2556 16609 2568 16643
rect 2602 16609 2614 16643
rect 2556 16603 2614 16609
rect 4430 16600 4436 16652
rect 4488 16640 4494 16652
rect 4617 16643 4675 16649
rect 4617 16640 4629 16643
rect 4488 16612 4629 16640
rect 4488 16600 4494 16612
rect 4617 16609 4629 16612
rect 4663 16609 4675 16643
rect 5166 16640 5172 16652
rect 5127 16612 5172 16640
rect 4617 16603 4675 16609
rect 5166 16600 5172 16612
rect 5224 16600 5230 16652
rect 5442 16640 5448 16652
rect 5403 16612 5448 16640
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 5997 16643 6055 16649
rect 5997 16609 6009 16643
rect 6043 16640 6055 16643
rect 6178 16640 6184 16652
rect 6043 16612 6184 16640
rect 6043 16609 6055 16612
rect 5997 16603 6055 16609
rect 6178 16600 6184 16612
rect 6236 16600 6242 16652
rect 7926 16640 7932 16652
rect 7887 16612 7932 16640
rect 7926 16600 7932 16612
rect 7984 16600 7990 16652
rect 13630 16640 13636 16652
rect 13591 16612 13636 16640
rect 13630 16600 13636 16612
rect 13688 16600 13694 16652
rect 14185 16643 14243 16649
rect 14185 16609 14197 16643
rect 14231 16609 14243 16643
rect 17310 16640 17316 16652
rect 17271 16612 17316 16640
rect 14185 16603 14243 16609
rect 2777 16575 2835 16581
rect 2777 16541 2789 16575
rect 2823 16572 2835 16575
rect 3510 16572 3516 16584
rect 2823 16544 3516 16572
rect 2823 16541 2835 16544
rect 2777 16535 2835 16541
rect 3510 16532 3516 16544
rect 3568 16532 3574 16584
rect 6086 16572 6092 16584
rect 6047 16544 6092 16572
rect 6086 16532 6092 16544
rect 6144 16532 6150 16584
rect 9766 16532 9772 16584
rect 9824 16572 9830 16584
rect 10137 16575 10195 16581
rect 10137 16572 10149 16575
rect 9824 16544 10149 16572
rect 9824 16532 9830 16544
rect 10137 16541 10149 16544
rect 10183 16541 10195 16575
rect 10137 16535 10195 16541
rect 11885 16575 11943 16581
rect 11885 16541 11897 16575
rect 11931 16541 11943 16575
rect 11885 16535 11943 16541
rect 2682 16504 2688 16516
rect 2643 16476 2688 16504
rect 2682 16464 2688 16476
rect 2740 16464 2746 16516
rect 1949 16439 2007 16445
rect 1949 16405 1961 16439
rect 1995 16436 2007 16439
rect 2406 16436 2412 16448
rect 1995 16408 2412 16436
rect 1995 16405 2007 16408
rect 1949 16399 2007 16405
rect 2406 16396 2412 16408
rect 2464 16396 2470 16448
rect 3050 16436 3056 16448
rect 3011 16408 3056 16436
rect 3050 16396 3056 16408
rect 3108 16396 3114 16448
rect 8294 16436 8300 16448
rect 8255 16408 8300 16436
rect 8294 16396 8300 16408
rect 8352 16396 8358 16448
rect 8478 16396 8484 16448
rect 8536 16436 8542 16448
rect 8849 16439 8907 16445
rect 8849 16436 8861 16439
rect 8536 16408 8861 16436
rect 8536 16396 8542 16408
rect 8849 16405 8861 16408
rect 8895 16405 8907 16439
rect 8849 16399 8907 16405
rect 11793 16439 11851 16445
rect 11793 16405 11805 16439
rect 11839 16436 11851 16439
rect 11900 16436 11928 16535
rect 14090 16464 14096 16516
rect 14148 16504 14154 16516
rect 14200 16504 14228 16603
rect 17310 16600 17316 16612
rect 17368 16600 17374 16652
rect 17862 16640 17868 16652
rect 17823 16612 17868 16640
rect 17862 16600 17868 16612
rect 17920 16600 17926 16652
rect 18874 16640 18880 16652
rect 18835 16612 18880 16640
rect 18874 16600 18880 16612
rect 18932 16600 18938 16652
rect 19429 16643 19487 16649
rect 19429 16609 19441 16643
rect 19475 16640 19487 16643
rect 19702 16640 19708 16652
rect 19475 16612 19708 16640
rect 19475 16609 19487 16612
rect 19429 16603 19487 16609
rect 15473 16575 15531 16581
rect 15473 16541 15485 16575
rect 15519 16572 15531 16575
rect 15654 16572 15660 16584
rect 15519 16544 15660 16572
rect 15519 16541 15531 16544
rect 15473 16535 15531 16541
rect 15654 16532 15660 16544
rect 15712 16572 15718 16584
rect 16393 16575 16451 16581
rect 16393 16572 16405 16575
rect 15712 16544 16405 16572
rect 15712 16532 15718 16544
rect 16393 16541 16405 16544
rect 16439 16541 16451 16575
rect 16393 16535 16451 16541
rect 19444 16504 19472 16603
rect 19702 16600 19708 16612
rect 19760 16600 19766 16652
rect 20901 16643 20959 16649
rect 20901 16609 20913 16643
rect 20947 16640 20959 16643
rect 21266 16640 21272 16652
rect 20947 16612 21272 16640
rect 20947 16609 20959 16612
rect 20901 16603 20959 16609
rect 21266 16600 21272 16612
rect 21324 16600 21330 16652
rect 21818 16600 21824 16652
rect 21876 16640 21882 16652
rect 21948 16643 22006 16649
rect 21948 16640 21960 16643
rect 21876 16612 21960 16640
rect 21876 16600 21882 16612
rect 21948 16609 21960 16612
rect 21994 16609 22006 16643
rect 21948 16603 22006 16609
rect 24581 16643 24639 16649
rect 24581 16609 24593 16643
rect 24627 16640 24639 16643
rect 24670 16640 24676 16652
rect 24627 16612 24676 16640
rect 24627 16609 24639 16612
rect 24581 16603 24639 16609
rect 24670 16600 24676 16612
rect 24728 16600 24734 16652
rect 14148 16476 19472 16504
rect 14148 16464 14154 16476
rect 12526 16436 12532 16448
rect 11839 16408 12532 16436
rect 11839 16405 11851 16408
rect 11793 16399 11851 16405
rect 12526 16396 12532 16408
rect 12584 16396 12590 16448
rect 17862 16396 17868 16448
rect 17920 16436 17926 16448
rect 18325 16439 18383 16445
rect 18325 16436 18337 16439
rect 17920 16408 18337 16436
rect 17920 16396 17926 16408
rect 18325 16405 18337 16408
rect 18371 16405 18383 16439
rect 18325 16399 18383 16405
rect 19702 16396 19708 16448
rect 19760 16436 19766 16448
rect 21085 16439 21143 16445
rect 21085 16436 21097 16439
rect 19760 16408 21097 16436
rect 19760 16396 19766 16408
rect 21085 16405 21097 16408
rect 21131 16405 21143 16439
rect 21085 16399 21143 16405
rect 21910 16396 21916 16448
rect 21968 16436 21974 16448
rect 22051 16439 22109 16445
rect 22051 16436 22063 16439
rect 21968 16408 22063 16436
rect 21968 16396 21974 16408
rect 22051 16405 22063 16408
rect 22097 16405 22109 16439
rect 22051 16399 22109 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2682 16192 2688 16244
rect 2740 16232 2746 16244
rect 3145 16235 3203 16241
rect 3145 16232 3157 16235
rect 2740 16204 3157 16232
rect 2740 16192 2746 16204
rect 3145 16201 3157 16204
rect 3191 16232 3203 16235
rect 3234 16232 3240 16244
rect 3191 16204 3240 16232
rect 3191 16201 3203 16204
rect 3145 16195 3203 16201
rect 3234 16192 3240 16204
rect 3292 16192 3298 16244
rect 3510 16232 3516 16244
rect 3471 16204 3516 16232
rect 3510 16192 3516 16204
rect 3568 16192 3574 16244
rect 3973 16235 4031 16241
rect 3973 16201 3985 16235
rect 4019 16232 4031 16235
rect 4341 16235 4399 16241
rect 4341 16232 4353 16235
rect 4019 16204 4353 16232
rect 4019 16201 4031 16204
rect 3973 16195 4031 16201
rect 4341 16201 4353 16204
rect 4387 16232 4399 16235
rect 4430 16232 4436 16244
rect 4387 16204 4436 16232
rect 4387 16201 4399 16204
rect 4341 16195 4399 16201
rect 4430 16192 4436 16204
rect 4488 16192 4494 16244
rect 7745 16235 7803 16241
rect 7745 16201 7757 16235
rect 7791 16232 7803 16235
rect 7926 16232 7932 16244
rect 7791 16204 7932 16232
rect 7791 16201 7803 16204
rect 7745 16195 7803 16201
rect 7926 16192 7932 16204
rect 7984 16192 7990 16244
rect 8294 16192 8300 16244
rect 8352 16232 8358 16244
rect 8389 16235 8447 16241
rect 8389 16232 8401 16235
rect 8352 16204 8401 16232
rect 8352 16192 8358 16204
rect 8389 16201 8401 16204
rect 8435 16201 8447 16235
rect 10229 16235 10287 16241
rect 10229 16232 10241 16235
rect 8389 16195 8447 16201
rect 9646 16204 10241 16232
rect 3528 16164 3556 16192
rect 4246 16164 4252 16176
rect 3528 16136 4252 16164
rect 4246 16124 4252 16136
rect 4304 16124 4310 16176
rect 5534 16096 5540 16108
rect 2332 16068 5540 16096
rect 1946 16028 1952 16040
rect 1907 16000 1952 16028
rect 1946 15988 1952 16000
rect 2004 15988 2010 16040
rect 2332 16037 2360 16068
rect 5534 16056 5540 16068
rect 5592 16056 5598 16108
rect 6086 16056 6092 16108
rect 6144 16096 6150 16108
rect 6825 16099 6883 16105
rect 6825 16096 6837 16099
rect 6144 16068 6837 16096
rect 6144 16056 6150 16068
rect 6825 16065 6837 16068
rect 6871 16096 6883 16099
rect 7282 16096 7288 16108
rect 6871 16068 7288 16096
rect 6871 16065 6883 16068
rect 6825 16059 6883 16065
rect 7282 16056 7288 16068
rect 7340 16056 7346 16108
rect 7742 16056 7748 16108
rect 7800 16096 7806 16108
rect 9646 16096 9674 16204
rect 10229 16201 10241 16204
rect 10275 16232 10287 16235
rect 11698 16232 11704 16244
rect 10275 16204 11704 16232
rect 10275 16201 10287 16204
rect 10229 16195 10287 16201
rect 11698 16192 11704 16204
rect 11756 16232 11762 16244
rect 11885 16235 11943 16241
rect 11885 16232 11897 16235
rect 11756 16204 11897 16232
rect 11756 16192 11762 16204
rect 11885 16201 11897 16204
rect 11931 16201 11943 16235
rect 14090 16232 14096 16244
rect 14051 16204 14096 16232
rect 11885 16195 11943 16201
rect 14090 16192 14096 16204
rect 14148 16192 14154 16244
rect 15838 16232 15844 16244
rect 15799 16204 15844 16232
rect 15838 16192 15844 16204
rect 15896 16192 15902 16244
rect 17497 16235 17555 16241
rect 17497 16201 17509 16235
rect 17543 16232 17555 16235
rect 17770 16232 17776 16244
rect 17543 16204 17776 16232
rect 17543 16201 17555 16204
rect 17497 16195 17555 16201
rect 17770 16192 17776 16204
rect 17828 16192 17834 16244
rect 17865 16235 17923 16241
rect 17865 16201 17877 16235
rect 17911 16232 17923 16235
rect 18046 16232 18052 16244
rect 17911 16204 18052 16232
rect 17911 16201 17923 16204
rect 17865 16195 17923 16201
rect 18046 16192 18052 16204
rect 18104 16192 18110 16244
rect 18874 16192 18880 16244
rect 18932 16232 18938 16244
rect 19245 16235 19303 16241
rect 19245 16232 19257 16235
rect 18932 16204 19257 16232
rect 18932 16192 18938 16204
rect 19245 16201 19257 16204
rect 19291 16201 19303 16235
rect 19702 16232 19708 16244
rect 19663 16204 19708 16232
rect 19245 16195 19303 16201
rect 19702 16192 19708 16204
rect 19760 16192 19766 16244
rect 21818 16192 21824 16244
rect 21876 16232 21882 16244
rect 22281 16235 22339 16241
rect 22281 16232 22293 16235
rect 21876 16204 22293 16232
rect 21876 16192 21882 16204
rect 22281 16201 22293 16204
rect 22327 16232 22339 16235
rect 23658 16232 23664 16244
rect 22327 16204 23664 16232
rect 22327 16201 22339 16204
rect 22281 16195 22339 16201
rect 23658 16192 23664 16204
rect 23716 16192 23722 16244
rect 23799 16235 23857 16241
rect 23799 16201 23811 16235
rect 23845 16232 23857 16235
rect 24670 16232 24676 16244
rect 23845 16204 24676 16232
rect 23845 16201 23857 16204
rect 23799 16195 23857 16201
rect 24670 16192 24676 16204
rect 24728 16192 24734 16244
rect 13538 16164 13544 16176
rect 7800 16068 9674 16096
rect 10796 16136 13544 16164
rect 7800 16056 7806 16068
rect 2317 16031 2375 16037
rect 2317 15997 2329 16031
rect 2363 15997 2375 16031
rect 2317 15991 2375 15997
rect 2406 15988 2412 16040
rect 2464 16028 2470 16040
rect 2866 16028 2872 16040
rect 2464 16000 2509 16028
rect 2827 16000 2872 16028
rect 2464 15988 2470 16000
rect 2866 15988 2872 16000
rect 2924 16028 2930 16040
rect 3510 16028 3516 16040
rect 2924 16000 3516 16028
rect 2924 15988 2930 16000
rect 3510 15988 3516 16000
rect 3568 15988 3574 16040
rect 4430 16028 4436 16040
rect 4391 16000 4436 16028
rect 4430 15988 4436 16000
rect 4488 15988 4494 16040
rect 5166 16028 5172 16040
rect 5127 16000 5172 16028
rect 5166 15988 5172 16000
rect 5224 15988 5230 16040
rect 5442 16028 5448 16040
rect 5403 16000 5448 16028
rect 5442 15988 5448 16000
rect 5500 15988 5506 16040
rect 5813 16031 5871 16037
rect 5813 15997 5825 16031
rect 5859 16028 5871 16031
rect 5994 16028 6000 16040
rect 5859 16000 6000 16028
rect 5859 15997 5871 16000
rect 5813 15991 5871 15997
rect 5994 15988 6000 16000
rect 6052 16028 6058 16040
rect 10796 16037 10824 16136
rect 13538 16124 13544 16136
rect 13596 16124 13602 16176
rect 15473 16167 15531 16173
rect 15473 16133 15485 16167
rect 15519 16164 15531 16167
rect 15654 16164 15660 16176
rect 15519 16136 15660 16164
rect 15519 16133 15531 16136
rect 15473 16127 15531 16133
rect 15654 16124 15660 16136
rect 15712 16124 15718 16176
rect 15746 16124 15752 16176
rect 15804 16164 15810 16176
rect 21959 16167 22017 16173
rect 21959 16164 21971 16167
rect 15804 16136 21971 16164
rect 15804 16124 15810 16136
rect 21959 16133 21971 16136
rect 22005 16133 22017 16167
rect 21959 16127 22017 16133
rect 11330 16096 11336 16108
rect 11291 16068 11336 16096
rect 11330 16056 11336 16068
rect 11388 16056 11394 16108
rect 14737 16099 14795 16105
rect 11440 16068 12940 16096
rect 8021 16031 8079 16037
rect 8021 16028 8033 16031
rect 6052 16000 8033 16028
rect 6052 15988 6058 16000
rect 8021 15997 8033 16000
rect 8067 15997 8079 16031
rect 8021 15991 8079 15997
rect 10689 16031 10747 16037
rect 10689 15997 10701 16031
rect 10735 16028 10747 16031
rect 10781 16031 10839 16037
rect 10781 16028 10793 16031
rect 10735 16000 10793 16028
rect 10735 15997 10747 16000
rect 10689 15991 10747 15997
rect 10781 15997 10793 16000
rect 10827 15997 10839 16031
rect 10781 15991 10839 15997
rect 10870 15988 10876 16040
rect 10928 16028 10934 16040
rect 11241 16031 11299 16037
rect 11241 16028 11253 16031
rect 10928 16000 11253 16028
rect 10928 15988 10934 16000
rect 11241 15997 11253 16000
rect 11287 16028 11299 16031
rect 11440 16028 11468 16068
rect 12618 16028 12624 16040
rect 11287 16000 11468 16028
rect 12579 16000 12624 16028
rect 11287 15997 11299 16000
rect 11241 15991 11299 15997
rect 12618 15988 12624 16000
rect 12676 15988 12682 16040
rect 12912 16037 12940 16068
rect 14737 16065 14749 16099
rect 14783 16096 14795 16099
rect 15010 16096 15016 16108
rect 14783 16068 15016 16096
rect 14783 16065 14795 16068
rect 14737 16059 14795 16065
rect 15010 16056 15016 16068
rect 15068 16096 15074 16108
rect 15562 16096 15568 16108
rect 15068 16068 15568 16096
rect 15068 16056 15074 16068
rect 15562 16056 15568 16068
rect 15620 16056 15626 16108
rect 20349 16099 20407 16105
rect 20349 16065 20361 16099
rect 20395 16096 20407 16099
rect 20438 16096 20444 16108
rect 20395 16068 20444 16096
rect 20395 16065 20407 16068
rect 20349 16059 20407 16065
rect 20438 16056 20444 16068
rect 20496 16056 20502 16108
rect 20622 16096 20628 16108
rect 20583 16068 20628 16096
rect 20622 16056 20628 16068
rect 20680 16056 20686 16108
rect 12897 16031 12955 16037
rect 12897 15997 12909 16031
rect 12943 16028 12955 16031
rect 12986 16028 12992 16040
rect 12943 16000 12992 16028
rect 12943 15997 12955 16000
rect 12897 15991 12955 15997
rect 12986 15988 12992 16000
rect 13044 15988 13050 16040
rect 15930 15988 15936 16040
rect 15988 16028 15994 16040
rect 16301 16031 16359 16037
rect 16301 16028 16313 16031
rect 15988 16000 16313 16028
rect 15988 15988 15994 16000
rect 16301 15997 16313 16000
rect 16347 16028 16359 16031
rect 16393 16031 16451 16037
rect 16393 16028 16405 16031
rect 16347 16000 16405 16028
rect 16347 15997 16359 16000
rect 16301 15991 16359 15997
rect 16393 15997 16405 16000
rect 16439 15997 16451 16031
rect 16393 15991 16451 15997
rect 5905 15963 5963 15969
rect 5905 15929 5917 15963
rect 5951 15960 5963 15963
rect 6086 15960 6092 15972
rect 5951 15932 6092 15960
rect 5951 15929 5963 15932
rect 5905 15923 5963 15929
rect 6086 15920 6092 15932
rect 6144 15920 6150 15972
rect 6638 15960 6644 15972
rect 6551 15932 6644 15960
rect 6638 15920 6644 15932
rect 6696 15960 6702 15972
rect 7187 15963 7245 15969
rect 7187 15960 7199 15963
rect 6696 15932 7199 15960
rect 6696 15920 6702 15932
rect 7187 15929 7199 15932
rect 7233 15960 7245 15963
rect 7742 15960 7748 15972
rect 7233 15932 7748 15960
rect 7233 15929 7245 15932
rect 7187 15923 7245 15929
rect 7742 15920 7748 15932
rect 7800 15920 7806 15972
rect 8478 15920 8484 15972
rect 8536 15960 8542 15972
rect 8665 15963 8723 15969
rect 8665 15960 8677 15963
rect 8536 15932 8677 15960
rect 8536 15920 8542 15932
rect 8665 15929 8677 15932
rect 8711 15929 8723 15963
rect 8665 15923 8723 15929
rect 8757 15963 8815 15969
rect 8757 15929 8769 15963
rect 8803 15929 8815 15963
rect 9306 15960 9312 15972
rect 9267 15932 9312 15960
rect 8757 15923 8815 15929
rect 2314 15852 2320 15904
rect 2372 15892 2378 15904
rect 3878 15892 3884 15904
rect 2372 15864 3884 15892
rect 2372 15852 2378 15864
rect 3878 15852 3884 15864
rect 3936 15852 3942 15904
rect 5994 15852 6000 15904
rect 6052 15892 6058 15904
rect 6178 15892 6184 15904
rect 6052 15864 6184 15892
rect 6052 15852 6058 15864
rect 6178 15852 6184 15864
rect 6236 15852 6242 15904
rect 8294 15852 8300 15904
rect 8352 15892 8358 15904
rect 8772 15892 8800 15923
rect 9306 15920 9312 15932
rect 9364 15920 9370 15972
rect 12636 15960 12664 15988
rect 13630 15960 13636 15972
rect 12636 15932 13636 15960
rect 13630 15920 13636 15932
rect 13688 15920 13694 15972
rect 14921 15963 14979 15969
rect 14921 15929 14933 15963
rect 14967 15929 14979 15963
rect 14921 15923 14979 15929
rect 9766 15892 9772 15904
rect 8352 15864 8800 15892
rect 9727 15864 9772 15892
rect 8352 15852 8358 15864
rect 9766 15852 9772 15864
rect 9824 15852 9830 15904
rect 12526 15892 12532 15904
rect 12487 15864 12532 15892
rect 12526 15852 12532 15864
rect 12584 15852 12590 15904
rect 14826 15852 14832 15904
rect 14884 15892 14890 15904
rect 14936 15892 14964 15923
rect 15010 15920 15016 15972
rect 15068 15960 15074 15972
rect 16408 15960 16436 15991
rect 16482 15988 16488 16040
rect 16540 16028 16546 16040
rect 16853 16031 16911 16037
rect 16853 16028 16865 16031
rect 16540 16000 16865 16028
rect 16540 15988 16546 16000
rect 16853 15997 16865 16000
rect 16899 15997 16911 16031
rect 16853 15991 16911 15997
rect 17862 15988 17868 16040
rect 17920 16028 17926 16040
rect 18049 16031 18107 16037
rect 18049 16028 18061 16031
rect 17920 16000 18061 16028
rect 17920 15988 17926 16000
rect 18049 15997 18061 16000
rect 18095 15997 18107 16031
rect 18049 15991 18107 15997
rect 21726 15988 21732 16040
rect 21784 16028 21790 16040
rect 21856 16031 21914 16037
rect 21856 16028 21868 16031
rect 21784 16000 21868 16028
rect 21784 15988 21790 16000
rect 21856 15997 21868 16000
rect 21902 16028 21914 16031
rect 22649 16031 22707 16037
rect 22649 16028 22661 16031
rect 21902 16000 22661 16028
rect 21902 15997 21914 16000
rect 21856 15991 21914 15997
rect 22649 15997 22661 16000
rect 22695 15997 22707 16031
rect 22649 15991 22707 15997
rect 23728 16031 23786 16037
rect 23728 15997 23740 16031
rect 23774 16028 23786 16031
rect 24118 16028 24124 16040
rect 23774 16000 24124 16028
rect 23774 15997 23786 16000
rect 23728 15991 23786 15997
rect 24118 15988 24124 16000
rect 24176 15988 24182 16040
rect 16758 15960 16764 15972
rect 15068 15932 15113 15960
rect 16408 15932 16764 15960
rect 15068 15920 15074 15932
rect 16758 15920 16764 15932
rect 16816 15920 16822 15972
rect 17126 15960 17132 15972
rect 17087 15932 17132 15960
rect 17126 15920 17132 15932
rect 17184 15920 17190 15972
rect 18138 15920 18144 15972
rect 18196 15960 18202 15972
rect 18370 15963 18428 15969
rect 18370 15960 18382 15963
rect 18196 15932 18382 15960
rect 18196 15920 18202 15932
rect 18370 15929 18382 15932
rect 18416 15929 18428 15963
rect 20073 15963 20131 15969
rect 20073 15960 20085 15963
rect 18370 15923 18428 15929
rect 18984 15932 20085 15960
rect 14884 15864 14964 15892
rect 14884 15852 14890 15864
rect 18874 15852 18880 15904
rect 18932 15892 18938 15904
rect 18984 15901 19012 15932
rect 20073 15929 20085 15932
rect 20119 15929 20131 15963
rect 20073 15923 20131 15929
rect 20441 15963 20499 15969
rect 20441 15929 20453 15963
rect 20487 15960 20499 15963
rect 21358 15960 21364 15972
rect 20487 15932 21364 15960
rect 20487 15929 20499 15932
rect 20441 15923 20499 15929
rect 18969 15895 19027 15901
rect 18969 15892 18981 15895
rect 18932 15864 18981 15892
rect 18932 15852 18938 15864
rect 18969 15861 18981 15864
rect 19015 15861 19027 15895
rect 20088 15892 20116 15923
rect 20456 15892 20484 15923
rect 21358 15920 21364 15932
rect 21416 15920 21422 15972
rect 21266 15892 21272 15904
rect 20088 15864 20484 15892
rect 21227 15864 21272 15892
rect 18969 15855 19027 15861
rect 21266 15852 21272 15864
rect 21324 15852 21330 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 2774 15648 2780 15700
rect 2832 15688 2838 15700
rect 3053 15691 3111 15697
rect 3053 15688 3065 15691
rect 2832 15660 3065 15688
rect 2832 15648 2838 15660
rect 3053 15657 3065 15660
rect 3099 15688 3111 15691
rect 3329 15691 3387 15697
rect 3329 15688 3341 15691
rect 3099 15660 3341 15688
rect 3099 15657 3111 15660
rect 3053 15651 3111 15657
rect 3329 15657 3341 15660
rect 3375 15657 3387 15691
rect 3329 15651 3387 15657
rect 3513 15691 3571 15697
rect 3513 15657 3525 15691
rect 3559 15688 3571 15691
rect 3694 15688 3700 15700
rect 3559 15660 3700 15688
rect 3559 15657 3571 15660
rect 3513 15651 3571 15657
rect 1765 15623 1823 15629
rect 1765 15589 1777 15623
rect 1811 15620 1823 15623
rect 1946 15620 1952 15632
rect 1811 15592 1952 15620
rect 1811 15589 1823 15592
rect 1765 15583 1823 15589
rect 1946 15580 1952 15592
rect 2004 15620 2010 15632
rect 2792 15620 2820 15648
rect 2004 15592 2820 15620
rect 2004 15580 2010 15592
rect 2056 15561 2084 15592
rect 2041 15555 2099 15561
rect 2041 15521 2053 15555
rect 2087 15521 2099 15555
rect 2314 15552 2320 15564
rect 2227 15524 2320 15552
rect 2041 15515 2099 15521
rect 2314 15512 2320 15524
rect 2372 15552 2378 15564
rect 3528 15552 3556 15651
rect 3694 15648 3700 15660
rect 3752 15648 3758 15700
rect 5442 15688 5448 15700
rect 5403 15660 5448 15688
rect 5442 15648 5448 15660
rect 5500 15648 5506 15700
rect 7282 15688 7288 15700
rect 7243 15660 7288 15688
rect 7282 15648 7288 15660
rect 7340 15648 7346 15700
rect 7926 15688 7932 15700
rect 7887 15660 7932 15688
rect 7926 15648 7932 15660
rect 7984 15688 7990 15700
rect 9766 15688 9772 15700
rect 7984 15660 8248 15688
rect 9727 15660 9772 15688
rect 7984 15648 7990 15660
rect 5166 15580 5172 15632
rect 5224 15620 5230 15632
rect 5350 15620 5356 15632
rect 5224 15592 5356 15620
rect 5224 15580 5230 15592
rect 5350 15580 5356 15592
rect 5408 15620 5414 15632
rect 5813 15623 5871 15629
rect 5813 15620 5825 15623
rect 5408 15592 5825 15620
rect 5408 15580 5414 15592
rect 5813 15589 5825 15592
rect 5859 15589 5871 15623
rect 5813 15583 5871 15589
rect 6451 15623 6509 15629
rect 6451 15589 6463 15623
rect 6497 15620 6509 15623
rect 6638 15620 6644 15632
rect 6497 15592 6644 15620
rect 6497 15589 6509 15592
rect 6451 15583 6509 15589
rect 6638 15580 6644 15592
rect 6696 15580 6702 15632
rect 8220 15629 8248 15660
rect 9766 15648 9772 15660
rect 9824 15648 9830 15700
rect 10778 15688 10784 15700
rect 10739 15660 10784 15688
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 11698 15688 11704 15700
rect 11659 15660 11704 15688
rect 11698 15648 11704 15660
rect 11756 15648 11762 15700
rect 11882 15648 11888 15700
rect 11940 15688 11946 15700
rect 12253 15691 12311 15697
rect 12253 15688 12265 15691
rect 11940 15660 12265 15688
rect 11940 15648 11946 15660
rect 12253 15657 12265 15660
rect 12299 15657 12311 15691
rect 12986 15688 12992 15700
rect 12947 15660 12992 15688
rect 12253 15651 12311 15657
rect 12986 15648 12992 15660
rect 13044 15648 13050 15700
rect 17310 15648 17316 15700
rect 17368 15688 17374 15700
rect 17405 15691 17463 15697
rect 17405 15688 17417 15691
rect 17368 15660 17417 15688
rect 17368 15648 17374 15660
rect 17405 15657 17417 15660
rect 17451 15688 17463 15691
rect 17678 15688 17684 15700
rect 17451 15660 17684 15688
rect 17451 15657 17463 15660
rect 17405 15651 17463 15657
rect 17678 15648 17684 15660
rect 17736 15648 17742 15700
rect 18969 15691 19027 15697
rect 18969 15657 18981 15691
rect 19015 15688 19027 15691
rect 20070 15688 20076 15700
rect 19015 15660 20076 15688
rect 19015 15657 19027 15660
rect 18969 15651 19027 15657
rect 20070 15648 20076 15660
rect 20128 15648 20134 15700
rect 20349 15691 20407 15697
rect 20349 15657 20361 15691
rect 20395 15688 20407 15691
rect 20438 15688 20444 15700
rect 20395 15660 20444 15688
rect 20395 15657 20407 15660
rect 20349 15651 20407 15657
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 21910 15688 21916 15700
rect 21871 15660 21916 15688
rect 21910 15648 21916 15660
rect 21968 15648 21974 15700
rect 24762 15688 24768 15700
rect 24723 15660 24768 15688
rect 24762 15648 24768 15660
rect 24820 15648 24826 15700
rect 8205 15623 8263 15629
rect 8205 15589 8217 15623
rect 8251 15589 8263 15623
rect 8205 15583 8263 15589
rect 8757 15623 8815 15629
rect 8757 15589 8769 15623
rect 8803 15620 8815 15623
rect 9306 15620 9312 15632
rect 8803 15592 9312 15620
rect 8803 15589 8815 15592
rect 8757 15583 8815 15589
rect 9306 15580 9312 15592
rect 9364 15580 9370 15632
rect 10686 15620 10692 15632
rect 9968 15592 10692 15620
rect 2372 15524 3556 15552
rect 3697 15555 3755 15561
rect 2372 15512 2378 15524
rect 3697 15521 3709 15555
rect 3743 15552 3755 15555
rect 4053 15555 4111 15561
rect 4053 15552 4065 15555
rect 3743 15524 4065 15552
rect 3743 15521 3755 15524
rect 3697 15515 3755 15521
rect 4053 15521 4065 15524
rect 4099 15521 4111 15555
rect 4053 15515 4111 15521
rect 4246 15512 4252 15564
rect 4304 15552 4310 15564
rect 9968 15561 9996 15592
rect 10686 15580 10692 15592
rect 10744 15580 10750 15632
rect 4341 15555 4399 15561
rect 4341 15552 4353 15555
rect 4304 15524 4353 15552
rect 4304 15512 4310 15524
rect 4341 15521 4353 15524
rect 4387 15521 4399 15555
rect 4341 15515 4399 15521
rect 9953 15555 10011 15561
rect 9953 15521 9965 15555
rect 9999 15521 10011 15555
rect 9953 15515 10011 15521
rect 10042 15512 10048 15564
rect 10100 15552 10106 15564
rect 10229 15555 10287 15561
rect 10229 15552 10241 15555
rect 10100 15524 10241 15552
rect 10100 15512 10106 15524
rect 10229 15521 10241 15524
rect 10275 15552 10287 15555
rect 10796 15552 10824 15648
rect 13817 15623 13875 15629
rect 13817 15589 13829 15623
rect 13863 15620 13875 15623
rect 14182 15620 14188 15632
rect 13863 15592 14188 15620
rect 13863 15589 13875 15592
rect 13817 15583 13875 15589
rect 14182 15580 14188 15592
rect 14240 15580 14246 15632
rect 15378 15580 15384 15632
rect 15436 15620 15442 15632
rect 15473 15623 15531 15629
rect 15473 15620 15485 15623
rect 15436 15592 15485 15620
rect 15436 15580 15442 15592
rect 15473 15589 15485 15592
rect 15519 15589 15531 15623
rect 15473 15583 15531 15589
rect 18138 15580 18144 15632
rect 18196 15620 18202 15632
rect 18370 15623 18428 15629
rect 18370 15620 18382 15623
rect 18196 15592 18382 15620
rect 18196 15580 18202 15592
rect 18370 15589 18382 15592
rect 18416 15589 18428 15623
rect 21082 15620 21088 15632
rect 21043 15592 21088 15620
rect 18370 15583 18428 15589
rect 21082 15580 21088 15592
rect 21140 15580 21146 15632
rect 21174 15580 21180 15632
rect 21232 15620 21238 15632
rect 22465 15623 22523 15629
rect 22465 15620 22477 15623
rect 21232 15592 22477 15620
rect 21232 15580 21238 15592
rect 22465 15589 22477 15592
rect 22511 15589 22523 15623
rect 22465 15583 22523 15589
rect 16850 15552 16856 15564
rect 10275 15524 10824 15552
rect 16811 15524 16856 15552
rect 10275 15521 10287 15524
rect 10229 15515 10287 15521
rect 16850 15512 16856 15524
rect 16908 15512 16914 15564
rect 17126 15512 17132 15564
rect 17184 15552 17190 15564
rect 17770 15552 17776 15564
rect 17184 15524 17776 15552
rect 17184 15512 17190 15524
rect 17770 15512 17776 15524
rect 17828 15552 17834 15564
rect 18049 15555 18107 15561
rect 18049 15552 18061 15555
rect 17828 15524 18061 15552
rect 17828 15512 17834 15524
rect 18049 15521 18061 15524
rect 18095 15521 18107 15555
rect 18049 15515 18107 15521
rect 19864 15555 19922 15561
rect 19864 15521 19876 15555
rect 19910 15552 19922 15555
rect 20162 15552 20168 15564
rect 19910 15524 20168 15552
rect 19910 15521 19922 15524
rect 19864 15515 19922 15521
rect 20162 15512 20168 15524
rect 20220 15512 20226 15564
rect 23658 15512 23664 15564
rect 23716 15552 23722 15564
rect 24210 15552 24216 15564
rect 23716 15524 24216 15552
rect 23716 15512 23722 15524
rect 24210 15512 24216 15524
rect 24268 15552 24274 15564
rect 24581 15555 24639 15561
rect 24581 15552 24593 15555
rect 24268 15524 24593 15552
rect 24268 15512 24274 15524
rect 24581 15521 24593 15524
rect 24627 15552 24639 15555
rect 24670 15552 24676 15564
rect 24627 15524 24676 15552
rect 24627 15521 24639 15524
rect 24581 15515 24639 15521
rect 24670 15512 24676 15524
rect 24728 15512 24734 15564
rect 2777 15487 2835 15493
rect 2777 15453 2789 15487
rect 2823 15484 2835 15487
rect 3142 15484 3148 15496
rect 2823 15456 3148 15484
rect 2823 15453 2835 15456
rect 2777 15447 2835 15453
rect 3142 15444 3148 15456
rect 3200 15444 3206 15496
rect 3234 15444 3240 15496
rect 3292 15484 3298 15496
rect 4157 15487 4215 15493
rect 4157 15484 4169 15487
rect 3292 15456 4169 15484
rect 3292 15444 3298 15456
rect 4157 15453 4169 15456
rect 4203 15453 4215 15487
rect 4157 15447 4215 15453
rect 4801 15487 4859 15493
rect 4801 15453 4813 15487
rect 4847 15484 4859 15487
rect 4890 15484 4896 15496
rect 4847 15456 4896 15484
rect 4847 15453 4859 15456
rect 4801 15447 4859 15453
rect 4890 15444 4896 15456
rect 4948 15444 4954 15496
rect 6086 15484 6092 15496
rect 6047 15456 6092 15484
rect 6086 15444 6092 15456
rect 6144 15444 6150 15496
rect 8110 15484 8116 15496
rect 8071 15456 8116 15484
rect 8110 15444 8116 15456
rect 8168 15444 8174 15496
rect 11330 15484 11336 15496
rect 11291 15456 11336 15484
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 12250 15444 12256 15496
rect 12308 15484 12314 15496
rect 13170 15484 13176 15496
rect 12308 15456 13176 15484
rect 12308 15444 12314 15456
rect 13170 15444 13176 15456
rect 13228 15444 13234 15496
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15484 13783 15487
rect 13906 15484 13912 15496
rect 13771 15456 13912 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 13906 15444 13912 15456
rect 13964 15444 13970 15496
rect 15378 15484 15384 15496
rect 15339 15456 15384 15484
rect 15378 15444 15384 15456
rect 15436 15444 15442 15496
rect 15657 15487 15715 15493
rect 15657 15453 15669 15487
rect 15703 15453 15715 15487
rect 15657 15447 15715 15453
rect 20993 15487 21051 15493
rect 20993 15453 21005 15487
rect 21039 15453 21051 15487
rect 20993 15447 21051 15453
rect 21637 15487 21695 15493
rect 21637 15453 21649 15487
rect 21683 15484 21695 15487
rect 22002 15484 22008 15496
rect 21683 15456 22008 15484
rect 21683 15453 21695 15456
rect 21637 15447 21695 15453
rect 2130 15416 2136 15428
rect 2091 15388 2136 15416
rect 2130 15376 2136 15388
rect 2188 15376 2194 15428
rect 3160 15348 3188 15444
rect 3329 15419 3387 15425
rect 3329 15385 3341 15419
rect 3375 15416 3387 15419
rect 14277 15419 14335 15425
rect 14277 15416 14289 15419
rect 3375 15388 4154 15416
rect 3375 15385 3387 15388
rect 3329 15379 3387 15385
rect 3697 15351 3755 15357
rect 3697 15348 3709 15351
rect 3160 15320 3709 15348
rect 3697 15317 3709 15320
rect 3743 15348 3755 15351
rect 3789 15351 3847 15357
rect 3789 15348 3801 15351
rect 3743 15320 3801 15348
rect 3743 15317 3755 15320
rect 3697 15311 3755 15317
rect 3789 15317 3801 15320
rect 3835 15317 3847 15351
rect 4126 15348 4154 15388
rect 13786 15388 14289 15416
rect 13786 15360 13814 15388
rect 14277 15385 14289 15388
rect 14323 15416 14335 15419
rect 15672 15416 15700 15447
rect 14323 15388 15700 15416
rect 14323 15385 14335 15388
rect 14277 15379 14335 15385
rect 15838 15376 15844 15428
rect 15896 15416 15902 15428
rect 17037 15419 17095 15425
rect 17037 15416 17049 15419
rect 15896 15388 17049 15416
rect 15896 15376 15902 15388
rect 17037 15385 17049 15388
rect 17083 15385 17095 15419
rect 17037 15379 17095 15385
rect 19058 15376 19064 15428
rect 19116 15416 19122 15428
rect 19935 15419 19993 15425
rect 19935 15416 19947 15419
rect 19116 15388 19947 15416
rect 19116 15376 19122 15388
rect 19935 15385 19947 15388
rect 19981 15385 19993 15419
rect 21008 15416 21036 15447
rect 22002 15444 22008 15456
rect 22060 15444 22066 15496
rect 22646 15416 22652 15428
rect 21008 15388 22652 15416
rect 19935 15379 19993 15385
rect 22646 15376 22652 15388
rect 22704 15376 22710 15428
rect 5074 15348 5080 15360
rect 4126 15320 5080 15348
rect 3789 15311 3847 15317
rect 5074 15308 5080 15320
rect 5132 15308 5138 15360
rect 7006 15348 7012 15360
rect 6967 15320 7012 15348
rect 7006 15308 7012 15320
rect 7064 15308 7070 15360
rect 11146 15348 11152 15360
rect 11107 15320 11152 15348
rect 11146 15308 11152 15320
rect 11204 15308 11210 15360
rect 12618 15348 12624 15360
rect 12579 15320 12624 15348
rect 12618 15308 12624 15320
rect 12676 15308 12682 15360
rect 13722 15308 13728 15360
rect 13780 15320 13814 15360
rect 14826 15348 14832 15360
rect 14787 15320 14832 15348
rect 13780 15308 13786 15320
rect 14826 15308 14832 15320
rect 14884 15308 14890 15360
rect 16482 15348 16488 15360
rect 16443 15320 16488 15348
rect 16482 15308 16488 15320
rect 16540 15308 16546 15360
rect 18506 15308 18512 15360
rect 18564 15348 18570 15360
rect 19337 15351 19395 15357
rect 19337 15348 19349 15351
rect 18564 15320 19349 15348
rect 18564 15308 18570 15320
rect 19337 15317 19349 15320
rect 19383 15348 19395 15351
rect 20162 15348 20168 15360
rect 19383 15320 20168 15348
rect 19383 15317 19395 15320
rect 19337 15311 19395 15317
rect 20162 15308 20168 15320
rect 20220 15308 20226 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 2501 15147 2559 15153
rect 2501 15113 2513 15147
rect 2547 15144 2559 15147
rect 2774 15144 2780 15156
rect 2547 15116 2780 15144
rect 2547 15113 2559 15116
rect 2501 15107 2559 15113
rect 2774 15104 2780 15116
rect 2832 15104 2838 15156
rect 3234 15104 3240 15156
rect 3292 15144 3298 15156
rect 3329 15147 3387 15153
rect 3329 15144 3341 15147
rect 3292 15116 3341 15144
rect 3292 15104 3298 15116
rect 3329 15113 3341 15116
rect 3375 15144 3387 15147
rect 4525 15147 4583 15153
rect 4525 15144 4537 15147
rect 3375 15116 4537 15144
rect 3375 15113 3387 15116
rect 3329 15107 3387 15113
rect 3620 15085 3648 15116
rect 4525 15113 4537 15116
rect 4571 15113 4583 15147
rect 4525 15107 4583 15113
rect 5074 15104 5080 15156
rect 5132 15144 5138 15156
rect 5215 15147 5273 15153
rect 5215 15144 5227 15147
rect 5132 15116 5227 15144
rect 5132 15104 5138 15116
rect 5215 15113 5227 15116
rect 5261 15113 5273 15147
rect 5350 15144 5356 15156
rect 5311 15116 5356 15144
rect 5215 15107 5273 15113
rect 5350 15104 5356 15116
rect 5408 15144 5414 15156
rect 6457 15147 6515 15153
rect 6457 15144 6469 15147
rect 5408 15116 6469 15144
rect 5408 15104 5414 15116
rect 6457 15113 6469 15116
rect 6503 15113 6515 15147
rect 6457 15107 6515 15113
rect 7926 15104 7932 15156
rect 7984 15144 7990 15156
rect 8389 15147 8447 15153
rect 8389 15144 8401 15147
rect 7984 15116 8401 15144
rect 7984 15104 7990 15116
rect 8389 15113 8401 15116
rect 8435 15113 8447 15147
rect 10042 15144 10048 15156
rect 10003 15116 10048 15144
rect 8389 15107 8447 15113
rect 10042 15104 10048 15116
rect 10100 15104 10106 15156
rect 10413 15147 10471 15153
rect 10413 15113 10425 15147
rect 10459 15144 10471 15147
rect 10686 15144 10692 15156
rect 10459 15116 10692 15144
rect 10459 15113 10471 15116
rect 10413 15107 10471 15113
rect 10686 15104 10692 15116
rect 10744 15104 10750 15156
rect 11330 15104 11336 15156
rect 11388 15144 11394 15156
rect 12161 15147 12219 15153
rect 12161 15144 12173 15147
rect 11388 15116 12173 15144
rect 11388 15104 11394 15116
rect 12161 15113 12173 15116
rect 12207 15113 12219 15147
rect 12161 15107 12219 15113
rect 12894 15104 12900 15156
rect 12952 15144 12958 15156
rect 14507 15147 14565 15153
rect 14507 15144 14519 15147
rect 12952 15116 14519 15144
rect 12952 15104 12958 15116
rect 14507 15113 14519 15116
rect 14553 15113 14565 15147
rect 15562 15144 15568 15156
rect 14507 15107 14565 15113
rect 15304 15116 15568 15144
rect 3605 15079 3663 15085
rect 3605 15076 3617 15079
rect 3583 15048 3617 15076
rect 3605 15045 3617 15048
rect 3651 15045 3663 15079
rect 3605 15039 3663 15045
rect 6181 15079 6239 15085
rect 6181 15045 6193 15079
rect 6227 15076 6239 15079
rect 6638 15076 6644 15088
rect 6227 15048 6644 15076
rect 6227 15045 6239 15048
rect 6181 15039 6239 15045
rect 6638 15036 6644 15048
rect 6696 15036 6702 15088
rect 6914 15036 6920 15088
rect 6972 15076 6978 15088
rect 11146 15076 11152 15088
rect 6972 15048 11152 15076
rect 6972 15036 6978 15048
rect 2130 14968 2136 15020
rect 2188 15008 2194 15020
rect 2869 15011 2927 15017
rect 2869 15008 2881 15011
rect 2188 14980 2881 15008
rect 2188 14968 2194 14980
rect 2869 14977 2881 14980
rect 2915 15008 2927 15011
rect 4062 15008 4068 15020
rect 2915 14980 4068 15008
rect 2915 14977 2927 14980
rect 2869 14971 2927 14977
rect 4062 14968 4068 14980
rect 4120 14968 4126 15020
rect 5442 15008 5448 15020
rect 5403 14980 5448 15008
rect 5442 14968 5448 14980
rect 5500 14968 5506 15020
rect 7190 14968 7196 15020
rect 7248 15008 7254 15020
rect 7469 15011 7527 15017
rect 7469 15008 7481 15011
rect 7248 14980 7481 15008
rect 7248 14968 7254 14980
rect 7469 14977 7481 14980
rect 7515 14977 7527 15011
rect 8110 15008 8116 15020
rect 8071 14980 8116 15008
rect 7469 14971 7527 14977
rect 8110 14968 8116 14980
rect 8168 14968 8174 15020
rect 10888 15017 10916 15048
rect 11146 15036 11152 15048
rect 11204 15036 11210 15088
rect 14182 15076 14188 15088
rect 12912 15048 13814 15076
rect 14143 15048 14188 15076
rect 12912 15020 12940 15048
rect 10873 15011 10931 15017
rect 10873 14977 10885 15011
rect 10919 14977 10931 15011
rect 12894 15008 12900 15020
rect 12807 14980 12900 15008
rect 10873 14971 10931 14977
rect 12894 14968 12900 14980
rect 12952 14968 12958 15020
rect 13170 15008 13176 15020
rect 13131 14980 13176 15008
rect 13170 14968 13176 14980
rect 13228 14968 13234 15020
rect 13786 15008 13814 15048
rect 14182 15036 14188 15048
rect 14240 15036 14246 15088
rect 15102 15036 15108 15088
rect 15160 15076 15166 15088
rect 15304 15076 15332 15116
rect 15562 15104 15568 15116
rect 15620 15104 15626 15156
rect 16666 15104 16672 15156
rect 16724 15144 16730 15156
rect 16761 15147 16819 15153
rect 16761 15144 16773 15147
rect 16724 15116 16773 15144
rect 16724 15104 16730 15116
rect 16761 15113 16773 15116
rect 16807 15113 16819 15147
rect 16761 15107 16819 15113
rect 16850 15104 16856 15156
rect 16908 15144 16914 15156
rect 17405 15147 17463 15153
rect 17405 15144 17417 15147
rect 16908 15116 17417 15144
rect 16908 15104 16914 15116
rect 17405 15113 17417 15116
rect 17451 15113 17463 15147
rect 17770 15144 17776 15156
rect 17731 15116 17776 15144
rect 17405 15107 17463 15113
rect 17770 15104 17776 15116
rect 17828 15104 17834 15156
rect 18138 15104 18144 15156
rect 18196 15144 18202 15156
rect 18233 15147 18291 15153
rect 18233 15144 18245 15147
rect 18196 15116 18245 15144
rect 18196 15104 18202 15116
rect 18233 15113 18245 15116
rect 18279 15113 18291 15147
rect 21082 15144 21088 15156
rect 21043 15116 21088 15144
rect 18233 15107 18291 15113
rect 21082 15104 21088 15116
rect 21140 15104 21146 15156
rect 21358 15144 21364 15156
rect 21319 15116 21364 15144
rect 21358 15104 21364 15116
rect 21416 15104 21422 15156
rect 22646 15144 22652 15156
rect 22607 15116 22652 15144
rect 22646 15104 22652 15116
rect 22704 15104 22710 15156
rect 24670 15144 24676 15156
rect 24631 15116 24676 15144
rect 24670 15104 24676 15116
rect 24728 15104 24734 15156
rect 24946 15144 24952 15156
rect 24907 15116 24952 15144
rect 24946 15104 24952 15116
rect 25004 15104 25010 15156
rect 15746 15076 15752 15088
rect 15160 15048 15332 15076
rect 15396 15048 15752 15076
rect 15160 15036 15166 15048
rect 15396 15008 15424 15048
rect 15746 15036 15752 15048
rect 15804 15076 15810 15088
rect 16025 15079 16083 15085
rect 16025 15076 16037 15079
rect 15804 15048 16037 15076
rect 15804 15036 15810 15048
rect 16025 15045 16037 15048
rect 16071 15045 16083 15079
rect 20622 15076 20628 15088
rect 20583 15048 20628 15076
rect 16025 15039 16083 15045
rect 20622 15036 20628 15048
rect 20680 15036 20686 15088
rect 13786 14980 15424 15008
rect 15473 15011 15531 15017
rect 15473 14977 15485 15011
rect 15519 15008 15531 15011
rect 15562 15008 15568 15020
rect 15519 14980 15568 15008
rect 15519 14977 15531 14980
rect 15473 14971 15531 14977
rect 15562 14968 15568 14980
rect 15620 14968 15626 15020
rect 15654 14968 15660 15020
rect 15712 15008 15718 15020
rect 17083 15011 17141 15017
rect 17083 15008 17095 15011
rect 15712 14980 17095 15008
rect 15712 14968 15718 14980
rect 17083 14977 17095 14980
rect 17129 14977 17141 15011
rect 18506 15008 18512 15020
rect 18467 14980 18512 15008
rect 17083 14971 17141 14977
rect 18506 14968 18512 14980
rect 18564 14968 18570 15020
rect 18598 14968 18604 15020
rect 18656 15008 18662 15020
rect 19889 15011 19947 15017
rect 18656 14980 19334 15008
rect 18656 14968 18662 14980
rect 658 14900 664 14952
rect 716 14940 722 14952
rect 1489 14943 1547 14949
rect 1489 14940 1501 14943
rect 716 14912 1501 14940
rect 716 14900 722 14912
rect 1489 14909 1501 14912
rect 1535 14940 1547 14943
rect 2406 14940 2412 14952
rect 1535 14912 2412 14940
rect 1535 14909 1547 14912
rect 1489 14903 1547 14909
rect 2406 14900 2412 14912
rect 2464 14940 2470 14952
rect 3050 14940 3056 14952
rect 2464 14912 3056 14940
rect 2464 14900 2470 14912
rect 3050 14900 3056 14912
rect 3108 14900 3114 14952
rect 3510 14940 3516 14952
rect 3471 14912 3516 14940
rect 3510 14900 3516 14912
rect 3568 14900 3574 14952
rect 3789 14943 3847 14949
rect 3789 14909 3801 14943
rect 3835 14940 3847 14943
rect 4246 14940 4252 14952
rect 3835 14912 4252 14940
rect 3835 14909 3847 14912
rect 3789 14903 3847 14909
rect 4246 14900 4252 14912
rect 4304 14940 4310 14952
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4304 14912 4905 14940
rect 4304 14900 4310 14912
rect 4893 14909 4905 14912
rect 4939 14909 4951 14943
rect 4893 14903 4951 14909
rect 4982 14900 4988 14952
rect 5040 14940 5046 14952
rect 5077 14943 5135 14949
rect 5077 14940 5089 14943
rect 5040 14912 5089 14940
rect 5040 14900 5046 14912
rect 5077 14909 5089 14912
rect 5123 14909 5135 14943
rect 8849 14943 8907 14949
rect 8849 14940 8861 14943
rect 5077 14903 5135 14909
rect 8128 14912 8861 14940
rect 2133 14875 2191 14881
rect 2133 14841 2145 14875
rect 2179 14872 2191 14875
rect 2314 14872 2320 14884
rect 2179 14844 2320 14872
rect 2179 14841 2191 14844
rect 2133 14835 2191 14841
rect 2314 14832 2320 14844
rect 2372 14832 2378 14884
rect 5813 14875 5871 14881
rect 5813 14841 5825 14875
rect 5859 14872 5871 14875
rect 7466 14872 7472 14884
rect 5859 14844 7472 14872
rect 5859 14841 5871 14844
rect 5813 14835 5871 14841
rect 7466 14832 7472 14844
rect 7524 14832 7530 14884
rect 7561 14875 7619 14881
rect 7561 14841 7573 14875
rect 7607 14872 7619 14875
rect 8128 14872 8156 14912
rect 8849 14909 8861 14912
rect 8895 14940 8907 14943
rect 9033 14943 9091 14949
rect 9033 14940 9045 14943
rect 8895 14912 9045 14940
rect 8895 14909 8907 14912
rect 8849 14903 8907 14909
rect 9033 14909 9045 14912
rect 9079 14909 9091 14943
rect 9033 14903 9091 14909
rect 14436 14943 14494 14949
rect 14436 14909 14448 14943
rect 14482 14940 14494 14943
rect 14918 14940 14924 14952
rect 14482 14912 14924 14940
rect 14482 14909 14494 14912
rect 14436 14903 14494 14909
rect 14918 14900 14924 14912
rect 14976 14900 14982 14952
rect 16666 14900 16672 14952
rect 16724 14940 16730 14952
rect 16980 14943 17038 14949
rect 16980 14940 16992 14943
rect 16724 14912 16992 14940
rect 16724 14900 16730 14912
rect 16980 14909 16992 14912
rect 17026 14909 17038 14943
rect 16980 14903 17038 14909
rect 7607 14844 8156 14872
rect 7607 14841 7619 14844
rect 7561 14835 7619 14841
rect 2866 14764 2872 14816
rect 2924 14804 2930 14816
rect 3973 14807 4031 14813
rect 3973 14804 3985 14807
rect 2924 14776 3985 14804
rect 2924 14764 2930 14776
rect 3973 14773 3985 14776
rect 4019 14773 4031 14807
rect 3973 14767 4031 14773
rect 7006 14764 7012 14816
rect 7064 14804 7070 14816
rect 7285 14807 7343 14813
rect 7285 14804 7297 14807
rect 7064 14776 7297 14804
rect 7064 14764 7070 14776
rect 7285 14773 7297 14776
rect 7331 14804 7343 14807
rect 7576 14804 7604 14835
rect 8570 14832 8576 14884
rect 8628 14872 8634 14884
rect 8941 14875 8999 14881
rect 8941 14872 8953 14875
rect 8628 14844 8953 14872
rect 8628 14832 8634 14844
rect 8941 14841 8953 14844
rect 8987 14841 8999 14875
rect 8941 14835 8999 14841
rect 10965 14875 11023 14881
rect 10965 14841 10977 14875
rect 11011 14872 11023 14875
rect 11238 14872 11244 14884
rect 11011 14844 11244 14872
rect 11011 14841 11023 14844
rect 10965 14835 11023 14841
rect 11238 14832 11244 14844
rect 11296 14832 11302 14884
rect 11514 14872 11520 14884
rect 11475 14844 11520 14872
rect 11514 14832 11520 14844
rect 11572 14832 11578 14884
rect 12713 14875 12771 14881
rect 12713 14841 12725 14875
rect 12759 14872 12771 14875
rect 12989 14875 13047 14881
rect 12989 14872 13001 14875
rect 12759 14844 13001 14872
rect 12759 14841 12771 14844
rect 12713 14835 12771 14841
rect 12989 14841 13001 14844
rect 13035 14872 13047 14875
rect 13170 14872 13176 14884
rect 13035 14844 13176 14872
rect 13035 14841 13047 14844
rect 12989 14835 13047 14841
rect 13170 14832 13176 14844
rect 13228 14832 13234 14884
rect 15574 14875 15632 14881
rect 15574 14841 15586 14875
rect 15620 14872 15632 14875
rect 16206 14872 16212 14884
rect 15620 14844 16212 14872
rect 15620 14841 15632 14844
rect 15574 14835 15632 14841
rect 16206 14832 16212 14844
rect 16264 14872 16270 14884
rect 16393 14875 16451 14881
rect 16393 14872 16405 14875
rect 16264 14844 16405 14872
rect 16264 14832 16270 14844
rect 16393 14841 16405 14844
rect 16439 14841 16451 14875
rect 18598 14872 18604 14884
rect 18559 14844 18604 14872
rect 16393 14835 16451 14841
rect 18598 14832 18604 14844
rect 18656 14832 18662 14884
rect 19150 14872 19156 14884
rect 19111 14844 19156 14872
rect 19150 14832 19156 14844
rect 19208 14832 19214 14884
rect 19306 14872 19334 14980
rect 19889 14977 19901 15011
rect 19935 15008 19947 15011
rect 20073 15011 20131 15017
rect 20073 15008 20085 15011
rect 19935 14980 20085 15008
rect 19935 14977 19947 14980
rect 19889 14971 19947 14977
rect 20073 14977 20085 14980
rect 20119 15008 20131 15011
rect 21174 15008 21180 15020
rect 20119 14980 21180 15008
rect 20119 14977 20131 14980
rect 20073 14971 20131 14977
rect 21174 14968 21180 14980
rect 21232 14968 21238 15020
rect 21637 15011 21695 15017
rect 21637 14977 21649 15011
rect 21683 15008 21695 15011
rect 21910 15008 21916 15020
rect 21683 14980 21916 15008
rect 21683 14977 21695 14980
rect 21637 14971 21695 14977
rect 21910 14968 21916 14980
rect 21968 14968 21974 15020
rect 22002 14968 22008 15020
rect 22060 15008 22066 15020
rect 22060 14980 22105 15008
rect 22060 14968 22066 14980
rect 24172 14943 24230 14949
rect 24172 14909 24184 14943
rect 24218 14940 24230 14943
rect 24946 14940 24952 14952
rect 24218 14912 24952 14940
rect 24218 14909 24230 14912
rect 24172 14903 24230 14909
rect 24946 14900 24952 14912
rect 25004 14900 25010 14952
rect 20070 14872 20076 14884
rect 19306 14844 20076 14872
rect 20070 14832 20076 14844
rect 20128 14872 20134 14884
rect 20165 14875 20223 14881
rect 20165 14872 20177 14875
rect 20128 14844 20177 14872
rect 20128 14832 20134 14844
rect 20165 14841 20177 14844
rect 20211 14872 20223 14875
rect 21082 14872 21088 14884
rect 20211 14844 21088 14872
rect 20211 14841 20223 14844
rect 20165 14835 20223 14841
rect 21082 14832 21088 14844
rect 21140 14832 21146 14884
rect 21358 14832 21364 14884
rect 21416 14872 21422 14884
rect 21729 14875 21787 14881
rect 21729 14872 21741 14875
rect 21416 14844 21741 14872
rect 21416 14832 21422 14844
rect 21729 14841 21741 14844
rect 21775 14841 21787 14875
rect 24259 14875 24317 14881
rect 24259 14872 24271 14875
rect 21729 14835 21787 14841
rect 21836 14844 24271 14872
rect 7331 14776 7604 14804
rect 11885 14807 11943 14813
rect 7331 14773 7343 14776
rect 7285 14767 7343 14773
rect 11885 14773 11897 14807
rect 11931 14804 11943 14807
rect 11974 14804 11980 14816
rect 11931 14776 11980 14804
rect 11931 14773 11943 14776
rect 11885 14767 11943 14773
rect 11974 14764 11980 14776
rect 12032 14764 12038 14816
rect 13906 14804 13912 14816
rect 13867 14776 13912 14804
rect 13906 14764 13912 14776
rect 13964 14764 13970 14816
rect 14918 14804 14924 14816
rect 14879 14776 14924 14804
rect 14918 14764 14924 14776
rect 14976 14764 14982 14816
rect 15286 14804 15292 14816
rect 15247 14776 15292 14804
rect 15286 14764 15292 14776
rect 15344 14764 15350 14816
rect 19518 14804 19524 14816
rect 19479 14776 19524 14804
rect 19518 14764 19524 14776
rect 19576 14764 19582 14816
rect 21634 14764 21640 14816
rect 21692 14804 21698 14816
rect 21836 14804 21864 14844
rect 24259 14841 24271 14844
rect 24305 14841 24317 14875
rect 24259 14835 24317 14841
rect 21692 14776 21864 14804
rect 21692 14764 21698 14776
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1486 14560 1492 14612
rect 1544 14600 1550 14612
rect 1581 14603 1639 14609
rect 1581 14600 1593 14603
rect 1544 14572 1593 14600
rect 1544 14560 1550 14572
rect 1581 14569 1593 14572
rect 1627 14569 1639 14603
rect 3050 14600 3056 14612
rect 3011 14572 3056 14600
rect 1581 14563 1639 14569
rect 3050 14560 3056 14572
rect 3108 14560 3114 14612
rect 4341 14603 4399 14609
rect 4341 14569 4353 14603
rect 4387 14600 4399 14603
rect 4430 14600 4436 14612
rect 4387 14572 4436 14600
rect 4387 14569 4399 14572
rect 4341 14563 4399 14569
rect 4430 14560 4436 14572
rect 4488 14560 4494 14612
rect 4982 14560 4988 14612
rect 5040 14600 5046 14612
rect 5445 14603 5503 14609
rect 5445 14600 5457 14603
rect 5040 14572 5457 14600
rect 5040 14560 5046 14572
rect 5445 14569 5457 14572
rect 5491 14569 5503 14603
rect 5445 14563 5503 14569
rect 6086 14560 6092 14612
rect 6144 14600 6150 14612
rect 6641 14603 6699 14609
rect 6641 14600 6653 14603
rect 6144 14572 6653 14600
rect 6144 14560 6150 14572
rect 6641 14569 6653 14572
rect 6687 14569 6699 14603
rect 6641 14563 6699 14569
rect 7190 14560 7196 14612
rect 7248 14600 7254 14612
rect 7377 14603 7435 14609
rect 7377 14600 7389 14603
rect 7248 14572 7389 14600
rect 7248 14560 7254 14572
rect 7377 14569 7389 14572
rect 7423 14569 7435 14603
rect 10686 14600 10692 14612
rect 7377 14563 7435 14569
rect 10428 14572 10692 14600
rect 566 14492 572 14544
rect 624 14532 630 14544
rect 1946 14532 1952 14544
rect 624 14504 1952 14532
rect 624 14492 630 14504
rect 1946 14492 1952 14504
rect 2004 14532 2010 14544
rect 2004 14504 2360 14532
rect 2004 14492 2010 14504
rect 2038 14464 2044 14476
rect 1999 14436 2044 14464
rect 2038 14424 2044 14436
rect 2096 14424 2102 14476
rect 2332 14473 2360 14504
rect 4062 14492 4068 14544
rect 4120 14532 4126 14544
rect 7929 14535 7987 14541
rect 4120 14504 5764 14532
rect 4120 14492 4126 14504
rect 2317 14467 2375 14473
rect 2317 14433 2329 14467
rect 2363 14433 2375 14467
rect 4246 14464 4252 14476
rect 4207 14436 4252 14464
rect 2317 14427 2375 14433
rect 4246 14424 4252 14436
rect 4304 14464 4310 14476
rect 5077 14467 5135 14473
rect 5077 14464 5089 14467
rect 4304 14436 5089 14464
rect 4304 14424 4310 14436
rect 5077 14433 5089 14436
rect 5123 14464 5135 14467
rect 5166 14464 5172 14476
rect 5123 14436 5172 14464
rect 5123 14433 5135 14436
rect 5077 14427 5135 14433
rect 5166 14424 5172 14436
rect 5224 14464 5230 14476
rect 5442 14464 5448 14476
rect 5224 14436 5448 14464
rect 5224 14424 5230 14436
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 5736 14473 5764 14504
rect 7929 14501 7941 14535
rect 7975 14532 7987 14535
rect 8570 14532 8576 14544
rect 7975 14504 8576 14532
rect 7975 14501 7987 14504
rect 7929 14495 7987 14501
rect 8570 14492 8576 14504
rect 8628 14492 8634 14544
rect 5721 14467 5779 14473
rect 5721 14433 5733 14467
rect 5767 14464 5779 14467
rect 6178 14464 6184 14476
rect 5767 14436 6184 14464
rect 5767 14433 5779 14436
rect 5721 14427 5779 14433
rect 6178 14424 6184 14436
rect 6236 14424 6242 14476
rect 10226 14424 10232 14476
rect 10284 14464 10290 14476
rect 10428 14473 10456 14572
rect 10686 14560 10692 14572
rect 10744 14560 10750 14612
rect 11974 14560 11980 14612
rect 12032 14600 12038 14612
rect 12069 14603 12127 14609
rect 12069 14600 12081 14603
rect 12032 14572 12081 14600
rect 12032 14560 12038 14572
rect 12069 14569 12081 14572
rect 12115 14569 12127 14603
rect 12069 14563 12127 14569
rect 12621 14603 12679 14609
rect 12621 14569 12633 14603
rect 12667 14600 12679 14603
rect 13446 14600 13452 14612
rect 12667 14572 13452 14600
rect 12667 14569 12679 14572
rect 12621 14563 12679 14569
rect 13446 14560 13452 14572
rect 13504 14600 13510 14612
rect 14737 14603 14795 14609
rect 13504 14572 13676 14600
rect 13504 14560 13510 14572
rect 12894 14532 12900 14544
rect 12855 14504 12900 14532
rect 12894 14492 12900 14504
rect 12952 14492 12958 14544
rect 13648 14541 13676 14572
rect 14737 14569 14749 14603
rect 14783 14600 14795 14603
rect 15378 14600 15384 14612
rect 14783 14572 15384 14600
rect 14783 14569 14795 14572
rect 14737 14563 14795 14569
rect 15378 14560 15384 14572
rect 15436 14600 15442 14612
rect 18598 14600 18604 14612
rect 15436 14572 18368 14600
rect 18559 14572 18604 14600
rect 15436 14560 15442 14572
rect 13633 14535 13691 14541
rect 13633 14501 13645 14535
rect 13679 14501 13691 14535
rect 15102 14532 15108 14544
rect 15063 14504 15108 14532
rect 13633 14495 13691 14501
rect 15102 14492 15108 14504
rect 15160 14492 15166 14544
rect 15286 14492 15292 14544
rect 15344 14532 15350 14544
rect 15657 14535 15715 14541
rect 15657 14532 15669 14535
rect 15344 14504 15669 14532
rect 15344 14492 15350 14504
rect 15657 14501 15669 14504
rect 15703 14532 15715 14535
rect 16022 14532 16028 14544
rect 15703 14504 16028 14532
rect 15703 14501 15715 14504
rect 15657 14495 15715 14501
rect 16022 14492 16028 14504
rect 16080 14492 16086 14544
rect 17862 14532 17868 14544
rect 17823 14504 17868 14532
rect 17862 14492 17868 14504
rect 17920 14492 17926 14544
rect 10413 14467 10471 14473
rect 10413 14464 10425 14467
rect 10284 14436 10425 14464
rect 10284 14424 10290 14436
rect 10413 14433 10425 14436
rect 10459 14433 10471 14467
rect 10686 14464 10692 14476
rect 10647 14436 10692 14464
rect 10413 14427 10471 14433
rect 10686 14424 10692 14436
rect 10744 14424 10750 14476
rect 16390 14424 16396 14476
rect 16448 14464 16454 14476
rect 16574 14464 16580 14476
rect 16448 14436 16580 14464
rect 16448 14424 16454 14436
rect 16574 14424 16580 14436
rect 16632 14464 16638 14476
rect 17126 14464 17132 14476
rect 16632 14436 17132 14464
rect 16632 14424 16638 14436
rect 17126 14424 17132 14436
rect 17184 14424 17190 14476
rect 17681 14467 17739 14473
rect 17681 14433 17693 14467
rect 17727 14464 17739 14467
rect 17727 14436 18276 14464
rect 17727 14433 17739 14436
rect 17681 14427 17739 14433
rect 1394 14356 1400 14408
rect 1452 14396 1458 14408
rect 2501 14399 2559 14405
rect 2501 14396 2513 14399
rect 1452 14368 2513 14396
rect 1452 14356 1458 14368
rect 2501 14365 2513 14368
rect 2547 14365 2559 14399
rect 2501 14359 2559 14365
rect 5534 14356 5540 14408
rect 5592 14396 5598 14408
rect 5629 14399 5687 14405
rect 5629 14396 5641 14399
rect 5592 14368 5641 14396
rect 5592 14356 5598 14368
rect 5629 14365 5641 14368
rect 5675 14365 5687 14399
rect 5629 14359 5687 14365
rect 7101 14399 7159 14405
rect 7101 14365 7113 14399
rect 7147 14396 7159 14399
rect 7837 14399 7895 14405
rect 7837 14396 7849 14399
rect 7147 14368 7849 14396
rect 7147 14365 7159 14368
rect 7101 14359 7159 14365
rect 7837 14365 7849 14368
rect 7883 14365 7895 14399
rect 8110 14396 8116 14408
rect 8071 14368 8116 14396
rect 7837 14359 7895 14365
rect 2130 14328 2136 14340
rect 2091 14300 2136 14328
rect 2130 14288 2136 14300
rect 2188 14288 2194 14340
rect 3605 14263 3663 14269
rect 3605 14229 3617 14263
rect 3651 14260 3663 14263
rect 4246 14260 4252 14272
rect 3651 14232 4252 14260
rect 3651 14229 3663 14232
rect 3605 14223 3663 14229
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 7852 14260 7880 14359
rect 8110 14356 8116 14368
rect 8168 14396 8174 14408
rect 8757 14399 8815 14405
rect 8757 14396 8769 14399
rect 8168 14368 8769 14396
rect 8168 14356 8174 14368
rect 8757 14365 8769 14368
rect 8803 14365 8815 14399
rect 8757 14359 8815 14365
rect 10873 14399 10931 14405
rect 10873 14365 10885 14399
rect 10919 14396 10931 14399
rect 11701 14399 11759 14405
rect 11701 14396 11713 14399
rect 10919 14368 11713 14396
rect 10919 14365 10931 14368
rect 10873 14359 10931 14365
rect 11701 14365 11713 14368
rect 11747 14396 11759 14399
rect 12250 14396 12256 14408
rect 11747 14368 12256 14396
rect 11747 14365 11759 14368
rect 11701 14359 11759 14365
rect 12250 14356 12256 14368
rect 12308 14356 12314 14408
rect 13541 14399 13599 14405
rect 13541 14365 13553 14399
rect 13587 14396 13599 14399
rect 13630 14396 13636 14408
rect 13587 14368 13636 14396
rect 13587 14365 13599 14368
rect 13541 14359 13599 14365
rect 13630 14356 13636 14368
rect 13688 14356 13694 14408
rect 15562 14396 15568 14408
rect 13786 14368 15424 14396
rect 15523 14368 15568 14396
rect 12526 14288 12532 14340
rect 12584 14328 12590 14340
rect 13786 14328 13814 14368
rect 14093 14331 14151 14337
rect 14093 14328 14105 14331
rect 12584 14300 13814 14328
rect 14016 14300 14105 14328
rect 12584 14288 12590 14300
rect 8110 14260 8116 14272
rect 7852 14232 8116 14260
rect 8110 14220 8116 14232
rect 8168 14220 8174 14272
rect 11238 14260 11244 14272
rect 11199 14232 11244 14260
rect 11238 14220 11244 14232
rect 11296 14220 11302 14272
rect 13262 14220 13268 14272
rect 13320 14260 13326 14272
rect 14016 14260 14044 14300
rect 14093 14297 14105 14300
rect 14139 14297 14151 14331
rect 15396 14328 15424 14368
rect 15562 14356 15568 14368
rect 15620 14356 15626 14408
rect 15841 14399 15899 14405
rect 15841 14365 15853 14399
rect 15887 14365 15899 14399
rect 15841 14359 15899 14365
rect 15856 14328 15884 14359
rect 16114 14328 16120 14340
rect 15396 14300 16120 14328
rect 14093 14291 14151 14297
rect 16114 14288 16120 14300
rect 16172 14288 16178 14340
rect 18248 14269 18276 14436
rect 18340 14328 18368 14572
rect 18598 14560 18604 14572
rect 18656 14560 18662 14612
rect 19518 14600 19524 14612
rect 18800 14572 19524 14600
rect 18800 14541 18828 14572
rect 19518 14560 19524 14572
rect 19576 14600 19582 14612
rect 21039 14603 21097 14609
rect 21039 14600 21051 14603
rect 19576 14572 21051 14600
rect 19576 14560 19582 14572
rect 21039 14569 21051 14572
rect 21085 14569 21097 14603
rect 21039 14563 21097 14569
rect 24765 14603 24823 14609
rect 24765 14569 24777 14603
rect 24811 14600 24823 14603
rect 25406 14600 25412 14612
rect 24811 14572 25412 14600
rect 24811 14569 24823 14572
rect 24765 14563 24823 14569
rect 25406 14560 25412 14572
rect 25464 14560 25470 14612
rect 18785 14535 18843 14541
rect 18785 14501 18797 14535
rect 18831 14501 18843 14535
rect 18785 14495 18843 14501
rect 18874 14492 18880 14544
rect 18932 14532 18938 14544
rect 20070 14532 20076 14544
rect 18932 14504 18977 14532
rect 20031 14504 20076 14532
rect 18932 14492 18938 14504
rect 20070 14492 20076 14504
rect 20128 14492 20134 14544
rect 20162 14492 20168 14544
rect 20220 14532 20226 14544
rect 23063 14535 23121 14541
rect 23063 14532 23075 14535
rect 20220 14504 23075 14532
rect 20220 14492 20226 14504
rect 23063 14501 23075 14504
rect 23109 14501 23121 14535
rect 23063 14495 23121 14501
rect 20254 14424 20260 14476
rect 20312 14464 20318 14476
rect 20990 14473 20996 14476
rect 20349 14467 20407 14473
rect 20349 14464 20361 14467
rect 20312 14436 20361 14464
rect 20312 14424 20318 14436
rect 20349 14433 20361 14436
rect 20395 14433 20407 14467
rect 20968 14467 20996 14473
rect 20968 14464 20980 14467
rect 20903 14436 20980 14464
rect 20349 14427 20407 14433
rect 20968 14433 20980 14436
rect 21048 14464 21054 14476
rect 21726 14464 21732 14476
rect 21048 14436 21732 14464
rect 20968 14427 20996 14433
rect 20990 14424 20996 14427
rect 21048 14424 21054 14436
rect 21726 14424 21732 14436
rect 21784 14424 21790 14476
rect 21980 14467 22038 14473
rect 21980 14433 21992 14467
rect 22026 14464 22038 14467
rect 22094 14464 22100 14476
rect 22026 14436 22100 14464
rect 22026 14433 22038 14436
rect 21980 14427 22038 14433
rect 22094 14424 22100 14436
rect 22152 14424 22158 14476
rect 22922 14464 22928 14476
rect 22883 14436 22928 14464
rect 22922 14424 22928 14436
rect 22980 14424 22986 14476
rect 24118 14424 24124 14476
rect 24176 14464 24182 14476
rect 24581 14467 24639 14473
rect 24581 14464 24593 14467
rect 24176 14436 24593 14464
rect 24176 14424 24182 14436
rect 24581 14433 24593 14436
rect 24627 14433 24639 14467
rect 24581 14427 24639 14433
rect 19150 14396 19156 14408
rect 19111 14368 19156 14396
rect 19150 14356 19156 14368
rect 19208 14356 19214 14408
rect 22051 14331 22109 14337
rect 22051 14328 22063 14331
rect 18340 14300 22063 14328
rect 22051 14297 22063 14300
rect 22097 14297 22109 14331
rect 22051 14291 22109 14297
rect 13320 14232 14044 14260
rect 18233 14263 18291 14269
rect 13320 14220 13326 14232
rect 18233 14229 18245 14263
rect 18279 14260 18291 14263
rect 18414 14260 18420 14272
rect 18279 14232 18420 14260
rect 18279 14229 18291 14232
rect 18233 14223 18291 14229
rect 18414 14220 18420 14232
rect 18472 14220 18478 14272
rect 18506 14220 18512 14272
rect 18564 14260 18570 14272
rect 19334 14260 19340 14272
rect 18564 14232 19340 14260
rect 18564 14220 18570 14232
rect 19334 14220 19340 14232
rect 19392 14220 19398 14272
rect 21453 14263 21511 14269
rect 21453 14229 21465 14263
rect 21499 14260 21511 14263
rect 21542 14260 21548 14272
rect 21499 14232 21548 14260
rect 21499 14229 21511 14232
rect 21453 14223 21511 14229
rect 21542 14220 21548 14232
rect 21600 14220 21606 14272
rect 21726 14260 21732 14272
rect 21687 14232 21732 14260
rect 21726 14220 21732 14232
rect 21784 14220 21790 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1578 14056 1584 14068
rect 1539 14028 1584 14056
rect 1578 14016 1584 14028
rect 1636 14016 1642 14068
rect 1946 14016 1952 14068
rect 2004 14056 2010 14068
rect 2041 14059 2099 14065
rect 2041 14056 2053 14059
rect 2004 14028 2053 14056
rect 2004 14016 2010 14028
rect 2041 14025 2053 14028
rect 2087 14056 2099 14059
rect 2314 14056 2320 14068
rect 2087 14028 2320 14056
rect 2087 14025 2099 14028
rect 2041 14019 2099 14025
rect 2314 14016 2320 14028
rect 2372 14056 2378 14068
rect 2409 14059 2467 14065
rect 2409 14056 2421 14059
rect 2372 14028 2421 14056
rect 2372 14016 2378 14028
rect 2409 14025 2421 14028
rect 2455 14056 2467 14059
rect 2958 14056 2964 14068
rect 2455 14028 2964 14056
rect 2455 14025 2467 14028
rect 2409 14019 2467 14025
rect 2958 14016 2964 14028
rect 3016 14016 3022 14068
rect 5166 14056 5172 14068
rect 5127 14028 5172 14056
rect 5166 14016 5172 14028
rect 5224 14016 5230 14068
rect 6178 14056 6184 14068
rect 6139 14028 6184 14056
rect 6178 14016 6184 14028
rect 6236 14016 6242 14068
rect 8570 14056 8576 14068
rect 8531 14028 8576 14056
rect 8570 14016 8576 14028
rect 8628 14016 8634 14068
rect 9306 14016 9312 14068
rect 9364 14056 9370 14068
rect 10137 14059 10195 14065
rect 10137 14056 10149 14059
rect 9364 14028 10149 14056
rect 9364 14016 9370 14028
rect 10137 14025 10149 14028
rect 10183 14056 10195 14059
rect 10226 14056 10232 14068
rect 10183 14028 10232 14056
rect 10183 14025 10195 14028
rect 10137 14019 10195 14025
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 11238 14016 11244 14068
rect 11296 14056 11302 14068
rect 11517 14059 11575 14065
rect 11517 14056 11529 14059
rect 11296 14028 11529 14056
rect 11296 14016 11302 14028
rect 11517 14025 11529 14028
rect 11563 14056 11575 14059
rect 13446 14056 13452 14068
rect 11563 14028 13124 14056
rect 13407 14028 13452 14056
rect 11563 14025 11575 14028
rect 11517 14019 11575 14025
rect 2130 13948 2136 14000
rect 2188 13988 2194 14000
rect 2682 13988 2688 14000
rect 2188 13960 2688 13988
rect 2188 13948 2194 13960
rect 2682 13948 2688 13960
rect 2740 13948 2746 14000
rect 3694 13948 3700 14000
rect 3752 13988 3758 14000
rect 5905 13991 5963 13997
rect 5905 13988 5917 13991
rect 3752 13960 5917 13988
rect 3752 13948 3758 13960
rect 5905 13957 5917 13960
rect 5951 13988 5963 13991
rect 9030 13988 9036 14000
rect 5951 13960 9036 13988
rect 5951 13957 5963 13960
rect 5905 13951 5963 13957
rect 9030 13948 9036 13960
rect 9088 13948 9094 14000
rect 11885 13991 11943 13997
rect 11885 13957 11897 13991
rect 11931 13988 11943 13991
rect 11974 13988 11980 14000
rect 11931 13960 11980 13988
rect 11931 13957 11943 13960
rect 11885 13951 11943 13957
rect 11974 13948 11980 13960
rect 12032 13948 12038 14000
rect 13096 13988 13124 14028
rect 13446 14016 13452 14028
rect 13504 14016 13510 14068
rect 13722 14016 13728 14068
rect 13780 14056 13786 14068
rect 13817 14059 13875 14065
rect 13817 14056 13829 14059
rect 13780 14028 13829 14056
rect 13780 14016 13786 14028
rect 13817 14025 13829 14028
rect 13863 14025 13875 14059
rect 17126 14056 17132 14068
rect 17087 14028 17132 14056
rect 13817 14019 13875 14025
rect 17126 14016 17132 14028
rect 17184 14016 17190 14068
rect 17865 14059 17923 14065
rect 17865 14025 17877 14059
rect 17911 14056 17923 14059
rect 18782 14056 18788 14068
rect 17911 14028 18788 14056
rect 17911 14025 17923 14028
rect 17865 14019 17923 14025
rect 14182 13988 14188 14000
rect 13096 13960 14188 13988
rect 14182 13948 14188 13960
rect 14240 13988 14246 14000
rect 14921 13991 14979 13997
rect 14921 13988 14933 13991
rect 14240 13960 14933 13988
rect 14240 13948 14246 13960
rect 14921 13957 14933 13960
rect 14967 13988 14979 13991
rect 15286 13988 15292 14000
rect 14967 13960 15292 13988
rect 14967 13957 14979 13960
rect 14921 13951 14979 13957
rect 15286 13948 15292 13960
rect 15344 13948 15350 14000
rect 15746 13988 15752 14000
rect 15707 13960 15752 13988
rect 15746 13948 15752 13960
rect 15804 13948 15810 14000
rect 1946 13880 1952 13932
rect 2004 13920 2010 13932
rect 3053 13923 3111 13929
rect 3053 13920 3065 13923
rect 2004 13892 3065 13920
rect 2004 13880 2010 13892
rect 3053 13889 3065 13892
rect 3099 13889 3111 13923
rect 3053 13883 3111 13889
rect 3881 13923 3939 13929
rect 3881 13889 3893 13923
rect 3927 13920 3939 13923
rect 4249 13923 4307 13929
rect 4249 13920 4261 13923
rect 3927 13892 4261 13920
rect 3927 13889 3939 13892
rect 3881 13883 3939 13889
rect 4249 13889 4261 13892
rect 4295 13889 4307 13923
rect 5537 13923 5595 13929
rect 5537 13920 5549 13923
rect 4249 13883 4307 13889
rect 4448 13892 5549 13920
rect 4448 13864 4476 13892
rect 5537 13889 5549 13892
rect 5583 13889 5595 13923
rect 6549 13923 6607 13929
rect 6549 13920 6561 13923
rect 5537 13883 5595 13889
rect 5736 13892 6561 13920
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 1486 13852 1492 13864
rect 1443 13824 1492 13852
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 1486 13812 1492 13824
rect 1544 13812 1550 13864
rect 2590 13812 2596 13864
rect 2648 13852 2654 13864
rect 2869 13855 2927 13861
rect 2648 13824 2693 13852
rect 2648 13812 2654 13824
rect 2869 13821 2881 13855
rect 2915 13852 2927 13855
rect 2958 13852 2964 13864
rect 2915 13824 2964 13852
rect 2915 13821 2927 13824
rect 2869 13815 2927 13821
rect 2958 13812 2964 13824
rect 3016 13812 3022 13864
rect 4062 13812 4068 13864
rect 4120 13852 4126 13864
rect 4157 13855 4215 13861
rect 4157 13852 4169 13855
rect 4120 13824 4169 13852
rect 4120 13812 4126 13824
rect 4157 13821 4169 13824
rect 4203 13821 4215 13855
rect 4157 13815 4215 13821
rect 4430 13812 4436 13864
rect 4488 13852 4494 13864
rect 4488 13824 4581 13852
rect 4488 13812 4494 13824
rect 5442 13812 5448 13864
rect 5500 13852 5506 13864
rect 5736 13861 5764 13892
rect 6549 13889 6561 13892
rect 6595 13889 6607 13923
rect 9048 13920 9076 13948
rect 9769 13923 9827 13929
rect 9048 13892 9536 13920
rect 6549 13883 6607 13889
rect 5721 13855 5779 13861
rect 5721 13852 5733 13855
rect 5500 13824 5733 13852
rect 5500 13812 5506 13824
rect 5721 13821 5733 13824
rect 5767 13821 5779 13855
rect 5721 13815 5779 13821
rect 7745 13855 7803 13861
rect 7745 13821 7757 13855
rect 7791 13821 7803 13855
rect 7926 13852 7932 13864
rect 7887 13824 7932 13852
rect 7745 13815 7803 13821
rect 3050 13744 3056 13796
rect 3108 13784 3114 13796
rect 3108 13756 4108 13784
rect 3108 13744 3114 13756
rect 2682 13676 2688 13728
rect 2740 13716 2746 13728
rect 3605 13719 3663 13725
rect 3605 13716 3617 13719
rect 2740 13688 3617 13716
rect 2740 13676 2746 13688
rect 3605 13685 3617 13688
rect 3651 13716 3663 13719
rect 3881 13719 3939 13725
rect 3881 13716 3893 13719
rect 3651 13688 3893 13716
rect 3651 13685 3663 13688
rect 3605 13679 3663 13685
rect 3881 13685 3893 13688
rect 3927 13716 3939 13719
rect 3973 13719 4031 13725
rect 3973 13716 3985 13719
rect 3927 13688 3985 13716
rect 3927 13685 3939 13688
rect 3881 13679 3939 13685
rect 3973 13685 3985 13688
rect 4019 13685 4031 13719
rect 4080 13716 4108 13756
rect 4430 13716 4436 13728
rect 4080 13688 4436 13716
rect 3973 13679 4031 13685
rect 4430 13676 4436 13688
rect 4488 13676 4494 13728
rect 4614 13716 4620 13728
rect 4575 13688 4620 13716
rect 4614 13676 4620 13688
rect 4672 13676 4678 13728
rect 7377 13719 7435 13725
rect 7377 13685 7389 13719
rect 7423 13716 7435 13719
rect 7760 13716 7788 13815
rect 7926 13812 7932 13824
rect 7984 13812 7990 13864
rect 9508 13861 9536 13892
rect 9769 13889 9781 13923
rect 9815 13920 9827 13923
rect 10597 13923 10655 13929
rect 10597 13920 10609 13923
rect 9815 13892 10609 13920
rect 9815 13889 9827 13892
rect 9769 13883 9827 13889
rect 10597 13889 10609 13892
rect 10643 13920 10655 13923
rect 10778 13920 10784 13932
rect 10643 13892 10784 13920
rect 10643 13889 10655 13892
rect 10597 13883 10655 13889
rect 10778 13880 10784 13892
rect 10836 13880 10842 13932
rect 11514 13880 11520 13932
rect 11572 13920 11578 13932
rect 12526 13920 12532 13932
rect 11572 13892 12532 13920
rect 11572 13880 11578 13892
rect 12526 13880 12532 13892
rect 12584 13880 12590 13932
rect 13173 13923 13231 13929
rect 13173 13889 13185 13923
rect 13219 13920 13231 13923
rect 13262 13920 13268 13932
rect 13219 13892 13268 13920
rect 13219 13889 13231 13892
rect 13173 13883 13231 13889
rect 13262 13880 13268 13892
rect 13320 13880 13326 13932
rect 13906 13880 13912 13932
rect 13964 13920 13970 13932
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 13964 13892 16681 13920
rect 13964 13880 13970 13892
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 18064 13864 18092 14028
rect 18782 14016 18788 14028
rect 18840 14016 18846 14068
rect 18874 14016 18880 14068
rect 18932 14056 18938 14068
rect 19061 14059 19119 14065
rect 19061 14056 19073 14059
rect 18932 14028 19073 14056
rect 18932 14016 18938 14028
rect 19061 14025 19073 14028
rect 19107 14025 19119 14059
rect 20990 14056 20996 14068
rect 20951 14028 20996 14056
rect 19061 14019 19119 14025
rect 20990 14016 20996 14028
rect 21048 14016 21054 14068
rect 21542 13988 21548 14000
rect 20272 13960 21548 13988
rect 20272 13920 20300 13960
rect 21542 13948 21548 13960
rect 21600 13948 21606 14000
rect 18616 13892 20300 13920
rect 9033 13855 9091 13861
rect 9033 13852 9045 13855
rect 8864 13824 9045 13852
rect 8202 13784 8208 13796
rect 8163 13756 8208 13784
rect 8202 13744 8208 13756
rect 8260 13744 8266 13796
rect 8294 13744 8300 13796
rect 8352 13784 8358 13796
rect 8570 13784 8576 13796
rect 8352 13756 8576 13784
rect 8352 13744 8358 13756
rect 8570 13744 8576 13756
rect 8628 13744 8634 13796
rect 8864 13716 8892 13824
rect 9033 13821 9045 13824
rect 9079 13821 9091 13855
rect 9033 13815 9091 13821
rect 9493 13855 9551 13861
rect 9493 13821 9505 13855
rect 9539 13821 9551 13855
rect 13998 13852 14004 13864
rect 13959 13824 14004 13852
rect 9493 13815 9551 13821
rect 13998 13812 14004 13824
rect 14056 13852 14062 13864
rect 14461 13855 14519 13861
rect 14461 13852 14473 13855
rect 14056 13824 14473 13852
rect 14056 13812 14062 13824
rect 14461 13821 14473 13824
rect 14507 13821 14519 13855
rect 18046 13852 18052 13864
rect 17959 13824 18052 13852
rect 14461 13815 14519 13821
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 18414 13852 18420 13864
rect 18327 13824 18420 13852
rect 18414 13812 18420 13824
rect 18472 13852 18478 13864
rect 18616 13861 18644 13892
rect 20806 13880 20812 13932
rect 20864 13920 20870 13932
rect 22922 13920 22928 13932
rect 20864 13892 22928 13920
rect 20864 13880 20870 13892
rect 22922 13880 22928 13892
rect 22980 13880 22986 13932
rect 18601 13855 18659 13861
rect 18601 13852 18613 13855
rect 18472 13824 18613 13852
rect 18472 13812 18478 13824
rect 18601 13821 18613 13824
rect 18647 13821 18659 13855
rect 18601 13815 18659 13821
rect 21361 13855 21419 13861
rect 21361 13821 21373 13855
rect 21407 13852 21419 13855
rect 21407 13824 21441 13852
rect 21407 13821 21419 13824
rect 21361 13815 21419 13821
rect 10505 13787 10563 13793
rect 10505 13753 10517 13787
rect 10551 13784 10563 13787
rect 10959 13787 11017 13793
rect 10959 13784 10971 13787
rect 10551 13756 10971 13784
rect 10551 13753 10563 13756
rect 10505 13747 10563 13753
rect 10959 13753 10971 13756
rect 11005 13784 11017 13787
rect 11974 13784 11980 13796
rect 11005 13756 11980 13784
rect 11005 13753 11017 13756
rect 10959 13747 11017 13753
rect 11974 13744 11980 13756
rect 12032 13744 12038 13796
rect 12621 13787 12679 13793
rect 12621 13753 12633 13787
rect 12667 13753 12679 13787
rect 12621 13747 12679 13753
rect 15197 13787 15255 13793
rect 15197 13753 15209 13787
rect 15243 13753 15255 13787
rect 15197 13747 15255 13753
rect 8941 13719 8999 13725
rect 8941 13716 8953 13719
rect 7423 13688 8953 13716
rect 7423 13685 7435 13688
rect 7377 13679 7435 13685
rect 8941 13685 8953 13688
rect 8987 13716 8999 13719
rect 9122 13716 9128 13728
rect 8987 13688 9128 13716
rect 8987 13685 8999 13688
rect 8941 13679 8999 13685
rect 9122 13676 9128 13688
rect 9180 13676 9186 13728
rect 11882 13676 11888 13728
rect 11940 13716 11946 13728
rect 12161 13719 12219 13725
rect 12161 13716 12173 13719
rect 11940 13688 12173 13716
rect 11940 13676 11946 13688
rect 12161 13685 12173 13688
rect 12207 13716 12219 13719
rect 12636 13716 12664 13747
rect 12207 13688 12664 13716
rect 12207 13685 12219 13688
rect 12161 13679 12219 13685
rect 12710 13676 12716 13728
rect 12768 13716 12774 13728
rect 14185 13719 14243 13725
rect 14185 13716 14197 13719
rect 12768 13688 14197 13716
rect 12768 13676 12774 13688
rect 14185 13685 14197 13688
rect 14231 13685 14243 13719
rect 15212 13716 15240 13747
rect 15286 13744 15292 13796
rect 15344 13784 15350 13796
rect 18432 13784 18460 13812
rect 15344 13756 15389 13784
rect 16500 13756 18460 13784
rect 15344 13744 15350 13756
rect 16500 13728 16528 13756
rect 19150 13744 19156 13796
rect 19208 13784 19214 13796
rect 19705 13787 19763 13793
rect 19705 13784 19717 13787
rect 19208 13756 19717 13784
rect 19208 13744 19214 13756
rect 19705 13753 19717 13756
rect 19751 13753 19763 13787
rect 19705 13747 19763 13753
rect 19797 13787 19855 13793
rect 19797 13753 19809 13787
rect 19843 13753 19855 13787
rect 19797 13747 19855 13753
rect 20349 13787 20407 13793
rect 20349 13753 20361 13787
rect 20395 13784 20407 13787
rect 21174 13784 21180 13796
rect 20395 13756 21180 13784
rect 20395 13753 20407 13756
rect 20349 13747 20407 13753
rect 15378 13716 15384 13728
rect 15212 13688 15384 13716
rect 14185 13679 14243 13685
rect 15378 13676 15384 13688
rect 15436 13676 15442 13728
rect 16022 13676 16028 13728
rect 16080 13716 16086 13728
rect 16117 13719 16175 13725
rect 16117 13716 16129 13719
rect 16080 13688 16129 13716
rect 16080 13676 16086 13688
rect 16117 13685 16129 13688
rect 16163 13685 16175 13719
rect 16117 13679 16175 13685
rect 16298 13676 16304 13728
rect 16356 13716 16362 13728
rect 16482 13716 16488 13728
rect 16356 13688 16488 13716
rect 16356 13676 16362 13688
rect 16482 13676 16488 13688
rect 16540 13676 16546 13728
rect 18138 13716 18144 13728
rect 18099 13688 18144 13716
rect 18138 13676 18144 13688
rect 18196 13676 18202 13728
rect 19426 13716 19432 13728
rect 19387 13688 19432 13716
rect 19426 13676 19432 13688
rect 19484 13716 19490 13728
rect 19812 13716 19840 13747
rect 21174 13744 21180 13756
rect 21232 13744 21238 13796
rect 21376 13784 21404 13815
rect 21542 13812 21548 13864
rect 21600 13852 21606 13864
rect 21637 13855 21695 13861
rect 21637 13852 21649 13855
rect 21600 13824 21649 13852
rect 21600 13812 21606 13824
rect 21637 13821 21649 13824
rect 21683 13821 21695 13855
rect 21637 13815 21695 13821
rect 21726 13784 21732 13796
rect 21376 13756 21732 13784
rect 21726 13744 21732 13756
rect 21784 13744 21790 13796
rect 19484 13688 19840 13716
rect 19484 13676 19490 13688
rect 19978 13676 19984 13728
rect 20036 13716 20042 13728
rect 21269 13719 21327 13725
rect 21269 13716 21281 13719
rect 20036 13688 21281 13716
rect 20036 13676 20042 13688
rect 21269 13685 21281 13688
rect 21315 13685 21327 13719
rect 21269 13679 21327 13685
rect 22094 13676 22100 13728
rect 22152 13716 22158 13728
rect 22189 13719 22247 13725
rect 22189 13716 22201 13719
rect 22152 13688 22201 13716
rect 22152 13676 22158 13688
rect 22189 13685 22201 13688
rect 22235 13685 22247 13719
rect 22189 13679 22247 13685
rect 24118 13676 24124 13728
rect 24176 13716 24182 13728
rect 24581 13719 24639 13725
rect 24581 13716 24593 13719
rect 24176 13688 24593 13716
rect 24176 13676 24182 13688
rect 24581 13685 24593 13688
rect 24627 13685 24639 13719
rect 24581 13679 24639 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 3602 13472 3608 13524
rect 3660 13512 3666 13524
rect 3789 13515 3847 13521
rect 3789 13512 3801 13515
rect 3660 13484 3801 13512
rect 3660 13472 3666 13484
rect 3789 13481 3801 13484
rect 3835 13481 3847 13515
rect 5534 13512 5540 13524
rect 3789 13475 3847 13481
rect 3896 13484 5540 13512
rect 2406 13444 2412 13456
rect 2319 13416 2412 13444
rect 2406 13404 2412 13416
rect 2464 13444 2470 13456
rect 3050 13444 3056 13456
rect 2464 13416 3056 13444
rect 2464 13404 2470 13416
rect 3050 13404 3056 13416
rect 3108 13404 3114 13456
rect 3513 13447 3571 13453
rect 3513 13413 3525 13447
rect 3559 13444 3571 13447
rect 3896 13444 3924 13484
rect 5534 13472 5540 13484
rect 5592 13472 5598 13524
rect 10134 13512 10140 13524
rect 10095 13484 10140 13512
rect 10134 13472 10140 13484
rect 10192 13472 10198 13524
rect 10778 13512 10784 13524
rect 10739 13484 10784 13512
rect 10778 13472 10784 13484
rect 10836 13472 10842 13524
rect 11882 13512 11888 13524
rect 11843 13484 11888 13512
rect 11882 13472 11888 13484
rect 11940 13472 11946 13524
rect 12250 13512 12256 13524
rect 12211 13484 12256 13512
rect 12250 13472 12256 13484
rect 12308 13472 12314 13524
rect 12526 13512 12532 13524
rect 12487 13484 12532 13512
rect 12526 13472 12532 13484
rect 12584 13472 12590 13524
rect 13170 13472 13176 13524
rect 13228 13512 13234 13524
rect 13633 13515 13691 13521
rect 13633 13512 13645 13515
rect 13228 13484 13645 13512
rect 13228 13472 13234 13484
rect 13633 13481 13645 13484
rect 13679 13481 13691 13515
rect 13633 13475 13691 13481
rect 15286 13472 15292 13524
rect 15344 13512 15350 13524
rect 17129 13515 17187 13521
rect 17129 13512 17141 13515
rect 15344 13484 17141 13512
rect 15344 13472 15350 13484
rect 17129 13481 17141 13484
rect 17175 13481 17187 13515
rect 17129 13475 17187 13481
rect 18230 13472 18236 13524
rect 18288 13512 18294 13524
rect 18325 13515 18383 13521
rect 18325 13512 18337 13515
rect 18288 13484 18337 13512
rect 18288 13472 18294 13484
rect 18325 13481 18337 13484
rect 18371 13481 18383 13515
rect 18325 13475 18383 13481
rect 19705 13515 19763 13521
rect 19705 13481 19717 13515
rect 19751 13512 19763 13515
rect 19751 13484 21128 13512
rect 19751 13481 19763 13484
rect 19705 13475 19763 13481
rect 3559 13416 3924 13444
rect 4065 13447 4123 13453
rect 3559 13413 3571 13416
rect 3513 13407 3571 13413
rect 4065 13413 4077 13447
rect 4111 13444 4123 13447
rect 4706 13444 4712 13456
rect 4111 13416 4712 13444
rect 4111 13413 4123 13416
rect 4065 13407 4123 13413
rect 4706 13404 4712 13416
rect 4764 13444 4770 13456
rect 5350 13444 5356 13456
rect 4764 13416 5356 13444
rect 4764 13404 4770 13416
rect 5350 13404 5356 13416
rect 5408 13404 5414 13456
rect 5899 13447 5957 13453
rect 5899 13413 5911 13447
rect 5945 13444 5957 13447
rect 6086 13444 6092 13456
rect 5945 13416 6092 13444
rect 5945 13413 5957 13416
rect 5899 13407 5957 13413
rect 6086 13404 6092 13416
rect 6144 13404 6150 13456
rect 8199 13447 8257 13453
rect 8199 13413 8211 13447
rect 8245 13444 8257 13447
rect 8294 13444 8300 13456
rect 8245 13416 8300 13444
rect 8245 13413 8257 13416
rect 8199 13407 8257 13413
rect 8294 13404 8300 13416
rect 8352 13444 8358 13456
rect 11327 13447 11385 13453
rect 11327 13444 11339 13447
rect 8352 13416 11339 13444
rect 8352 13404 8358 13416
rect 11327 13413 11339 13416
rect 11373 13444 11385 13447
rect 11974 13444 11980 13456
rect 11373 13416 11980 13444
rect 11373 13413 11385 13416
rect 11327 13407 11385 13413
rect 11974 13404 11980 13416
rect 12032 13444 12038 13456
rect 13075 13447 13133 13453
rect 13075 13444 13087 13447
rect 12032 13416 13087 13444
rect 12032 13404 12038 13416
rect 13075 13413 13087 13416
rect 13121 13444 13133 13447
rect 13446 13444 13452 13456
rect 13121 13416 13452 13444
rect 13121 13413 13133 13416
rect 13075 13407 13133 13413
rect 13446 13404 13452 13416
rect 13504 13404 13510 13456
rect 14734 13404 14740 13456
rect 14792 13444 14798 13456
rect 15657 13447 15715 13453
rect 15657 13444 15669 13447
rect 14792 13416 15669 13444
rect 14792 13404 14798 13416
rect 15657 13413 15669 13416
rect 15703 13444 15715 13447
rect 16022 13444 16028 13456
rect 15703 13416 16028 13444
rect 15703 13413 15715 13416
rect 15657 13407 15715 13413
rect 16022 13404 16028 13416
rect 16080 13404 16086 13456
rect 18046 13444 18052 13456
rect 17328 13416 18052 13444
rect 2314 13376 2320 13388
rect 2275 13348 2320 13376
rect 2314 13336 2320 13348
rect 2372 13336 2378 13388
rect 4154 13336 4160 13388
rect 4212 13376 4218 13388
rect 4249 13379 4307 13385
rect 4249 13376 4261 13379
rect 4212 13348 4261 13376
rect 4212 13336 4218 13348
rect 4249 13345 4261 13348
rect 4295 13345 4307 13379
rect 4249 13339 4307 13345
rect 4985 13379 5043 13385
rect 4985 13345 4997 13379
rect 5031 13376 5043 13379
rect 5994 13376 6000 13388
rect 5031 13348 6000 13376
rect 5031 13345 5043 13348
rect 4985 13339 5043 13345
rect 2222 13268 2228 13320
rect 2280 13308 2286 13320
rect 4801 13311 4859 13317
rect 4801 13308 4813 13311
rect 2280 13280 4813 13308
rect 2280 13268 2286 13280
rect 4801 13277 4813 13280
rect 4847 13277 4859 13311
rect 4801 13271 4859 13277
rect 2038 13200 2044 13252
rect 2096 13240 2102 13252
rect 4062 13240 4068 13252
rect 2096 13212 4068 13240
rect 2096 13200 2102 13212
rect 2884 13184 2912 13212
rect 4062 13200 4068 13212
rect 4120 13240 4126 13252
rect 5000 13240 5028 13339
rect 5994 13336 6000 13348
rect 6052 13336 6058 13388
rect 8757 13379 8815 13385
rect 8757 13345 8769 13379
rect 8803 13376 8815 13379
rect 9858 13376 9864 13388
rect 8803 13348 9864 13376
rect 8803 13345 8815 13348
rect 8757 13339 8815 13345
rect 9858 13336 9864 13348
rect 9916 13336 9922 13388
rect 9953 13379 10011 13385
rect 9953 13345 9965 13379
rect 9999 13376 10011 13379
rect 10778 13376 10784 13388
rect 9999 13348 10784 13376
rect 9999 13345 10011 13348
rect 9953 13339 10011 13345
rect 5534 13308 5540 13320
rect 5495 13280 5540 13308
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 7834 13308 7840 13320
rect 7795 13280 7840 13308
rect 7834 13268 7840 13280
rect 7892 13268 7898 13320
rect 9030 13268 9036 13320
rect 9088 13308 9094 13320
rect 9125 13311 9183 13317
rect 9125 13308 9137 13311
rect 9088 13280 9137 13308
rect 9088 13268 9094 13280
rect 9125 13277 9137 13280
rect 9171 13308 9183 13311
rect 9968 13308 9996 13339
rect 10778 13336 10784 13348
rect 10836 13336 10842 13388
rect 14645 13379 14703 13385
rect 14645 13345 14657 13379
rect 14691 13376 14703 13379
rect 14918 13376 14924 13388
rect 14691 13348 14924 13376
rect 14691 13345 14703 13348
rect 14645 13339 14703 13345
rect 14918 13336 14924 13348
rect 14976 13336 14982 13388
rect 17126 13336 17132 13388
rect 17184 13376 17190 13388
rect 17328 13385 17356 13416
rect 18046 13404 18052 13416
rect 18104 13404 18110 13456
rect 18340 13444 18368 13475
rect 18690 13444 18696 13456
rect 18340 13416 18696 13444
rect 18690 13404 18696 13416
rect 18748 13444 18754 13456
rect 19106 13447 19164 13453
rect 19106 13444 19118 13447
rect 18748 13416 19118 13444
rect 18748 13404 18754 13416
rect 19106 13413 19118 13416
rect 19152 13413 19164 13447
rect 19106 13407 19164 13413
rect 20622 13404 20628 13456
rect 20680 13444 20686 13456
rect 21100 13453 21128 13484
rect 20993 13447 21051 13453
rect 20993 13444 21005 13447
rect 20680 13416 21005 13444
rect 20680 13404 20686 13416
rect 20993 13413 21005 13416
rect 21039 13413 21051 13447
rect 20993 13407 21051 13413
rect 21085 13447 21143 13453
rect 21085 13413 21097 13447
rect 21131 13444 21143 13447
rect 21266 13444 21272 13456
rect 21131 13416 21272 13444
rect 21131 13413 21143 13416
rect 21085 13407 21143 13413
rect 21266 13404 21272 13416
rect 21324 13404 21330 13456
rect 21450 13404 21456 13456
rect 21508 13444 21514 13456
rect 22094 13444 22100 13456
rect 21508 13416 22100 13444
rect 21508 13404 21514 13416
rect 22094 13404 22100 13416
rect 22152 13404 22158 13456
rect 17313 13379 17371 13385
rect 17313 13376 17325 13379
rect 17184 13348 17325 13376
rect 17184 13336 17190 13348
rect 17313 13345 17325 13348
rect 17359 13345 17371 13379
rect 17494 13376 17500 13388
rect 17455 13348 17500 13376
rect 17313 13339 17371 13345
rect 17494 13336 17500 13348
rect 17552 13336 17558 13388
rect 18785 13379 18843 13385
rect 18785 13345 18797 13379
rect 18831 13376 18843 13379
rect 19518 13376 19524 13388
rect 18831 13348 19524 13376
rect 18831 13345 18843 13348
rect 18785 13339 18843 13345
rect 19518 13336 19524 13348
rect 19576 13376 19582 13388
rect 19978 13376 19984 13388
rect 19576 13348 19984 13376
rect 19576 13336 19582 13348
rect 19978 13336 19984 13348
rect 20036 13336 20042 13388
rect 10962 13308 10968 13320
rect 9171 13280 9996 13308
rect 10923 13280 10968 13308
rect 9171 13277 9183 13280
rect 9125 13271 9183 13277
rect 10962 13268 10968 13280
rect 11020 13268 11026 13320
rect 12710 13308 12716 13320
rect 12671 13280 12716 13308
rect 12710 13268 12716 13280
rect 12768 13268 12774 13320
rect 15105 13311 15163 13317
rect 15105 13277 15117 13311
rect 15151 13308 15163 13311
rect 15378 13308 15384 13320
rect 15151 13280 15384 13308
rect 15151 13277 15163 13280
rect 15105 13271 15163 13277
rect 15378 13268 15384 13280
rect 15436 13268 15442 13320
rect 15565 13311 15623 13317
rect 15565 13277 15577 13311
rect 15611 13277 15623 13311
rect 15565 13271 15623 13277
rect 4120 13212 5028 13240
rect 4120 13200 4126 13212
rect 11698 13200 11704 13252
rect 11756 13240 11762 13252
rect 15580 13240 15608 13271
rect 15746 13268 15752 13320
rect 15804 13308 15810 13320
rect 15841 13311 15899 13317
rect 15841 13308 15853 13311
rect 15804 13280 15853 13308
rect 15804 13268 15810 13280
rect 15841 13277 15853 13280
rect 15887 13277 15899 13311
rect 15841 13271 15899 13277
rect 18414 13268 18420 13320
rect 18472 13308 18478 13320
rect 19334 13308 19340 13320
rect 18472 13280 19340 13308
rect 18472 13268 18478 13280
rect 19334 13268 19340 13280
rect 19392 13268 19398 13320
rect 21174 13268 21180 13320
rect 21232 13308 21238 13320
rect 21269 13311 21327 13317
rect 21269 13308 21281 13311
rect 21232 13280 21281 13308
rect 21232 13268 21238 13280
rect 21269 13277 21281 13280
rect 21315 13277 21327 13311
rect 21269 13271 21327 13277
rect 15930 13240 15936 13252
rect 11756 13212 15240 13240
rect 15580 13212 15936 13240
rect 11756 13200 11762 13212
rect 2130 13132 2136 13184
rect 2188 13172 2194 13184
rect 2682 13172 2688 13184
rect 2188 13144 2688 13172
rect 2188 13132 2194 13144
rect 2682 13132 2688 13144
rect 2740 13132 2746 13184
rect 2866 13132 2872 13184
rect 2924 13172 2930 13184
rect 3053 13175 3111 13181
rect 3053 13172 3065 13175
rect 2924 13144 3065 13172
rect 2924 13132 2930 13144
rect 3053 13141 3065 13144
rect 3099 13141 3111 13175
rect 3053 13135 3111 13141
rect 3786 13132 3792 13184
rect 3844 13172 3850 13184
rect 4341 13175 4399 13181
rect 4341 13172 4353 13175
rect 3844 13144 4353 13172
rect 3844 13132 3850 13144
rect 4341 13141 4353 13144
rect 4387 13141 4399 13175
rect 4341 13135 4399 13141
rect 4801 13175 4859 13181
rect 4801 13141 4813 13175
rect 4847 13172 4859 13175
rect 5261 13175 5319 13181
rect 5261 13172 5273 13175
rect 4847 13144 5273 13172
rect 4847 13141 4859 13144
rect 4801 13135 4859 13141
rect 5261 13141 5273 13144
rect 5307 13172 5319 13175
rect 6362 13172 6368 13184
rect 5307 13144 6368 13172
rect 5307 13141 5319 13144
rect 5261 13135 5319 13141
rect 6362 13132 6368 13144
rect 6420 13132 6426 13184
rect 6457 13175 6515 13181
rect 6457 13141 6469 13175
rect 6503 13172 6515 13175
rect 6825 13175 6883 13181
rect 6825 13172 6837 13175
rect 6503 13144 6837 13172
rect 6503 13141 6515 13144
rect 6457 13135 6515 13141
rect 6825 13141 6837 13144
rect 6871 13172 6883 13175
rect 7006 13172 7012 13184
rect 6871 13144 7012 13172
rect 6871 13141 6883 13144
rect 6825 13135 6883 13141
rect 7006 13132 7012 13144
rect 7064 13132 7070 13184
rect 7098 13132 7104 13184
rect 7156 13172 7162 13184
rect 7469 13175 7527 13181
rect 7469 13172 7481 13175
rect 7156 13144 7481 13172
rect 7156 13132 7162 13144
rect 7469 13141 7481 13144
rect 7515 13172 7527 13175
rect 7926 13172 7932 13184
rect 7515 13144 7932 13172
rect 7515 13141 7527 13144
rect 7469 13135 7527 13141
rect 7926 13132 7932 13144
rect 7984 13132 7990 13184
rect 10410 13172 10416 13184
rect 10371 13144 10416 13172
rect 10410 13132 10416 13144
rect 10468 13172 10474 13184
rect 10686 13172 10692 13184
rect 10468 13144 10692 13172
rect 10468 13132 10474 13144
rect 10686 13132 10692 13144
rect 10744 13132 10750 13184
rect 13906 13172 13912 13184
rect 13867 13144 13912 13172
rect 13906 13132 13912 13144
rect 13964 13132 13970 13184
rect 15212 13172 15240 13212
rect 15930 13200 15936 13212
rect 15988 13200 15994 13252
rect 16390 13172 16396 13184
rect 15212 13144 16396 13172
rect 16390 13132 16396 13144
rect 16448 13132 16454 13184
rect 19150 13132 19156 13184
rect 19208 13172 19214 13184
rect 19981 13175 20039 13181
rect 19981 13172 19993 13175
rect 19208 13144 19993 13172
rect 19208 13132 19214 13144
rect 19981 13141 19993 13144
rect 20027 13141 20039 13175
rect 19981 13135 20039 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1118 12928 1124 12980
rect 1176 12968 1182 12980
rect 1581 12971 1639 12977
rect 1581 12968 1593 12971
rect 1176 12940 1593 12968
rect 1176 12928 1182 12940
rect 1581 12937 1593 12940
rect 1627 12937 1639 12971
rect 1581 12931 1639 12937
rect 2041 12971 2099 12977
rect 2041 12937 2053 12971
rect 2087 12968 2099 12971
rect 2314 12968 2320 12980
rect 2087 12940 2320 12968
rect 2087 12937 2099 12940
rect 2041 12931 2099 12937
rect 2314 12928 2320 12940
rect 2372 12968 2378 12980
rect 2682 12968 2688 12980
rect 2372 12940 2688 12968
rect 2372 12928 2378 12940
rect 2682 12928 2688 12940
rect 2740 12968 2746 12980
rect 3142 12968 3148 12980
rect 2740 12940 3148 12968
rect 2740 12928 2746 12940
rect 3142 12928 3148 12940
rect 3200 12928 3206 12980
rect 6086 12928 6092 12980
rect 6144 12968 6150 12980
rect 6638 12968 6644 12980
rect 6144 12940 6644 12968
rect 6144 12928 6150 12940
rect 6638 12928 6644 12940
rect 6696 12968 6702 12980
rect 7837 12971 7895 12977
rect 7837 12968 7849 12971
rect 6696 12940 7849 12968
rect 6696 12928 6702 12940
rect 7837 12937 7849 12940
rect 7883 12968 7895 12971
rect 8294 12968 8300 12980
rect 7883 12940 8300 12968
rect 7883 12937 7895 12940
rect 7837 12931 7895 12937
rect 8294 12928 8300 12940
rect 8352 12968 8358 12980
rect 8389 12971 8447 12977
rect 8389 12968 8401 12971
rect 8352 12940 8401 12968
rect 8352 12928 8358 12940
rect 8389 12937 8401 12940
rect 8435 12937 8447 12971
rect 8389 12931 8447 12937
rect 9493 12971 9551 12977
rect 9493 12937 9505 12971
rect 9539 12968 9551 12971
rect 13633 12971 13691 12977
rect 13633 12968 13645 12971
rect 9539 12940 13645 12968
rect 9539 12937 9551 12940
rect 9493 12931 9551 12937
rect 13633 12937 13645 12940
rect 13679 12968 13691 12971
rect 13998 12968 14004 12980
rect 13679 12940 14004 12968
rect 13679 12937 13691 12940
rect 13633 12931 13691 12937
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 14734 12928 14740 12980
rect 14792 12968 14798 12980
rect 15289 12971 15347 12977
rect 15289 12968 15301 12971
rect 14792 12940 15301 12968
rect 14792 12928 14798 12940
rect 15289 12937 15301 12940
rect 15335 12937 15347 12971
rect 17126 12968 17132 12980
rect 17087 12940 17132 12968
rect 15289 12931 15347 12937
rect 17126 12928 17132 12940
rect 17184 12928 17190 12980
rect 19245 12971 19303 12977
rect 19245 12937 19257 12971
rect 19291 12968 19303 12971
rect 19426 12968 19432 12980
rect 19291 12940 19432 12968
rect 19291 12937 19303 12940
rect 19245 12931 19303 12937
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 21266 12968 21272 12980
rect 21227 12940 21272 12968
rect 21266 12928 21272 12940
rect 21324 12928 21330 12980
rect 5074 12900 5080 12912
rect 1412 12872 5080 12900
rect 1412 12773 1440 12872
rect 5074 12860 5080 12872
rect 5132 12860 5138 12912
rect 5350 12860 5356 12912
rect 5408 12900 5414 12912
rect 9769 12903 9827 12909
rect 9769 12900 9781 12903
rect 5408 12872 9781 12900
rect 5408 12860 5414 12872
rect 9769 12869 9781 12872
rect 9815 12869 9827 12903
rect 9769 12863 9827 12869
rect 11425 12903 11483 12909
rect 11425 12869 11437 12903
rect 11471 12900 11483 12903
rect 11974 12900 11980 12912
rect 11471 12872 11980 12900
rect 11471 12869 11483 12872
rect 11425 12863 11483 12869
rect 2409 12835 2467 12841
rect 2409 12801 2421 12835
rect 2455 12832 2467 12835
rect 2498 12832 2504 12844
rect 2455 12804 2504 12832
rect 2455 12801 2467 12804
rect 2409 12795 2467 12801
rect 2498 12792 2504 12804
rect 2556 12832 2562 12844
rect 2961 12835 3019 12841
rect 2961 12832 2973 12835
rect 2556 12804 2973 12832
rect 2556 12792 2562 12804
rect 2961 12801 2973 12804
rect 3007 12801 3019 12835
rect 2961 12795 3019 12801
rect 6362 12792 6368 12844
rect 6420 12832 6426 12844
rect 7193 12835 7251 12841
rect 7193 12832 7205 12835
rect 6420 12804 7205 12832
rect 6420 12792 6426 12804
rect 7193 12801 7205 12804
rect 7239 12801 7251 12835
rect 7193 12795 7251 12801
rect 8202 12792 8208 12844
rect 8260 12832 8266 12844
rect 8573 12835 8631 12841
rect 8573 12832 8585 12835
rect 8260 12804 8585 12832
rect 8260 12792 8266 12804
rect 8573 12801 8585 12804
rect 8619 12832 8631 12835
rect 9030 12832 9036 12844
rect 8619 12804 9036 12832
rect 8619 12801 8631 12804
rect 8573 12795 8631 12801
rect 9030 12792 9036 12804
rect 9088 12792 9094 12844
rect 9784 12832 9812 12863
rect 11974 12860 11980 12872
rect 12032 12860 12038 12912
rect 13538 12860 13544 12912
rect 13596 12900 13602 12912
rect 16114 12900 16120 12912
rect 13596 12872 14228 12900
rect 16075 12872 16120 12900
rect 13596 12860 13602 12872
rect 9784 12804 10824 12832
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12733 1455 12767
rect 1397 12727 1455 12733
rect 2590 12724 2596 12776
rect 2648 12764 2654 12776
rect 2869 12767 2927 12773
rect 2869 12764 2881 12767
rect 2648 12736 2881 12764
rect 2648 12724 2654 12736
rect 2869 12733 2881 12736
rect 2915 12733 2927 12767
rect 3142 12764 3148 12776
rect 3103 12736 3148 12764
rect 2869 12727 2927 12733
rect 2884 12696 2912 12727
rect 3142 12724 3148 12736
rect 3200 12724 3206 12776
rect 5077 12767 5135 12773
rect 5077 12764 5089 12767
rect 4540 12736 5089 12764
rect 2958 12696 2964 12708
rect 2884 12668 2964 12696
rect 2958 12656 2964 12668
rect 3016 12656 3022 12708
rect 3329 12631 3387 12637
rect 3329 12597 3341 12631
rect 3375 12628 3387 12631
rect 3418 12628 3424 12640
rect 3375 12600 3424 12628
rect 3375 12597 3387 12600
rect 3329 12591 3387 12597
rect 3418 12588 3424 12600
rect 3476 12588 3482 12640
rect 3602 12588 3608 12640
rect 3660 12628 3666 12640
rect 4065 12631 4123 12637
rect 4065 12628 4077 12631
rect 3660 12600 4077 12628
rect 3660 12588 3666 12600
rect 4065 12597 4077 12600
rect 4111 12628 4123 12631
rect 4154 12628 4160 12640
rect 4111 12600 4160 12628
rect 4111 12597 4123 12600
rect 4065 12591 4123 12597
rect 4154 12588 4160 12600
rect 4212 12588 4218 12640
rect 4430 12588 4436 12640
rect 4488 12628 4494 12640
rect 4540 12637 4568 12736
rect 5077 12733 5089 12736
rect 5123 12733 5135 12767
rect 5077 12727 5135 12733
rect 5537 12767 5595 12773
rect 5537 12733 5549 12767
rect 5583 12733 5595 12767
rect 5537 12727 5595 12733
rect 5552 12696 5580 12727
rect 9122 12724 9128 12776
rect 9180 12764 9186 12776
rect 9766 12764 9772 12776
rect 9180 12736 9772 12764
rect 9180 12724 9186 12736
rect 9766 12724 9772 12736
rect 9824 12764 9830 12776
rect 10137 12767 10195 12773
rect 10137 12764 10149 12767
rect 9824 12736 10149 12764
rect 9824 12724 9830 12736
rect 10137 12733 10149 12736
rect 10183 12764 10195 12767
rect 10321 12767 10379 12773
rect 10321 12764 10333 12767
rect 10183 12736 10333 12764
rect 10183 12733 10195 12736
rect 10137 12727 10195 12733
rect 10321 12733 10333 12736
rect 10367 12764 10379 12767
rect 10410 12764 10416 12776
rect 10367 12736 10416 12764
rect 10367 12733 10379 12736
rect 10321 12727 10379 12733
rect 10410 12724 10416 12736
rect 10468 12724 10474 12776
rect 10796 12773 10824 12804
rect 10962 12792 10968 12844
rect 11020 12832 11026 12844
rect 14200 12841 14228 12872
rect 16114 12860 16120 12872
rect 16172 12860 16178 12912
rect 21174 12860 21180 12912
rect 21232 12900 21238 12912
rect 22002 12900 22008 12912
rect 21232 12872 22008 12900
rect 21232 12860 21238 12872
rect 22002 12860 22008 12872
rect 22060 12900 22066 12912
rect 22465 12903 22523 12909
rect 22465 12900 22477 12903
rect 22060 12872 22477 12900
rect 22060 12860 22066 12872
rect 22465 12869 22477 12872
rect 22511 12869 22523 12903
rect 22465 12863 22523 12869
rect 11057 12835 11115 12841
rect 11057 12832 11069 12835
rect 11020 12804 11069 12832
rect 11020 12792 11026 12804
rect 11057 12801 11069 12804
rect 11103 12832 11115 12835
rect 11701 12835 11759 12841
rect 11701 12832 11713 12835
rect 11103 12804 11713 12832
rect 11103 12801 11115 12804
rect 11057 12795 11115 12801
rect 11701 12801 11713 12804
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 14185 12835 14243 12841
rect 14185 12801 14197 12835
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 15565 12835 15623 12841
rect 15565 12801 15577 12835
rect 15611 12832 15623 12835
rect 16577 12835 16635 12841
rect 16577 12832 16589 12835
rect 15611 12804 16589 12832
rect 15611 12801 15623 12804
rect 15565 12795 15623 12801
rect 16577 12801 16589 12804
rect 16623 12832 16635 12835
rect 24719 12835 24777 12841
rect 24719 12832 24731 12835
rect 16623 12804 24731 12832
rect 16623 12801 16635 12804
rect 16577 12795 16635 12801
rect 24719 12801 24731 12804
rect 24765 12801 24777 12835
rect 24719 12795 24777 12801
rect 10781 12767 10839 12773
rect 10781 12733 10793 12767
rect 10827 12764 10839 12767
rect 12437 12767 12495 12773
rect 12437 12764 12449 12767
rect 10827 12736 12449 12764
rect 10827 12733 10839 12736
rect 10781 12727 10839 12733
rect 12437 12733 12449 12736
rect 12483 12764 12495 12767
rect 13265 12767 13323 12773
rect 13265 12764 13277 12767
rect 12483 12736 13277 12764
rect 12483 12733 12495 12736
rect 12437 12727 12495 12733
rect 13265 12733 13277 12736
rect 13311 12733 13323 12767
rect 13265 12727 13323 12733
rect 17865 12767 17923 12773
rect 17865 12733 17877 12767
rect 17911 12764 17923 12767
rect 18322 12764 18328 12776
rect 17911 12736 18328 12764
rect 17911 12733 17923 12736
rect 17865 12727 17923 12733
rect 18322 12724 18328 12736
rect 18380 12724 18386 12776
rect 20070 12764 20076 12776
rect 20031 12736 20076 12764
rect 20070 12724 20076 12736
rect 20128 12724 20134 12776
rect 20993 12767 21051 12773
rect 20993 12733 21005 12767
rect 21039 12764 21051 12767
rect 21637 12767 21695 12773
rect 21637 12764 21649 12767
rect 21039 12736 21649 12764
rect 21039 12733 21051 12736
rect 20993 12727 21051 12733
rect 21637 12733 21649 12736
rect 21683 12733 21695 12767
rect 21637 12727 21695 12733
rect 24632 12767 24690 12773
rect 24632 12733 24644 12767
rect 24678 12764 24690 12767
rect 24678 12736 25176 12764
rect 24678 12733 24690 12736
rect 24632 12727 24690 12733
rect 5810 12696 5816 12708
rect 5000 12668 5580 12696
rect 5771 12668 5816 12696
rect 5000 12640 5028 12668
rect 5810 12656 5816 12668
rect 5868 12656 5874 12708
rect 6917 12699 6975 12705
rect 6917 12696 6929 12699
rect 6656 12668 6929 12696
rect 6656 12640 6684 12668
rect 6917 12665 6929 12668
rect 6963 12665 6975 12699
rect 6917 12659 6975 12665
rect 7006 12656 7012 12708
rect 7064 12696 7070 12708
rect 7064 12668 7109 12696
rect 7064 12656 7070 12668
rect 8294 12656 8300 12708
rect 8352 12696 8358 12708
rect 8894 12699 8952 12705
rect 8894 12696 8906 12699
rect 8352 12668 8906 12696
rect 8352 12656 8358 12668
rect 8894 12665 8906 12668
rect 8940 12665 8952 12699
rect 13906 12696 13912 12708
rect 13867 12668 13912 12696
rect 8894 12659 8952 12665
rect 13906 12656 13912 12668
rect 13964 12656 13970 12708
rect 13998 12656 14004 12708
rect 14056 12696 14062 12708
rect 14921 12699 14979 12705
rect 14921 12696 14933 12699
rect 14056 12668 14933 12696
rect 14056 12656 14062 12668
rect 14921 12665 14933 12668
rect 14967 12696 14979 12699
rect 15657 12699 15715 12705
rect 15657 12696 15669 12699
rect 14967 12668 15669 12696
rect 14967 12665 14979 12668
rect 14921 12659 14979 12665
rect 15657 12665 15669 12668
rect 15703 12696 15715 12699
rect 16206 12696 16212 12708
rect 15703 12668 16212 12696
rect 15703 12665 15715 12668
rect 15657 12659 15715 12665
rect 16206 12656 16212 12668
rect 16264 12656 16270 12708
rect 20394 12699 20452 12705
rect 20394 12696 20406 12699
rect 19904 12668 20406 12696
rect 4525 12631 4583 12637
rect 4525 12628 4537 12631
rect 4488 12600 4537 12628
rect 4488 12588 4494 12600
rect 4525 12597 4537 12600
rect 4571 12597 4583 12631
rect 4982 12628 4988 12640
rect 4943 12600 4988 12628
rect 4525 12591 4583 12597
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 6086 12628 6092 12640
rect 6047 12600 6092 12628
rect 6086 12588 6092 12600
rect 6144 12588 6150 12640
rect 6638 12628 6644 12640
rect 6599 12600 6644 12628
rect 6638 12588 6644 12600
rect 6696 12588 6702 12640
rect 12618 12628 12624 12640
rect 12579 12600 12624 12628
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 12989 12631 13047 12637
rect 12989 12597 13001 12631
rect 13035 12628 13047 12631
rect 13446 12628 13452 12640
rect 13035 12600 13452 12628
rect 13035 12597 13047 12600
rect 12989 12591 13047 12597
rect 13446 12588 13452 12600
rect 13504 12588 13510 12640
rect 17494 12628 17500 12640
rect 17407 12600 17500 12628
rect 17494 12588 17500 12600
rect 17552 12628 17558 12640
rect 17954 12628 17960 12640
rect 17552 12600 17960 12628
rect 17552 12588 17558 12600
rect 17954 12588 17960 12600
rect 18012 12588 18018 12640
rect 18690 12628 18696 12640
rect 18651 12600 18696 12628
rect 18690 12588 18696 12600
rect 18748 12628 18754 12640
rect 19904 12637 19932 12668
rect 20394 12665 20406 12668
rect 20440 12665 20452 12699
rect 20394 12659 20452 12665
rect 19521 12631 19579 12637
rect 19521 12628 19533 12631
rect 18748 12600 19533 12628
rect 18748 12588 18754 12600
rect 19521 12597 19533 12600
rect 19567 12628 19579 12631
rect 19889 12631 19947 12637
rect 19889 12628 19901 12631
rect 19567 12600 19901 12628
rect 19567 12597 19579 12600
rect 19521 12591 19579 12597
rect 19889 12597 19901 12600
rect 19935 12597 19947 12631
rect 21652 12628 21680 12727
rect 21910 12696 21916 12708
rect 21871 12668 21916 12696
rect 21910 12656 21916 12668
rect 21968 12656 21974 12708
rect 22005 12699 22063 12705
rect 22005 12665 22017 12699
rect 22051 12665 22063 12699
rect 22005 12659 22063 12665
rect 22020 12628 22048 12659
rect 25148 12637 25176 12736
rect 21652 12600 22048 12628
rect 25133 12631 25191 12637
rect 19889 12591 19947 12597
rect 25133 12597 25145 12631
rect 25179 12628 25191 12631
rect 26418 12628 26424 12640
rect 25179 12600 26424 12628
rect 25179 12597 25191 12600
rect 25133 12591 25191 12597
rect 26418 12588 26424 12600
rect 26476 12588 26482 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 3694 12384 3700 12436
rect 3752 12424 3758 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 3752 12396 3801 12424
rect 3752 12384 3758 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 4246 12424 4252 12436
rect 4207 12396 4252 12424
rect 3789 12387 3847 12393
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 4706 12424 4712 12436
rect 4667 12396 4712 12424
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 5074 12424 5080 12436
rect 5035 12396 5080 12424
rect 5074 12384 5080 12396
rect 5132 12384 5138 12436
rect 5810 12384 5816 12436
rect 5868 12424 5874 12436
rect 6181 12427 6239 12433
rect 6181 12424 6193 12427
rect 5868 12396 6193 12424
rect 5868 12384 5874 12396
rect 6181 12393 6193 12396
rect 6227 12393 6239 12427
rect 7190 12424 7196 12436
rect 7151 12396 7196 12424
rect 6181 12387 6239 12393
rect 7190 12384 7196 12396
rect 7248 12384 7254 12436
rect 7834 12424 7840 12436
rect 7795 12396 7840 12424
rect 7834 12384 7840 12396
rect 7892 12384 7898 12436
rect 9030 12424 9036 12436
rect 8991 12396 9036 12424
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 10778 12424 10784 12436
rect 10739 12396 10784 12424
rect 10778 12384 10784 12396
rect 10836 12384 10842 12436
rect 11422 12424 11428 12436
rect 11383 12396 11428 12424
rect 11422 12384 11428 12396
rect 11480 12384 11486 12436
rect 15473 12427 15531 12433
rect 15473 12393 15485 12427
rect 15519 12424 15531 12427
rect 16298 12424 16304 12436
rect 15519 12396 16304 12424
rect 15519 12393 15531 12396
rect 15473 12387 15531 12393
rect 16298 12384 16304 12396
rect 16356 12384 16362 12436
rect 19518 12424 19524 12436
rect 19479 12396 19524 12424
rect 19518 12384 19524 12396
rect 19576 12384 19582 12436
rect 20622 12424 20628 12436
rect 20583 12396 20628 12424
rect 20622 12384 20628 12396
rect 20680 12424 20686 12436
rect 20680 12396 21680 12424
rect 20680 12384 20686 12396
rect 3970 12356 3976 12368
rect 2976 12328 3976 12356
rect 1302 12248 1308 12300
rect 1360 12288 1366 12300
rect 2976 12297 3004 12328
rect 3970 12316 3976 12328
rect 4028 12356 4034 12368
rect 4614 12356 4620 12368
rect 4028 12328 4620 12356
rect 4028 12316 4034 12328
rect 4614 12316 4620 12328
rect 4672 12316 4678 12368
rect 6270 12356 6276 12368
rect 5092 12328 6276 12356
rect 1489 12291 1547 12297
rect 1489 12288 1501 12291
rect 1360 12260 1501 12288
rect 1360 12248 1366 12260
rect 1489 12257 1501 12260
rect 1535 12257 1547 12291
rect 1489 12251 1547 12257
rect 2961 12291 3019 12297
rect 2961 12257 2973 12291
rect 3007 12257 3019 12291
rect 4062 12288 4068 12300
rect 4023 12260 4068 12288
rect 2961 12251 3019 12257
rect 4062 12248 4068 12260
rect 4120 12248 4126 12300
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12220 2191 12223
rect 2314 12220 2320 12232
rect 2179 12192 2320 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 2314 12180 2320 12192
rect 2372 12220 2378 12232
rect 2866 12220 2872 12232
rect 2372 12192 2872 12220
rect 2372 12180 2378 12192
rect 2866 12180 2872 12192
rect 2924 12180 2930 12232
rect 5092 12220 5120 12328
rect 5368 12297 5396 12328
rect 6270 12316 6276 12328
rect 6328 12316 6334 12368
rect 7208 12356 7236 12384
rect 10505 12359 10563 12365
rect 7208 12328 10364 12356
rect 5353 12291 5411 12297
rect 5353 12257 5365 12291
rect 5399 12257 5411 12291
rect 5353 12251 5411 12257
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 5629 12291 5687 12297
rect 5629 12288 5641 12291
rect 5592 12260 5641 12288
rect 5592 12248 5598 12260
rect 5629 12257 5641 12260
rect 5675 12257 5687 12291
rect 7006 12288 7012 12300
rect 6967 12260 7012 12288
rect 5629 12251 5687 12257
rect 7006 12248 7012 12260
rect 7064 12248 7070 12300
rect 8021 12291 8079 12297
rect 8021 12288 8033 12291
rect 7116 12260 8033 12288
rect 4126 12192 5120 12220
rect 5905 12223 5963 12229
rect 2958 12152 2964 12164
rect 2608 12124 2964 12152
rect 2038 12044 2044 12096
rect 2096 12084 2102 12096
rect 2608 12093 2636 12124
rect 2958 12112 2964 12124
rect 3016 12152 3022 12164
rect 3421 12155 3479 12161
rect 3421 12152 3433 12155
rect 3016 12124 3433 12152
rect 3016 12112 3022 12124
rect 3421 12121 3433 12124
rect 3467 12121 3479 12155
rect 3421 12115 3479 12121
rect 2593 12087 2651 12093
rect 2593 12084 2605 12087
rect 2096 12056 2605 12084
rect 2096 12044 2102 12056
rect 2593 12053 2605 12056
rect 2639 12053 2651 12087
rect 2593 12047 2651 12053
rect 3145 12087 3203 12093
rect 3145 12053 3157 12087
rect 3191 12084 3203 12087
rect 4126 12084 4154 12192
rect 5905 12189 5917 12223
rect 5951 12220 5963 12223
rect 5994 12220 6000 12232
rect 5951 12192 6000 12220
rect 5951 12189 5963 12192
rect 5905 12183 5963 12189
rect 5994 12180 6000 12192
rect 6052 12180 6058 12232
rect 4430 12112 4436 12164
rect 4488 12152 4494 12164
rect 7116 12152 7144 12260
rect 8021 12257 8033 12260
rect 8067 12288 8079 12291
rect 8202 12288 8208 12300
rect 8067 12260 8208 12288
rect 8067 12257 8079 12260
rect 8021 12251 8079 12257
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 8386 12248 8392 12300
rect 8444 12288 8450 12300
rect 8481 12291 8539 12297
rect 8481 12288 8493 12291
rect 8444 12260 8493 12288
rect 8444 12248 8450 12260
rect 8481 12257 8493 12260
rect 8527 12257 8539 12291
rect 9766 12288 9772 12300
rect 9727 12260 9772 12288
rect 8481 12251 8539 12257
rect 9766 12248 9772 12260
rect 9824 12248 9830 12300
rect 10229 12291 10287 12297
rect 10229 12257 10241 12291
rect 10275 12257 10287 12291
rect 10336 12288 10364 12328
rect 10505 12325 10517 12359
rect 10551 12356 10563 12359
rect 12710 12356 12716 12368
rect 10551 12328 12716 12356
rect 10551 12325 10563 12328
rect 10505 12319 10563 12325
rect 12710 12316 12716 12328
rect 12768 12316 12774 12368
rect 13814 12316 13820 12368
rect 13872 12356 13878 12368
rect 16482 12356 16488 12368
rect 13872 12328 13917 12356
rect 16443 12328 16488 12356
rect 13872 12316 13878 12328
rect 16482 12316 16488 12328
rect 16540 12316 16546 12368
rect 18595 12359 18653 12365
rect 18595 12325 18607 12359
rect 18641 12356 18653 12359
rect 18690 12356 18696 12368
rect 18641 12328 18696 12356
rect 18641 12325 18653 12328
rect 18595 12319 18653 12325
rect 18690 12316 18696 12328
rect 18748 12316 18754 12368
rect 21082 12356 21088 12368
rect 21043 12328 21088 12356
rect 21082 12316 21088 12328
rect 21140 12316 21146 12368
rect 21652 12365 21680 12396
rect 21637 12359 21695 12365
rect 21637 12325 21649 12359
rect 21683 12325 21695 12359
rect 21637 12319 21695 12325
rect 11333 12291 11391 12297
rect 11333 12288 11345 12291
rect 10336 12260 11345 12288
rect 10229 12251 10287 12257
rect 11333 12257 11345 12260
rect 11379 12288 11391 12291
rect 11698 12288 11704 12300
rect 11379 12260 11704 12288
rect 11379 12257 11391 12260
rect 11333 12251 11391 12257
rect 8754 12220 8760 12232
rect 8715 12192 8760 12220
rect 8754 12180 8760 12192
rect 8812 12180 8818 12232
rect 9398 12180 9404 12232
rect 9456 12220 9462 12232
rect 10244 12220 10272 12251
rect 11698 12248 11704 12260
rect 11756 12248 11762 12300
rect 11790 12248 11796 12300
rect 11848 12288 11854 12300
rect 11848 12260 11893 12288
rect 11848 12248 11854 12260
rect 14642 12248 14648 12300
rect 14700 12288 14706 12300
rect 15289 12291 15347 12297
rect 15289 12288 15301 12291
rect 14700 12260 15301 12288
rect 14700 12248 14706 12260
rect 15289 12257 15301 12260
rect 15335 12257 15347 12291
rect 15289 12251 15347 12257
rect 18138 12248 18144 12300
rect 18196 12288 18202 12300
rect 18233 12291 18291 12297
rect 18233 12288 18245 12291
rect 18196 12260 18245 12288
rect 18196 12248 18202 12260
rect 18233 12257 18245 12260
rect 18279 12257 18291 12291
rect 18233 12251 18291 12257
rect 13722 12220 13728 12232
rect 9456 12192 10272 12220
rect 13683 12192 13728 12220
rect 9456 12180 9462 12192
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 14090 12220 14096 12232
rect 14051 12192 14096 12220
rect 14090 12180 14096 12192
rect 14148 12180 14154 12232
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12220 16451 12223
rect 16850 12220 16856 12232
rect 16439 12192 16856 12220
rect 16439 12189 16451 12192
rect 16393 12183 16451 12189
rect 16850 12180 16856 12192
rect 16908 12220 16914 12232
rect 20993 12223 21051 12229
rect 16908 12192 18638 12220
rect 16908 12180 16914 12192
rect 4488 12124 7144 12152
rect 4488 12112 4494 12124
rect 12618 12112 12624 12164
rect 12676 12152 12682 12164
rect 16942 12152 16948 12164
rect 12676 12124 16804 12152
rect 16903 12124 16948 12152
rect 12676 12112 12682 12124
rect 6914 12084 6920 12096
rect 3191 12056 4154 12084
rect 6875 12056 6920 12084
rect 3191 12053 3203 12056
rect 3145 12047 3203 12053
rect 6914 12044 6920 12056
rect 6972 12044 6978 12096
rect 13078 12084 13084 12096
rect 13039 12056 13084 12084
rect 13078 12044 13084 12056
rect 13136 12044 13142 12096
rect 15841 12087 15899 12093
rect 15841 12053 15853 12087
rect 15887 12084 15899 12087
rect 15930 12084 15936 12096
rect 15887 12056 15936 12084
rect 15887 12053 15899 12056
rect 15841 12047 15899 12053
rect 15930 12044 15936 12056
rect 15988 12044 15994 12096
rect 16776 12084 16804 12124
rect 16942 12112 16948 12124
rect 17000 12112 17006 12164
rect 18610 12152 18638 12192
rect 20993 12189 21005 12223
rect 21039 12220 21051 12223
rect 21358 12220 21364 12232
rect 21039 12192 21364 12220
rect 21039 12189 21051 12192
rect 20993 12183 21051 12189
rect 21358 12180 21364 12192
rect 21416 12180 21422 12232
rect 22738 12152 22744 12164
rect 18610 12124 22744 12152
rect 22738 12112 22744 12124
rect 22796 12112 22802 12164
rect 19058 12084 19064 12096
rect 16776 12056 19064 12084
rect 19058 12044 19064 12056
rect 19116 12044 19122 12096
rect 19153 12087 19211 12093
rect 19153 12053 19165 12087
rect 19199 12084 19211 12087
rect 19242 12084 19248 12096
rect 19199 12056 19248 12084
rect 19199 12053 19211 12056
rect 19153 12047 19211 12053
rect 19242 12044 19248 12056
rect 19300 12044 19306 12096
rect 20070 12084 20076 12096
rect 20031 12056 20076 12084
rect 20070 12044 20076 12056
rect 20128 12044 20134 12096
rect 21910 12084 21916 12096
rect 21871 12056 21916 12084
rect 21910 12044 21916 12056
rect 21968 12044 21974 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2038 11840 2044 11892
rect 2096 11880 2102 11892
rect 3053 11883 3111 11889
rect 3053 11880 3065 11883
rect 2096 11852 3065 11880
rect 2096 11840 2102 11852
rect 3053 11849 3065 11852
rect 3099 11849 3111 11883
rect 3053 11843 3111 11849
rect 4062 11840 4068 11892
rect 4120 11880 4126 11892
rect 4522 11880 4528 11892
rect 4120 11852 4528 11880
rect 4120 11840 4126 11852
rect 4522 11840 4528 11852
rect 4580 11880 4586 11892
rect 4617 11883 4675 11889
rect 4617 11880 4629 11883
rect 4580 11852 4629 11880
rect 4580 11840 4586 11852
rect 4617 11849 4629 11852
rect 4663 11849 4675 11883
rect 6270 11880 6276 11892
rect 6231 11852 6276 11880
rect 4617 11843 4675 11849
rect 6270 11840 6276 11852
rect 6328 11840 6334 11892
rect 11698 11840 11704 11892
rect 11756 11880 11762 11892
rect 11793 11883 11851 11889
rect 11793 11880 11805 11883
rect 11756 11852 11805 11880
rect 11756 11840 11762 11852
rect 11793 11849 11805 11852
rect 11839 11849 11851 11883
rect 11793 11843 11851 11849
rect 13814 11840 13820 11892
rect 13872 11880 13878 11892
rect 13909 11883 13967 11889
rect 13909 11880 13921 11883
rect 13872 11852 13921 11880
rect 13872 11840 13878 11852
rect 13909 11849 13921 11852
rect 13955 11849 13967 11883
rect 14642 11880 14648 11892
rect 14603 11852 14648 11880
rect 13909 11843 13967 11849
rect 14642 11840 14648 11852
rect 14700 11840 14706 11892
rect 15562 11840 15568 11892
rect 15620 11880 15626 11892
rect 16117 11883 16175 11889
rect 16117 11880 16129 11883
rect 15620 11852 16129 11880
rect 15620 11840 15626 11852
rect 16117 11849 16129 11852
rect 16163 11880 16175 11883
rect 16482 11880 16488 11892
rect 16163 11852 16488 11880
rect 16163 11849 16175 11852
rect 16117 11843 16175 11849
rect 16482 11840 16488 11852
rect 16540 11840 16546 11892
rect 16850 11880 16856 11892
rect 16811 11852 16856 11880
rect 16850 11840 16856 11852
rect 16908 11840 16914 11892
rect 17865 11883 17923 11889
rect 17865 11849 17877 11883
rect 17911 11880 17923 11883
rect 18138 11880 18144 11892
rect 17911 11852 18144 11880
rect 17911 11849 17923 11852
rect 17865 11843 17923 11849
rect 18138 11840 18144 11852
rect 18196 11840 18202 11892
rect 18325 11883 18383 11889
rect 18325 11849 18337 11883
rect 18371 11880 18383 11883
rect 18690 11880 18696 11892
rect 18371 11852 18696 11880
rect 18371 11849 18383 11852
rect 18325 11843 18383 11849
rect 4982 11772 4988 11824
rect 5040 11812 5046 11824
rect 5077 11815 5135 11821
rect 5077 11812 5089 11815
rect 5040 11784 5089 11812
rect 5040 11772 5046 11784
rect 5077 11781 5089 11784
rect 5123 11812 5135 11815
rect 5123 11784 5580 11812
rect 5123 11781 5135 11784
rect 5077 11775 5135 11781
rect 5552 11756 5580 11784
rect 8294 11772 8300 11824
rect 8352 11812 8358 11824
rect 8573 11815 8631 11821
rect 8573 11812 8585 11815
rect 8352 11784 8585 11812
rect 8352 11772 8358 11784
rect 8573 11781 8585 11784
rect 8619 11781 8631 11815
rect 12618 11812 12624 11824
rect 8573 11775 8631 11781
rect 10796 11784 12624 11812
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11744 2835 11747
rect 5442 11744 5448 11756
rect 2823 11716 5448 11744
rect 2823 11713 2835 11716
rect 2777 11707 2835 11713
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 5534 11704 5540 11756
rect 5592 11744 5598 11756
rect 5592 11716 6960 11744
rect 5592 11704 5598 11716
rect 1578 11636 1584 11688
rect 1636 11676 1642 11688
rect 2038 11676 2044 11688
rect 1636 11648 2044 11676
rect 1636 11636 1642 11648
rect 2038 11636 2044 11648
rect 2096 11636 2102 11688
rect 2130 11636 2136 11688
rect 2188 11676 2194 11688
rect 2317 11679 2375 11685
rect 2188 11648 2233 11676
rect 2188 11636 2194 11648
rect 2317 11645 2329 11679
rect 2363 11676 2375 11679
rect 2406 11676 2412 11688
rect 2363 11648 2412 11676
rect 2363 11645 2375 11648
rect 2317 11639 2375 11645
rect 2406 11636 2412 11648
rect 2464 11636 2470 11688
rect 3694 11676 3700 11688
rect 3655 11648 3700 11676
rect 3694 11636 3700 11648
rect 3752 11636 3758 11688
rect 5736 11685 5764 11716
rect 6932 11688 6960 11716
rect 4065 11679 4123 11685
rect 4065 11645 4077 11679
rect 4111 11645 4123 11679
rect 4065 11639 4123 11645
rect 5353 11679 5411 11685
rect 5353 11645 5365 11679
rect 5399 11645 5411 11679
rect 5353 11639 5411 11645
rect 5721 11679 5779 11685
rect 5721 11645 5733 11679
rect 5767 11645 5779 11679
rect 5721 11639 5779 11645
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11645 6883 11679
rect 6825 11639 6883 11645
rect 2866 11568 2872 11620
rect 2924 11608 2930 11620
rect 3421 11611 3479 11617
rect 3421 11608 3433 11611
rect 2924 11580 3433 11608
rect 2924 11568 2930 11580
rect 3421 11577 3433 11580
rect 3467 11608 3479 11611
rect 4080 11608 4108 11639
rect 4982 11608 4988 11620
rect 3467 11580 4988 11608
rect 3467 11577 3479 11580
rect 3421 11571 3479 11577
rect 4982 11568 4988 11580
rect 5040 11568 5046 11620
rect 5368 11608 5396 11639
rect 5442 11608 5448 11620
rect 5368 11580 5448 11608
rect 5442 11568 5448 11580
rect 5500 11568 5506 11620
rect 5902 11608 5908 11620
rect 5863 11580 5908 11608
rect 5902 11568 5908 11580
rect 5960 11568 5966 11620
rect 6641 11611 6699 11617
rect 6641 11577 6653 11611
rect 6687 11608 6699 11611
rect 6840 11608 6868 11639
rect 6914 11636 6920 11688
rect 6972 11676 6978 11688
rect 7285 11679 7343 11685
rect 7285 11676 7297 11679
rect 6972 11648 7297 11676
rect 6972 11636 6978 11648
rect 7285 11645 7297 11648
rect 7331 11645 7343 11679
rect 7285 11639 7343 11645
rect 7926 11608 7932 11620
rect 6687 11580 7932 11608
rect 6687 11577 6699 11580
rect 6641 11571 6699 11577
rect 7926 11568 7932 11580
rect 7984 11568 7990 11620
rect 8588 11608 8616 11775
rect 8754 11744 8760 11756
rect 8715 11716 8760 11744
rect 8754 11704 8760 11716
rect 8812 11704 8818 11756
rect 10796 11685 10824 11784
rect 12618 11772 12624 11784
rect 12676 11772 12682 11824
rect 13722 11772 13728 11824
rect 13780 11812 13786 11824
rect 14369 11815 14427 11821
rect 14369 11812 14381 11815
rect 13780 11784 14381 11812
rect 13780 11772 13786 11784
rect 14369 11781 14381 11784
rect 14415 11812 14427 11815
rect 16942 11812 16948 11824
rect 14415 11784 16948 11812
rect 14415 11781 14427 11784
rect 14369 11775 14427 11781
rect 16942 11772 16948 11784
rect 17000 11772 17006 11824
rect 17221 11815 17279 11821
rect 17221 11781 17233 11815
rect 17267 11812 17279 11815
rect 18340 11812 18368 11843
rect 18690 11840 18696 11852
rect 18748 11840 18754 11892
rect 19242 11840 19248 11892
rect 19300 11880 19306 11892
rect 19889 11883 19947 11889
rect 19889 11880 19901 11883
rect 19300 11852 19901 11880
rect 19300 11840 19306 11852
rect 19889 11849 19901 11852
rect 19935 11880 19947 11883
rect 21082 11880 21088 11892
rect 19935 11852 21088 11880
rect 19935 11849 19947 11852
rect 19889 11843 19947 11849
rect 21082 11840 21088 11852
rect 21140 11840 21146 11892
rect 22002 11880 22008 11892
rect 21963 11852 22008 11880
rect 22002 11840 22008 11852
rect 22060 11840 22066 11892
rect 17267 11784 18368 11812
rect 17267 11781 17279 11784
rect 17221 11775 17279 11781
rect 11517 11747 11575 11753
rect 11517 11713 11529 11747
rect 11563 11744 11575 11747
rect 12713 11747 12771 11753
rect 12713 11744 12725 11747
rect 11563 11716 12725 11744
rect 11563 11713 11575 11716
rect 11517 11707 11575 11713
rect 12713 11713 12725 11716
rect 12759 11744 12771 11747
rect 13078 11744 13084 11756
rect 12759 11716 13084 11744
rect 12759 11713 12771 11716
rect 12713 11707 12771 11713
rect 13078 11704 13084 11716
rect 13136 11704 13142 11756
rect 13906 11704 13912 11756
rect 13964 11744 13970 11756
rect 17083 11747 17141 11753
rect 17083 11744 17095 11747
rect 13964 11716 17095 11744
rect 13964 11704 13970 11716
rect 17083 11713 17095 11716
rect 17129 11713 17141 11747
rect 18506 11744 18512 11756
rect 17083 11707 17141 11713
rect 17420 11716 18512 11744
rect 10689 11679 10747 11685
rect 10689 11645 10701 11679
rect 10735 11676 10747 11679
rect 10781 11679 10839 11685
rect 10781 11676 10793 11679
rect 10735 11648 10793 11676
rect 10735 11645 10747 11648
rect 10689 11639 10747 11645
rect 10781 11645 10793 11648
rect 10827 11645 10839 11679
rect 10781 11639 10839 11645
rect 10870 11636 10876 11688
rect 10928 11676 10934 11688
rect 11241 11679 11299 11685
rect 11241 11676 11253 11679
rect 10928 11648 11253 11676
rect 10928 11636 10934 11648
rect 11241 11645 11253 11648
rect 11287 11676 11299 11679
rect 11790 11676 11796 11688
rect 11287 11648 11796 11676
rect 11287 11645 11299 11648
rect 11241 11639 11299 11645
rect 11790 11636 11796 11648
rect 11848 11676 11854 11688
rect 12161 11679 12219 11685
rect 12161 11676 12173 11679
rect 11848 11648 12173 11676
rect 11848 11636 11854 11648
rect 12161 11645 12173 11648
rect 12207 11676 12219 11679
rect 14734 11676 14740 11688
rect 12207 11648 14740 11676
rect 12207 11645 12219 11648
rect 12161 11639 12219 11645
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 15197 11679 15255 11685
rect 15197 11645 15209 11679
rect 15243 11676 15255 11679
rect 15286 11676 15292 11688
rect 15243 11648 15292 11676
rect 15243 11645 15255 11648
rect 15197 11639 15255 11645
rect 15286 11636 15292 11648
rect 15344 11636 15350 11688
rect 16850 11636 16856 11688
rect 16908 11676 16914 11688
rect 17420 11685 17448 11716
rect 18506 11704 18512 11716
rect 18564 11704 18570 11756
rect 19150 11744 19156 11756
rect 19111 11716 19156 11744
rect 19150 11704 19156 11716
rect 19208 11704 19214 11756
rect 20717 11747 20775 11753
rect 20717 11713 20729 11747
rect 20763 11744 20775 11747
rect 21910 11744 21916 11756
rect 20763 11716 21916 11744
rect 20763 11713 20775 11716
rect 20717 11707 20775 11713
rect 21910 11704 21916 11716
rect 21968 11704 21974 11756
rect 16980 11679 17038 11685
rect 16980 11676 16992 11679
rect 16908 11648 16992 11676
rect 16908 11636 16914 11648
rect 16980 11645 16992 11648
rect 17026 11676 17038 11679
rect 17405 11679 17463 11685
rect 17405 11676 17417 11679
rect 17026 11648 17417 11676
rect 17026 11645 17038 11648
rect 16980 11639 17038 11645
rect 17405 11645 17417 11648
rect 17451 11645 17463 11679
rect 17405 11639 17463 11645
rect 21612 11679 21670 11685
rect 21612 11645 21624 11679
rect 21658 11676 21670 11679
rect 22002 11676 22008 11688
rect 21658 11648 22008 11676
rect 21658 11645 21670 11648
rect 21612 11639 21670 11645
rect 22002 11636 22008 11648
rect 22060 11636 22066 11688
rect 9078 11611 9136 11617
rect 9078 11608 9090 11611
rect 8588 11580 9090 11608
rect 9078 11577 9090 11580
rect 9124 11577 9136 11611
rect 9078 11571 9136 11577
rect 9214 11568 9220 11620
rect 9272 11608 9278 11620
rect 9766 11608 9772 11620
rect 9272 11580 9772 11608
rect 9272 11568 9278 11580
rect 9766 11568 9772 11580
rect 9824 11608 9830 11620
rect 9953 11611 10011 11617
rect 9953 11608 9965 11611
rect 9824 11580 9965 11608
rect 9824 11568 9830 11580
rect 9953 11577 9965 11580
rect 9999 11577 10011 11611
rect 9953 11571 10011 11577
rect 13446 11568 13452 11620
rect 13504 11608 13510 11620
rect 15105 11611 15163 11617
rect 15105 11608 15117 11611
rect 13504 11580 15117 11608
rect 13504 11568 13510 11580
rect 15105 11577 15117 11580
rect 15151 11608 15163 11611
rect 15559 11611 15617 11617
rect 15559 11608 15571 11611
rect 15151 11580 15571 11608
rect 15151 11577 15163 11580
rect 15105 11571 15163 11577
rect 15559 11577 15571 11580
rect 15605 11608 15617 11611
rect 16390 11608 16396 11620
rect 15605 11580 16396 11608
rect 15605 11577 15617 11580
rect 15559 11571 15617 11577
rect 16390 11568 16396 11580
rect 16448 11608 16454 11620
rect 17221 11611 17279 11617
rect 17221 11608 17233 11611
rect 16448 11580 17233 11608
rect 16448 11568 16454 11580
rect 17221 11577 17233 11580
rect 17267 11577 17279 11611
rect 18506 11608 18512 11620
rect 18467 11580 18512 11608
rect 17221 11571 17279 11577
rect 18506 11568 18512 11580
rect 18564 11568 18570 11620
rect 18598 11568 18604 11620
rect 18656 11608 18662 11620
rect 19242 11608 19248 11620
rect 18656 11580 19248 11608
rect 18656 11568 18662 11580
rect 19242 11568 19248 11580
rect 19300 11568 19306 11620
rect 19521 11611 19579 11617
rect 19521 11577 19533 11611
rect 19567 11608 19579 11611
rect 20073 11611 20131 11617
rect 20073 11608 20085 11611
rect 19567 11580 20085 11608
rect 19567 11577 19579 11580
rect 19521 11571 19579 11577
rect 20073 11577 20085 11580
rect 20119 11577 20131 11611
rect 20073 11571 20131 11577
rect 20165 11611 20223 11617
rect 20165 11577 20177 11611
rect 20211 11608 20223 11611
rect 21082 11608 21088 11620
rect 20211 11580 21088 11608
rect 20211 11577 20223 11580
rect 20165 11571 20223 11577
rect 1302 11500 1308 11552
rect 1360 11540 1366 11552
rect 1581 11543 1639 11549
rect 1581 11540 1593 11543
rect 1360 11512 1593 11540
rect 1360 11500 1366 11512
rect 1581 11509 1593 11512
rect 1627 11509 1639 11543
rect 3878 11540 3884 11552
rect 3839 11512 3884 11540
rect 1581 11503 1639 11509
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 6730 11500 6736 11552
rect 6788 11540 6794 11552
rect 6917 11543 6975 11549
rect 6917 11540 6929 11543
rect 6788 11512 6929 11540
rect 6788 11500 6794 11512
rect 6917 11509 6929 11512
rect 6963 11509 6975 11543
rect 6917 11503 6975 11509
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 8021 11543 8079 11549
rect 8021 11540 8033 11543
rect 7524 11512 8033 11540
rect 7524 11500 7530 11512
rect 8021 11509 8033 11512
rect 8067 11540 8079 11543
rect 8386 11540 8392 11552
rect 8067 11512 8392 11540
rect 8067 11509 8079 11512
rect 8021 11503 8079 11509
rect 8386 11500 8392 11512
rect 8444 11500 8450 11552
rect 9677 11543 9735 11549
rect 9677 11509 9689 11543
rect 9723 11540 9735 11543
rect 9858 11540 9864 11552
rect 9723 11512 9864 11540
rect 9723 11509 9735 11512
rect 9677 11503 9735 11509
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 13081 11543 13139 11549
rect 13081 11509 13093 11543
rect 13127 11540 13139 11543
rect 13464 11540 13492 11568
rect 13630 11540 13636 11552
rect 13127 11512 13492 11540
rect 13591 11512 13636 11540
rect 13127 11509 13139 11512
rect 13081 11503 13139 11509
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 20088 11540 20116 11571
rect 21082 11568 21088 11580
rect 21140 11568 21146 11620
rect 20898 11540 20904 11552
rect 20088 11512 20904 11540
rect 20898 11500 20904 11512
rect 20956 11500 20962 11552
rect 21358 11540 21364 11552
rect 21319 11512 21364 11540
rect 21358 11500 21364 11512
rect 21416 11500 21422 11552
rect 21683 11543 21741 11549
rect 21683 11509 21695 11543
rect 21729 11540 21741 11543
rect 21910 11540 21916 11552
rect 21729 11512 21916 11540
rect 21729 11509 21741 11512
rect 21683 11503 21741 11509
rect 21910 11500 21916 11512
rect 21968 11500 21974 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 3881 11339 3939 11345
rect 1627 11308 2452 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 1394 11200 1400 11212
rect 1355 11172 1400 11200
rect 1394 11160 1400 11172
rect 1452 11160 1458 11212
rect 2424 11209 2452 11308
rect 3881 11305 3893 11339
rect 3927 11336 3939 11339
rect 3970 11336 3976 11348
rect 3927 11308 3976 11336
rect 3927 11305 3939 11308
rect 3881 11299 3939 11305
rect 3970 11296 3976 11308
rect 4028 11296 4034 11348
rect 5261 11339 5319 11345
rect 5261 11305 5273 11339
rect 5307 11336 5319 11339
rect 5534 11336 5540 11348
rect 5307 11308 5540 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 5902 11296 5908 11348
rect 5960 11336 5966 11348
rect 6822 11336 6828 11348
rect 5960 11308 6828 11336
rect 5960 11296 5966 11308
rect 6822 11296 6828 11308
rect 6880 11336 6886 11348
rect 7377 11339 7435 11345
rect 7377 11336 7389 11339
rect 6880 11308 7389 11336
rect 6880 11296 6886 11308
rect 7377 11305 7389 11308
rect 7423 11305 7435 11339
rect 7834 11336 7840 11348
rect 7795 11308 7840 11336
rect 7377 11299 7435 11305
rect 7834 11296 7840 11308
rect 7892 11296 7898 11348
rect 8754 11296 8760 11348
rect 8812 11336 8818 11348
rect 8941 11339 8999 11345
rect 8941 11336 8953 11339
rect 8812 11308 8953 11336
rect 8812 11296 8818 11308
rect 8941 11305 8953 11308
rect 8987 11305 8999 11339
rect 12805 11339 12863 11345
rect 12805 11336 12817 11339
rect 8941 11299 8999 11305
rect 11710 11308 12817 11336
rect 4246 11268 4252 11280
rect 4207 11240 4252 11268
rect 4246 11228 4252 11240
rect 4304 11228 4310 11280
rect 6086 11268 6092 11280
rect 6047 11240 6092 11268
rect 6086 11228 6092 11240
rect 6144 11228 6150 11280
rect 6270 11228 6276 11280
rect 6328 11268 6334 11280
rect 9398 11268 9404 11280
rect 6328 11240 9404 11268
rect 6328 11228 6334 11240
rect 9398 11228 9404 11240
rect 9456 11228 9462 11280
rect 9858 11268 9864 11280
rect 9819 11240 9864 11268
rect 9858 11228 9864 11240
rect 9916 11228 9922 11280
rect 11710 11277 11738 11308
rect 12805 11305 12817 11308
rect 12851 11336 12863 11339
rect 13446 11336 13452 11348
rect 12851 11308 13452 11336
rect 12851 11305 12863 11308
rect 12805 11299 12863 11305
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 13814 11296 13820 11348
rect 13872 11336 13878 11348
rect 14001 11339 14059 11345
rect 14001 11336 14013 11339
rect 13872 11308 14013 11336
rect 13872 11296 13878 11308
rect 14001 11305 14013 11308
rect 14047 11305 14059 11339
rect 14001 11299 14059 11305
rect 15286 11296 15292 11348
rect 15344 11336 15350 11348
rect 15473 11339 15531 11345
rect 15473 11336 15485 11339
rect 15344 11308 15485 11336
rect 15344 11296 15350 11308
rect 15473 11305 15485 11308
rect 15519 11305 15531 11339
rect 17589 11339 17647 11345
rect 17589 11336 17601 11339
rect 15473 11299 15531 11305
rect 15764 11308 17601 11336
rect 11695 11271 11753 11277
rect 11695 11237 11707 11271
rect 11741 11237 11753 11271
rect 11695 11231 11753 11237
rect 15764 11212 15792 11308
rect 17589 11305 17601 11308
rect 17635 11305 17647 11339
rect 17589 11299 17647 11305
rect 18506 11296 18512 11348
rect 18564 11336 18570 11348
rect 18877 11339 18935 11345
rect 18877 11336 18889 11339
rect 18564 11308 18889 11336
rect 18564 11296 18570 11308
rect 18877 11305 18889 11308
rect 18923 11336 18935 11339
rect 19518 11336 19524 11348
rect 18923 11308 19524 11336
rect 18923 11305 18935 11308
rect 18877 11299 18935 11305
rect 19518 11296 19524 11308
rect 19576 11296 19582 11348
rect 20898 11296 20904 11348
rect 20956 11336 20962 11348
rect 21039 11339 21097 11345
rect 21039 11336 21051 11339
rect 20956 11308 21051 11336
rect 20956 11296 20962 11308
rect 21039 11305 21051 11308
rect 21085 11305 21097 11339
rect 21039 11299 21097 11305
rect 16111 11271 16169 11277
rect 16111 11237 16123 11271
rect 16157 11268 16169 11271
rect 16390 11268 16396 11280
rect 16157 11240 16396 11268
rect 16157 11237 16169 11240
rect 16111 11231 16169 11237
rect 16390 11228 16396 11240
rect 16448 11228 16454 11280
rect 18598 11268 18604 11280
rect 18559 11240 18604 11268
rect 18598 11228 18604 11240
rect 18656 11228 18662 11280
rect 19797 11271 19855 11277
rect 19797 11237 19809 11271
rect 19843 11268 19855 11271
rect 20070 11268 20076 11280
rect 19843 11240 20076 11268
rect 19843 11237 19855 11240
rect 19797 11231 19855 11237
rect 20070 11228 20076 11240
rect 20128 11228 20134 11280
rect 2409 11203 2467 11209
rect 2409 11169 2421 11203
rect 2455 11169 2467 11203
rect 2866 11200 2872 11212
rect 2827 11172 2872 11200
rect 2409 11163 2467 11169
rect 2424 11064 2452 11163
rect 2866 11160 2872 11172
rect 2924 11160 2930 11212
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11200 5871 11203
rect 5994 11200 6000 11212
rect 5859 11172 6000 11200
rect 5859 11169 5871 11172
rect 5813 11163 5871 11169
rect 5994 11160 6000 11172
rect 6052 11160 6058 11212
rect 7834 11200 7840 11212
rect 7795 11172 7840 11200
rect 7834 11160 7840 11172
rect 7892 11160 7898 11212
rect 8018 11200 8024 11212
rect 7979 11172 8024 11200
rect 8018 11160 8024 11172
rect 8076 11160 8082 11212
rect 11333 11203 11391 11209
rect 11333 11169 11345 11203
rect 11379 11200 11391 11203
rect 11422 11200 11428 11212
rect 11379 11172 11428 11200
rect 11379 11169 11391 11172
rect 11333 11163 11391 11169
rect 11422 11160 11428 11172
rect 11480 11160 11486 11212
rect 15746 11200 15752 11212
rect 15659 11172 15752 11200
rect 15746 11160 15752 11172
rect 15804 11160 15810 11212
rect 16758 11160 16764 11212
rect 16816 11200 16822 11212
rect 17497 11203 17555 11209
rect 17497 11200 17509 11203
rect 16816 11172 17509 11200
rect 16816 11160 16822 11172
rect 17497 11169 17509 11172
rect 17543 11200 17555 11203
rect 17586 11200 17592 11212
rect 17543 11172 17592 11200
rect 17543 11169 17555 11172
rect 17497 11163 17555 11169
rect 17586 11160 17592 11172
rect 17644 11160 17650 11212
rect 17954 11200 17960 11212
rect 17915 11172 17960 11200
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 19058 11200 19064 11212
rect 19019 11172 19064 11200
rect 19058 11160 19064 11172
rect 19116 11160 19122 11212
rect 19334 11160 19340 11212
rect 19392 11200 19398 11212
rect 19521 11203 19579 11209
rect 19521 11200 19533 11203
rect 19392 11172 19533 11200
rect 19392 11160 19398 11172
rect 19521 11169 19533 11172
rect 19567 11169 19579 11203
rect 19521 11163 19579 11169
rect 20809 11203 20867 11209
rect 20809 11169 20821 11203
rect 20855 11200 20867 11203
rect 20898 11200 20904 11212
rect 20855 11172 20904 11200
rect 20855 11169 20867 11172
rect 20809 11163 20867 11169
rect 20898 11160 20904 11172
rect 20956 11160 20962 11212
rect 21910 11160 21916 11212
rect 21968 11200 21974 11212
rect 24210 11200 24216 11212
rect 21968 11172 24216 11200
rect 21968 11160 21974 11172
rect 24210 11160 24216 11172
rect 24268 11200 24274 11212
rect 24581 11203 24639 11209
rect 24581 11200 24593 11203
rect 24268 11172 24593 11200
rect 24268 11160 24274 11172
rect 24581 11169 24593 11172
rect 24627 11169 24639 11203
rect 24581 11163 24639 11169
rect 3142 11132 3148 11144
rect 3103 11104 3148 11132
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 4154 11092 4160 11144
rect 4212 11132 4218 11144
rect 4801 11135 4859 11141
rect 4212 11104 4257 11132
rect 4212 11092 4218 11104
rect 4801 11101 4813 11135
rect 4847 11132 4859 11135
rect 5258 11132 5264 11144
rect 4847 11104 5264 11132
rect 4847 11101 4859 11104
rect 4801 11095 4859 11101
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 5445 11135 5503 11141
rect 5445 11101 5457 11135
rect 5491 11132 5503 11135
rect 7006 11132 7012 11144
rect 5491 11104 7012 11132
rect 5491 11101 5503 11104
rect 5445 11095 5503 11101
rect 7006 11092 7012 11104
rect 7064 11092 7070 11144
rect 9398 11092 9404 11144
rect 9456 11132 9462 11144
rect 9769 11135 9827 11141
rect 9769 11132 9781 11135
rect 9456 11104 9781 11132
rect 9456 11092 9462 11104
rect 9769 11101 9781 11104
rect 9815 11101 9827 11135
rect 9769 11095 9827 11101
rect 13081 11135 13139 11141
rect 13081 11101 13093 11135
rect 13127 11132 13139 11135
rect 13538 11132 13544 11144
rect 13127 11104 13544 11132
rect 13127 11101 13139 11104
rect 13081 11095 13139 11101
rect 13538 11092 13544 11104
rect 13596 11092 13602 11144
rect 3326 11064 3332 11076
rect 2424 11036 3332 11064
rect 3326 11024 3332 11036
rect 3384 11064 3390 11076
rect 3384 11036 4154 11064
rect 3384 11024 3390 11036
rect 2038 10996 2044 11008
rect 1999 10968 2044 10996
rect 2038 10956 2044 10968
rect 2096 10956 2102 11008
rect 2406 10956 2412 11008
rect 2464 10996 2470 11008
rect 3421 10999 3479 11005
rect 3421 10996 3433 10999
rect 2464 10968 3433 10996
rect 2464 10956 2470 10968
rect 3421 10965 3433 10968
rect 3467 10965 3479 10999
rect 4126 10996 4154 11036
rect 5350 11024 5356 11076
rect 5408 11064 5414 11076
rect 6733 11067 6791 11073
rect 6733 11064 6745 11067
rect 5408 11036 6745 11064
rect 5408 11024 5414 11036
rect 6733 11033 6745 11036
rect 6779 11033 6791 11067
rect 6733 11027 6791 11033
rect 9490 11024 9496 11076
rect 9548 11064 9554 11076
rect 10321 11067 10379 11073
rect 10321 11064 10333 11067
rect 9548 11036 10333 11064
rect 9548 11024 9554 11036
rect 10321 11033 10333 11036
rect 10367 11064 10379 11067
rect 14090 11064 14096 11076
rect 10367 11036 14096 11064
rect 10367 11033 10379 11036
rect 10321 11027 10379 11033
rect 14090 11024 14096 11036
rect 14148 11024 14154 11076
rect 5445 10999 5503 11005
rect 5445 10996 5457 10999
rect 4126 10968 5457 10996
rect 3421 10959 3479 10965
rect 5445 10965 5457 10968
rect 5491 10965 5503 10999
rect 5445 10959 5503 10965
rect 5534 10956 5540 11008
rect 5592 10996 5598 11008
rect 5592 10968 5637 10996
rect 5592 10956 5598 10968
rect 8202 10956 8208 11008
rect 8260 10996 8266 11008
rect 8573 10999 8631 11005
rect 8573 10996 8585 10999
rect 8260 10968 8585 10996
rect 8260 10956 8266 10968
rect 8573 10965 8585 10968
rect 8619 10965 8631 10999
rect 10778 10996 10784 11008
rect 10739 10968 10784 10996
rect 8573 10959 8631 10965
rect 10778 10956 10784 10968
rect 10836 10956 10842 11008
rect 12250 10996 12256 11008
rect 12211 10968 12256 10996
rect 12250 10956 12256 10968
rect 12308 10956 12314 11008
rect 16666 10996 16672 11008
rect 16627 10968 16672 10996
rect 16666 10956 16672 10968
rect 16724 10956 16730 11008
rect 24765 10999 24823 11005
rect 24765 10965 24777 10999
rect 24811 10996 24823 10999
rect 27706 10996 27712 11008
rect 24811 10968 27712 10996
rect 24811 10965 24823 10968
rect 24765 10959 24823 10965
rect 27706 10956 27712 10968
rect 27764 10956 27770 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 4246 10792 4252 10804
rect 4207 10764 4252 10792
rect 4246 10752 4252 10764
rect 4304 10792 4310 10804
rect 4525 10795 4583 10801
rect 4525 10792 4537 10795
rect 4304 10764 4537 10792
rect 4304 10752 4310 10764
rect 4525 10761 4537 10764
rect 4571 10761 4583 10795
rect 4525 10755 4583 10761
rect 7834 10752 7840 10804
rect 7892 10792 7898 10804
rect 8389 10795 8447 10801
rect 8389 10792 8401 10795
rect 7892 10764 8401 10792
rect 7892 10752 7898 10764
rect 8389 10761 8401 10764
rect 8435 10792 8447 10795
rect 9214 10792 9220 10804
rect 8435 10764 9220 10792
rect 8435 10761 8447 10764
rect 8389 10755 8447 10761
rect 9214 10752 9220 10764
rect 9272 10752 9278 10804
rect 9401 10795 9459 10801
rect 9401 10761 9413 10795
rect 9447 10792 9459 10795
rect 9490 10792 9496 10804
rect 9447 10764 9496 10792
rect 9447 10761 9459 10764
rect 9401 10755 9459 10761
rect 3786 10684 3792 10736
rect 3844 10724 3850 10736
rect 8987 10727 9045 10733
rect 8987 10724 8999 10727
rect 3844 10696 8999 10724
rect 3844 10684 3850 10696
rect 8987 10693 8999 10696
rect 9033 10693 9045 10727
rect 8987 10687 9045 10693
rect 2498 10656 2504 10668
rect 2459 10628 2504 10656
rect 2498 10616 2504 10628
rect 2556 10616 2562 10668
rect 3142 10616 3148 10668
rect 3200 10656 3206 10668
rect 3329 10659 3387 10665
rect 3329 10656 3341 10659
rect 3200 10628 3341 10656
rect 3200 10616 3206 10628
rect 3329 10625 3341 10628
rect 3375 10625 3387 10659
rect 3329 10619 3387 10625
rect 5905 10659 5963 10665
rect 5905 10625 5917 10659
rect 5951 10656 5963 10659
rect 6362 10656 6368 10668
rect 5951 10628 6368 10656
rect 5951 10625 5963 10628
rect 5905 10619 5963 10625
rect 6362 10616 6368 10628
rect 6420 10616 6426 10668
rect 6822 10656 6828 10668
rect 6783 10628 6828 10656
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10588 1731 10591
rect 2038 10588 2044 10600
rect 1719 10560 2044 10588
rect 1719 10557 1731 10560
rect 1673 10551 1731 10557
rect 2038 10548 2044 10560
rect 2096 10548 2102 10600
rect 8916 10591 8974 10597
rect 8916 10557 8928 10591
rect 8962 10588 8974 10591
rect 9416 10588 9444 10755
rect 9490 10752 9496 10764
rect 9548 10752 9554 10804
rect 9858 10752 9864 10804
rect 9916 10792 9922 10804
rect 10045 10795 10103 10801
rect 10045 10792 10057 10795
rect 9916 10764 10057 10792
rect 9916 10752 9922 10764
rect 10045 10761 10057 10764
rect 10091 10761 10103 10795
rect 10045 10755 10103 10761
rect 11422 10752 11428 10804
rect 11480 10792 11486 10804
rect 12161 10795 12219 10801
rect 12161 10792 12173 10795
rect 11480 10764 12173 10792
rect 11480 10752 11486 10764
rect 12161 10761 12173 10764
rect 12207 10761 12219 10795
rect 12161 10755 12219 10761
rect 13357 10795 13415 10801
rect 13357 10761 13369 10795
rect 13403 10792 13415 10795
rect 13446 10792 13452 10804
rect 13403 10764 13452 10792
rect 13403 10761 13415 10764
rect 13357 10755 13415 10761
rect 11885 10727 11943 10733
rect 11885 10693 11897 10727
rect 11931 10724 11943 10727
rect 13372 10724 13400 10755
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 15378 10752 15384 10804
rect 15436 10792 15442 10804
rect 17083 10795 17141 10801
rect 17083 10792 17095 10795
rect 15436 10764 17095 10792
rect 15436 10752 15442 10764
rect 17083 10761 17095 10764
rect 17129 10761 17141 10795
rect 17770 10792 17776 10804
rect 17731 10764 17776 10792
rect 17083 10755 17141 10761
rect 17770 10752 17776 10764
rect 17828 10752 17834 10804
rect 19058 10792 19064 10804
rect 19019 10764 19064 10792
rect 19058 10752 19064 10764
rect 19116 10752 19122 10804
rect 19334 10752 19340 10804
rect 19392 10792 19398 10804
rect 19429 10795 19487 10801
rect 19429 10792 19441 10795
rect 19392 10764 19441 10792
rect 19392 10752 19398 10764
rect 19429 10761 19441 10764
rect 19475 10761 19487 10795
rect 19429 10755 19487 10761
rect 19518 10752 19524 10804
rect 19576 10792 19582 10804
rect 19751 10795 19809 10801
rect 19751 10792 19763 10795
rect 19576 10764 19763 10792
rect 19576 10752 19582 10764
rect 19751 10761 19763 10764
rect 19797 10761 19809 10795
rect 19751 10755 19809 10761
rect 20165 10795 20223 10801
rect 20165 10761 20177 10795
rect 20211 10792 20223 10795
rect 20254 10792 20260 10804
rect 20211 10764 20260 10792
rect 20211 10761 20223 10764
rect 20165 10755 20223 10761
rect 14090 10724 14096 10736
rect 11931 10696 13400 10724
rect 14051 10696 14096 10724
rect 11931 10693 11943 10696
rect 11885 10687 11943 10693
rect 14090 10684 14096 10696
rect 14148 10684 14154 10736
rect 14734 10684 14740 10736
rect 14792 10724 14798 10736
rect 16761 10727 16819 10733
rect 16761 10724 16773 10727
rect 14792 10696 16773 10724
rect 14792 10684 14798 10696
rect 16761 10693 16773 10696
rect 16807 10724 16819 10727
rect 17954 10724 17960 10736
rect 16807 10696 17960 10724
rect 16807 10693 16819 10696
rect 16761 10687 16819 10693
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 13541 10659 13599 10665
rect 13541 10625 13553 10659
rect 13587 10656 13599 10659
rect 13906 10656 13912 10668
rect 13587 10628 13912 10656
rect 13587 10625 13599 10628
rect 13541 10619 13599 10625
rect 13906 10616 13912 10628
rect 13964 10656 13970 10668
rect 15749 10659 15807 10665
rect 15749 10656 15761 10659
rect 13964 10628 15761 10656
rect 13964 10616 13970 10628
rect 15749 10625 15761 10628
rect 15795 10625 15807 10659
rect 16390 10656 16396 10668
rect 16351 10628 16396 10656
rect 15749 10619 15807 10625
rect 16390 10616 16396 10628
rect 16448 10616 16454 10668
rect 10686 10588 10692 10600
rect 8962 10560 9444 10588
rect 10599 10560 10692 10588
rect 8962 10557 8974 10560
rect 8916 10551 8974 10557
rect 10686 10548 10692 10560
rect 10744 10588 10750 10600
rect 11054 10588 11060 10600
rect 10744 10560 11060 10588
rect 10744 10548 10750 10560
rect 11054 10548 11060 10560
rect 11112 10548 11118 10600
rect 11241 10591 11299 10597
rect 11241 10557 11253 10591
rect 11287 10557 11299 10591
rect 11241 10551 11299 10557
rect 12504 10591 12562 10597
rect 12504 10557 12516 10591
rect 12550 10588 12562 10591
rect 12986 10588 12992 10600
rect 12550 10560 12992 10588
rect 12550 10557 12562 10560
rect 12504 10551 12562 10557
rect 3237 10523 3295 10529
rect 3237 10489 3249 10523
rect 3283 10520 3295 10523
rect 3650 10523 3708 10529
rect 3650 10520 3662 10523
rect 3283 10492 3662 10520
rect 3283 10489 3295 10492
rect 3237 10483 3295 10489
rect 3650 10489 3662 10492
rect 3696 10520 3708 10523
rect 4246 10520 4252 10532
rect 3696 10492 4252 10520
rect 3696 10489 3708 10492
rect 3650 10483 3708 10489
rect 4246 10480 4252 10492
rect 4304 10480 4310 10532
rect 5258 10520 5264 10532
rect 5219 10492 5264 10520
rect 5258 10480 5264 10492
rect 5316 10480 5322 10532
rect 5350 10480 5356 10532
rect 5408 10520 5414 10532
rect 7146 10523 7204 10529
rect 7146 10520 7158 10523
rect 5408 10492 5453 10520
rect 6564 10492 7158 10520
rect 5408 10480 5414 10492
rect 2866 10452 2872 10464
rect 2827 10424 2872 10452
rect 2866 10412 2872 10424
rect 2924 10412 2930 10464
rect 5077 10455 5135 10461
rect 5077 10421 5089 10455
rect 5123 10452 5135 10455
rect 5368 10452 5396 10480
rect 5123 10424 5396 10452
rect 5123 10421 5135 10424
rect 5077 10415 5135 10421
rect 5442 10412 5448 10464
rect 5500 10452 5506 10464
rect 6086 10452 6092 10464
rect 5500 10424 6092 10452
rect 5500 10412 5506 10424
rect 6086 10412 6092 10424
rect 6144 10452 6150 10464
rect 6564 10461 6592 10492
rect 7146 10489 7158 10492
rect 7192 10489 7204 10523
rect 7146 10483 7204 10489
rect 7558 10480 7564 10532
rect 7616 10520 7622 10532
rect 8018 10520 8024 10532
rect 7616 10492 8024 10520
rect 7616 10480 7622 10492
rect 8018 10480 8024 10492
rect 8076 10480 8082 10532
rect 10778 10480 10784 10532
rect 10836 10520 10842 10532
rect 11256 10520 11284 10551
rect 12986 10548 12992 10560
rect 13044 10548 13050 10600
rect 17012 10591 17070 10597
rect 17012 10557 17024 10591
rect 17058 10588 17070 10591
rect 17058 10560 17540 10588
rect 17058 10557 17070 10560
rect 17012 10551 17070 10557
rect 10836 10492 11284 10520
rect 11517 10523 11575 10529
rect 10836 10480 10842 10492
rect 11517 10489 11529 10523
rect 11563 10520 11575 10523
rect 13630 10520 13636 10532
rect 11563 10492 13486 10520
rect 13591 10492 13636 10520
rect 11563 10489 11575 10492
rect 11517 10483 11575 10489
rect 6181 10455 6239 10461
rect 6181 10452 6193 10455
rect 6144 10424 6193 10452
rect 6144 10412 6150 10424
rect 6181 10421 6193 10424
rect 6227 10452 6239 10455
rect 6549 10455 6607 10461
rect 6549 10452 6561 10455
rect 6227 10424 6561 10452
rect 6227 10421 6239 10424
rect 6181 10415 6239 10421
rect 6549 10421 6561 10424
rect 6595 10421 6607 10455
rect 7742 10452 7748 10464
rect 7703 10424 7748 10452
rect 6549 10415 6607 10421
rect 7742 10412 7748 10424
rect 7800 10412 7806 10464
rect 9398 10412 9404 10464
rect 9456 10452 9462 10464
rect 9677 10455 9735 10461
rect 9677 10452 9689 10455
rect 9456 10424 9689 10452
rect 9456 10412 9462 10424
rect 9677 10421 9689 10424
rect 9723 10421 9735 10455
rect 9677 10415 9735 10421
rect 12575 10455 12633 10461
rect 12575 10421 12587 10455
rect 12621 10452 12633 10455
rect 12802 10452 12808 10464
rect 12621 10424 12808 10452
rect 12621 10421 12633 10424
rect 12575 10415 12633 10421
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 12986 10452 12992 10464
rect 12947 10424 12992 10452
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 13458 10452 13486 10492
rect 13630 10480 13636 10492
rect 13688 10520 13694 10532
rect 14921 10523 14979 10529
rect 13688 10492 13814 10520
rect 13688 10480 13694 10492
rect 13538 10452 13544 10464
rect 13458 10424 13544 10452
rect 13538 10412 13544 10424
rect 13596 10412 13602 10464
rect 13786 10452 13814 10492
rect 14921 10489 14933 10523
rect 14967 10520 14979 10523
rect 15470 10520 15476 10532
rect 14967 10492 15476 10520
rect 14967 10489 14979 10492
rect 14921 10483 14979 10489
rect 15470 10480 15476 10492
rect 15528 10480 15534 10532
rect 15562 10480 15568 10532
rect 15620 10520 15626 10532
rect 17512 10529 17540 10560
rect 17770 10548 17776 10600
rect 17828 10588 17834 10600
rect 18049 10591 18107 10597
rect 18049 10588 18061 10591
rect 17828 10560 18061 10588
rect 17828 10548 17834 10560
rect 18049 10557 18061 10560
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 18138 10548 18144 10600
rect 18196 10588 18202 10600
rect 18601 10591 18659 10597
rect 18601 10588 18613 10591
rect 18196 10560 18613 10588
rect 18196 10548 18202 10560
rect 18601 10557 18613 10560
rect 18647 10588 18659 10591
rect 19334 10588 19340 10600
rect 18647 10560 19340 10588
rect 18647 10557 18659 10560
rect 18601 10551 18659 10557
rect 19334 10548 19340 10560
rect 19392 10548 19398 10600
rect 19426 10548 19432 10600
rect 19484 10588 19490 10600
rect 19680 10591 19738 10597
rect 19680 10588 19692 10591
rect 19484 10560 19692 10588
rect 19484 10548 19490 10560
rect 19680 10557 19692 10560
rect 19726 10588 19738 10591
rect 20180 10588 20208 10755
rect 20254 10752 20260 10764
rect 20312 10752 20318 10804
rect 24210 10752 24216 10804
rect 24268 10792 24274 10804
rect 24397 10795 24455 10801
rect 24397 10792 24409 10795
rect 24268 10764 24409 10792
rect 24268 10752 24274 10764
rect 24397 10761 24409 10764
rect 24443 10761 24455 10795
rect 24397 10755 24455 10761
rect 24762 10724 24768 10736
rect 24723 10696 24768 10724
rect 24762 10684 24768 10696
rect 24820 10684 24826 10736
rect 19726 10560 20208 10588
rect 19726 10557 19738 10560
rect 19680 10551 19738 10557
rect 24026 10548 24032 10600
rect 24084 10588 24090 10600
rect 24581 10591 24639 10597
rect 24581 10588 24593 10591
rect 24084 10560 24593 10588
rect 24084 10548 24090 10560
rect 24581 10557 24593 10560
rect 24627 10588 24639 10591
rect 25133 10591 25191 10597
rect 25133 10588 25145 10591
rect 24627 10560 25145 10588
rect 24627 10557 24639 10560
rect 24581 10551 24639 10557
rect 25133 10557 25145 10560
rect 25179 10557 25191 10591
rect 25133 10551 25191 10557
rect 17497 10523 17555 10529
rect 15620 10492 15665 10520
rect 15620 10480 15626 10492
rect 17497 10489 17509 10523
rect 17543 10520 17555 10523
rect 17954 10520 17960 10532
rect 17543 10492 17960 10520
rect 17543 10489 17555 10492
rect 17497 10483 17555 10489
rect 17954 10480 17960 10492
rect 18012 10520 18018 10532
rect 20806 10520 20812 10532
rect 18012 10492 20812 10520
rect 18012 10480 18018 10492
rect 20806 10480 20812 10492
rect 20864 10480 20870 10532
rect 14461 10455 14519 10461
rect 14461 10452 14473 10455
rect 13786 10424 14473 10452
rect 14461 10421 14473 10424
rect 14507 10421 14519 10455
rect 14461 10415 14519 10421
rect 15289 10455 15347 10461
rect 15289 10421 15301 10455
rect 15335 10452 15347 10455
rect 15580 10452 15608 10480
rect 18322 10452 18328 10464
rect 15335 10424 15608 10452
rect 18283 10424 18328 10452
rect 15335 10421 15347 10424
rect 15289 10415 15347 10421
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 20898 10452 20904 10464
rect 20859 10424 20904 10452
rect 20898 10412 20904 10424
rect 20956 10412 20962 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1394 10208 1400 10260
rect 1452 10248 1458 10260
rect 2225 10251 2283 10257
rect 2225 10248 2237 10251
rect 1452 10220 2237 10248
rect 1452 10208 1458 10220
rect 2225 10217 2237 10220
rect 2271 10217 2283 10251
rect 2225 10211 2283 10217
rect 3142 10208 3148 10260
rect 3200 10248 3206 10260
rect 3789 10251 3847 10257
rect 3789 10248 3801 10251
rect 3200 10220 3801 10248
rect 3200 10208 3206 10220
rect 3789 10217 3801 10220
rect 3835 10217 3847 10251
rect 4154 10248 4160 10260
rect 3789 10211 3847 10217
rect 4126 10208 4160 10248
rect 4212 10248 4218 10260
rect 4249 10251 4307 10257
rect 4249 10248 4261 10251
rect 4212 10220 4261 10248
rect 4212 10208 4218 10220
rect 4249 10217 4261 10220
rect 4295 10217 4307 10251
rect 4249 10211 4307 10217
rect 5994 10208 6000 10260
rect 6052 10248 6058 10260
rect 6089 10251 6147 10257
rect 6089 10248 6101 10251
rect 6052 10220 6101 10248
rect 6052 10208 6058 10220
rect 6089 10217 6101 10220
rect 6135 10217 6147 10251
rect 6089 10211 6147 10217
rect 8757 10251 8815 10257
rect 8757 10217 8769 10251
rect 8803 10248 8815 10251
rect 9306 10248 9312 10260
rect 8803 10220 9312 10248
rect 8803 10217 8815 10220
rect 8757 10211 8815 10217
rect 9306 10208 9312 10220
rect 9364 10208 9370 10260
rect 10505 10251 10563 10257
rect 10505 10217 10517 10251
rect 10551 10248 10563 10251
rect 10686 10248 10692 10260
rect 10551 10220 10692 10248
rect 10551 10217 10563 10220
rect 10505 10211 10563 10217
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 13906 10248 13912 10260
rect 13458 10220 13912 10248
rect 1673 10183 1731 10189
rect 1673 10149 1685 10183
rect 1719 10180 1731 10183
rect 4126 10180 4154 10208
rect 1719 10152 4154 10180
rect 5255 10183 5313 10189
rect 1719 10149 1731 10152
rect 1673 10143 1731 10149
rect 5255 10149 5267 10183
rect 5301 10180 5313 10183
rect 5350 10180 5356 10192
rect 5301 10152 5356 10180
rect 5301 10149 5313 10152
rect 5255 10143 5313 10149
rect 5350 10140 5356 10152
rect 5408 10140 5414 10192
rect 6270 10140 6276 10192
rect 6328 10180 6334 10192
rect 6825 10183 6883 10189
rect 6825 10180 6837 10183
rect 6328 10152 6837 10180
rect 6328 10140 6334 10152
rect 6825 10149 6837 10152
rect 6871 10180 6883 10183
rect 7742 10180 7748 10192
rect 6871 10152 7748 10180
rect 6871 10149 6883 10152
rect 6825 10143 6883 10149
rect 7742 10140 7748 10152
rect 7800 10140 7806 10192
rect 12250 10140 12256 10192
rect 12308 10180 12314 10192
rect 12710 10180 12716 10192
rect 12308 10152 12716 10180
rect 12308 10140 12314 10152
rect 12710 10140 12716 10152
rect 12768 10180 12774 10192
rect 12805 10183 12863 10189
rect 12805 10180 12817 10183
rect 12768 10152 12817 10180
rect 12768 10140 12774 10152
rect 12805 10149 12817 10152
rect 12851 10149 12863 10183
rect 12805 10143 12863 10149
rect 13357 10183 13415 10189
rect 13357 10149 13369 10183
rect 13403 10180 13415 10183
rect 13458 10180 13486 10220
rect 13906 10208 13912 10220
rect 13964 10248 13970 10260
rect 14001 10251 14059 10257
rect 14001 10248 14013 10251
rect 13964 10220 14013 10248
rect 13964 10208 13970 10220
rect 14001 10217 14013 10220
rect 14047 10217 14059 10251
rect 14001 10211 14059 10217
rect 14323 10251 14381 10257
rect 14323 10217 14335 10251
rect 14369 10248 14381 10251
rect 14826 10248 14832 10260
rect 14369 10220 14832 10248
rect 14369 10217 14381 10220
rect 14323 10211 14381 10217
rect 14826 10208 14832 10220
rect 14884 10208 14890 10260
rect 15470 10208 15476 10260
rect 15528 10248 15534 10260
rect 15565 10251 15623 10257
rect 15565 10248 15577 10251
rect 15528 10220 15577 10248
rect 15528 10208 15534 10220
rect 15565 10217 15577 10220
rect 15611 10217 15623 10251
rect 15746 10248 15752 10260
rect 15707 10220 15752 10248
rect 15565 10211 15623 10217
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 17586 10248 17592 10260
rect 17547 10220 17592 10248
rect 17586 10208 17592 10220
rect 17644 10208 17650 10260
rect 18138 10248 18144 10260
rect 18099 10220 18144 10248
rect 18138 10208 18144 10220
rect 18196 10208 18202 10260
rect 13403 10152 13486 10180
rect 13403 10149 13415 10152
rect 13357 10143 13415 10149
rect 13538 10140 13544 10192
rect 13596 10180 13602 10192
rect 13633 10183 13691 10189
rect 13633 10180 13645 10183
rect 13596 10152 13645 10180
rect 13596 10140 13602 10152
rect 13633 10149 13645 10152
rect 13679 10149 13691 10183
rect 13633 10143 13691 10149
rect 13722 10140 13728 10192
rect 13780 10180 13786 10192
rect 13814 10180 13820 10192
rect 13780 10152 13820 10180
rect 13780 10140 13786 10152
rect 13814 10140 13820 10152
rect 13872 10140 13878 10192
rect 16666 10140 16672 10192
rect 16724 10180 16730 10192
rect 16761 10183 16819 10189
rect 16761 10180 16773 10183
rect 16724 10152 16773 10180
rect 16724 10140 16730 10152
rect 16761 10149 16773 10152
rect 16807 10149 16819 10183
rect 16761 10143 16819 10149
rect 1464 10115 1522 10121
rect 1464 10081 1476 10115
rect 1510 10112 1522 10115
rect 1854 10112 1860 10124
rect 1510 10084 1860 10112
rect 1510 10081 1522 10084
rect 1464 10075 1522 10081
rect 1854 10072 1860 10084
rect 1912 10072 1918 10124
rect 2406 10112 2412 10124
rect 2367 10084 2412 10112
rect 2406 10072 2412 10084
rect 2464 10072 2470 10124
rect 2498 10072 2504 10124
rect 2556 10112 2562 10124
rect 2682 10112 2688 10124
rect 2556 10084 2601 10112
rect 2643 10084 2688 10112
rect 2556 10072 2562 10084
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 3326 10072 3332 10124
rect 3384 10112 3390 10124
rect 3421 10115 3479 10121
rect 3421 10112 3433 10115
rect 3384 10084 3433 10112
rect 3384 10072 3390 10084
rect 3421 10081 3433 10084
rect 3467 10081 3479 10115
rect 3421 10075 3479 10081
rect 8202 10072 8208 10124
rect 8260 10112 8266 10124
rect 8573 10115 8631 10121
rect 8573 10112 8585 10115
rect 8260 10084 8585 10112
rect 8260 10072 8266 10084
rect 8573 10081 8585 10084
rect 8619 10112 8631 10115
rect 8846 10112 8852 10124
rect 8619 10084 8852 10112
rect 8619 10081 8631 10084
rect 8573 10075 8631 10081
rect 8846 10072 8852 10084
rect 8904 10072 8910 10124
rect 9582 10072 9588 10124
rect 9640 10112 9646 10124
rect 10318 10112 10324 10124
rect 9640 10084 10324 10112
rect 9640 10072 9646 10084
rect 10318 10072 10324 10084
rect 10376 10072 10382 10124
rect 14182 10112 14188 10124
rect 14143 10084 14188 10112
rect 14182 10072 14188 10084
rect 14240 10072 14246 10124
rect 15197 10115 15255 10121
rect 15197 10081 15209 10115
rect 15243 10112 15255 10115
rect 15378 10112 15384 10124
rect 15243 10084 15384 10112
rect 15243 10081 15255 10084
rect 15197 10075 15255 10081
rect 15378 10072 15384 10084
rect 15436 10072 15442 10124
rect 3142 10044 3148 10056
rect 3103 10016 3148 10044
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10044 4951 10047
rect 5074 10044 5080 10056
rect 4939 10016 5080 10044
rect 4939 10013 4951 10016
rect 4893 10007 4951 10013
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 6733 10047 6791 10053
rect 6733 10013 6745 10047
rect 6779 10044 6791 10047
rect 7834 10044 7840 10056
rect 6779 10016 7840 10044
rect 6779 10013 6791 10016
rect 6733 10007 6791 10013
rect 7834 10004 7840 10016
rect 7892 10004 7898 10056
rect 12158 10004 12164 10056
rect 12216 10044 12222 10056
rect 12713 10047 12771 10053
rect 12713 10044 12725 10047
rect 12216 10016 12725 10044
rect 12216 10004 12222 10016
rect 12713 10013 12725 10016
rect 12759 10013 12771 10047
rect 12713 10007 12771 10013
rect 16669 10047 16727 10053
rect 16669 10013 16681 10047
rect 16715 10044 16727 10047
rect 16758 10044 16764 10056
rect 16715 10016 16764 10044
rect 16715 10013 16727 10016
rect 16669 10007 16727 10013
rect 16758 10004 16764 10016
rect 16816 10004 16822 10056
rect 16942 10044 16948 10056
rect 16903 10016 16948 10044
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 6362 9936 6368 9988
rect 6420 9976 6426 9988
rect 7285 9979 7343 9985
rect 7285 9976 7297 9979
rect 6420 9948 7297 9976
rect 6420 9936 6426 9948
rect 7285 9945 7297 9948
rect 7331 9945 7343 9979
rect 7285 9939 7343 9945
rect 7466 9936 7472 9988
rect 7524 9976 7530 9988
rect 10778 9976 10784 9988
rect 7524 9948 10784 9976
rect 7524 9936 7530 9948
rect 10778 9936 10784 9948
rect 10836 9936 10842 9988
rect 1854 9868 1860 9920
rect 1912 9908 1918 9920
rect 3602 9908 3608 9920
rect 1912 9880 3608 9908
rect 1912 9868 1918 9880
rect 3602 9868 3608 9880
rect 3660 9868 3666 9920
rect 4801 9911 4859 9917
rect 4801 9877 4813 9911
rect 4847 9908 4859 9911
rect 5258 9908 5264 9920
rect 4847 9880 5264 9908
rect 4847 9877 4859 9880
rect 4801 9871 4859 9877
rect 5258 9868 5264 9880
rect 5316 9868 5322 9920
rect 5813 9911 5871 9917
rect 5813 9877 5825 9911
rect 5859 9908 5871 9911
rect 6546 9908 6552 9920
rect 5859 9880 6552 9908
rect 5859 9877 5871 9880
rect 5813 9871 5871 9877
rect 6546 9868 6552 9880
rect 6604 9868 6610 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 1578 9704 1584 9716
rect 1539 9676 1584 9704
rect 1578 9664 1584 9676
rect 1636 9664 1642 9716
rect 2498 9664 2504 9716
rect 2556 9704 2562 9716
rect 2777 9707 2835 9713
rect 2777 9704 2789 9707
rect 2556 9676 2789 9704
rect 2556 9664 2562 9676
rect 2777 9673 2789 9676
rect 2823 9673 2835 9707
rect 6270 9704 6276 9716
rect 6231 9676 6276 9704
rect 2777 9667 2835 9673
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 6546 9704 6552 9716
rect 6507 9676 6552 9704
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 8846 9704 8852 9716
rect 8807 9676 8852 9704
rect 8846 9664 8852 9676
rect 8904 9664 8910 9716
rect 10318 9704 10324 9716
rect 10279 9676 10324 9704
rect 10318 9664 10324 9676
rect 10376 9664 10382 9716
rect 12710 9704 12716 9716
rect 12671 9676 12716 9704
rect 12710 9664 12716 9676
rect 12768 9704 12774 9716
rect 13081 9707 13139 9713
rect 13081 9704 13093 9707
rect 12768 9676 13093 9704
rect 12768 9664 12774 9676
rect 13081 9673 13093 9676
rect 13127 9704 13139 9707
rect 13446 9704 13452 9716
rect 13127 9676 13452 9704
rect 13127 9673 13139 9676
rect 13081 9667 13139 9673
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 13538 9664 13544 9716
rect 13596 9704 13602 9716
rect 14182 9704 14188 9716
rect 13596 9676 14188 9704
rect 13596 9664 13602 9676
rect 14182 9664 14188 9676
rect 14240 9704 14246 9716
rect 14277 9707 14335 9713
rect 14277 9704 14289 9707
rect 14240 9676 14289 9704
rect 14240 9664 14246 9676
rect 14277 9673 14289 9676
rect 14323 9673 14335 9707
rect 14277 9667 14335 9673
rect 15930 9664 15936 9716
rect 15988 9704 15994 9716
rect 16071 9707 16129 9713
rect 16071 9704 16083 9707
rect 15988 9676 16083 9704
rect 15988 9664 15994 9676
rect 16071 9673 16083 9676
rect 16117 9673 16129 9707
rect 16071 9667 16129 9673
rect 16666 9664 16672 9716
rect 16724 9704 16730 9716
rect 16761 9707 16819 9713
rect 16761 9704 16773 9707
rect 16724 9676 16773 9704
rect 16724 9664 16730 9676
rect 16761 9673 16773 9676
rect 16807 9673 16819 9707
rect 16761 9667 16819 9673
rect 5074 9596 5080 9648
rect 5132 9636 5138 9648
rect 5905 9639 5963 9645
rect 5905 9636 5917 9639
rect 5132 9608 5917 9636
rect 5132 9596 5138 9608
rect 5905 9605 5917 9608
rect 5951 9636 5963 9639
rect 6730 9636 6736 9648
rect 5951 9608 6736 9636
rect 5951 9605 5963 9608
rect 5905 9599 5963 9605
rect 6730 9596 6736 9608
rect 6788 9596 6794 9648
rect 16485 9639 16543 9645
rect 16485 9605 16497 9639
rect 16531 9636 16543 9639
rect 19426 9636 19432 9648
rect 16531 9608 19432 9636
rect 16531 9605 16543 9608
rect 16485 9599 16543 9605
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2682 9568 2688 9580
rect 2547 9540 2688 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 3050 9528 3056 9580
rect 3108 9568 3114 9580
rect 3510 9568 3516 9580
rect 3108 9540 3516 9568
rect 3108 9528 3114 9540
rect 3510 9528 3516 9540
rect 3568 9528 3574 9580
rect 3878 9528 3884 9580
rect 3936 9568 3942 9580
rect 4249 9571 4307 9577
rect 4249 9568 4261 9571
rect 3936 9540 4261 9568
rect 3936 9528 3942 9540
rect 4249 9537 4261 9540
rect 4295 9537 4307 9571
rect 4249 9531 4307 9537
rect 6917 9571 6975 9577
rect 6917 9537 6929 9571
rect 6963 9568 6975 9571
rect 7006 9568 7012 9580
rect 6963 9540 7012 9568
rect 6963 9537 6975 9540
rect 6917 9531 6975 9537
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 7190 9568 7196 9580
rect 7151 9540 7196 9568
rect 7190 9528 7196 9540
rect 7248 9528 7254 9580
rect 8389 9571 8447 9577
rect 8389 9537 8401 9571
rect 8435 9568 8447 9571
rect 8478 9568 8484 9580
rect 8435 9540 8484 9568
rect 8435 9537 8447 9540
rect 8389 9531 8447 9537
rect 8478 9528 8484 9540
rect 8536 9528 8542 9580
rect 9398 9568 9404 9580
rect 9359 9540 9404 9568
rect 9398 9528 9404 9540
rect 9456 9528 9462 9580
rect 12802 9528 12808 9580
rect 12860 9568 12866 9580
rect 13354 9568 13360 9580
rect 12860 9540 13360 9568
rect 12860 9528 12866 9540
rect 13354 9528 13360 9540
rect 13412 9528 13418 9580
rect 13814 9528 13820 9580
rect 13872 9568 13878 9580
rect 13872 9540 13917 9568
rect 13872 9528 13878 9540
rect 1302 9460 1308 9512
rect 1360 9500 1366 9512
rect 1397 9503 1455 9509
rect 1397 9500 1409 9503
rect 1360 9472 1409 9500
rect 1360 9460 1366 9472
rect 1397 9469 1409 9472
rect 1443 9500 1455 9503
rect 1857 9503 1915 9509
rect 1857 9500 1869 9503
rect 1443 9472 1869 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1857 9469 1869 9472
rect 1903 9469 1915 9503
rect 1857 9463 1915 9469
rect 3304 9503 3362 9509
rect 3304 9469 3316 9503
rect 3350 9500 3362 9503
rect 3694 9500 3700 9512
rect 3350 9472 3700 9500
rect 3350 9469 3362 9472
rect 3304 9463 3362 9469
rect 106 9392 112 9444
rect 164 9432 170 9444
rect 3319 9432 3347 9463
rect 3694 9460 3700 9472
rect 3752 9460 3758 9512
rect 16000 9503 16058 9509
rect 16000 9469 16012 9503
rect 16046 9500 16058 9503
rect 16500 9500 16528 9599
rect 19426 9596 19432 9608
rect 19484 9596 19490 9648
rect 16046 9472 16528 9500
rect 24648 9503 24706 9509
rect 16046 9469 16058 9472
rect 16000 9463 16058 9469
rect 24648 9469 24660 9503
rect 24694 9500 24706 9503
rect 24694 9472 25176 9500
rect 24694 9469 24706 9472
rect 24648 9463 24706 9469
rect 164 9404 3347 9432
rect 164 9392 170 9404
rect 3510 9392 3516 9444
rect 3568 9432 3574 9444
rect 4157 9435 4215 9441
rect 4157 9432 4169 9435
rect 3568 9404 4169 9432
rect 3568 9392 3574 9404
rect 4157 9401 4169 9404
rect 4203 9432 4215 9435
rect 4246 9432 4252 9444
rect 4203 9404 4252 9432
rect 4203 9401 4215 9404
rect 4157 9395 4215 9401
rect 4246 9392 4252 9404
rect 4304 9432 4310 9444
rect 4570 9435 4628 9441
rect 4570 9432 4582 9435
rect 4304 9404 4582 9432
rect 4304 9392 4310 9404
rect 4570 9401 4582 9404
rect 4616 9432 4628 9435
rect 5350 9432 5356 9444
rect 4616 9404 5356 9432
rect 4616 9401 4628 9404
rect 4570 9395 4628 9401
rect 5350 9392 5356 9404
rect 5408 9432 5414 9444
rect 5445 9435 5503 9441
rect 5445 9432 5457 9435
rect 5408 9404 5457 9432
rect 5408 9392 5414 9404
rect 5445 9401 5457 9404
rect 5491 9401 5503 9435
rect 5445 9395 5503 9401
rect 7009 9435 7067 9441
rect 7009 9401 7021 9435
rect 7055 9401 7067 9435
rect 13446 9432 13452 9444
rect 13407 9404 13452 9432
rect 7009 9395 7067 9401
rect 3375 9367 3433 9373
rect 3375 9333 3387 9367
rect 3421 9364 3433 9367
rect 3602 9364 3608 9376
rect 3421 9336 3608 9364
rect 3421 9333 3433 9336
rect 3375 9327 3433 9333
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 5166 9364 5172 9376
rect 5127 9336 5172 9364
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 6546 9324 6552 9376
rect 6604 9364 6610 9376
rect 7024 9364 7052 9395
rect 13446 9392 13452 9404
rect 13504 9392 13510 9444
rect 15378 9432 15384 9444
rect 15291 9404 15384 9432
rect 15378 9392 15384 9404
rect 15436 9432 15442 9444
rect 21450 9432 21456 9444
rect 15436 9404 21456 9432
rect 15436 9392 15442 9404
rect 21450 9392 21456 9404
rect 21508 9392 21514 9444
rect 25148 9376 25176 9472
rect 7834 9364 7840 9376
rect 6604 9336 7052 9364
rect 7795 9336 7840 9364
rect 6604 9324 6610 9336
rect 7834 9324 7840 9336
rect 7892 9324 7898 9376
rect 12158 9364 12164 9376
rect 12119 9336 12164 9364
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 16758 9324 16764 9376
rect 16816 9364 16822 9376
rect 17221 9367 17279 9373
rect 17221 9364 17233 9367
rect 16816 9336 17233 9364
rect 16816 9324 16822 9336
rect 17221 9333 17233 9336
rect 17267 9364 17279 9367
rect 24719 9367 24777 9373
rect 24719 9364 24731 9367
rect 17267 9336 24731 9364
rect 17267 9333 17279 9336
rect 17221 9327 17279 9333
rect 24719 9333 24731 9336
rect 24765 9333 24777 9367
rect 25130 9364 25136 9376
rect 25091 9336 25136 9364
rect 24719 9327 24777 9333
rect 25130 9324 25136 9336
rect 25188 9324 25194 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1578 9160 1584 9172
rect 1539 9132 1584 9160
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 2406 9160 2412 9172
rect 2367 9132 2412 9160
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 3878 9120 3884 9172
rect 3936 9160 3942 9172
rect 4249 9163 4307 9169
rect 4249 9160 4261 9163
rect 3936 9132 4261 9160
rect 3936 9120 3942 9132
rect 4249 9129 4261 9132
rect 4295 9129 4307 9163
rect 4249 9123 4307 9129
rect 6549 9163 6607 9169
rect 6549 9129 6561 9163
rect 6595 9160 6607 9163
rect 6638 9160 6644 9172
rect 6595 9132 6644 9160
rect 6595 9129 6607 9132
rect 6549 9123 6607 9129
rect 6638 9120 6644 9132
rect 6696 9120 6702 9172
rect 7650 9120 7656 9172
rect 7708 9160 7714 9172
rect 7745 9163 7803 9169
rect 7745 9160 7757 9163
rect 7708 9132 7757 9160
rect 7708 9120 7714 9132
rect 7745 9129 7757 9132
rect 7791 9129 7803 9163
rect 13354 9160 13360 9172
rect 13315 9132 13360 9160
rect 7745 9123 7803 9129
rect 13354 9120 13360 9132
rect 13412 9120 13418 9172
rect 24762 9160 24768 9172
rect 24723 9132 24768 9160
rect 24762 9120 24768 9132
rect 24820 9120 24826 9172
rect 1946 9052 1952 9104
rect 2004 9092 2010 9104
rect 5166 9092 5172 9104
rect 2004 9064 3004 9092
rect 5127 9064 5172 9092
rect 2004 9052 2010 9064
rect 2976 9036 3004 9064
rect 5166 9052 5172 9064
rect 5224 9052 5230 9104
rect 5258 9052 5264 9104
rect 5316 9092 5322 9104
rect 5721 9095 5779 9101
rect 5721 9092 5733 9095
rect 5316 9064 5733 9092
rect 5316 9052 5322 9064
rect 5721 9061 5733 9064
rect 5767 9092 5779 9095
rect 7190 9092 7196 9104
rect 5767 9064 7196 9092
rect 5767 9061 5779 9064
rect 5721 9055 5779 9061
rect 7190 9052 7196 9064
rect 7248 9052 7254 9104
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2314 9024 2320 9036
rect 1443 8996 2320 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2314 8984 2320 8996
rect 2372 8984 2378 9036
rect 2958 9024 2964 9036
rect 2871 8996 2964 9024
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 7561 9027 7619 9033
rect 7561 8993 7573 9027
rect 7607 8993 7619 9027
rect 7561 8987 7619 8993
rect 3602 8916 3608 8968
rect 3660 8956 3666 8968
rect 5077 8959 5135 8965
rect 5077 8956 5089 8959
rect 3660 8928 5089 8956
rect 3660 8916 3666 8928
rect 5077 8925 5089 8928
rect 5123 8956 5135 8959
rect 5994 8956 6000 8968
rect 5123 8928 6000 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5994 8916 6000 8928
rect 6052 8916 6058 8968
rect 7576 8900 7604 8987
rect 21726 8984 21732 9036
rect 21784 9024 21790 9036
rect 24581 9027 24639 9033
rect 24581 9024 24593 9027
rect 21784 8996 24593 9024
rect 21784 8984 21790 8996
rect 24581 8993 24593 8996
rect 24627 9024 24639 9027
rect 24670 9024 24676 9036
rect 24627 8996 24676 9024
rect 24627 8993 24639 8996
rect 24581 8987 24639 8993
rect 24670 8984 24676 8996
rect 24728 8984 24734 9036
rect 3145 8891 3203 8897
rect 3145 8857 3157 8891
rect 3191 8888 3203 8891
rect 7558 8888 7564 8900
rect 3191 8860 7564 8888
rect 3191 8857 3203 8860
rect 3145 8851 3203 8857
rect 7558 8848 7564 8860
rect 7616 8848 7622 8900
rect 7006 8820 7012 8832
rect 6967 8792 7012 8820
rect 7006 8780 7012 8792
rect 7064 8780 7070 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1535 8619 1593 8625
rect 1535 8585 1547 8619
rect 1581 8616 1593 8619
rect 1670 8616 1676 8628
rect 1581 8588 1676 8616
rect 1581 8585 1593 8588
rect 1535 8579 1593 8585
rect 1670 8576 1676 8588
rect 1728 8576 1734 8628
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 3329 8619 3387 8625
rect 3329 8616 3341 8619
rect 2924 8588 3341 8616
rect 2924 8576 2930 8588
rect 3329 8585 3341 8588
rect 3375 8585 3387 8619
rect 3329 8579 3387 8585
rect 5077 8619 5135 8625
rect 5077 8585 5089 8619
rect 5123 8616 5135 8619
rect 5166 8616 5172 8628
rect 5123 8588 5172 8616
rect 5123 8585 5135 8588
rect 5077 8579 5135 8585
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 5307 8619 5365 8625
rect 5307 8585 5319 8619
rect 5353 8616 5365 8619
rect 7006 8616 7012 8628
rect 5353 8588 7012 8616
rect 5353 8585 5365 8588
rect 5307 8579 5365 8585
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 7558 8616 7564 8628
rect 7519 8588 7564 8616
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 24670 8616 24676 8628
rect 24631 8588 24676 8616
rect 24670 8576 24676 8588
rect 24728 8576 24734 8628
rect 2958 8548 2964 8560
rect 2919 8520 2964 8548
rect 2958 8508 2964 8520
rect 3016 8508 3022 8560
rect 3418 8508 3424 8560
rect 3476 8548 3482 8560
rect 4341 8551 4399 8557
rect 3476 8520 4200 8548
rect 3476 8508 3482 8520
rect 2314 8480 2320 8492
rect 2275 8452 2320 8480
rect 2314 8440 2320 8452
rect 2372 8440 2378 8492
rect 1464 8415 1522 8421
rect 1464 8381 1476 8415
rect 1510 8412 1522 8415
rect 1762 8412 1768 8424
rect 1510 8384 1768 8412
rect 1510 8381 1522 8384
rect 1464 8375 1522 8381
rect 1762 8372 1768 8384
rect 1820 8412 1826 8424
rect 1857 8415 1915 8421
rect 1857 8412 1869 8415
rect 1820 8384 1869 8412
rect 1820 8372 1826 8384
rect 1857 8381 1869 8384
rect 1903 8381 1915 8415
rect 1857 8375 1915 8381
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 4172 8421 4200 8520
rect 4341 8517 4353 8551
rect 4387 8548 4399 8551
rect 5534 8548 5540 8560
rect 4387 8520 5540 8548
rect 4387 8517 4399 8520
rect 4341 8511 4399 8517
rect 5534 8508 5540 8520
rect 5592 8508 5598 8560
rect 5994 8548 6000 8560
rect 5955 8520 6000 8548
rect 5994 8508 6000 8520
rect 6052 8508 6058 8560
rect 5721 8483 5779 8489
rect 5721 8480 5733 8483
rect 5251 8452 5733 8480
rect 5251 8421 5279 8452
rect 5721 8449 5733 8452
rect 5767 8480 5779 8483
rect 13538 8480 13544 8492
rect 5767 8452 13544 8480
rect 5767 8449 5779 8452
rect 5721 8443 5779 8449
rect 13538 8440 13544 8452
rect 13596 8440 13602 8492
rect 3145 8415 3203 8421
rect 3145 8412 3157 8415
rect 2832 8384 3157 8412
rect 2832 8372 2838 8384
rect 3145 8381 3157 8384
rect 3191 8412 3203 8415
rect 3605 8415 3663 8421
rect 3605 8412 3617 8415
rect 3191 8384 3617 8412
rect 3191 8381 3203 8384
rect 3145 8375 3203 8381
rect 3605 8381 3617 8384
rect 3651 8381 3663 8415
rect 3605 8375 3663 8381
rect 4166 8415 4224 8421
rect 4166 8381 4178 8415
rect 4212 8412 4224 8415
rect 4617 8415 4675 8421
rect 4617 8412 4629 8415
rect 4212 8384 4629 8412
rect 4212 8381 4224 8384
rect 4166 8375 4224 8381
rect 4617 8381 4629 8384
rect 4663 8381 4675 8415
rect 4617 8375 4675 8381
rect 5236 8415 5294 8421
rect 5236 8381 5248 8415
rect 5282 8381 5294 8415
rect 5236 8375 5294 8381
rect 5251 8344 5279 8375
rect 4126 8316 5279 8344
rect 1394 8236 1400 8288
rect 1452 8276 1458 8288
rect 4126 8276 4154 8316
rect 1452 8248 4154 8276
rect 1452 8236 1458 8248
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 842 8032 848 8084
rect 900 8072 906 8084
rect 1581 8075 1639 8081
rect 1581 8072 1593 8075
rect 900 8044 1593 8072
rect 900 8032 906 8044
rect 1581 8041 1593 8044
rect 1627 8041 1639 8075
rect 1581 8035 1639 8041
rect 4249 8075 4307 8081
rect 4249 8041 4261 8075
rect 4295 8072 4307 8075
rect 4430 8072 4436 8084
rect 4295 8044 4436 8072
rect 4295 8041 4307 8044
rect 4249 8035 4307 8041
rect 4430 8032 4436 8044
rect 4488 8032 4494 8084
rect 5261 8075 5319 8081
rect 5261 8041 5273 8075
rect 5307 8072 5319 8075
rect 7466 8072 7472 8084
rect 5307 8044 7472 8072
rect 5307 8041 5319 8044
rect 5261 8035 5319 8041
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7905 1455 7939
rect 1397 7899 1455 7905
rect 1412 7868 1440 7899
rect 3142 7896 3148 7948
rect 3200 7936 3206 7948
rect 4062 7936 4068 7948
rect 3200 7908 4068 7936
rect 3200 7896 3206 7908
rect 4062 7896 4068 7908
rect 4120 7896 4126 7948
rect 4890 7896 4896 7948
rect 4948 7936 4954 7948
rect 5077 7939 5135 7945
rect 5077 7936 5089 7939
rect 4948 7908 5089 7936
rect 4948 7896 4954 7908
rect 5077 7905 5089 7908
rect 5123 7905 5135 7939
rect 5077 7899 5135 7905
rect 1486 7868 1492 7880
rect 1412 7840 1492 7868
rect 1486 7828 1492 7840
rect 1544 7828 1550 7880
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1486 7488 1492 7540
rect 1544 7528 1550 7540
rect 1581 7531 1639 7537
rect 1581 7528 1593 7531
rect 1544 7500 1593 7528
rect 1544 7488 1550 7500
rect 1581 7497 1593 7500
rect 1627 7497 1639 7531
rect 4062 7528 4068 7540
rect 4023 7500 4068 7528
rect 1581 7491 1639 7497
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 4890 7488 4896 7540
rect 4948 7528 4954 7540
rect 5077 7531 5135 7537
rect 5077 7528 5089 7531
rect 4948 7500 5089 7528
rect 4948 7488 4954 7500
rect 5077 7497 5089 7500
rect 5123 7497 5135 7531
rect 5077 7491 5135 7497
rect 24765 7463 24823 7469
rect 24765 7429 24777 7463
rect 24811 7460 24823 7463
rect 27614 7460 27620 7472
rect 24811 7432 27620 7460
rect 24811 7429 24823 7432
rect 24765 7423 24823 7429
rect 27614 7420 27620 7432
rect 27672 7420 27678 7472
rect 24210 7284 24216 7336
rect 24268 7324 24274 7336
rect 24581 7327 24639 7333
rect 24581 7324 24593 7327
rect 24268 7296 24593 7324
rect 24268 7284 24274 7296
rect 24581 7293 24593 7296
rect 24627 7324 24639 7327
rect 25133 7327 25191 7333
rect 25133 7324 25145 7327
rect 24627 7296 25145 7324
rect 24627 7293 24639 7296
rect 24581 7287 24639 7293
rect 25133 7293 25145 7296
rect 25179 7293 25191 7327
rect 25133 7287 25191 7293
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1578 6984 1584 6996
rect 1539 6956 1584 6984
rect 1578 6944 1584 6956
rect 1636 6944 1642 6996
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1394 6400 1400 6452
rect 1452 6440 1458 6452
rect 1581 6443 1639 6449
rect 1581 6440 1593 6443
rect 1452 6412 1593 6440
rect 1452 6400 1458 6412
rect 1581 6409 1593 6412
rect 1627 6409 1639 6443
rect 1581 6403 1639 6409
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 24765 5899 24823 5905
rect 24765 5865 24777 5899
rect 24811 5896 24823 5899
rect 27522 5896 27528 5908
rect 24811 5868 27528 5896
rect 24811 5865 24823 5868
rect 24765 5859 24823 5865
rect 27522 5856 27528 5868
rect 27580 5856 27586 5908
rect 24118 5720 24124 5772
rect 24176 5760 24182 5772
rect 24581 5763 24639 5769
rect 24581 5760 24593 5763
rect 24176 5732 24593 5760
rect 24176 5720 24182 5732
rect 24581 5729 24593 5732
rect 24627 5760 24639 5763
rect 24670 5760 24676 5772
rect 24627 5732 24676 5760
rect 24627 5729 24639 5732
rect 24581 5723 24639 5729
rect 24670 5720 24676 5732
rect 24728 5720 24734 5772
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 24670 5352 24676 5364
rect 24631 5324 24676 5352
rect 24670 5312 24676 5324
rect 24728 5312 24734 5364
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 3050 2932 3056 2984
rect 3108 2972 3114 2984
rect 3916 2975 3974 2981
rect 3916 2972 3928 2975
rect 3108 2944 3928 2972
rect 3108 2932 3114 2944
rect 3916 2941 3928 2944
rect 3962 2972 3974 2975
rect 4341 2975 4399 2981
rect 4341 2972 4353 2975
rect 3962 2944 4353 2972
rect 3962 2941 3974 2944
rect 3916 2935 3974 2941
rect 4341 2941 4353 2944
rect 4387 2941 4399 2975
rect 4341 2935 4399 2941
rect 4019 2839 4077 2845
rect 4019 2805 4031 2839
rect 4065 2836 4077 2839
rect 8938 2836 8944 2848
rect 4065 2808 8944 2836
rect 4065 2805 4077 2808
rect 4019 2799 4077 2805
rect 8938 2796 8944 2808
rect 8996 2796 9002 2848
rect 14274 2796 14280 2848
rect 14332 2836 14338 2848
rect 19242 2836 19248 2848
rect 14332 2808 19248 2836
rect 14332 2796 14338 2808
rect 19242 2796 19248 2808
rect 19300 2796 19306 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 7055 2635 7113 2641
rect 7055 2601 7067 2635
rect 7101 2632 7113 2635
rect 7834 2632 7840 2644
rect 7101 2604 7840 2632
rect 7101 2601 7113 2604
rect 7055 2595 7113 2601
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 8110 2592 8116 2644
rect 8168 2632 8174 2644
rect 8205 2635 8263 2641
rect 8205 2632 8217 2635
rect 8168 2604 8217 2632
rect 8168 2592 8174 2604
rect 8205 2601 8217 2604
rect 8251 2601 8263 2635
rect 8205 2595 8263 2601
rect 11655 2635 11713 2641
rect 11655 2601 11667 2635
rect 11701 2632 11713 2635
rect 12158 2632 12164 2644
rect 11701 2604 12164 2632
rect 11701 2601 11713 2604
rect 11655 2595 11713 2601
rect 12158 2592 12164 2604
rect 12216 2592 12222 2644
rect 21358 2592 21364 2644
rect 21416 2632 21422 2644
rect 21453 2635 21511 2641
rect 21453 2632 21465 2635
rect 21416 2604 21465 2632
rect 21416 2592 21422 2604
rect 21453 2601 21465 2604
rect 21499 2601 21511 2635
rect 21453 2595 21511 2601
rect 24765 2635 24823 2641
rect 24765 2601 24777 2635
rect 24811 2632 24823 2635
rect 24946 2632 24952 2644
rect 24811 2604 24952 2632
rect 24811 2601 24823 2604
rect 24765 2595 24823 2601
rect 24946 2592 24952 2604
rect 25004 2592 25010 2644
rect 5534 2524 5540 2576
rect 5592 2564 5598 2576
rect 5592 2536 11627 2564
rect 5592 2524 5598 2536
rect 6984 2499 7042 2505
rect 6984 2465 6996 2499
rect 7030 2496 7042 2499
rect 7374 2496 7380 2508
rect 7030 2468 7380 2496
rect 7030 2465 7042 2468
rect 6984 2459 7042 2465
rect 7374 2456 7380 2468
rect 7432 2456 7438 2508
rect 11599 2505 11627 2536
rect 19242 2524 19248 2576
rect 19300 2564 19306 2576
rect 19300 2536 24624 2564
rect 19300 2524 19306 2536
rect 7996 2499 8054 2505
rect 7996 2465 8008 2499
rect 8042 2496 8054 2499
rect 11584 2499 11642 2505
rect 8042 2468 8524 2496
rect 8042 2465 8054 2468
rect 7996 2459 8054 2465
rect 7374 2292 7380 2304
rect 7335 2264 7380 2292
rect 7374 2252 7380 2264
rect 7432 2252 7438 2304
rect 8496 2301 8524 2468
rect 11584 2465 11596 2499
rect 11630 2496 11642 2499
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11630 2468 11989 2496
rect 11630 2465 11642 2468
rect 11584 2459 11642 2465
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 14090 2496 14096 2508
rect 14051 2468 14096 2496
rect 11977 2459 12035 2465
rect 14090 2456 14096 2468
rect 14148 2496 14154 2508
rect 24596 2505 24624 2536
rect 14645 2499 14703 2505
rect 14645 2496 14657 2499
rect 14148 2468 14657 2496
rect 14148 2456 14154 2468
rect 14645 2465 14657 2468
rect 14691 2465 14703 2499
rect 14645 2459 14703 2465
rect 18325 2499 18383 2505
rect 18325 2465 18337 2499
rect 18371 2465 18383 2499
rect 18325 2459 18383 2465
rect 21244 2499 21302 2505
rect 21244 2465 21256 2499
rect 21290 2496 21302 2499
rect 22808 2499 22866 2505
rect 21290 2468 21772 2496
rect 21290 2465 21302 2468
rect 21244 2459 21302 2465
rect 18340 2428 18368 2459
rect 18874 2428 18880 2440
rect 18340 2400 18880 2428
rect 18874 2388 18880 2400
rect 18932 2388 18938 2440
rect 14277 2363 14335 2369
rect 14277 2329 14289 2363
rect 14323 2360 14335 2363
rect 16114 2360 16120 2372
rect 14323 2332 16120 2360
rect 14323 2329 14335 2332
rect 14277 2323 14335 2329
rect 16114 2320 16120 2332
rect 16172 2320 16178 2372
rect 18509 2363 18567 2369
rect 18509 2329 18521 2363
rect 18555 2360 18567 2363
rect 20070 2360 20076 2372
rect 18555 2332 20076 2360
rect 18555 2329 18567 2332
rect 18509 2323 18567 2329
rect 20070 2320 20076 2332
rect 20128 2320 20134 2372
rect 8481 2295 8539 2301
rect 8481 2261 8493 2295
rect 8527 2292 8539 2295
rect 9214 2292 9220 2304
rect 8527 2264 9220 2292
rect 8527 2261 8539 2264
rect 8481 2255 8539 2261
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 21744 2301 21772 2468
rect 22808 2465 22820 2499
rect 22854 2496 22866 2499
rect 23201 2499 23259 2505
rect 23201 2496 23213 2499
rect 22854 2468 23213 2496
rect 22854 2465 22866 2468
rect 22808 2459 22866 2465
rect 23201 2465 23213 2468
rect 23247 2496 23259 2499
rect 24581 2499 24639 2505
rect 23247 2468 23474 2496
rect 23247 2465 23259 2468
rect 23201 2459 23259 2465
rect 23446 2428 23474 2468
rect 24581 2465 24593 2499
rect 24627 2496 24639 2499
rect 25133 2499 25191 2505
rect 25133 2496 25145 2499
rect 24627 2468 25145 2496
rect 24627 2465 24639 2468
rect 24581 2459 24639 2465
rect 25133 2465 25145 2468
rect 25179 2465 25191 2499
rect 25133 2459 25191 2465
rect 24762 2428 24768 2440
rect 23446 2400 24768 2428
rect 24762 2388 24768 2400
rect 24820 2388 24826 2440
rect 21729 2295 21787 2301
rect 21729 2261 21741 2295
rect 21775 2292 21787 2295
rect 22094 2292 22100 2304
rect 21775 2264 22100 2292
rect 21775 2261 21787 2264
rect 21729 2255 21787 2261
rect 22094 2252 22100 2264
rect 22152 2252 22158 2304
rect 22186 2252 22192 2304
rect 22244 2292 22250 2304
rect 22879 2295 22937 2301
rect 22879 2292 22891 2295
rect 22244 2264 22891 2292
rect 22244 2252 22250 2264
rect 22879 2261 22891 2264
rect 22925 2261 22937 2295
rect 22879 2255 22937 2261
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 15838 184 15844 196
rect 11716 156 15844 184
rect 11716 128 11744 156
rect 15838 144 15844 156
rect 15896 144 15902 196
rect 11698 76 11704 128
rect 11756 76 11762 128
<< via1 >>
rect 24952 27480 25004 27532
rect 25964 27480 26016 27532
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 12164 25304 12216 25356
rect 12716 25347 12768 25356
rect 12716 25313 12734 25347
rect 12734 25313 12768 25347
rect 12716 25304 12768 25313
rect 27620 25304 27672 25356
rect 5632 25168 5684 25220
rect 6552 25168 6604 25220
rect 9404 25168 9456 25220
rect 13544 25168 13596 25220
rect 12440 25100 12492 25152
rect 12532 25100 12584 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 12716 24939 12768 24948
rect 12716 24905 12725 24939
rect 12725 24905 12759 24939
rect 12759 24905 12768 24939
rect 12716 24896 12768 24905
rect 13268 24896 13320 24948
rect 1860 24735 1912 24744
rect 1860 24701 1869 24735
rect 1869 24701 1903 24735
rect 1903 24701 1912 24735
rect 1860 24692 1912 24701
rect 8668 24624 8720 24676
rect 14096 24692 14148 24744
rect 15200 24735 15252 24744
rect 15200 24701 15209 24735
rect 15209 24701 15243 24735
rect 15243 24701 15252 24735
rect 15200 24692 15252 24701
rect 12256 24624 12308 24676
rect 15384 24624 15436 24676
rect 11336 24556 11388 24608
rect 12164 24599 12216 24608
rect 12164 24565 12173 24599
rect 12173 24565 12207 24599
rect 12207 24565 12216 24599
rect 12164 24556 12216 24565
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 11612 24395 11664 24404
rect 11612 24361 11621 24395
rect 11621 24361 11655 24395
rect 11655 24361 11664 24395
rect 11612 24352 11664 24361
rect 14556 24352 14608 24404
rect 112 24148 164 24200
rect 6092 24216 6144 24268
rect 6920 24259 6972 24268
rect 6920 24225 6929 24259
rect 6929 24225 6963 24259
rect 6963 24225 6972 24259
rect 6920 24216 6972 24225
rect 11336 24216 11388 24268
rect 12440 24216 12492 24268
rect 13452 24216 13504 24268
rect 15752 24216 15804 24268
rect 16948 24216 17000 24268
rect 18604 24216 18656 24268
rect 21456 24216 21508 24268
rect 1952 24148 2004 24200
rect 2044 24148 2096 24200
rect 6828 24080 6880 24132
rect 15936 24123 15988 24132
rect 15936 24089 15945 24123
rect 15945 24089 15979 24123
rect 15979 24089 15988 24123
rect 15936 24080 15988 24089
rect 6000 24012 6052 24064
rect 6460 24012 6512 24064
rect 10600 24055 10652 24064
rect 10600 24021 10609 24055
rect 10609 24021 10643 24055
rect 10643 24021 10652 24055
rect 10600 24012 10652 24021
rect 14188 24055 14240 24064
rect 14188 24021 14197 24055
rect 14197 24021 14231 24055
rect 14231 24021 14240 24055
rect 14188 24012 14240 24021
rect 16212 24012 16264 24064
rect 16304 24012 16356 24064
rect 18880 24012 18932 24064
rect 20352 24012 20404 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1952 23808 2004 23860
rect 6644 23808 6696 23860
rect 11336 23808 11388 23860
rect 13452 23851 13504 23860
rect 13452 23817 13461 23851
rect 13461 23817 13495 23851
rect 13495 23817 13504 23851
rect 13452 23808 13504 23817
rect 15752 23808 15804 23860
rect 17316 23808 17368 23860
rect 19340 23808 19392 23860
rect 20904 23808 20956 23860
rect 21456 23851 21508 23860
rect 21456 23817 21465 23851
rect 21465 23817 21499 23851
rect 21499 23817 21508 23851
rect 21456 23808 21508 23817
rect 8208 23740 8260 23792
rect 18604 23783 18656 23792
rect 18604 23749 18613 23783
rect 18613 23749 18647 23783
rect 18647 23749 18656 23783
rect 18604 23740 18656 23749
rect 4804 23672 4856 23724
rect 6092 23672 6144 23724
rect 12532 23715 12584 23724
rect 12532 23681 12541 23715
rect 12541 23681 12575 23715
rect 12575 23681 12584 23715
rect 12532 23672 12584 23681
rect 12808 23715 12860 23724
rect 12808 23681 12817 23715
rect 12817 23681 12851 23715
rect 12851 23681 12860 23715
rect 12808 23672 12860 23681
rect 14648 23715 14700 23724
rect 14648 23681 14657 23715
rect 14657 23681 14691 23715
rect 14691 23681 14700 23715
rect 14648 23672 14700 23681
rect 15936 23715 15988 23724
rect 15936 23681 15945 23715
rect 15945 23681 15979 23715
rect 15979 23681 15988 23715
rect 15936 23672 15988 23681
rect 16120 23672 16172 23724
rect 1492 23604 1544 23656
rect 2228 23604 2280 23656
rect 3148 23604 3200 23656
rect 6644 23604 6696 23656
rect 8484 23647 8536 23656
rect 8484 23613 8502 23647
rect 8502 23613 8536 23647
rect 8484 23604 8536 23613
rect 10600 23647 10652 23656
rect 10600 23613 10609 23647
rect 10609 23613 10643 23647
rect 10643 23613 10652 23647
rect 10600 23604 10652 23613
rect 10968 23647 11020 23656
rect 10968 23613 10977 23647
rect 10977 23613 11011 23647
rect 11011 23613 11020 23647
rect 10968 23604 11020 23613
rect 13820 23604 13872 23656
rect 14188 23604 14240 23656
rect 17776 23604 17828 23656
rect 19340 23604 19392 23656
rect 24676 23808 24728 23860
rect 27252 23808 27304 23860
rect 6276 23536 6328 23588
rect 6920 23536 6972 23588
rect 11060 23536 11112 23588
rect 16948 23579 17000 23588
rect 112 23468 164 23520
rect 3516 23468 3568 23520
rect 3792 23468 3844 23520
rect 7748 23468 7800 23520
rect 8392 23468 8444 23520
rect 10968 23468 11020 23520
rect 11336 23468 11388 23520
rect 12716 23468 12768 23520
rect 15752 23511 15804 23520
rect 15752 23477 15761 23511
rect 15761 23477 15795 23511
rect 15795 23477 15804 23511
rect 16948 23545 16957 23579
rect 16957 23545 16991 23579
rect 16991 23545 17000 23579
rect 16948 23536 17000 23545
rect 23388 23536 23440 23588
rect 15752 23468 15804 23477
rect 20904 23468 20956 23520
rect 22744 23468 22796 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 8668 23307 8720 23316
rect 8668 23273 8677 23307
rect 8677 23273 8711 23307
rect 8711 23273 8720 23307
rect 8668 23264 8720 23273
rect 12532 23307 12584 23316
rect 12532 23273 12541 23307
rect 12541 23273 12575 23307
rect 12575 23273 12584 23307
rect 12532 23264 12584 23273
rect 16304 23307 16356 23316
rect 16304 23273 16313 23307
rect 16313 23273 16347 23307
rect 16347 23273 16356 23307
rect 16304 23264 16356 23273
rect 18880 23307 18932 23316
rect 18880 23273 18889 23307
rect 18889 23273 18923 23307
rect 18923 23273 18932 23307
rect 18880 23264 18932 23273
rect 10416 23196 10468 23248
rect 12716 23196 12768 23248
rect 15476 23239 15528 23248
rect 15476 23205 15485 23239
rect 15485 23205 15519 23239
rect 15519 23205 15528 23239
rect 15476 23196 15528 23205
rect 16212 23196 16264 23248
rect 16948 23239 17000 23248
rect 16948 23205 16957 23239
rect 16957 23205 16991 23239
rect 16991 23205 17000 23239
rect 16948 23196 17000 23205
rect 17040 23239 17092 23248
rect 17040 23205 17049 23239
rect 17049 23205 17083 23239
rect 17083 23205 17092 23239
rect 17040 23196 17092 23205
rect 17316 23196 17368 23248
rect 18236 23196 18288 23248
rect 20 22924 72 22976
rect 2320 23128 2372 23180
rect 2780 23128 2832 23180
rect 4896 23128 4948 23180
rect 8024 23128 8076 23180
rect 13728 23171 13780 23180
rect 13728 23137 13737 23171
rect 13737 23137 13771 23171
rect 13771 23137 13780 23171
rect 13728 23128 13780 23137
rect 14188 23171 14240 23180
rect 14188 23137 14197 23171
rect 14197 23137 14231 23171
rect 14231 23137 14240 23171
rect 14188 23128 14240 23137
rect 21364 23196 21416 23248
rect 22560 23128 22612 23180
rect 6092 23060 6144 23112
rect 11704 23060 11756 23112
rect 14832 23060 14884 23112
rect 15384 23103 15436 23112
rect 15384 23069 15393 23103
rect 15393 23069 15427 23103
rect 15427 23069 15436 23103
rect 15384 23060 15436 23069
rect 15660 23103 15712 23112
rect 15660 23069 15669 23103
rect 15669 23069 15703 23103
rect 15703 23069 15712 23103
rect 15660 23060 15712 23069
rect 16120 23060 16172 23112
rect 20996 23103 21048 23112
rect 20996 23069 21005 23103
rect 21005 23069 21039 23103
rect 21039 23069 21048 23103
rect 20996 23060 21048 23069
rect 21272 23103 21324 23112
rect 21272 23069 21281 23103
rect 21281 23069 21315 23103
rect 21315 23069 21324 23103
rect 21272 23060 21324 23069
rect 9496 22992 9548 23044
rect 12072 23035 12124 23044
rect 12072 23001 12081 23035
rect 12081 23001 12115 23035
rect 12115 23001 12124 23035
rect 12072 22992 12124 23001
rect 2320 22924 2372 22976
rect 3240 22924 3292 22976
rect 4988 22924 5040 22976
rect 5264 22967 5316 22976
rect 5264 22933 5273 22967
rect 5273 22933 5307 22967
rect 5307 22933 5316 22967
rect 5264 22924 5316 22933
rect 6736 22967 6788 22976
rect 6736 22933 6745 22967
rect 6745 22933 6779 22967
rect 6779 22933 6788 22967
rect 6736 22924 6788 22933
rect 8576 22924 8628 22976
rect 12532 22924 12584 22976
rect 12808 22967 12860 22976
rect 12808 22933 12817 22967
rect 12817 22933 12851 22967
rect 12851 22933 12860 22967
rect 12808 22924 12860 22933
rect 18328 22924 18380 22976
rect 21088 22924 21140 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 2780 22763 2832 22772
rect 2780 22729 2789 22763
rect 2789 22729 2823 22763
rect 2823 22729 2832 22763
rect 2780 22720 2832 22729
rect 11704 22763 11756 22772
rect 11704 22729 11713 22763
rect 11713 22729 11747 22763
rect 11747 22729 11756 22763
rect 11704 22720 11756 22729
rect 13728 22763 13780 22772
rect 13728 22729 13737 22763
rect 13737 22729 13771 22763
rect 13771 22729 13780 22763
rect 13728 22720 13780 22729
rect 16948 22720 17000 22772
rect 18236 22763 18288 22772
rect 18236 22729 18245 22763
rect 18245 22729 18279 22763
rect 18279 22729 18288 22763
rect 18236 22720 18288 22729
rect 20996 22720 21048 22772
rect 22560 22763 22612 22772
rect 22560 22729 22569 22763
rect 22569 22729 22603 22763
rect 22603 22729 22612 22763
rect 22560 22720 22612 22729
rect 4896 22652 4948 22704
rect 8484 22652 8536 22704
rect 12164 22652 12216 22704
rect 13268 22652 13320 22704
rect 8668 22584 8720 22636
rect 1768 22491 1820 22500
rect 1768 22457 1777 22491
rect 1777 22457 1811 22491
rect 1811 22457 1820 22491
rect 1768 22448 1820 22457
rect 3148 22516 3200 22568
rect 5264 22559 5316 22568
rect 5264 22525 5273 22559
rect 5273 22525 5307 22559
rect 5307 22525 5316 22559
rect 5264 22516 5316 22525
rect 13912 22584 13964 22636
rect 14372 22627 14424 22636
rect 14372 22593 14381 22627
rect 14381 22593 14415 22627
rect 14415 22593 14424 22627
rect 14372 22584 14424 22593
rect 15660 22584 15712 22636
rect 16304 22652 16356 22704
rect 16212 22627 16264 22636
rect 16212 22593 16221 22627
rect 16221 22593 16255 22627
rect 16255 22593 16264 22627
rect 16212 22584 16264 22593
rect 6184 22448 6236 22500
rect 1952 22380 2004 22432
rect 3056 22380 3108 22432
rect 6368 22380 6420 22432
rect 6736 22380 6788 22432
rect 7564 22380 7616 22432
rect 11336 22516 11388 22568
rect 8576 22448 8628 22500
rect 8944 22491 8996 22500
rect 8944 22457 8953 22491
rect 8953 22457 8987 22491
rect 8987 22457 8996 22491
rect 12532 22491 12584 22500
rect 8944 22448 8996 22457
rect 12532 22457 12541 22491
rect 12541 22457 12575 22491
rect 12575 22457 12584 22491
rect 12532 22448 12584 22457
rect 12624 22491 12676 22500
rect 12624 22457 12633 22491
rect 12633 22457 12667 22491
rect 12667 22457 12676 22491
rect 14464 22491 14516 22500
rect 12624 22448 12676 22457
rect 14464 22457 14473 22491
rect 14473 22457 14507 22491
rect 14507 22457 14516 22491
rect 14464 22448 14516 22457
rect 15476 22448 15528 22500
rect 7840 22380 7892 22432
rect 8024 22423 8076 22432
rect 8024 22389 8033 22423
rect 8033 22389 8067 22423
rect 8067 22389 8076 22423
rect 8024 22380 8076 22389
rect 11152 22380 11204 22432
rect 12716 22380 12768 22432
rect 14188 22380 14240 22432
rect 17040 22584 17092 22636
rect 18880 22652 18932 22704
rect 18972 22652 19024 22704
rect 21364 22695 21416 22704
rect 21364 22661 21373 22695
rect 21373 22661 21407 22695
rect 21407 22661 21416 22695
rect 21364 22652 21416 22661
rect 20352 22627 20404 22636
rect 20352 22593 20361 22627
rect 20361 22593 20395 22627
rect 20395 22593 20404 22627
rect 20352 22584 20404 22593
rect 21272 22584 21324 22636
rect 19984 22448 20036 22500
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 7748 22176 7800 22228
rect 1952 22108 2004 22160
rect 6092 22151 6144 22160
rect 6092 22117 6101 22151
rect 6101 22117 6135 22151
rect 6135 22117 6144 22151
rect 6092 22108 6144 22117
rect 6184 22151 6236 22160
rect 6184 22117 6193 22151
rect 6193 22117 6227 22151
rect 6227 22117 6236 22151
rect 7932 22176 7984 22228
rect 12624 22176 12676 22228
rect 14372 22176 14424 22228
rect 15384 22176 15436 22228
rect 20352 22219 20404 22228
rect 20352 22185 20361 22219
rect 20361 22185 20395 22219
rect 20395 22185 20404 22219
rect 20352 22176 20404 22185
rect 6184 22108 6236 22117
rect 11244 22108 11296 22160
rect 13452 22108 13504 22160
rect 14464 22108 14516 22160
rect 15292 22108 15344 22160
rect 15752 22108 15804 22160
rect 16212 22108 16264 22160
rect 18328 22151 18380 22160
rect 18328 22117 18337 22151
rect 18337 22117 18371 22151
rect 18371 22117 18380 22151
rect 18328 22108 18380 22117
rect 18420 22151 18472 22160
rect 18420 22117 18429 22151
rect 18429 22117 18463 22151
rect 18463 22117 18472 22151
rect 18420 22108 18472 22117
rect 20996 22108 21048 22160
rect 4620 22083 4672 22092
rect 4620 22049 4629 22083
rect 4629 22049 4663 22083
rect 4663 22049 4672 22083
rect 4620 22040 4672 22049
rect 9588 22083 9640 22092
rect 9588 22049 9597 22083
rect 9597 22049 9631 22083
rect 9631 22049 9640 22083
rect 9588 22040 9640 22049
rect 1860 21972 1912 22024
rect 2504 21972 2556 22024
rect 6368 22015 6420 22024
rect 6368 21981 6377 22015
rect 6377 21981 6411 22015
rect 6411 21981 6420 22015
rect 6368 21972 6420 21981
rect 8760 22015 8812 22024
rect 8760 21981 8769 22015
rect 8769 21981 8803 22015
rect 8803 21981 8812 22015
rect 8760 21972 8812 21981
rect 11152 22015 11204 22024
rect 11152 21981 11161 22015
rect 11161 21981 11195 22015
rect 11195 21981 11204 22015
rect 11152 21972 11204 21981
rect 12992 22015 13044 22024
rect 12992 21981 13001 22015
rect 13001 21981 13035 22015
rect 13035 21981 13044 22015
rect 12992 21972 13044 21981
rect 13268 22015 13320 22024
rect 13268 21981 13277 22015
rect 13277 21981 13311 22015
rect 13311 21981 13320 22015
rect 13268 21972 13320 21981
rect 15936 21972 15988 22024
rect 18972 22015 19024 22024
rect 18972 21981 18981 22015
rect 18981 21981 19015 22015
rect 19015 21981 19024 22015
rect 18972 21972 19024 21981
rect 21088 21972 21140 22024
rect 21272 22015 21324 22024
rect 21272 21981 21281 22015
rect 21281 21981 21315 22015
rect 21315 21981 21324 22015
rect 21272 21972 21324 21981
rect 6828 21904 6880 21956
rect 11336 21904 11388 21956
rect 12072 21904 12124 21956
rect 19892 21947 19944 21956
rect 19892 21913 19901 21947
rect 19901 21913 19935 21947
rect 19935 21913 19944 21947
rect 19892 21904 19944 21913
rect 3608 21879 3660 21888
rect 3608 21845 3617 21879
rect 3617 21845 3651 21879
rect 3651 21845 3660 21879
rect 3608 21836 3660 21845
rect 4712 21879 4764 21888
rect 4712 21845 4721 21879
rect 4721 21845 4755 21879
rect 4755 21845 4764 21879
rect 4712 21836 4764 21845
rect 5540 21879 5592 21888
rect 5540 21845 5549 21879
rect 5549 21845 5583 21879
rect 5583 21845 5592 21879
rect 5540 21836 5592 21845
rect 9404 21836 9456 21888
rect 10048 21836 10100 21888
rect 10784 21879 10836 21888
rect 10784 21845 10793 21879
rect 10793 21845 10827 21879
rect 10827 21845 10836 21879
rect 10784 21836 10836 21845
rect 13820 21836 13872 21888
rect 16488 21836 16540 21888
rect 18052 21879 18104 21888
rect 18052 21845 18061 21879
rect 18061 21845 18095 21879
rect 18095 21845 18104 21879
rect 18052 21836 18104 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1768 21675 1820 21684
rect 1768 21641 1777 21675
rect 1777 21641 1811 21675
rect 1811 21641 1820 21675
rect 1768 21632 1820 21641
rect 4620 21675 4672 21684
rect 4620 21641 4629 21675
rect 4629 21641 4663 21675
rect 4663 21641 4672 21675
rect 4620 21632 4672 21641
rect 5264 21632 5316 21684
rect 6184 21675 6236 21684
rect 6184 21641 6193 21675
rect 6193 21641 6227 21675
rect 6227 21641 6236 21675
rect 6184 21632 6236 21641
rect 11152 21632 11204 21684
rect 12440 21632 12492 21684
rect 13544 21632 13596 21684
rect 15476 21632 15528 21684
rect 15936 21675 15988 21684
rect 15936 21641 15945 21675
rect 15945 21641 15979 21675
rect 15979 21641 15988 21675
rect 15936 21632 15988 21641
rect 18328 21632 18380 21684
rect 18420 21632 18472 21684
rect 20996 21632 21048 21684
rect 21916 21675 21968 21684
rect 21916 21641 21925 21675
rect 21925 21641 21959 21675
rect 21959 21641 21968 21675
rect 21916 21632 21968 21641
rect 25136 21675 25188 21684
rect 25136 21641 25145 21675
rect 25145 21641 25179 21675
rect 25179 21641 25188 21675
rect 25136 21632 25188 21641
rect 8392 21564 8444 21616
rect 2044 21539 2096 21548
rect 2044 21505 2053 21539
rect 2053 21505 2087 21539
rect 2087 21505 2096 21539
rect 2044 21496 2096 21505
rect 2504 21539 2556 21548
rect 2504 21505 2513 21539
rect 2513 21505 2547 21539
rect 2547 21505 2556 21539
rect 2504 21496 2556 21505
rect 3884 21539 3936 21548
rect 3884 21505 3893 21539
rect 3893 21505 3927 21539
rect 3927 21505 3936 21539
rect 3884 21496 3936 21505
rect 5540 21496 5592 21548
rect 6368 21496 6420 21548
rect 12072 21564 12124 21616
rect 8760 21539 8812 21548
rect 8760 21505 8769 21539
rect 8769 21505 8803 21539
rect 8803 21505 8812 21539
rect 8760 21496 8812 21505
rect 8944 21496 8996 21548
rect 16580 21564 16632 21616
rect 13268 21496 13320 21548
rect 14648 21539 14700 21548
rect 14648 21505 14657 21539
rect 14657 21505 14691 21539
rect 14691 21505 14700 21539
rect 14648 21496 14700 21505
rect 18052 21539 18104 21548
rect 18052 21505 18061 21539
rect 18061 21505 18095 21539
rect 18095 21505 18104 21539
rect 18052 21496 18104 21505
rect 19892 21539 19944 21548
rect 19892 21505 19901 21539
rect 19901 21505 19935 21539
rect 19935 21505 19944 21539
rect 19892 21496 19944 21505
rect 6000 21428 6052 21480
rect 6920 21428 6972 21480
rect 13544 21428 13596 21480
rect 16488 21471 16540 21480
rect 1768 21360 1820 21412
rect 3608 21403 3660 21412
rect 3608 21369 3617 21403
rect 3617 21369 3651 21403
rect 3651 21369 3660 21403
rect 3608 21360 3660 21369
rect 5356 21403 5408 21412
rect 5356 21369 5365 21403
rect 5365 21369 5399 21403
rect 5399 21369 5408 21403
rect 5356 21360 5408 21369
rect 7472 21360 7524 21412
rect 8576 21403 8628 21412
rect 8576 21369 8585 21403
rect 8585 21369 8619 21403
rect 8619 21369 8628 21403
rect 8576 21360 8628 21369
rect 9772 21360 9824 21412
rect 10048 21403 10100 21412
rect 10048 21369 10057 21403
rect 10057 21369 10091 21403
rect 10091 21369 10100 21403
rect 10048 21360 10100 21369
rect 10140 21403 10192 21412
rect 10140 21369 10149 21403
rect 10149 21369 10183 21403
rect 10183 21369 10192 21403
rect 10140 21360 10192 21369
rect 7932 21292 7984 21344
rect 8668 21292 8720 21344
rect 9588 21292 9640 21344
rect 11244 21335 11296 21344
rect 11244 21301 11253 21335
rect 11253 21301 11287 21335
rect 11287 21301 11296 21335
rect 11244 21292 11296 21301
rect 12164 21335 12216 21344
rect 12164 21301 12173 21335
rect 12173 21301 12207 21335
rect 12207 21301 12216 21335
rect 12992 21360 13044 21412
rect 13452 21335 13504 21344
rect 12164 21292 12216 21301
rect 13452 21301 13461 21335
rect 13461 21301 13495 21335
rect 13495 21301 13504 21335
rect 13452 21292 13504 21301
rect 16488 21437 16497 21471
rect 16497 21437 16531 21471
rect 16531 21437 16540 21471
rect 16488 21428 16540 21437
rect 21916 21428 21968 21480
rect 25136 21428 25188 21480
rect 17132 21360 17184 21412
rect 20536 21403 20588 21412
rect 15384 21292 15436 21344
rect 17776 21335 17828 21344
rect 17776 21301 17785 21335
rect 17785 21301 17819 21335
rect 17819 21301 17828 21335
rect 17776 21292 17828 21301
rect 19524 21292 19576 21344
rect 20536 21369 20545 21403
rect 20545 21369 20579 21403
rect 20579 21369 20588 21403
rect 20536 21360 20588 21369
rect 20444 21292 20496 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 2044 21063 2096 21072
rect 2044 21029 2053 21063
rect 2053 21029 2087 21063
rect 2087 21029 2096 21063
rect 2044 21020 2096 21029
rect 2872 21088 2924 21140
rect 3884 21088 3936 21140
rect 5356 21088 5408 21140
rect 6092 21131 6144 21140
rect 6092 21097 6101 21131
rect 6101 21097 6135 21131
rect 6135 21097 6144 21131
rect 6092 21088 6144 21097
rect 6828 21131 6880 21140
rect 6828 21097 6837 21131
rect 6837 21097 6871 21131
rect 6871 21097 6880 21131
rect 6828 21088 6880 21097
rect 7748 21088 7800 21140
rect 8392 21088 8444 21140
rect 12164 21088 12216 21140
rect 14648 21131 14700 21140
rect 14648 21097 14657 21131
rect 14657 21097 14691 21131
rect 14691 21097 14700 21131
rect 14648 21088 14700 21097
rect 15292 21088 15344 21140
rect 16580 21131 16632 21140
rect 16580 21097 16589 21131
rect 16589 21097 16623 21131
rect 16623 21097 16632 21131
rect 16580 21088 16632 21097
rect 18420 21088 18472 21140
rect 19064 21131 19116 21140
rect 19064 21097 19073 21131
rect 19073 21097 19107 21131
rect 19107 21097 19116 21131
rect 19064 21088 19116 21097
rect 19524 21088 19576 21140
rect 19984 21131 20036 21140
rect 19984 21097 19993 21131
rect 19993 21097 20027 21131
rect 20027 21097 20036 21131
rect 19984 21088 20036 21097
rect 21088 21088 21140 21140
rect 3240 21063 3292 21072
rect 3240 21029 3249 21063
rect 3249 21029 3283 21063
rect 3283 21029 3292 21063
rect 3240 21020 3292 21029
rect 3516 21020 3568 21072
rect 4896 21020 4948 21072
rect 7932 21020 7984 21072
rect 10140 21063 10192 21072
rect 10140 21029 10149 21063
rect 10149 21029 10183 21063
rect 10183 21029 10192 21063
rect 10140 21020 10192 21029
rect 11244 21020 11296 21072
rect 13544 21020 13596 21072
rect 15384 21020 15436 21072
rect 8116 20952 8168 21004
rect 8208 20952 8260 21004
rect 9312 20952 9364 21004
rect 11060 20995 11112 21004
rect 11060 20961 11069 20995
rect 11069 20961 11103 20995
rect 11103 20961 11112 20995
rect 11060 20952 11112 20961
rect 14832 20952 14884 21004
rect 16764 20952 16816 21004
rect 17224 20952 17276 21004
rect 4528 20884 4580 20936
rect 7472 20927 7524 20936
rect 7472 20893 7481 20927
rect 7481 20893 7515 20927
rect 7515 20893 7524 20927
rect 7472 20884 7524 20893
rect 12808 20927 12860 20936
rect 12808 20893 12817 20927
rect 12817 20893 12851 20927
rect 12851 20893 12860 20927
rect 12808 20884 12860 20893
rect 17868 20927 17920 20936
rect 17868 20893 17877 20927
rect 17877 20893 17911 20927
rect 17911 20893 17920 20927
rect 17868 20884 17920 20893
rect 18696 20927 18748 20936
rect 18696 20893 18705 20927
rect 18705 20893 18739 20927
rect 18739 20893 18748 20927
rect 18696 20884 18748 20893
rect 19984 20884 20036 20936
rect 2964 20791 3016 20800
rect 2964 20757 2973 20791
rect 2973 20757 3007 20791
rect 3007 20757 3016 20791
rect 2964 20748 3016 20757
rect 8576 20748 8628 20800
rect 9588 20748 9640 20800
rect 9680 20748 9732 20800
rect 12532 20791 12584 20800
rect 12532 20757 12541 20791
rect 12541 20757 12575 20791
rect 12575 20757 12584 20791
rect 12532 20748 12584 20757
rect 12624 20748 12676 20800
rect 14372 20748 14424 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1584 20587 1636 20596
rect 1584 20553 1593 20587
rect 1593 20553 1627 20587
rect 1627 20553 1636 20587
rect 1584 20544 1636 20553
rect 4712 20544 4764 20596
rect 5264 20544 5316 20596
rect 8024 20544 8076 20596
rect 11244 20544 11296 20596
rect 13728 20544 13780 20596
rect 16764 20587 16816 20596
rect 2872 20451 2924 20460
rect 2872 20417 2881 20451
rect 2881 20417 2915 20451
rect 2915 20417 2924 20451
rect 2872 20408 2924 20417
rect 3332 20451 3384 20460
rect 3332 20417 3341 20451
rect 3341 20417 3375 20451
rect 3375 20417 3384 20451
rect 3332 20408 3384 20417
rect 4988 20408 5040 20460
rect 8760 20476 8812 20528
rect 5540 20451 5592 20460
rect 5540 20417 5549 20451
rect 5549 20417 5583 20451
rect 5583 20417 5592 20451
rect 5540 20408 5592 20417
rect 1400 20383 1452 20392
rect 1400 20349 1409 20383
rect 1409 20349 1443 20383
rect 1443 20349 1452 20383
rect 1400 20340 1452 20349
rect 8668 20408 8720 20460
rect 9220 20408 9272 20460
rect 12532 20451 12584 20460
rect 12532 20417 12541 20451
rect 12541 20417 12575 20451
rect 12575 20417 12584 20451
rect 12532 20408 12584 20417
rect 12992 20476 13044 20528
rect 16764 20553 16773 20587
rect 16773 20553 16807 20587
rect 16807 20553 16816 20587
rect 16764 20544 16816 20553
rect 17132 20587 17184 20596
rect 17132 20553 17141 20587
rect 17141 20553 17175 20587
rect 17175 20553 17184 20587
rect 17132 20544 17184 20553
rect 19892 20544 19944 20596
rect 20996 20544 21048 20596
rect 21640 20544 21692 20596
rect 16212 20476 16264 20528
rect 14004 20408 14056 20460
rect 16580 20408 16632 20460
rect 17868 20408 17920 20460
rect 19984 20451 20036 20460
rect 19984 20417 19993 20451
rect 19993 20417 20027 20451
rect 20027 20417 20036 20451
rect 19984 20408 20036 20417
rect 20260 20408 20312 20460
rect 2964 20315 3016 20324
rect 2964 20281 2973 20315
rect 2973 20281 3007 20315
rect 3007 20281 3016 20315
rect 2964 20272 3016 20281
rect 3700 20272 3752 20324
rect 4896 20315 4948 20324
rect 4896 20281 4905 20315
rect 4905 20281 4939 20315
rect 4939 20281 4948 20315
rect 4896 20272 4948 20281
rect 5264 20315 5316 20324
rect 5264 20281 5273 20315
rect 5273 20281 5307 20315
rect 5307 20281 5316 20315
rect 5264 20272 5316 20281
rect 1952 20247 2004 20256
rect 1952 20213 1961 20247
rect 1961 20213 1995 20247
rect 1995 20213 2004 20247
rect 1952 20204 2004 20213
rect 2044 20204 2096 20256
rect 2596 20204 2648 20256
rect 4528 20204 4580 20256
rect 7748 20272 7800 20324
rect 14372 20340 14424 20392
rect 9496 20272 9548 20324
rect 12624 20315 12676 20324
rect 6184 20204 6236 20256
rect 7932 20204 7984 20256
rect 9128 20247 9180 20256
rect 9128 20213 9137 20247
rect 9137 20213 9171 20247
rect 9171 20213 9180 20247
rect 9128 20204 9180 20213
rect 9312 20204 9364 20256
rect 9588 20204 9640 20256
rect 12624 20281 12633 20315
rect 12633 20281 12667 20315
rect 12667 20281 12676 20315
rect 12624 20272 12676 20281
rect 13544 20247 13596 20256
rect 13544 20213 13553 20247
rect 13553 20213 13587 20247
rect 13587 20213 13596 20247
rect 13544 20204 13596 20213
rect 14096 20247 14148 20256
rect 14096 20213 14105 20247
rect 14105 20213 14139 20247
rect 14139 20213 14148 20247
rect 14096 20204 14148 20213
rect 15384 20247 15436 20256
rect 15384 20213 15393 20247
rect 15393 20213 15427 20247
rect 15427 20213 15436 20247
rect 15384 20204 15436 20213
rect 15752 20204 15804 20256
rect 19064 20272 19116 20324
rect 19984 20272 20036 20324
rect 21548 20315 21600 20324
rect 21548 20281 21557 20315
rect 21557 20281 21591 20315
rect 21591 20281 21600 20315
rect 21548 20272 21600 20281
rect 21640 20315 21692 20324
rect 21640 20281 21649 20315
rect 21649 20281 21683 20315
rect 21683 20281 21692 20315
rect 21640 20272 21692 20281
rect 17776 20247 17828 20256
rect 17776 20213 17785 20247
rect 17785 20213 17819 20247
rect 17819 20213 17828 20247
rect 17776 20204 17828 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 3608 20000 3660 20052
rect 4620 20000 4672 20052
rect 5356 20000 5408 20052
rect 7472 20043 7524 20052
rect 7472 20009 7481 20043
rect 7481 20009 7515 20043
rect 7515 20009 7524 20043
rect 7472 20000 7524 20009
rect 7748 20000 7800 20052
rect 7932 20000 7984 20052
rect 2504 19975 2556 19984
rect 2504 19941 2513 19975
rect 2513 19941 2547 19975
rect 2547 19941 2556 19975
rect 2504 19932 2556 19941
rect 3240 19932 3292 19984
rect 4896 19932 4948 19984
rect 6460 19932 6512 19984
rect 6736 19932 6788 19984
rect 7564 19932 7616 19984
rect 9128 20000 9180 20052
rect 11060 20043 11112 20052
rect 11060 20009 11069 20043
rect 11069 20009 11103 20043
rect 11103 20009 11112 20043
rect 11060 20000 11112 20009
rect 12808 20043 12860 20052
rect 12808 20009 12817 20043
rect 12817 20009 12851 20043
rect 12851 20009 12860 20043
rect 12808 20000 12860 20009
rect 14096 20000 14148 20052
rect 14832 20000 14884 20052
rect 15384 20000 15436 20052
rect 8760 19975 8812 19984
rect 8760 19941 8769 19975
rect 8769 19941 8803 19975
rect 8803 19941 8812 19975
rect 8760 19932 8812 19941
rect 9496 19975 9548 19984
rect 9496 19941 9505 19975
rect 9505 19941 9539 19975
rect 9539 19941 9548 19975
rect 9496 19932 9548 19941
rect 13544 19932 13596 19984
rect 17776 20000 17828 20052
rect 17868 20000 17920 20052
rect 19248 20043 19300 20052
rect 19248 20009 19257 20043
rect 19257 20009 19291 20043
rect 19291 20009 19300 20043
rect 19248 20000 19300 20009
rect 20260 20043 20312 20052
rect 20260 20009 20269 20043
rect 20269 20009 20303 20043
rect 20303 20009 20312 20043
rect 20260 20000 20312 20009
rect 21548 20043 21600 20052
rect 21548 20009 21557 20043
rect 21557 20009 21591 20043
rect 21591 20009 21600 20043
rect 21548 20000 21600 20009
rect 1768 19864 1820 19916
rect 3332 19796 3384 19848
rect 3516 19796 3568 19848
rect 3792 19796 3844 19848
rect 2964 19728 3016 19780
rect 6276 19864 6328 19916
rect 9588 19864 9640 19916
rect 10232 19907 10284 19916
rect 2136 19703 2188 19712
rect 2136 19669 2145 19703
rect 2145 19669 2179 19703
rect 2179 19669 2188 19703
rect 2136 19660 2188 19669
rect 3424 19703 3476 19712
rect 3424 19669 3433 19703
rect 3433 19669 3467 19703
rect 3467 19669 3476 19703
rect 3424 19660 3476 19669
rect 3608 19660 3660 19712
rect 4068 19660 4120 19712
rect 6460 19839 6512 19848
rect 6460 19805 6469 19839
rect 6469 19805 6503 19839
rect 6503 19805 6512 19839
rect 6460 19796 6512 19805
rect 10232 19873 10241 19907
rect 10241 19873 10275 19907
rect 10275 19873 10284 19907
rect 10232 19864 10284 19873
rect 10784 19864 10836 19916
rect 11612 19839 11664 19848
rect 11612 19805 11621 19839
rect 11621 19805 11655 19839
rect 11655 19805 11664 19839
rect 11612 19796 11664 19805
rect 13452 19864 13504 19916
rect 13636 19907 13688 19916
rect 13636 19873 13645 19907
rect 13645 19873 13679 19907
rect 13679 19873 13688 19907
rect 13636 19864 13688 19873
rect 14188 19907 14240 19916
rect 14188 19873 14197 19907
rect 14197 19873 14231 19907
rect 14231 19873 14240 19907
rect 14188 19864 14240 19873
rect 17592 19907 17644 19916
rect 13360 19796 13412 19848
rect 14832 19796 14884 19848
rect 17592 19873 17601 19907
rect 17601 19873 17635 19907
rect 17635 19873 17644 19907
rect 17592 19864 17644 19873
rect 18696 19932 18748 19984
rect 19156 19907 19208 19916
rect 17132 19796 17184 19848
rect 17868 19796 17920 19848
rect 19156 19873 19165 19907
rect 19165 19873 19199 19907
rect 19199 19873 19208 19907
rect 19156 19864 19208 19873
rect 20812 19907 20864 19916
rect 20812 19873 20821 19907
rect 20821 19873 20855 19907
rect 20855 19873 20864 19907
rect 20812 19864 20864 19873
rect 25504 19864 25556 19916
rect 15752 19728 15804 19780
rect 14740 19703 14792 19712
rect 14740 19669 14749 19703
rect 14749 19669 14783 19703
rect 14783 19669 14792 19703
rect 14740 19660 14792 19669
rect 16212 19703 16264 19712
rect 16212 19669 16221 19703
rect 16221 19669 16255 19703
rect 16255 19669 16264 19703
rect 16212 19660 16264 19669
rect 18604 19660 18656 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 2964 19499 3016 19508
rect 2964 19465 2973 19499
rect 2973 19465 3007 19499
rect 3007 19465 3016 19499
rect 2964 19456 3016 19465
rect 3240 19499 3292 19508
rect 3240 19465 3249 19499
rect 3249 19465 3283 19499
rect 3283 19465 3292 19499
rect 3240 19456 3292 19465
rect 3976 19456 4028 19508
rect 6276 19499 6328 19508
rect 6276 19465 6285 19499
rect 6285 19465 6319 19499
rect 6319 19465 6328 19499
rect 6276 19456 6328 19465
rect 10232 19456 10284 19508
rect 10692 19456 10744 19508
rect 13636 19456 13688 19508
rect 15384 19499 15436 19508
rect 15384 19465 15393 19499
rect 15393 19465 15427 19499
rect 15427 19465 15436 19499
rect 15384 19456 15436 19465
rect 16212 19456 16264 19508
rect 17132 19456 17184 19508
rect 18880 19456 18932 19508
rect 19156 19456 19208 19508
rect 25136 19499 25188 19508
rect 25136 19465 25145 19499
rect 25145 19465 25179 19499
rect 25179 19465 25188 19499
rect 25136 19456 25188 19465
rect 25504 19499 25556 19508
rect 25504 19465 25513 19499
rect 25513 19465 25547 19499
rect 25547 19465 25556 19499
rect 25504 19456 25556 19465
rect 6460 19388 6512 19440
rect 12348 19388 12400 19440
rect 13912 19388 13964 19440
rect 17592 19388 17644 19440
rect 18512 19388 18564 19440
rect 21364 19388 21416 19440
rect 1768 19320 1820 19372
rect 2688 19320 2740 19372
rect 3608 19320 3660 19372
rect 3884 19320 3936 19372
rect 3700 19252 3752 19304
rect 3976 19295 4028 19304
rect 3976 19261 3985 19295
rect 3985 19261 4019 19295
rect 4019 19261 4028 19295
rect 3976 19252 4028 19261
rect 4620 19320 4672 19372
rect 5264 19320 5316 19372
rect 5540 19363 5592 19372
rect 5540 19329 5549 19363
rect 5549 19329 5583 19363
rect 5583 19329 5592 19363
rect 5540 19320 5592 19329
rect 9220 19320 9272 19372
rect 10784 19320 10836 19372
rect 11612 19320 11664 19372
rect 4896 19252 4948 19304
rect 7380 19295 7432 19304
rect 7380 19261 7389 19295
rect 7389 19261 7423 19295
rect 7423 19261 7432 19295
rect 7380 19252 7432 19261
rect 2136 19184 2188 19236
rect 2964 19184 3016 19236
rect 3884 19184 3936 19236
rect 5356 19227 5408 19236
rect 5356 19193 5365 19227
rect 5365 19193 5399 19227
rect 5399 19193 5408 19227
rect 5356 19184 5408 19193
rect 5540 19184 5592 19236
rect 9036 19227 9088 19236
rect 6092 19116 6144 19168
rect 6276 19116 6328 19168
rect 8208 19159 8260 19168
rect 8208 19125 8217 19159
rect 8217 19125 8251 19159
rect 8251 19125 8260 19159
rect 9036 19193 9045 19227
rect 9045 19193 9079 19227
rect 9079 19193 9088 19227
rect 9036 19184 9088 19193
rect 8208 19116 8260 19125
rect 8576 19116 8628 19168
rect 9588 19116 9640 19168
rect 9864 19116 9916 19168
rect 11428 19184 11480 19236
rect 12532 19227 12584 19236
rect 12532 19193 12541 19227
rect 12541 19193 12575 19227
rect 12575 19193 12584 19227
rect 12532 19184 12584 19193
rect 12624 19227 12676 19236
rect 12624 19193 12633 19227
rect 12633 19193 12667 19227
rect 12667 19193 12676 19227
rect 13360 19320 13412 19372
rect 14372 19320 14424 19372
rect 14740 19320 14792 19372
rect 16120 19320 16172 19372
rect 20260 19320 20312 19372
rect 20536 19363 20588 19372
rect 20536 19329 20545 19363
rect 20545 19329 20579 19363
rect 20579 19329 20588 19363
rect 20536 19320 20588 19329
rect 21272 19320 21324 19372
rect 13728 19252 13780 19304
rect 14464 19295 14516 19304
rect 14464 19261 14473 19295
rect 14473 19261 14507 19295
rect 14507 19261 14516 19295
rect 14464 19252 14516 19261
rect 17776 19295 17828 19304
rect 17776 19261 17785 19295
rect 17785 19261 17819 19295
rect 17819 19261 17828 19295
rect 17776 19252 17828 19261
rect 18052 19295 18104 19304
rect 18052 19261 18061 19295
rect 18061 19261 18095 19295
rect 18095 19261 18104 19295
rect 18052 19252 18104 19261
rect 22100 19252 22152 19304
rect 25136 19252 25188 19304
rect 12624 19184 12676 19193
rect 11704 19159 11756 19168
rect 11704 19125 11713 19159
rect 11713 19125 11747 19159
rect 11747 19125 11756 19159
rect 11704 19116 11756 19125
rect 13728 19116 13780 19168
rect 16120 19184 16172 19236
rect 16764 19184 16816 19236
rect 18420 19184 18472 19236
rect 19984 19227 20036 19236
rect 19984 19193 19993 19227
rect 19993 19193 20027 19227
rect 20027 19193 20036 19227
rect 19984 19184 20036 19193
rect 17868 19116 17920 19168
rect 20076 19116 20128 19168
rect 20812 19116 20864 19168
rect 21916 19116 21968 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 2596 18955 2648 18964
rect 2596 18921 2605 18955
rect 2605 18921 2639 18955
rect 2639 18921 2648 18955
rect 2596 18912 2648 18921
rect 4068 18912 4120 18964
rect 6184 18955 6236 18964
rect 6184 18921 6193 18955
rect 6193 18921 6227 18955
rect 6227 18921 6236 18955
rect 6184 18912 6236 18921
rect 7564 18912 7616 18964
rect 9220 18912 9272 18964
rect 9680 18912 9732 18964
rect 11704 18955 11756 18964
rect 2136 18844 2188 18896
rect 3792 18844 3844 18896
rect 8208 18887 8260 18896
rect 2596 18776 2648 18828
rect 3424 18776 3476 18828
rect 4620 18819 4672 18828
rect 4620 18785 4629 18819
rect 4629 18785 4663 18819
rect 4663 18785 4672 18819
rect 4620 18776 4672 18785
rect 4712 18776 4764 18828
rect 2412 18708 2464 18760
rect 5080 18708 5132 18760
rect 5448 18776 5500 18828
rect 6276 18819 6328 18828
rect 6276 18785 6285 18819
rect 6285 18785 6319 18819
rect 6319 18785 6328 18819
rect 6276 18776 6328 18785
rect 8208 18853 8217 18887
rect 8217 18853 8251 18887
rect 8251 18853 8260 18887
rect 8208 18844 8260 18853
rect 11704 18921 11713 18955
rect 11713 18921 11747 18955
rect 11747 18921 11756 18955
rect 11704 18912 11756 18921
rect 14832 18912 14884 18964
rect 18052 18912 18104 18964
rect 19248 18912 19300 18964
rect 9864 18887 9916 18896
rect 9864 18853 9873 18887
rect 9873 18853 9907 18887
rect 9907 18853 9916 18887
rect 12624 18887 12676 18896
rect 9864 18844 9916 18853
rect 12624 18853 12633 18887
rect 12633 18853 12667 18887
rect 12667 18853 12676 18887
rect 12624 18844 12676 18853
rect 13820 18844 13872 18896
rect 15752 18887 15804 18896
rect 15752 18853 15761 18887
rect 15761 18853 15795 18887
rect 15795 18853 15804 18887
rect 15752 18844 15804 18853
rect 19156 18887 19208 18896
rect 19156 18853 19165 18887
rect 19165 18853 19199 18887
rect 19199 18853 19208 18887
rect 19156 18844 19208 18853
rect 20168 18844 20220 18896
rect 20536 18844 20588 18896
rect 6552 18776 6604 18828
rect 7932 18776 7984 18828
rect 10784 18819 10836 18828
rect 10784 18785 10793 18819
rect 10793 18785 10827 18819
rect 10827 18785 10836 18819
rect 10784 18776 10836 18785
rect 17868 18819 17920 18828
rect 6000 18708 6052 18760
rect 6828 18751 6880 18760
rect 6828 18717 6837 18751
rect 6837 18717 6871 18751
rect 6871 18717 6880 18751
rect 6828 18708 6880 18717
rect 8116 18751 8168 18760
rect 8116 18717 8125 18751
rect 8125 18717 8159 18751
rect 8159 18717 8168 18751
rect 8116 18708 8168 18717
rect 1952 18640 2004 18692
rect 4712 18640 4764 18692
rect 9128 18640 9180 18692
rect 10968 18708 11020 18760
rect 13544 18708 13596 18760
rect 15476 18708 15528 18760
rect 16028 18751 16080 18760
rect 16028 18717 16037 18751
rect 16037 18717 16071 18751
rect 16071 18717 16080 18751
rect 16028 18708 16080 18717
rect 17868 18785 17877 18819
rect 17877 18785 17911 18819
rect 17911 18785 17920 18819
rect 17868 18776 17920 18785
rect 3792 18572 3844 18624
rect 7656 18572 7708 18624
rect 11428 18640 11480 18692
rect 14556 18683 14608 18692
rect 14556 18649 14565 18683
rect 14565 18649 14599 18683
rect 14599 18649 14608 18683
rect 17960 18708 18012 18760
rect 18696 18708 18748 18760
rect 19064 18751 19116 18760
rect 19064 18717 19073 18751
rect 19073 18717 19107 18751
rect 19107 18717 19116 18751
rect 19064 18708 19116 18717
rect 19248 18708 19300 18760
rect 14556 18640 14608 18649
rect 16672 18640 16724 18692
rect 21732 18640 21784 18692
rect 12348 18572 12400 18624
rect 12532 18572 12584 18624
rect 12992 18615 13044 18624
rect 12992 18581 13001 18615
rect 13001 18581 13035 18615
rect 13035 18581 13044 18615
rect 12992 18572 13044 18581
rect 14188 18615 14240 18624
rect 14188 18581 14197 18615
rect 14197 18581 14231 18615
rect 14231 18581 14240 18615
rect 14188 18572 14240 18581
rect 19984 18615 20036 18624
rect 19984 18581 19993 18615
rect 19993 18581 20027 18615
rect 20027 18581 20036 18615
rect 19984 18572 20036 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 2688 18411 2740 18420
rect 2688 18377 2697 18411
rect 2697 18377 2731 18411
rect 2731 18377 2740 18411
rect 2964 18411 3016 18420
rect 2688 18368 2740 18377
rect 2964 18377 2973 18411
rect 2973 18377 3007 18411
rect 3007 18377 3016 18411
rect 2964 18368 3016 18377
rect 4620 18368 4672 18420
rect 6552 18411 6604 18420
rect 6552 18377 6561 18411
rect 6561 18377 6595 18411
rect 6595 18377 6604 18411
rect 6552 18368 6604 18377
rect 7748 18411 7800 18420
rect 7748 18377 7757 18411
rect 7757 18377 7791 18411
rect 7791 18377 7800 18411
rect 7748 18368 7800 18377
rect 9680 18368 9732 18420
rect 11704 18368 11756 18420
rect 13820 18411 13872 18420
rect 13820 18377 13829 18411
rect 13829 18377 13863 18411
rect 13863 18377 13872 18411
rect 13820 18368 13872 18377
rect 17224 18368 17276 18420
rect 17868 18368 17920 18420
rect 18420 18368 18472 18420
rect 19984 18368 20036 18420
rect 9036 18300 9088 18352
rect 11612 18300 11664 18352
rect 13636 18300 13688 18352
rect 13912 18300 13964 18352
rect 19064 18300 19116 18352
rect 3056 18232 3108 18284
rect 9956 18232 10008 18284
rect 12900 18232 12952 18284
rect 16028 18232 16080 18284
rect 16488 18275 16540 18284
rect 16488 18241 16497 18275
rect 16497 18241 16531 18275
rect 16531 18241 16540 18275
rect 16488 18232 16540 18241
rect 16764 18275 16816 18284
rect 16764 18241 16773 18275
rect 16773 18241 16807 18275
rect 16807 18241 16816 18275
rect 16764 18232 16816 18241
rect 18696 18275 18748 18284
rect 18696 18241 18705 18275
rect 18705 18241 18739 18275
rect 18739 18241 18748 18275
rect 18696 18232 18748 18241
rect 20260 18232 20312 18284
rect 2412 18207 2464 18216
rect 1768 18096 1820 18148
rect 2412 18173 2421 18207
rect 2421 18173 2455 18207
rect 2455 18173 2464 18207
rect 2412 18164 2464 18173
rect 4620 18207 4672 18216
rect 4620 18173 4629 18207
rect 4629 18173 4663 18207
rect 4663 18173 4672 18207
rect 4620 18164 4672 18173
rect 5080 18164 5132 18216
rect 5448 18207 5500 18216
rect 3792 18096 3844 18148
rect 5448 18173 5457 18207
rect 5457 18173 5491 18207
rect 5491 18173 5500 18207
rect 5448 18164 5500 18173
rect 6644 18164 6696 18216
rect 7656 18164 7708 18216
rect 7748 18096 7800 18148
rect 11520 18164 11572 18216
rect 14648 18207 14700 18216
rect 14648 18173 14657 18207
rect 14657 18173 14691 18207
rect 14691 18173 14700 18207
rect 14648 18164 14700 18173
rect 9864 18096 9916 18148
rect 12624 18139 12676 18148
rect 12624 18105 12633 18139
rect 12633 18105 12667 18139
rect 12667 18105 12676 18139
rect 14556 18139 14608 18148
rect 12624 18096 12676 18105
rect 14556 18105 14565 18139
rect 14565 18105 14599 18139
rect 14599 18105 14608 18139
rect 14556 18096 14608 18105
rect 4528 18071 4580 18080
rect 4528 18037 4537 18071
rect 4537 18037 4571 18071
rect 4571 18037 4580 18071
rect 4528 18028 4580 18037
rect 4620 18028 4672 18080
rect 6184 18071 6236 18080
rect 6184 18037 6193 18071
rect 6193 18037 6227 18071
rect 6227 18037 6236 18071
rect 6184 18028 6236 18037
rect 7196 18028 7248 18080
rect 10968 18071 11020 18080
rect 10968 18037 10977 18071
rect 10977 18037 11011 18071
rect 11011 18037 11020 18071
rect 10968 18028 11020 18037
rect 13544 18071 13596 18080
rect 13544 18037 13553 18071
rect 13553 18037 13587 18071
rect 13587 18037 13596 18071
rect 13544 18028 13596 18037
rect 15568 18071 15620 18080
rect 15568 18037 15577 18071
rect 15577 18037 15611 18071
rect 15611 18037 15620 18071
rect 15568 18028 15620 18037
rect 15752 18028 15804 18080
rect 16212 18071 16264 18080
rect 16212 18037 16221 18071
rect 16221 18037 16255 18071
rect 16255 18037 16264 18071
rect 18420 18096 18472 18148
rect 20536 18139 20588 18148
rect 20536 18105 20545 18139
rect 20545 18105 20579 18139
rect 20579 18105 20588 18139
rect 20536 18096 20588 18105
rect 16212 18028 16264 18037
rect 17960 18028 18012 18080
rect 21364 18096 21416 18148
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2596 17867 2648 17876
rect 2596 17833 2605 17867
rect 2605 17833 2639 17867
rect 2639 17833 2648 17867
rect 2596 17824 2648 17833
rect 3056 17824 3108 17876
rect 3976 17824 4028 17876
rect 4528 17824 4580 17876
rect 4804 17867 4856 17876
rect 4804 17833 4813 17867
rect 4813 17833 4847 17867
rect 4847 17833 4856 17867
rect 4804 17824 4856 17833
rect 8116 17824 8168 17876
rect 8208 17824 8260 17876
rect 9956 17867 10008 17876
rect 9956 17833 9965 17867
rect 9965 17833 9999 17867
rect 9999 17833 10008 17867
rect 9956 17824 10008 17833
rect 11428 17824 11480 17876
rect 11612 17867 11664 17876
rect 11612 17833 11621 17867
rect 11621 17833 11655 17867
rect 11655 17833 11664 17867
rect 11612 17824 11664 17833
rect 16212 17867 16264 17876
rect 16212 17833 16221 17867
rect 16221 17833 16255 17867
rect 16255 17833 16264 17867
rect 16212 17824 16264 17833
rect 16488 17867 16540 17876
rect 16488 17833 16497 17867
rect 16497 17833 16531 17867
rect 16531 17833 16540 17867
rect 16488 17824 16540 17833
rect 17224 17867 17276 17876
rect 17224 17833 17233 17867
rect 17233 17833 17267 17867
rect 17267 17833 17276 17867
rect 17224 17824 17276 17833
rect 18420 17824 18472 17876
rect 19156 17824 19208 17876
rect 20536 17867 20588 17876
rect 20536 17833 20545 17867
rect 20545 17833 20579 17867
rect 20579 17833 20588 17867
rect 20536 17824 20588 17833
rect 1768 17731 1820 17740
rect 1768 17697 1777 17731
rect 1777 17697 1811 17731
rect 1811 17697 1820 17731
rect 1768 17688 1820 17697
rect 1952 17688 2004 17740
rect 2504 17731 2556 17740
rect 2504 17697 2513 17731
rect 2513 17697 2547 17731
rect 2547 17697 2556 17731
rect 2504 17688 2556 17697
rect 2872 17688 2924 17740
rect 6276 17756 6328 17808
rect 7748 17799 7800 17808
rect 7748 17765 7757 17799
rect 7757 17765 7791 17799
rect 7791 17765 7800 17799
rect 7748 17756 7800 17765
rect 10968 17799 11020 17808
rect 10968 17765 10977 17799
rect 10977 17765 11011 17799
rect 11011 17765 11020 17799
rect 10968 17756 11020 17765
rect 11888 17756 11940 17808
rect 16028 17756 16080 17808
rect 4528 17688 4580 17740
rect 6092 17731 6144 17740
rect 6092 17697 6101 17731
rect 6101 17697 6135 17731
rect 6135 17697 6144 17731
rect 6092 17688 6144 17697
rect 6736 17688 6788 17740
rect 10140 17688 10192 17740
rect 2596 17620 2648 17672
rect 7472 17663 7524 17672
rect 7472 17629 7481 17663
rect 7481 17629 7515 17663
rect 7515 17629 7524 17663
rect 7472 17620 7524 17629
rect 3516 17552 3568 17604
rect 6920 17552 6972 17604
rect 10600 17688 10652 17740
rect 13544 17688 13596 17740
rect 13728 17688 13780 17740
rect 14096 17731 14148 17740
rect 14096 17697 14105 17731
rect 14105 17697 14139 17731
rect 14139 17697 14148 17731
rect 14096 17688 14148 17697
rect 15476 17688 15528 17740
rect 17040 17731 17092 17740
rect 17040 17697 17049 17731
rect 17049 17697 17083 17731
rect 17083 17697 17092 17731
rect 17040 17688 17092 17697
rect 20628 17688 20680 17740
rect 21364 17688 21416 17740
rect 11612 17620 11664 17672
rect 12164 17663 12216 17672
rect 12164 17629 12173 17663
rect 12173 17629 12207 17663
rect 12207 17629 12216 17663
rect 12164 17620 12216 17629
rect 16304 17620 16356 17672
rect 18144 17663 18196 17672
rect 18144 17629 18153 17663
rect 18153 17629 18187 17663
rect 18187 17629 18196 17663
rect 18144 17620 18196 17629
rect 3424 17527 3476 17536
rect 3424 17493 3433 17527
rect 3433 17493 3467 17527
rect 3467 17493 3476 17527
rect 3424 17484 3476 17493
rect 5540 17484 5592 17536
rect 12900 17527 12952 17536
rect 12900 17493 12909 17527
rect 12909 17493 12943 17527
rect 12943 17493 12952 17527
rect 12900 17484 12952 17493
rect 14648 17552 14700 17604
rect 18972 17552 19024 17604
rect 14004 17484 14056 17536
rect 15936 17484 15988 17536
rect 19432 17484 19484 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2504 17280 2556 17332
rect 4252 17280 4304 17332
rect 4988 17280 5040 17332
rect 6092 17280 6144 17332
rect 7104 17280 7156 17332
rect 7748 17280 7800 17332
rect 8208 17280 8260 17332
rect 1676 17144 1728 17196
rect 2688 17144 2740 17196
rect 9404 17280 9456 17332
rect 16304 17323 16356 17332
rect 16304 17289 16313 17323
rect 16313 17289 16347 17323
rect 16347 17289 16356 17323
rect 16304 17280 16356 17289
rect 17040 17323 17092 17332
rect 17040 17289 17049 17323
rect 17049 17289 17083 17323
rect 17083 17289 17092 17323
rect 17040 17280 17092 17289
rect 18144 17280 18196 17332
rect 9128 17255 9180 17264
rect 3884 17144 3936 17196
rect 4436 17144 4488 17196
rect 6368 17144 6420 17196
rect 6736 17144 6788 17196
rect 9128 17221 9137 17255
rect 9137 17221 9171 17255
rect 9171 17221 9180 17255
rect 9128 17212 9180 17221
rect 7656 17187 7708 17196
rect 3424 17076 3476 17128
rect 3700 17076 3752 17128
rect 7656 17153 7665 17187
rect 7665 17153 7699 17187
rect 7699 17153 7708 17187
rect 7656 17144 7708 17153
rect 10600 17212 10652 17264
rect 10784 17212 10836 17264
rect 11428 17212 11480 17264
rect 12164 17144 12216 17196
rect 16672 17212 16724 17264
rect 18052 17212 18104 17264
rect 18420 17280 18472 17332
rect 19432 17323 19484 17332
rect 19432 17289 19441 17323
rect 19441 17289 19475 17323
rect 19475 17289 19484 17323
rect 19432 17280 19484 17289
rect 20536 17280 20588 17332
rect 20628 17280 20680 17332
rect 25136 17323 25188 17332
rect 25136 17289 25145 17323
rect 25145 17289 25179 17323
rect 25179 17289 25188 17323
rect 25136 17280 25188 17289
rect 19064 17212 19116 17264
rect 10600 17119 10652 17128
rect 2412 17008 2464 17060
rect 4252 17008 4304 17060
rect 10600 17085 10609 17119
rect 10609 17085 10643 17119
rect 10643 17085 10652 17119
rect 10600 17076 10652 17085
rect 7656 17008 7708 17060
rect 8576 17008 8628 17060
rect 5540 16940 5592 16992
rect 8208 16940 8260 16992
rect 10140 16940 10192 16992
rect 12348 17008 12400 17060
rect 11060 16940 11112 16992
rect 11888 16983 11940 16992
rect 11888 16949 11897 16983
rect 11897 16949 11931 16983
rect 11931 16949 11940 16983
rect 11888 16940 11940 16949
rect 12808 16940 12860 16992
rect 13544 16940 13596 16992
rect 17316 17144 17368 17196
rect 14740 17119 14792 17128
rect 14740 17085 14749 17119
rect 14749 17085 14783 17119
rect 14783 17085 14792 17119
rect 14740 17076 14792 17085
rect 16764 17076 16816 17128
rect 14556 17008 14608 17060
rect 16028 17051 16080 17060
rect 16028 17017 16037 17051
rect 16037 17017 16071 17051
rect 16071 17017 16080 17051
rect 16028 17008 16080 17017
rect 18052 17008 18104 17060
rect 18512 17051 18564 17060
rect 18512 17017 18521 17051
rect 18521 17017 18555 17051
rect 18555 17017 18564 17051
rect 18512 17008 18564 17017
rect 21364 17119 21416 17128
rect 21364 17085 21373 17119
rect 21373 17085 21407 17119
rect 21407 17085 21416 17119
rect 21364 17076 21416 17085
rect 25136 17076 25188 17128
rect 14096 16983 14148 16992
rect 14096 16949 14105 16983
rect 14105 16949 14139 16983
rect 14139 16949 14148 16983
rect 14096 16940 14148 16949
rect 15844 16940 15896 16992
rect 16856 16940 16908 16992
rect 20352 16983 20404 16992
rect 20352 16949 20361 16983
rect 20361 16949 20395 16983
rect 20395 16949 20404 16983
rect 20352 16940 20404 16949
rect 22652 16940 22704 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1400 16736 1452 16788
rect 3424 16779 3476 16788
rect 3424 16745 3433 16779
rect 3433 16745 3467 16779
rect 3467 16745 3476 16779
rect 3424 16736 3476 16745
rect 5172 16736 5224 16788
rect 6736 16736 6788 16788
rect 7472 16779 7524 16788
rect 7472 16745 7481 16779
rect 7481 16745 7515 16779
rect 7515 16745 7524 16779
rect 7472 16736 7524 16745
rect 11060 16779 11112 16788
rect 11060 16745 11069 16779
rect 11069 16745 11103 16779
rect 11103 16745 11112 16779
rect 11060 16736 11112 16745
rect 12808 16779 12860 16788
rect 12808 16745 12817 16779
rect 12817 16745 12851 16779
rect 12851 16745 12860 16779
rect 12808 16736 12860 16745
rect 16764 16779 16816 16788
rect 2412 16711 2464 16720
rect 2412 16677 2421 16711
rect 2421 16677 2455 16711
rect 2455 16677 2464 16711
rect 2412 16668 2464 16677
rect 2228 16600 2280 16652
rect 2780 16668 2832 16720
rect 3884 16668 3936 16720
rect 11704 16668 11756 16720
rect 12348 16668 12400 16720
rect 14740 16711 14792 16720
rect 14740 16677 14749 16711
rect 14749 16677 14783 16711
rect 14783 16677 14792 16711
rect 14740 16668 14792 16677
rect 15844 16668 15896 16720
rect 16764 16745 16773 16779
rect 16773 16745 16807 16779
rect 16807 16745 16816 16779
rect 16764 16736 16816 16745
rect 18512 16736 18564 16788
rect 18972 16779 19024 16788
rect 18972 16745 18981 16779
rect 18981 16745 19015 16779
rect 19015 16745 19024 16779
rect 18972 16736 19024 16745
rect 24768 16779 24820 16788
rect 24768 16745 24777 16779
rect 24777 16745 24811 16779
rect 24811 16745 24820 16779
rect 24768 16736 24820 16745
rect 18144 16668 18196 16720
rect 4436 16600 4488 16652
rect 5172 16643 5224 16652
rect 5172 16609 5181 16643
rect 5181 16609 5215 16643
rect 5215 16609 5224 16643
rect 5172 16600 5224 16609
rect 5448 16643 5500 16652
rect 5448 16609 5457 16643
rect 5457 16609 5491 16643
rect 5491 16609 5500 16643
rect 5448 16600 5500 16609
rect 6184 16600 6236 16652
rect 7932 16643 7984 16652
rect 7932 16609 7941 16643
rect 7941 16609 7975 16643
rect 7975 16609 7984 16643
rect 7932 16600 7984 16609
rect 13636 16643 13688 16652
rect 13636 16609 13645 16643
rect 13645 16609 13679 16643
rect 13679 16609 13688 16643
rect 13636 16600 13688 16609
rect 17316 16643 17368 16652
rect 3516 16532 3568 16584
rect 6092 16575 6144 16584
rect 6092 16541 6101 16575
rect 6101 16541 6135 16575
rect 6135 16541 6144 16575
rect 6092 16532 6144 16541
rect 9772 16532 9824 16584
rect 2688 16507 2740 16516
rect 2688 16473 2697 16507
rect 2697 16473 2731 16507
rect 2731 16473 2740 16507
rect 2688 16464 2740 16473
rect 2412 16396 2464 16448
rect 3056 16439 3108 16448
rect 3056 16405 3065 16439
rect 3065 16405 3099 16439
rect 3099 16405 3108 16439
rect 3056 16396 3108 16405
rect 8300 16439 8352 16448
rect 8300 16405 8309 16439
rect 8309 16405 8343 16439
rect 8343 16405 8352 16439
rect 8300 16396 8352 16405
rect 8484 16396 8536 16448
rect 14096 16464 14148 16516
rect 17316 16609 17325 16643
rect 17325 16609 17359 16643
rect 17359 16609 17368 16643
rect 17316 16600 17368 16609
rect 17868 16643 17920 16652
rect 17868 16609 17877 16643
rect 17877 16609 17911 16643
rect 17911 16609 17920 16643
rect 17868 16600 17920 16609
rect 18880 16643 18932 16652
rect 18880 16609 18889 16643
rect 18889 16609 18923 16643
rect 18923 16609 18932 16643
rect 18880 16600 18932 16609
rect 15660 16532 15712 16584
rect 19708 16600 19760 16652
rect 21272 16600 21324 16652
rect 21824 16600 21876 16652
rect 24676 16600 24728 16652
rect 12532 16396 12584 16448
rect 17868 16396 17920 16448
rect 19708 16396 19760 16448
rect 21916 16396 21968 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2688 16192 2740 16244
rect 3240 16192 3292 16244
rect 3516 16235 3568 16244
rect 3516 16201 3525 16235
rect 3525 16201 3559 16235
rect 3559 16201 3568 16235
rect 3516 16192 3568 16201
rect 4436 16192 4488 16244
rect 7932 16192 7984 16244
rect 8300 16192 8352 16244
rect 4252 16124 4304 16176
rect 1952 16031 2004 16040
rect 1952 15997 1961 16031
rect 1961 15997 1995 16031
rect 1995 15997 2004 16031
rect 1952 15988 2004 15997
rect 5540 16056 5592 16108
rect 6092 16056 6144 16108
rect 7288 16056 7340 16108
rect 7748 16056 7800 16108
rect 11704 16192 11756 16244
rect 14096 16235 14148 16244
rect 14096 16201 14105 16235
rect 14105 16201 14139 16235
rect 14139 16201 14148 16235
rect 14096 16192 14148 16201
rect 15844 16235 15896 16244
rect 15844 16201 15853 16235
rect 15853 16201 15887 16235
rect 15887 16201 15896 16235
rect 15844 16192 15896 16201
rect 17776 16192 17828 16244
rect 18052 16192 18104 16244
rect 18880 16192 18932 16244
rect 19708 16235 19760 16244
rect 19708 16201 19717 16235
rect 19717 16201 19751 16235
rect 19751 16201 19760 16235
rect 19708 16192 19760 16201
rect 21824 16192 21876 16244
rect 23664 16192 23716 16244
rect 24676 16235 24728 16244
rect 24676 16201 24685 16235
rect 24685 16201 24719 16235
rect 24719 16201 24728 16235
rect 24676 16192 24728 16201
rect 2412 16031 2464 16040
rect 2412 15997 2421 16031
rect 2421 15997 2455 16031
rect 2455 15997 2464 16031
rect 2872 16031 2924 16040
rect 2412 15988 2464 15997
rect 2872 15997 2881 16031
rect 2881 15997 2915 16031
rect 2915 15997 2924 16031
rect 2872 15988 2924 15997
rect 3516 15988 3568 16040
rect 4436 16031 4488 16040
rect 4436 15997 4445 16031
rect 4445 15997 4479 16031
rect 4479 15997 4488 16031
rect 4436 15988 4488 15997
rect 5172 16031 5224 16040
rect 5172 15997 5181 16031
rect 5181 15997 5215 16031
rect 5215 15997 5224 16031
rect 5172 15988 5224 15997
rect 5448 16031 5500 16040
rect 5448 15997 5457 16031
rect 5457 15997 5491 16031
rect 5491 15997 5500 16031
rect 5448 15988 5500 15997
rect 6000 15988 6052 16040
rect 13544 16124 13596 16176
rect 15660 16124 15712 16176
rect 15752 16124 15804 16176
rect 11336 16099 11388 16108
rect 11336 16065 11345 16099
rect 11345 16065 11379 16099
rect 11379 16065 11388 16099
rect 11336 16056 11388 16065
rect 10876 15988 10928 16040
rect 12624 16031 12676 16040
rect 12624 15997 12633 16031
rect 12633 15997 12667 16031
rect 12667 15997 12676 16031
rect 12624 15988 12676 15997
rect 15016 16056 15068 16108
rect 15568 16056 15620 16108
rect 20444 16056 20496 16108
rect 20628 16099 20680 16108
rect 20628 16065 20637 16099
rect 20637 16065 20671 16099
rect 20671 16065 20680 16099
rect 20628 16056 20680 16065
rect 12992 15988 13044 16040
rect 15936 15988 15988 16040
rect 6092 15920 6144 15972
rect 6644 15963 6696 15972
rect 6644 15929 6653 15963
rect 6653 15929 6687 15963
rect 6687 15929 6696 15963
rect 6644 15920 6696 15929
rect 7748 15920 7800 15972
rect 8484 15920 8536 15972
rect 9312 15963 9364 15972
rect 2320 15852 2372 15904
rect 3884 15852 3936 15904
rect 6000 15852 6052 15904
rect 6184 15895 6236 15904
rect 6184 15861 6193 15895
rect 6193 15861 6227 15895
rect 6227 15861 6236 15895
rect 6184 15852 6236 15861
rect 8300 15852 8352 15904
rect 9312 15929 9321 15963
rect 9321 15929 9355 15963
rect 9355 15929 9364 15963
rect 9312 15920 9364 15929
rect 13636 15963 13688 15972
rect 13636 15929 13645 15963
rect 13645 15929 13679 15963
rect 13679 15929 13688 15963
rect 13636 15920 13688 15929
rect 9772 15895 9824 15904
rect 9772 15861 9781 15895
rect 9781 15861 9815 15895
rect 9815 15861 9824 15895
rect 9772 15852 9824 15861
rect 12532 15895 12584 15904
rect 12532 15861 12541 15895
rect 12541 15861 12575 15895
rect 12575 15861 12584 15895
rect 12532 15852 12584 15861
rect 14832 15852 14884 15904
rect 15016 15963 15068 15972
rect 15016 15929 15025 15963
rect 15025 15929 15059 15963
rect 15059 15929 15068 15963
rect 16488 15988 16540 16040
rect 17868 15988 17920 16040
rect 21732 15988 21784 16040
rect 24124 16031 24176 16040
rect 24124 15997 24133 16031
rect 24133 15997 24167 16031
rect 24167 15997 24176 16031
rect 24124 15988 24176 15997
rect 15016 15920 15068 15929
rect 16764 15920 16816 15972
rect 17132 15963 17184 15972
rect 17132 15929 17141 15963
rect 17141 15929 17175 15963
rect 17175 15929 17184 15963
rect 17132 15920 17184 15929
rect 18144 15920 18196 15972
rect 18880 15852 18932 15904
rect 21364 15920 21416 15972
rect 21272 15895 21324 15904
rect 21272 15861 21281 15895
rect 21281 15861 21315 15895
rect 21315 15861 21324 15895
rect 21272 15852 21324 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2780 15648 2832 15700
rect 1952 15580 2004 15632
rect 2320 15555 2372 15564
rect 2320 15521 2329 15555
rect 2329 15521 2363 15555
rect 2363 15521 2372 15555
rect 3700 15648 3752 15700
rect 5448 15691 5500 15700
rect 5448 15657 5457 15691
rect 5457 15657 5491 15691
rect 5491 15657 5500 15691
rect 5448 15648 5500 15657
rect 7288 15691 7340 15700
rect 7288 15657 7297 15691
rect 7297 15657 7331 15691
rect 7331 15657 7340 15691
rect 7288 15648 7340 15657
rect 7932 15691 7984 15700
rect 7932 15657 7941 15691
rect 7941 15657 7975 15691
rect 7975 15657 7984 15691
rect 9772 15691 9824 15700
rect 7932 15648 7984 15657
rect 5172 15580 5224 15632
rect 5356 15580 5408 15632
rect 6644 15580 6696 15632
rect 9772 15657 9781 15691
rect 9781 15657 9815 15691
rect 9815 15657 9824 15691
rect 9772 15648 9824 15657
rect 10784 15691 10836 15700
rect 10784 15657 10793 15691
rect 10793 15657 10827 15691
rect 10827 15657 10836 15691
rect 10784 15648 10836 15657
rect 11704 15691 11756 15700
rect 11704 15657 11713 15691
rect 11713 15657 11747 15691
rect 11747 15657 11756 15691
rect 11704 15648 11756 15657
rect 11888 15648 11940 15700
rect 12992 15691 13044 15700
rect 12992 15657 13001 15691
rect 13001 15657 13035 15691
rect 13035 15657 13044 15691
rect 12992 15648 13044 15657
rect 17316 15648 17368 15700
rect 17684 15648 17736 15700
rect 20076 15648 20128 15700
rect 20444 15648 20496 15700
rect 21916 15691 21968 15700
rect 21916 15657 21925 15691
rect 21925 15657 21959 15691
rect 21959 15657 21968 15691
rect 21916 15648 21968 15657
rect 24768 15691 24820 15700
rect 24768 15657 24777 15691
rect 24777 15657 24811 15691
rect 24811 15657 24820 15691
rect 24768 15648 24820 15657
rect 9312 15580 9364 15632
rect 2320 15512 2372 15521
rect 4252 15512 4304 15564
rect 10692 15580 10744 15632
rect 10048 15512 10100 15564
rect 14188 15580 14240 15632
rect 15384 15580 15436 15632
rect 18144 15580 18196 15632
rect 21088 15623 21140 15632
rect 21088 15589 21097 15623
rect 21097 15589 21131 15623
rect 21131 15589 21140 15623
rect 21088 15580 21140 15589
rect 21180 15580 21232 15632
rect 16856 15555 16908 15564
rect 16856 15521 16865 15555
rect 16865 15521 16899 15555
rect 16899 15521 16908 15555
rect 16856 15512 16908 15521
rect 17132 15512 17184 15564
rect 17776 15512 17828 15564
rect 20168 15512 20220 15564
rect 23664 15512 23716 15564
rect 24216 15512 24268 15564
rect 24676 15512 24728 15564
rect 3148 15444 3200 15496
rect 3240 15444 3292 15496
rect 4896 15444 4948 15496
rect 6092 15487 6144 15496
rect 6092 15453 6101 15487
rect 6101 15453 6135 15487
rect 6135 15453 6144 15487
rect 6092 15444 6144 15453
rect 8116 15487 8168 15496
rect 8116 15453 8125 15487
rect 8125 15453 8159 15487
rect 8159 15453 8168 15487
rect 8116 15444 8168 15453
rect 11336 15487 11388 15496
rect 11336 15453 11345 15487
rect 11345 15453 11379 15487
rect 11379 15453 11388 15487
rect 11336 15444 11388 15453
rect 12256 15444 12308 15496
rect 13176 15444 13228 15496
rect 13912 15444 13964 15496
rect 15384 15487 15436 15496
rect 15384 15453 15393 15487
rect 15393 15453 15427 15487
rect 15427 15453 15436 15487
rect 15384 15444 15436 15453
rect 2136 15419 2188 15428
rect 2136 15385 2145 15419
rect 2145 15385 2179 15419
rect 2179 15385 2188 15419
rect 2136 15376 2188 15385
rect 15844 15376 15896 15428
rect 19064 15376 19116 15428
rect 22008 15444 22060 15496
rect 22652 15376 22704 15428
rect 5080 15351 5132 15360
rect 5080 15317 5089 15351
rect 5089 15317 5123 15351
rect 5123 15317 5132 15351
rect 5080 15308 5132 15317
rect 7012 15351 7064 15360
rect 7012 15317 7021 15351
rect 7021 15317 7055 15351
rect 7055 15317 7064 15351
rect 7012 15308 7064 15317
rect 11152 15351 11204 15360
rect 11152 15317 11161 15351
rect 11161 15317 11195 15351
rect 11195 15317 11204 15351
rect 11152 15308 11204 15317
rect 12624 15351 12676 15360
rect 12624 15317 12633 15351
rect 12633 15317 12667 15351
rect 12667 15317 12676 15351
rect 12624 15308 12676 15317
rect 13728 15308 13780 15360
rect 14832 15351 14884 15360
rect 14832 15317 14841 15351
rect 14841 15317 14875 15351
rect 14875 15317 14884 15351
rect 14832 15308 14884 15317
rect 16488 15351 16540 15360
rect 16488 15317 16497 15351
rect 16497 15317 16531 15351
rect 16531 15317 16540 15351
rect 16488 15308 16540 15317
rect 18512 15308 18564 15360
rect 20168 15308 20220 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2780 15104 2832 15156
rect 3240 15104 3292 15156
rect 5080 15104 5132 15156
rect 5356 15147 5408 15156
rect 5356 15113 5365 15147
rect 5365 15113 5399 15147
rect 5399 15113 5408 15147
rect 5356 15104 5408 15113
rect 7932 15104 7984 15156
rect 10048 15147 10100 15156
rect 10048 15113 10057 15147
rect 10057 15113 10091 15147
rect 10091 15113 10100 15147
rect 10048 15104 10100 15113
rect 10692 15104 10744 15156
rect 11336 15104 11388 15156
rect 12900 15104 12952 15156
rect 6644 15036 6696 15088
rect 6920 15036 6972 15088
rect 2136 14968 2188 15020
rect 4068 14968 4120 15020
rect 5448 15011 5500 15020
rect 5448 14977 5457 15011
rect 5457 14977 5491 15011
rect 5491 14977 5500 15011
rect 5448 14968 5500 14977
rect 7196 14968 7248 15020
rect 8116 15011 8168 15020
rect 8116 14977 8125 15011
rect 8125 14977 8159 15011
rect 8159 14977 8168 15011
rect 8116 14968 8168 14977
rect 11152 15036 11204 15088
rect 14188 15079 14240 15088
rect 12900 15011 12952 15020
rect 12900 14977 12909 15011
rect 12909 14977 12943 15011
rect 12943 14977 12952 15011
rect 12900 14968 12952 14977
rect 13176 15011 13228 15020
rect 13176 14977 13185 15011
rect 13185 14977 13219 15011
rect 13219 14977 13228 15011
rect 13176 14968 13228 14977
rect 14188 15045 14197 15079
rect 14197 15045 14231 15079
rect 14231 15045 14240 15079
rect 14188 15036 14240 15045
rect 15108 15036 15160 15088
rect 15568 15104 15620 15156
rect 16672 15104 16724 15156
rect 16856 15104 16908 15156
rect 17776 15147 17828 15156
rect 17776 15113 17785 15147
rect 17785 15113 17819 15147
rect 17819 15113 17828 15147
rect 17776 15104 17828 15113
rect 18144 15104 18196 15156
rect 21088 15147 21140 15156
rect 21088 15113 21097 15147
rect 21097 15113 21131 15147
rect 21131 15113 21140 15147
rect 21088 15104 21140 15113
rect 21364 15147 21416 15156
rect 21364 15113 21373 15147
rect 21373 15113 21407 15147
rect 21407 15113 21416 15147
rect 21364 15104 21416 15113
rect 22652 15147 22704 15156
rect 22652 15113 22661 15147
rect 22661 15113 22695 15147
rect 22695 15113 22704 15147
rect 22652 15104 22704 15113
rect 24676 15147 24728 15156
rect 24676 15113 24685 15147
rect 24685 15113 24719 15147
rect 24719 15113 24728 15147
rect 24676 15104 24728 15113
rect 24952 15147 25004 15156
rect 24952 15113 24961 15147
rect 24961 15113 24995 15147
rect 24995 15113 25004 15147
rect 24952 15104 25004 15113
rect 15752 15036 15804 15088
rect 20628 15079 20680 15088
rect 20628 15045 20637 15079
rect 20637 15045 20671 15079
rect 20671 15045 20680 15079
rect 20628 15036 20680 15045
rect 15568 14968 15620 15020
rect 15660 14968 15712 15020
rect 18512 15011 18564 15020
rect 18512 14977 18521 15011
rect 18521 14977 18555 15011
rect 18555 14977 18564 15011
rect 18512 14968 18564 14977
rect 18604 14968 18656 15020
rect 664 14900 716 14952
rect 2412 14900 2464 14952
rect 3056 14900 3108 14952
rect 3516 14943 3568 14952
rect 3516 14909 3525 14943
rect 3525 14909 3559 14943
rect 3559 14909 3568 14943
rect 3516 14900 3568 14909
rect 4252 14900 4304 14952
rect 4988 14900 5040 14952
rect 2320 14832 2372 14884
rect 7472 14832 7524 14884
rect 14924 14900 14976 14952
rect 16672 14900 16724 14952
rect 2872 14764 2924 14816
rect 7012 14764 7064 14816
rect 8576 14832 8628 14884
rect 11244 14832 11296 14884
rect 11520 14875 11572 14884
rect 11520 14841 11529 14875
rect 11529 14841 11563 14875
rect 11563 14841 11572 14875
rect 11520 14832 11572 14841
rect 13176 14832 13228 14884
rect 16212 14832 16264 14884
rect 18604 14875 18656 14884
rect 18604 14841 18613 14875
rect 18613 14841 18647 14875
rect 18647 14841 18656 14875
rect 18604 14832 18656 14841
rect 19156 14875 19208 14884
rect 19156 14841 19165 14875
rect 19165 14841 19199 14875
rect 19199 14841 19208 14875
rect 19156 14832 19208 14841
rect 21180 14968 21232 15020
rect 21916 14968 21968 15020
rect 22008 15011 22060 15020
rect 22008 14977 22017 15011
rect 22017 14977 22051 15011
rect 22051 14977 22060 15011
rect 22008 14968 22060 14977
rect 24952 14900 25004 14952
rect 20076 14832 20128 14884
rect 21088 14832 21140 14884
rect 21364 14832 21416 14884
rect 11980 14764 12032 14816
rect 13912 14807 13964 14816
rect 13912 14773 13921 14807
rect 13921 14773 13955 14807
rect 13955 14773 13964 14807
rect 13912 14764 13964 14773
rect 14924 14807 14976 14816
rect 14924 14773 14933 14807
rect 14933 14773 14967 14807
rect 14967 14773 14976 14807
rect 14924 14764 14976 14773
rect 15292 14807 15344 14816
rect 15292 14773 15301 14807
rect 15301 14773 15335 14807
rect 15335 14773 15344 14807
rect 15292 14764 15344 14773
rect 19524 14807 19576 14816
rect 19524 14773 19533 14807
rect 19533 14773 19567 14807
rect 19567 14773 19576 14807
rect 19524 14764 19576 14773
rect 21640 14764 21692 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1492 14560 1544 14612
rect 3056 14603 3108 14612
rect 3056 14569 3065 14603
rect 3065 14569 3099 14603
rect 3099 14569 3108 14603
rect 3056 14560 3108 14569
rect 4436 14560 4488 14612
rect 4988 14560 5040 14612
rect 6092 14560 6144 14612
rect 7196 14560 7248 14612
rect 572 14492 624 14544
rect 1952 14492 2004 14544
rect 2044 14467 2096 14476
rect 2044 14433 2053 14467
rect 2053 14433 2087 14467
rect 2087 14433 2096 14467
rect 2044 14424 2096 14433
rect 4068 14492 4120 14544
rect 4252 14467 4304 14476
rect 4252 14433 4261 14467
rect 4261 14433 4295 14467
rect 4295 14433 4304 14467
rect 4252 14424 4304 14433
rect 5172 14424 5224 14476
rect 5448 14424 5500 14476
rect 8576 14492 8628 14544
rect 6184 14424 6236 14476
rect 10232 14424 10284 14476
rect 10692 14560 10744 14612
rect 11980 14560 12032 14612
rect 13452 14560 13504 14612
rect 12900 14535 12952 14544
rect 12900 14501 12909 14535
rect 12909 14501 12943 14535
rect 12943 14501 12952 14535
rect 12900 14492 12952 14501
rect 15384 14560 15436 14612
rect 18604 14603 18656 14612
rect 15108 14535 15160 14544
rect 15108 14501 15117 14535
rect 15117 14501 15151 14535
rect 15151 14501 15160 14535
rect 15108 14492 15160 14501
rect 15292 14492 15344 14544
rect 16028 14492 16080 14544
rect 17868 14535 17920 14544
rect 17868 14501 17877 14535
rect 17877 14501 17911 14535
rect 17911 14501 17920 14535
rect 17868 14492 17920 14501
rect 10692 14467 10744 14476
rect 10692 14433 10701 14467
rect 10701 14433 10735 14467
rect 10735 14433 10744 14467
rect 10692 14424 10744 14433
rect 16396 14424 16448 14476
rect 16580 14424 16632 14476
rect 17132 14467 17184 14476
rect 17132 14433 17141 14467
rect 17141 14433 17175 14467
rect 17175 14433 17184 14467
rect 17132 14424 17184 14433
rect 1400 14356 1452 14408
rect 5540 14356 5592 14408
rect 8116 14399 8168 14408
rect 2136 14331 2188 14340
rect 2136 14297 2145 14331
rect 2145 14297 2179 14331
rect 2179 14297 2188 14331
rect 2136 14288 2188 14297
rect 4252 14220 4304 14272
rect 8116 14365 8125 14399
rect 8125 14365 8159 14399
rect 8159 14365 8168 14399
rect 8116 14356 8168 14365
rect 12256 14356 12308 14408
rect 13636 14356 13688 14408
rect 15568 14399 15620 14408
rect 12532 14288 12584 14340
rect 8116 14220 8168 14272
rect 11244 14263 11296 14272
rect 11244 14229 11253 14263
rect 11253 14229 11287 14263
rect 11287 14229 11296 14263
rect 11244 14220 11296 14229
rect 13268 14220 13320 14272
rect 15568 14365 15577 14399
rect 15577 14365 15611 14399
rect 15611 14365 15620 14399
rect 15568 14356 15620 14365
rect 16120 14288 16172 14340
rect 18604 14569 18613 14603
rect 18613 14569 18647 14603
rect 18647 14569 18656 14603
rect 18604 14560 18656 14569
rect 19524 14560 19576 14612
rect 25412 14560 25464 14612
rect 18880 14535 18932 14544
rect 18880 14501 18889 14535
rect 18889 14501 18923 14535
rect 18923 14501 18932 14535
rect 20076 14535 20128 14544
rect 18880 14492 18932 14501
rect 20076 14501 20085 14535
rect 20085 14501 20119 14535
rect 20119 14501 20128 14535
rect 20076 14492 20128 14501
rect 20168 14492 20220 14544
rect 20260 14424 20312 14476
rect 20996 14467 21048 14476
rect 20996 14433 21014 14467
rect 21014 14433 21048 14467
rect 20996 14424 21048 14433
rect 21732 14424 21784 14476
rect 22100 14424 22152 14476
rect 22928 14467 22980 14476
rect 22928 14433 22937 14467
rect 22937 14433 22971 14467
rect 22971 14433 22980 14467
rect 22928 14424 22980 14433
rect 24124 14424 24176 14476
rect 19156 14399 19208 14408
rect 19156 14365 19165 14399
rect 19165 14365 19199 14399
rect 19199 14365 19208 14399
rect 19156 14356 19208 14365
rect 18420 14220 18472 14272
rect 18512 14220 18564 14272
rect 19340 14220 19392 14272
rect 21548 14220 21600 14272
rect 21732 14263 21784 14272
rect 21732 14229 21741 14263
rect 21741 14229 21775 14263
rect 21775 14229 21784 14263
rect 21732 14220 21784 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 1952 14016 2004 14068
rect 2320 14016 2372 14068
rect 2964 14016 3016 14068
rect 5172 14059 5224 14068
rect 5172 14025 5181 14059
rect 5181 14025 5215 14059
rect 5215 14025 5224 14059
rect 5172 14016 5224 14025
rect 6184 14059 6236 14068
rect 6184 14025 6193 14059
rect 6193 14025 6227 14059
rect 6227 14025 6236 14059
rect 6184 14016 6236 14025
rect 8576 14059 8628 14068
rect 8576 14025 8585 14059
rect 8585 14025 8619 14059
rect 8619 14025 8628 14059
rect 8576 14016 8628 14025
rect 9312 14016 9364 14068
rect 10232 14016 10284 14068
rect 11244 14016 11296 14068
rect 13452 14059 13504 14068
rect 2136 13948 2188 14000
rect 2688 13991 2740 14000
rect 2688 13957 2697 13991
rect 2697 13957 2731 13991
rect 2731 13957 2740 13991
rect 2688 13948 2740 13957
rect 3700 13948 3752 14000
rect 9036 13948 9088 14000
rect 11980 13948 12032 14000
rect 13452 14025 13461 14059
rect 13461 14025 13495 14059
rect 13495 14025 13504 14059
rect 13452 14016 13504 14025
rect 13728 14016 13780 14068
rect 17132 14059 17184 14068
rect 17132 14025 17141 14059
rect 17141 14025 17175 14059
rect 17175 14025 17184 14059
rect 17132 14016 17184 14025
rect 14188 13948 14240 14000
rect 15292 13948 15344 14000
rect 15752 13991 15804 14000
rect 15752 13957 15761 13991
rect 15761 13957 15795 13991
rect 15795 13957 15804 13991
rect 15752 13948 15804 13957
rect 1952 13880 2004 13932
rect 1492 13812 1544 13864
rect 2596 13855 2648 13864
rect 2596 13821 2605 13855
rect 2605 13821 2639 13855
rect 2639 13821 2648 13855
rect 2596 13812 2648 13821
rect 2964 13812 3016 13864
rect 4068 13812 4120 13864
rect 4436 13855 4488 13864
rect 4436 13821 4445 13855
rect 4445 13821 4479 13855
rect 4479 13821 4488 13855
rect 4436 13812 4488 13821
rect 5448 13812 5500 13864
rect 7932 13855 7984 13864
rect 3056 13744 3108 13796
rect 2688 13676 2740 13728
rect 4436 13676 4488 13728
rect 4620 13719 4672 13728
rect 4620 13685 4629 13719
rect 4629 13685 4663 13719
rect 4663 13685 4672 13719
rect 4620 13676 4672 13685
rect 7932 13821 7941 13855
rect 7941 13821 7975 13855
rect 7975 13821 7984 13855
rect 7932 13812 7984 13821
rect 10784 13880 10836 13932
rect 11520 13880 11572 13932
rect 12532 13923 12584 13932
rect 12532 13889 12541 13923
rect 12541 13889 12575 13923
rect 12575 13889 12584 13923
rect 12532 13880 12584 13889
rect 13268 13880 13320 13932
rect 13912 13880 13964 13932
rect 18788 14016 18840 14068
rect 18880 14016 18932 14068
rect 20996 14059 21048 14068
rect 20996 14025 21005 14059
rect 21005 14025 21039 14059
rect 21039 14025 21048 14059
rect 20996 14016 21048 14025
rect 21548 13948 21600 14000
rect 8208 13787 8260 13796
rect 8208 13753 8217 13787
rect 8217 13753 8251 13787
rect 8251 13753 8260 13787
rect 8208 13744 8260 13753
rect 8300 13744 8352 13796
rect 8576 13744 8628 13796
rect 14004 13855 14056 13864
rect 14004 13821 14013 13855
rect 14013 13821 14047 13855
rect 14047 13821 14056 13855
rect 14004 13812 14056 13821
rect 18052 13855 18104 13864
rect 18052 13821 18061 13855
rect 18061 13821 18095 13855
rect 18095 13821 18104 13855
rect 18052 13812 18104 13821
rect 18420 13812 18472 13864
rect 20812 13880 20864 13932
rect 22928 13923 22980 13932
rect 22928 13889 22937 13923
rect 22937 13889 22971 13923
rect 22971 13889 22980 13923
rect 22928 13880 22980 13889
rect 11980 13744 12032 13796
rect 9128 13676 9180 13728
rect 11888 13676 11940 13728
rect 12716 13676 12768 13728
rect 15292 13787 15344 13796
rect 15292 13753 15301 13787
rect 15301 13753 15335 13787
rect 15335 13753 15344 13787
rect 15292 13744 15344 13753
rect 19156 13744 19208 13796
rect 15384 13676 15436 13728
rect 16028 13676 16080 13728
rect 16304 13676 16356 13728
rect 16488 13719 16540 13728
rect 16488 13685 16497 13719
rect 16497 13685 16531 13719
rect 16531 13685 16540 13719
rect 16488 13676 16540 13685
rect 18144 13719 18196 13728
rect 18144 13685 18153 13719
rect 18153 13685 18187 13719
rect 18187 13685 18196 13719
rect 18144 13676 18196 13685
rect 19432 13719 19484 13728
rect 19432 13685 19441 13719
rect 19441 13685 19475 13719
rect 19475 13685 19484 13719
rect 21180 13744 21232 13796
rect 21548 13812 21600 13864
rect 21732 13744 21784 13796
rect 19432 13676 19484 13685
rect 19984 13676 20036 13728
rect 22100 13676 22152 13728
rect 24124 13676 24176 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 3608 13472 3660 13524
rect 2412 13447 2464 13456
rect 2412 13413 2421 13447
rect 2421 13413 2455 13447
rect 2455 13413 2464 13447
rect 2412 13404 2464 13413
rect 3056 13404 3108 13456
rect 5540 13472 5592 13524
rect 10140 13515 10192 13524
rect 10140 13481 10149 13515
rect 10149 13481 10183 13515
rect 10183 13481 10192 13515
rect 10140 13472 10192 13481
rect 10784 13515 10836 13524
rect 10784 13481 10793 13515
rect 10793 13481 10827 13515
rect 10827 13481 10836 13515
rect 10784 13472 10836 13481
rect 11888 13515 11940 13524
rect 11888 13481 11897 13515
rect 11897 13481 11931 13515
rect 11931 13481 11940 13515
rect 11888 13472 11940 13481
rect 12256 13515 12308 13524
rect 12256 13481 12265 13515
rect 12265 13481 12299 13515
rect 12299 13481 12308 13515
rect 12256 13472 12308 13481
rect 12532 13515 12584 13524
rect 12532 13481 12541 13515
rect 12541 13481 12575 13515
rect 12575 13481 12584 13515
rect 12532 13472 12584 13481
rect 13176 13472 13228 13524
rect 15292 13472 15344 13524
rect 18236 13472 18288 13524
rect 4712 13404 4764 13456
rect 5356 13404 5408 13456
rect 6092 13404 6144 13456
rect 8300 13404 8352 13456
rect 11980 13404 12032 13456
rect 13452 13404 13504 13456
rect 14740 13404 14792 13456
rect 16028 13404 16080 13456
rect 2320 13379 2372 13388
rect 2320 13345 2329 13379
rect 2329 13345 2363 13379
rect 2363 13345 2372 13379
rect 2320 13336 2372 13345
rect 4160 13336 4212 13388
rect 2228 13268 2280 13320
rect 2044 13200 2096 13252
rect 4068 13200 4120 13252
rect 6000 13336 6052 13388
rect 9864 13336 9916 13388
rect 5540 13311 5592 13320
rect 5540 13277 5549 13311
rect 5549 13277 5583 13311
rect 5583 13277 5592 13311
rect 5540 13268 5592 13277
rect 7840 13311 7892 13320
rect 7840 13277 7849 13311
rect 7849 13277 7883 13311
rect 7883 13277 7892 13311
rect 7840 13268 7892 13277
rect 9036 13268 9088 13320
rect 10784 13336 10836 13388
rect 14924 13336 14976 13388
rect 17132 13336 17184 13388
rect 18052 13404 18104 13456
rect 18696 13404 18748 13456
rect 20628 13404 20680 13456
rect 21272 13404 21324 13456
rect 21456 13404 21508 13456
rect 22100 13404 22152 13456
rect 17500 13379 17552 13388
rect 17500 13345 17509 13379
rect 17509 13345 17543 13379
rect 17543 13345 17552 13379
rect 17500 13336 17552 13345
rect 19524 13336 19576 13388
rect 19984 13336 20036 13388
rect 10968 13311 11020 13320
rect 10968 13277 10977 13311
rect 10977 13277 11011 13311
rect 11011 13277 11020 13311
rect 10968 13268 11020 13277
rect 12716 13311 12768 13320
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 15384 13268 15436 13320
rect 11704 13200 11756 13252
rect 15752 13268 15804 13320
rect 18420 13268 18472 13320
rect 19340 13268 19392 13320
rect 21180 13268 21232 13320
rect 2136 13132 2188 13184
rect 2688 13175 2740 13184
rect 2688 13141 2697 13175
rect 2697 13141 2731 13175
rect 2731 13141 2740 13175
rect 2688 13132 2740 13141
rect 2872 13132 2924 13184
rect 3792 13132 3844 13184
rect 6368 13132 6420 13184
rect 7012 13132 7064 13184
rect 7104 13132 7156 13184
rect 7932 13132 7984 13184
rect 10416 13175 10468 13184
rect 10416 13141 10425 13175
rect 10425 13141 10459 13175
rect 10459 13141 10468 13175
rect 10416 13132 10468 13141
rect 10692 13132 10744 13184
rect 13912 13175 13964 13184
rect 13912 13141 13921 13175
rect 13921 13141 13955 13175
rect 13955 13141 13964 13175
rect 13912 13132 13964 13141
rect 15936 13200 15988 13252
rect 16396 13132 16448 13184
rect 19156 13132 19208 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1124 12928 1176 12980
rect 2320 12928 2372 12980
rect 2688 12971 2740 12980
rect 2688 12937 2697 12971
rect 2697 12937 2731 12971
rect 2731 12937 2740 12971
rect 2688 12928 2740 12937
rect 3148 12928 3200 12980
rect 6092 12928 6144 12980
rect 6644 12928 6696 12980
rect 8300 12928 8352 12980
rect 14004 12928 14056 12980
rect 14740 12928 14792 12980
rect 17132 12971 17184 12980
rect 17132 12937 17141 12971
rect 17141 12937 17175 12971
rect 17175 12937 17184 12971
rect 17132 12928 17184 12937
rect 19432 12928 19484 12980
rect 21272 12971 21324 12980
rect 21272 12937 21281 12971
rect 21281 12937 21315 12971
rect 21315 12937 21324 12971
rect 21272 12928 21324 12937
rect 5080 12860 5132 12912
rect 5356 12860 5408 12912
rect 2504 12792 2556 12844
rect 6368 12792 6420 12844
rect 8208 12792 8260 12844
rect 9036 12792 9088 12844
rect 11980 12860 12032 12912
rect 13544 12860 13596 12912
rect 16120 12903 16172 12912
rect 2596 12724 2648 12776
rect 3148 12767 3200 12776
rect 3148 12733 3157 12767
rect 3157 12733 3191 12767
rect 3191 12733 3200 12767
rect 3148 12724 3200 12733
rect 2964 12656 3016 12708
rect 3424 12588 3476 12640
rect 3608 12588 3660 12640
rect 4160 12588 4212 12640
rect 4436 12588 4488 12640
rect 9128 12724 9180 12776
rect 9772 12724 9824 12776
rect 10416 12724 10468 12776
rect 10968 12792 11020 12844
rect 16120 12869 16129 12903
rect 16129 12869 16163 12903
rect 16163 12869 16172 12903
rect 16120 12860 16172 12869
rect 21180 12860 21232 12912
rect 22008 12860 22060 12912
rect 18328 12767 18380 12776
rect 18328 12733 18337 12767
rect 18337 12733 18371 12767
rect 18371 12733 18380 12767
rect 18328 12724 18380 12733
rect 20076 12767 20128 12776
rect 20076 12733 20085 12767
rect 20085 12733 20119 12767
rect 20119 12733 20128 12767
rect 20076 12724 20128 12733
rect 5816 12699 5868 12708
rect 5816 12665 5825 12699
rect 5825 12665 5859 12699
rect 5859 12665 5868 12699
rect 5816 12656 5868 12665
rect 7012 12699 7064 12708
rect 7012 12665 7021 12699
rect 7021 12665 7055 12699
rect 7055 12665 7064 12699
rect 7012 12656 7064 12665
rect 8300 12656 8352 12708
rect 13912 12699 13964 12708
rect 13912 12665 13921 12699
rect 13921 12665 13955 12699
rect 13955 12665 13964 12699
rect 13912 12656 13964 12665
rect 14004 12699 14056 12708
rect 14004 12665 14013 12699
rect 14013 12665 14047 12699
rect 14047 12665 14056 12699
rect 14004 12656 14056 12665
rect 16212 12656 16264 12708
rect 4988 12631 5040 12640
rect 4988 12597 4997 12631
rect 4997 12597 5031 12631
rect 5031 12597 5040 12631
rect 4988 12588 5040 12597
rect 6092 12631 6144 12640
rect 6092 12597 6101 12631
rect 6101 12597 6135 12631
rect 6135 12597 6144 12631
rect 6092 12588 6144 12597
rect 6644 12631 6696 12640
rect 6644 12597 6653 12631
rect 6653 12597 6687 12631
rect 6687 12597 6696 12631
rect 6644 12588 6696 12597
rect 12624 12631 12676 12640
rect 12624 12597 12633 12631
rect 12633 12597 12667 12631
rect 12667 12597 12676 12631
rect 12624 12588 12676 12597
rect 13452 12588 13504 12640
rect 17500 12631 17552 12640
rect 17500 12597 17509 12631
rect 17509 12597 17543 12631
rect 17543 12597 17552 12631
rect 17500 12588 17552 12597
rect 17960 12588 18012 12640
rect 18696 12631 18748 12640
rect 18696 12597 18705 12631
rect 18705 12597 18739 12631
rect 18739 12597 18748 12631
rect 18696 12588 18748 12597
rect 21916 12699 21968 12708
rect 21916 12665 21925 12699
rect 21925 12665 21959 12699
rect 21959 12665 21968 12699
rect 21916 12656 21968 12665
rect 26424 12588 26476 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 3700 12384 3752 12436
rect 4252 12427 4304 12436
rect 4252 12393 4261 12427
rect 4261 12393 4295 12427
rect 4295 12393 4304 12427
rect 4252 12384 4304 12393
rect 4712 12427 4764 12436
rect 4712 12393 4721 12427
rect 4721 12393 4755 12427
rect 4755 12393 4764 12427
rect 4712 12384 4764 12393
rect 5080 12427 5132 12436
rect 5080 12393 5089 12427
rect 5089 12393 5123 12427
rect 5123 12393 5132 12427
rect 5080 12384 5132 12393
rect 5816 12384 5868 12436
rect 7196 12427 7248 12436
rect 7196 12393 7205 12427
rect 7205 12393 7239 12427
rect 7239 12393 7248 12427
rect 7196 12384 7248 12393
rect 7840 12427 7892 12436
rect 7840 12393 7849 12427
rect 7849 12393 7883 12427
rect 7883 12393 7892 12427
rect 7840 12384 7892 12393
rect 9036 12427 9088 12436
rect 9036 12393 9045 12427
rect 9045 12393 9079 12427
rect 9079 12393 9088 12427
rect 9036 12384 9088 12393
rect 10784 12427 10836 12436
rect 10784 12393 10793 12427
rect 10793 12393 10827 12427
rect 10827 12393 10836 12427
rect 10784 12384 10836 12393
rect 11428 12427 11480 12436
rect 11428 12393 11437 12427
rect 11437 12393 11471 12427
rect 11471 12393 11480 12427
rect 11428 12384 11480 12393
rect 16304 12384 16356 12436
rect 19524 12427 19576 12436
rect 19524 12393 19533 12427
rect 19533 12393 19567 12427
rect 19567 12393 19576 12427
rect 19524 12384 19576 12393
rect 20628 12427 20680 12436
rect 20628 12393 20637 12427
rect 20637 12393 20671 12427
rect 20671 12393 20680 12427
rect 20628 12384 20680 12393
rect 1308 12248 1360 12300
rect 3976 12316 4028 12368
rect 4620 12316 4672 12368
rect 4068 12291 4120 12300
rect 4068 12257 4077 12291
rect 4077 12257 4111 12291
rect 4111 12257 4120 12291
rect 4068 12248 4120 12257
rect 2320 12180 2372 12232
rect 2872 12180 2924 12232
rect 6276 12316 6328 12368
rect 5540 12248 5592 12300
rect 7012 12291 7064 12300
rect 7012 12257 7021 12291
rect 7021 12257 7055 12291
rect 7055 12257 7064 12291
rect 7012 12248 7064 12257
rect 2044 12044 2096 12096
rect 2964 12112 3016 12164
rect 6000 12180 6052 12232
rect 4436 12112 4488 12164
rect 8208 12248 8260 12300
rect 8392 12248 8444 12300
rect 9772 12291 9824 12300
rect 9772 12257 9781 12291
rect 9781 12257 9815 12291
rect 9815 12257 9824 12291
rect 9772 12248 9824 12257
rect 12716 12359 12768 12368
rect 12716 12325 12725 12359
rect 12725 12325 12759 12359
rect 12759 12325 12768 12359
rect 12716 12316 12768 12325
rect 13820 12359 13872 12368
rect 13820 12325 13829 12359
rect 13829 12325 13863 12359
rect 13863 12325 13872 12359
rect 16488 12359 16540 12368
rect 13820 12316 13872 12325
rect 16488 12325 16497 12359
rect 16497 12325 16531 12359
rect 16531 12325 16540 12359
rect 16488 12316 16540 12325
rect 18696 12316 18748 12368
rect 21088 12359 21140 12368
rect 21088 12325 21097 12359
rect 21097 12325 21131 12359
rect 21131 12325 21140 12359
rect 21088 12316 21140 12325
rect 8760 12223 8812 12232
rect 8760 12189 8769 12223
rect 8769 12189 8803 12223
rect 8803 12189 8812 12223
rect 8760 12180 8812 12189
rect 9404 12180 9456 12232
rect 11704 12248 11756 12300
rect 11796 12291 11848 12300
rect 11796 12257 11805 12291
rect 11805 12257 11839 12291
rect 11839 12257 11848 12291
rect 11796 12248 11848 12257
rect 14648 12248 14700 12300
rect 18144 12248 18196 12300
rect 13728 12223 13780 12232
rect 13728 12189 13737 12223
rect 13737 12189 13771 12223
rect 13771 12189 13780 12223
rect 13728 12180 13780 12189
rect 14096 12223 14148 12232
rect 14096 12189 14105 12223
rect 14105 12189 14139 12223
rect 14139 12189 14148 12223
rect 14096 12180 14148 12189
rect 16856 12180 16908 12232
rect 12624 12112 12676 12164
rect 16948 12155 17000 12164
rect 6920 12087 6972 12096
rect 6920 12053 6929 12087
rect 6929 12053 6963 12087
rect 6963 12053 6972 12087
rect 6920 12044 6972 12053
rect 13084 12087 13136 12096
rect 13084 12053 13093 12087
rect 13093 12053 13127 12087
rect 13127 12053 13136 12087
rect 13084 12044 13136 12053
rect 15936 12044 15988 12096
rect 16948 12121 16957 12155
rect 16957 12121 16991 12155
rect 16991 12121 17000 12155
rect 16948 12112 17000 12121
rect 21364 12180 21416 12232
rect 22744 12112 22796 12164
rect 19064 12044 19116 12096
rect 19248 12044 19300 12096
rect 20076 12087 20128 12096
rect 20076 12053 20085 12087
rect 20085 12053 20119 12087
rect 20119 12053 20128 12087
rect 20076 12044 20128 12053
rect 21916 12087 21968 12096
rect 21916 12053 21925 12087
rect 21925 12053 21959 12087
rect 21959 12053 21968 12087
rect 21916 12044 21968 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2044 11840 2096 11892
rect 4068 11840 4120 11892
rect 4528 11840 4580 11892
rect 6276 11883 6328 11892
rect 6276 11849 6285 11883
rect 6285 11849 6319 11883
rect 6319 11849 6328 11883
rect 6276 11840 6328 11849
rect 11704 11840 11756 11892
rect 13820 11840 13872 11892
rect 14648 11883 14700 11892
rect 14648 11849 14657 11883
rect 14657 11849 14691 11883
rect 14691 11849 14700 11883
rect 14648 11840 14700 11849
rect 15568 11840 15620 11892
rect 16488 11883 16540 11892
rect 16488 11849 16497 11883
rect 16497 11849 16531 11883
rect 16531 11849 16540 11883
rect 16488 11840 16540 11849
rect 16856 11883 16908 11892
rect 16856 11849 16865 11883
rect 16865 11849 16899 11883
rect 16899 11849 16908 11883
rect 16856 11840 16908 11849
rect 18144 11840 18196 11892
rect 4988 11772 5040 11824
rect 8300 11772 8352 11824
rect 5448 11704 5500 11756
rect 5540 11704 5592 11756
rect 1584 11636 1636 11688
rect 2044 11679 2096 11688
rect 2044 11645 2053 11679
rect 2053 11645 2087 11679
rect 2087 11645 2096 11679
rect 2044 11636 2096 11645
rect 2136 11679 2188 11688
rect 2136 11645 2145 11679
rect 2145 11645 2179 11679
rect 2179 11645 2188 11679
rect 2136 11636 2188 11645
rect 2412 11636 2464 11688
rect 3700 11679 3752 11688
rect 3700 11645 3709 11679
rect 3709 11645 3743 11679
rect 3743 11645 3752 11679
rect 3700 11636 3752 11645
rect 2872 11568 2924 11620
rect 4988 11568 5040 11620
rect 5448 11568 5500 11620
rect 5908 11611 5960 11620
rect 5908 11577 5917 11611
rect 5917 11577 5951 11611
rect 5951 11577 5960 11611
rect 5908 11568 5960 11577
rect 6920 11636 6972 11688
rect 7932 11568 7984 11620
rect 8760 11747 8812 11756
rect 8760 11713 8769 11747
rect 8769 11713 8803 11747
rect 8803 11713 8812 11747
rect 8760 11704 8812 11713
rect 12624 11772 12676 11824
rect 13728 11772 13780 11824
rect 16948 11772 17000 11824
rect 18696 11840 18748 11892
rect 19248 11840 19300 11892
rect 21088 11883 21140 11892
rect 21088 11849 21097 11883
rect 21097 11849 21131 11883
rect 21131 11849 21140 11883
rect 21088 11840 21140 11849
rect 22008 11883 22060 11892
rect 22008 11849 22017 11883
rect 22017 11849 22051 11883
rect 22051 11849 22060 11883
rect 22008 11840 22060 11849
rect 13084 11704 13136 11756
rect 13912 11704 13964 11756
rect 10876 11636 10928 11688
rect 11796 11636 11848 11688
rect 14740 11636 14792 11688
rect 15292 11636 15344 11688
rect 16856 11636 16908 11688
rect 18512 11704 18564 11756
rect 19156 11747 19208 11756
rect 19156 11713 19165 11747
rect 19165 11713 19199 11747
rect 19199 11713 19208 11747
rect 19156 11704 19208 11713
rect 21916 11704 21968 11756
rect 22008 11636 22060 11688
rect 9220 11568 9272 11620
rect 9772 11568 9824 11620
rect 13452 11568 13504 11620
rect 16396 11568 16448 11620
rect 18512 11611 18564 11620
rect 18512 11577 18521 11611
rect 18521 11577 18555 11611
rect 18555 11577 18564 11611
rect 18512 11568 18564 11577
rect 18604 11611 18656 11620
rect 18604 11577 18613 11611
rect 18613 11577 18647 11611
rect 18647 11577 18656 11611
rect 18604 11568 18656 11577
rect 19248 11568 19300 11620
rect 1308 11500 1360 11552
rect 3884 11543 3936 11552
rect 3884 11509 3893 11543
rect 3893 11509 3927 11543
rect 3927 11509 3936 11543
rect 3884 11500 3936 11509
rect 6736 11500 6788 11552
rect 7472 11500 7524 11552
rect 8392 11500 8444 11552
rect 9864 11500 9916 11552
rect 13636 11543 13688 11552
rect 13636 11509 13645 11543
rect 13645 11509 13679 11543
rect 13679 11509 13688 11543
rect 13636 11500 13688 11509
rect 21088 11568 21140 11620
rect 20904 11500 20956 11552
rect 21364 11543 21416 11552
rect 21364 11509 21373 11543
rect 21373 11509 21407 11543
rect 21407 11509 21416 11543
rect 21364 11500 21416 11509
rect 21916 11500 21968 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 3976 11296 4028 11348
rect 5540 11296 5592 11348
rect 5908 11296 5960 11348
rect 6828 11296 6880 11348
rect 7840 11339 7892 11348
rect 7840 11305 7849 11339
rect 7849 11305 7883 11339
rect 7883 11305 7892 11339
rect 7840 11296 7892 11305
rect 8760 11296 8812 11348
rect 4252 11271 4304 11280
rect 4252 11237 4261 11271
rect 4261 11237 4295 11271
rect 4295 11237 4304 11271
rect 4252 11228 4304 11237
rect 6092 11271 6144 11280
rect 6092 11237 6101 11271
rect 6101 11237 6135 11271
rect 6135 11237 6144 11271
rect 6092 11228 6144 11237
rect 6276 11228 6328 11280
rect 9404 11271 9456 11280
rect 9404 11237 9413 11271
rect 9413 11237 9447 11271
rect 9447 11237 9456 11271
rect 9404 11228 9456 11237
rect 9864 11271 9916 11280
rect 9864 11237 9873 11271
rect 9873 11237 9907 11271
rect 9907 11237 9916 11271
rect 9864 11228 9916 11237
rect 13452 11339 13504 11348
rect 13452 11305 13461 11339
rect 13461 11305 13495 11339
rect 13495 11305 13504 11339
rect 13452 11296 13504 11305
rect 13820 11296 13872 11348
rect 15292 11296 15344 11348
rect 18512 11296 18564 11348
rect 19524 11296 19576 11348
rect 20904 11296 20956 11348
rect 16396 11228 16448 11280
rect 18604 11271 18656 11280
rect 18604 11237 18613 11271
rect 18613 11237 18647 11271
rect 18647 11237 18656 11271
rect 18604 11228 18656 11237
rect 20076 11228 20128 11280
rect 2872 11203 2924 11212
rect 2872 11169 2881 11203
rect 2881 11169 2915 11203
rect 2915 11169 2924 11203
rect 2872 11160 2924 11169
rect 6000 11160 6052 11212
rect 7840 11203 7892 11212
rect 7840 11169 7849 11203
rect 7849 11169 7883 11203
rect 7883 11169 7892 11203
rect 7840 11160 7892 11169
rect 8024 11203 8076 11212
rect 8024 11169 8033 11203
rect 8033 11169 8067 11203
rect 8067 11169 8076 11203
rect 8024 11160 8076 11169
rect 11428 11160 11480 11212
rect 15752 11203 15804 11212
rect 15752 11169 15761 11203
rect 15761 11169 15795 11203
rect 15795 11169 15804 11203
rect 15752 11160 15804 11169
rect 16764 11160 16816 11212
rect 17592 11160 17644 11212
rect 17960 11203 18012 11212
rect 17960 11169 17969 11203
rect 17969 11169 18003 11203
rect 18003 11169 18012 11203
rect 17960 11160 18012 11169
rect 19064 11203 19116 11212
rect 19064 11169 19073 11203
rect 19073 11169 19107 11203
rect 19107 11169 19116 11203
rect 19064 11160 19116 11169
rect 19340 11160 19392 11212
rect 20904 11160 20956 11212
rect 21916 11160 21968 11212
rect 24216 11160 24268 11212
rect 3148 11135 3200 11144
rect 3148 11101 3157 11135
rect 3157 11101 3191 11135
rect 3191 11101 3200 11135
rect 3148 11092 3200 11101
rect 4160 11135 4212 11144
rect 4160 11101 4169 11135
rect 4169 11101 4203 11135
rect 4203 11101 4212 11135
rect 4160 11092 4212 11101
rect 5264 11092 5316 11144
rect 7012 11135 7064 11144
rect 7012 11101 7021 11135
rect 7021 11101 7055 11135
rect 7055 11101 7064 11135
rect 7012 11092 7064 11101
rect 9404 11092 9456 11144
rect 13544 11092 13596 11144
rect 3332 11024 3384 11076
rect 2044 10999 2096 11008
rect 2044 10965 2053 10999
rect 2053 10965 2087 10999
rect 2087 10965 2096 10999
rect 2044 10956 2096 10965
rect 2412 10956 2464 11008
rect 5356 11024 5408 11076
rect 9496 11024 9548 11076
rect 14096 11024 14148 11076
rect 5540 10999 5592 11008
rect 5540 10965 5549 10999
rect 5549 10965 5583 10999
rect 5583 10965 5592 10999
rect 5540 10956 5592 10965
rect 8208 10956 8260 11008
rect 10784 10999 10836 11008
rect 10784 10965 10793 10999
rect 10793 10965 10827 10999
rect 10827 10965 10836 10999
rect 10784 10956 10836 10965
rect 12256 10999 12308 11008
rect 12256 10965 12265 10999
rect 12265 10965 12299 10999
rect 12299 10965 12308 10999
rect 12256 10956 12308 10965
rect 16672 10999 16724 11008
rect 16672 10965 16681 10999
rect 16681 10965 16715 10999
rect 16715 10965 16724 10999
rect 16672 10956 16724 10965
rect 27712 10956 27764 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 4252 10795 4304 10804
rect 4252 10761 4261 10795
rect 4261 10761 4295 10795
rect 4295 10761 4304 10795
rect 4252 10752 4304 10761
rect 7840 10752 7892 10804
rect 9220 10752 9272 10804
rect 3792 10684 3844 10736
rect 2504 10659 2556 10668
rect 2504 10625 2513 10659
rect 2513 10625 2547 10659
rect 2547 10625 2556 10659
rect 2504 10616 2556 10625
rect 3148 10616 3200 10668
rect 6368 10616 6420 10668
rect 6828 10659 6880 10668
rect 6828 10625 6837 10659
rect 6837 10625 6871 10659
rect 6871 10625 6880 10659
rect 6828 10616 6880 10625
rect 2044 10591 2096 10600
rect 2044 10557 2053 10591
rect 2053 10557 2087 10591
rect 2087 10557 2096 10591
rect 2044 10548 2096 10557
rect 9496 10752 9548 10804
rect 9864 10752 9916 10804
rect 11428 10752 11480 10804
rect 13452 10752 13504 10804
rect 15384 10752 15436 10804
rect 17776 10795 17828 10804
rect 17776 10761 17785 10795
rect 17785 10761 17819 10795
rect 17819 10761 17828 10795
rect 17776 10752 17828 10761
rect 19064 10795 19116 10804
rect 19064 10761 19073 10795
rect 19073 10761 19107 10795
rect 19107 10761 19116 10795
rect 19064 10752 19116 10761
rect 19340 10752 19392 10804
rect 19524 10752 19576 10804
rect 14096 10727 14148 10736
rect 14096 10693 14105 10727
rect 14105 10693 14139 10727
rect 14139 10693 14148 10727
rect 14096 10684 14148 10693
rect 14740 10684 14792 10736
rect 17960 10684 18012 10736
rect 13912 10616 13964 10668
rect 16396 10659 16448 10668
rect 16396 10625 16405 10659
rect 16405 10625 16439 10659
rect 16439 10625 16448 10659
rect 16396 10616 16448 10625
rect 10692 10591 10744 10600
rect 10692 10557 10701 10591
rect 10701 10557 10735 10591
rect 10735 10557 10744 10591
rect 11060 10591 11112 10600
rect 10692 10548 10744 10557
rect 11060 10557 11069 10591
rect 11069 10557 11103 10591
rect 11103 10557 11112 10591
rect 11060 10548 11112 10557
rect 4252 10480 4304 10532
rect 5264 10523 5316 10532
rect 5264 10489 5273 10523
rect 5273 10489 5307 10523
rect 5307 10489 5316 10523
rect 5264 10480 5316 10489
rect 5356 10523 5408 10532
rect 5356 10489 5365 10523
rect 5365 10489 5399 10523
rect 5399 10489 5408 10523
rect 5356 10480 5408 10489
rect 2872 10455 2924 10464
rect 2872 10421 2881 10455
rect 2881 10421 2915 10455
rect 2915 10421 2924 10455
rect 2872 10412 2924 10421
rect 5448 10412 5500 10464
rect 6092 10412 6144 10464
rect 7564 10480 7616 10532
rect 8024 10523 8076 10532
rect 8024 10489 8033 10523
rect 8033 10489 8067 10523
rect 8067 10489 8076 10523
rect 8024 10480 8076 10489
rect 10784 10480 10836 10532
rect 12992 10548 13044 10600
rect 13636 10523 13688 10532
rect 7748 10455 7800 10464
rect 7748 10421 7757 10455
rect 7757 10421 7791 10455
rect 7791 10421 7800 10455
rect 7748 10412 7800 10421
rect 9404 10412 9456 10464
rect 12808 10412 12860 10464
rect 12992 10455 13044 10464
rect 12992 10421 13001 10455
rect 13001 10421 13035 10455
rect 13035 10421 13044 10455
rect 12992 10412 13044 10421
rect 13636 10489 13645 10523
rect 13645 10489 13679 10523
rect 13679 10489 13688 10523
rect 13636 10480 13688 10489
rect 13544 10412 13596 10464
rect 15476 10523 15528 10532
rect 15476 10489 15485 10523
rect 15485 10489 15519 10523
rect 15519 10489 15528 10523
rect 15476 10480 15528 10489
rect 15568 10523 15620 10532
rect 15568 10489 15577 10523
rect 15577 10489 15611 10523
rect 15611 10489 15620 10523
rect 17776 10548 17828 10600
rect 18144 10548 18196 10600
rect 19340 10548 19392 10600
rect 19432 10548 19484 10600
rect 20260 10752 20312 10804
rect 24216 10752 24268 10804
rect 24768 10727 24820 10736
rect 24768 10693 24777 10727
rect 24777 10693 24811 10727
rect 24811 10693 24820 10727
rect 24768 10684 24820 10693
rect 24032 10548 24084 10600
rect 15568 10480 15620 10489
rect 17960 10480 18012 10532
rect 20812 10480 20864 10532
rect 18328 10455 18380 10464
rect 18328 10421 18337 10455
rect 18337 10421 18371 10455
rect 18371 10421 18380 10455
rect 18328 10412 18380 10421
rect 20904 10455 20956 10464
rect 20904 10421 20913 10455
rect 20913 10421 20947 10455
rect 20947 10421 20956 10455
rect 20904 10412 20956 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1400 10208 1452 10260
rect 3148 10208 3200 10260
rect 4160 10208 4212 10260
rect 6000 10208 6052 10260
rect 9312 10208 9364 10260
rect 10692 10208 10744 10260
rect 5356 10140 5408 10192
rect 6276 10140 6328 10192
rect 7748 10140 7800 10192
rect 12256 10140 12308 10192
rect 12716 10140 12768 10192
rect 13912 10208 13964 10260
rect 14832 10208 14884 10260
rect 15476 10208 15528 10260
rect 15752 10251 15804 10260
rect 15752 10217 15761 10251
rect 15761 10217 15795 10251
rect 15795 10217 15804 10251
rect 15752 10208 15804 10217
rect 17592 10251 17644 10260
rect 17592 10217 17601 10251
rect 17601 10217 17635 10251
rect 17635 10217 17644 10251
rect 17592 10208 17644 10217
rect 18144 10251 18196 10260
rect 18144 10217 18153 10251
rect 18153 10217 18187 10251
rect 18187 10217 18196 10251
rect 18144 10208 18196 10217
rect 13544 10140 13596 10192
rect 13728 10140 13780 10192
rect 13820 10140 13872 10192
rect 16672 10140 16724 10192
rect 1860 10115 1912 10124
rect 1860 10081 1869 10115
rect 1869 10081 1903 10115
rect 1903 10081 1912 10115
rect 1860 10072 1912 10081
rect 2412 10115 2464 10124
rect 2412 10081 2421 10115
rect 2421 10081 2455 10115
rect 2455 10081 2464 10115
rect 2412 10072 2464 10081
rect 2504 10115 2556 10124
rect 2504 10081 2513 10115
rect 2513 10081 2547 10115
rect 2547 10081 2556 10115
rect 2688 10115 2740 10124
rect 2504 10072 2556 10081
rect 2688 10081 2697 10115
rect 2697 10081 2731 10115
rect 2731 10081 2740 10115
rect 2688 10072 2740 10081
rect 3332 10072 3384 10124
rect 8208 10072 8260 10124
rect 8852 10072 8904 10124
rect 9588 10072 9640 10124
rect 10324 10115 10376 10124
rect 10324 10081 10333 10115
rect 10333 10081 10367 10115
rect 10367 10081 10376 10115
rect 10324 10072 10376 10081
rect 14188 10115 14240 10124
rect 14188 10081 14197 10115
rect 14197 10081 14231 10115
rect 14231 10081 14240 10115
rect 14188 10072 14240 10081
rect 15384 10072 15436 10124
rect 3148 10047 3200 10056
rect 3148 10013 3157 10047
rect 3157 10013 3191 10047
rect 3191 10013 3200 10047
rect 3148 10004 3200 10013
rect 5080 10004 5132 10056
rect 7840 10004 7892 10056
rect 12164 10004 12216 10056
rect 16764 10004 16816 10056
rect 16948 10047 17000 10056
rect 16948 10013 16957 10047
rect 16957 10013 16991 10047
rect 16991 10013 17000 10047
rect 16948 10004 17000 10013
rect 6368 9936 6420 9988
rect 7472 9936 7524 9988
rect 10784 9979 10836 9988
rect 10784 9945 10793 9979
rect 10793 9945 10827 9979
rect 10827 9945 10836 9979
rect 10784 9936 10836 9945
rect 1860 9868 1912 9920
rect 3608 9868 3660 9920
rect 5264 9868 5316 9920
rect 6552 9868 6604 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1584 9707 1636 9716
rect 1584 9673 1593 9707
rect 1593 9673 1627 9707
rect 1627 9673 1636 9707
rect 1584 9664 1636 9673
rect 2504 9664 2556 9716
rect 6276 9707 6328 9716
rect 6276 9673 6285 9707
rect 6285 9673 6319 9707
rect 6319 9673 6328 9707
rect 6276 9664 6328 9673
rect 6552 9707 6604 9716
rect 6552 9673 6561 9707
rect 6561 9673 6595 9707
rect 6595 9673 6604 9707
rect 6552 9664 6604 9673
rect 8852 9707 8904 9716
rect 8852 9673 8861 9707
rect 8861 9673 8895 9707
rect 8895 9673 8904 9707
rect 8852 9664 8904 9673
rect 10324 9707 10376 9716
rect 10324 9673 10333 9707
rect 10333 9673 10367 9707
rect 10367 9673 10376 9707
rect 10324 9664 10376 9673
rect 12716 9707 12768 9716
rect 12716 9673 12725 9707
rect 12725 9673 12759 9707
rect 12759 9673 12768 9707
rect 12716 9664 12768 9673
rect 13452 9664 13504 9716
rect 13544 9664 13596 9716
rect 14188 9664 14240 9716
rect 15936 9664 15988 9716
rect 16672 9664 16724 9716
rect 5080 9596 5132 9648
rect 6736 9596 6788 9648
rect 2688 9528 2740 9580
rect 3056 9528 3108 9580
rect 3516 9528 3568 9580
rect 3884 9528 3936 9580
rect 7012 9528 7064 9580
rect 7196 9571 7248 9580
rect 7196 9537 7205 9571
rect 7205 9537 7239 9571
rect 7239 9537 7248 9571
rect 7196 9528 7248 9537
rect 8484 9528 8536 9580
rect 9404 9571 9456 9580
rect 9404 9537 9413 9571
rect 9413 9537 9447 9571
rect 9447 9537 9456 9571
rect 9404 9528 9456 9537
rect 12808 9528 12860 9580
rect 13360 9571 13412 9580
rect 13360 9537 13369 9571
rect 13369 9537 13403 9571
rect 13403 9537 13412 9571
rect 13360 9528 13412 9537
rect 13820 9571 13872 9580
rect 13820 9537 13829 9571
rect 13829 9537 13863 9571
rect 13863 9537 13872 9571
rect 13820 9528 13872 9537
rect 1308 9460 1360 9512
rect 3700 9503 3752 9512
rect 112 9392 164 9444
rect 3700 9469 3709 9503
rect 3709 9469 3743 9503
rect 3743 9469 3752 9503
rect 3700 9460 3752 9469
rect 19432 9596 19484 9648
rect 3516 9392 3568 9444
rect 4252 9392 4304 9444
rect 5356 9392 5408 9444
rect 13452 9435 13504 9444
rect 3608 9324 3660 9376
rect 5172 9367 5224 9376
rect 5172 9333 5181 9367
rect 5181 9333 5215 9367
rect 5215 9333 5224 9367
rect 5172 9324 5224 9333
rect 6552 9324 6604 9376
rect 13452 9401 13461 9435
rect 13461 9401 13495 9435
rect 13495 9401 13504 9435
rect 13452 9392 13504 9401
rect 15384 9435 15436 9444
rect 15384 9401 15393 9435
rect 15393 9401 15427 9435
rect 15427 9401 15436 9435
rect 15384 9392 15436 9401
rect 21456 9392 21508 9444
rect 7840 9367 7892 9376
rect 7840 9333 7849 9367
rect 7849 9333 7883 9367
rect 7883 9333 7892 9367
rect 7840 9324 7892 9333
rect 12164 9367 12216 9376
rect 12164 9333 12173 9367
rect 12173 9333 12207 9367
rect 12207 9333 12216 9367
rect 12164 9324 12216 9333
rect 16764 9324 16816 9376
rect 25136 9367 25188 9376
rect 25136 9333 25145 9367
rect 25145 9333 25179 9367
rect 25179 9333 25188 9367
rect 25136 9324 25188 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1584 9163 1636 9172
rect 1584 9129 1593 9163
rect 1593 9129 1627 9163
rect 1627 9129 1636 9163
rect 1584 9120 1636 9129
rect 2412 9163 2464 9172
rect 2412 9129 2421 9163
rect 2421 9129 2455 9163
rect 2455 9129 2464 9163
rect 2412 9120 2464 9129
rect 3884 9120 3936 9172
rect 6644 9120 6696 9172
rect 7656 9120 7708 9172
rect 13360 9163 13412 9172
rect 13360 9129 13369 9163
rect 13369 9129 13403 9163
rect 13403 9129 13412 9163
rect 13360 9120 13412 9129
rect 24768 9163 24820 9172
rect 24768 9129 24777 9163
rect 24777 9129 24811 9163
rect 24811 9129 24820 9163
rect 24768 9120 24820 9129
rect 1952 9052 2004 9104
rect 5172 9095 5224 9104
rect 5172 9061 5181 9095
rect 5181 9061 5215 9095
rect 5215 9061 5224 9095
rect 5172 9052 5224 9061
rect 5264 9052 5316 9104
rect 7196 9052 7248 9104
rect 2320 8984 2372 9036
rect 2964 9027 3016 9036
rect 2964 8993 2973 9027
rect 2973 8993 3007 9027
rect 3007 8993 3016 9027
rect 2964 8984 3016 8993
rect 3608 8916 3660 8968
rect 6000 8916 6052 8968
rect 21732 8984 21784 9036
rect 24676 8984 24728 9036
rect 7564 8848 7616 8900
rect 7012 8823 7064 8832
rect 7012 8789 7021 8823
rect 7021 8789 7055 8823
rect 7055 8789 7064 8823
rect 7012 8780 7064 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1676 8576 1728 8628
rect 2872 8576 2924 8628
rect 5172 8576 5224 8628
rect 7012 8576 7064 8628
rect 7564 8619 7616 8628
rect 7564 8585 7573 8619
rect 7573 8585 7607 8619
rect 7607 8585 7616 8619
rect 7564 8576 7616 8585
rect 24676 8619 24728 8628
rect 24676 8585 24685 8619
rect 24685 8585 24719 8619
rect 24719 8585 24728 8619
rect 24676 8576 24728 8585
rect 2964 8551 3016 8560
rect 2964 8517 2973 8551
rect 2973 8517 3007 8551
rect 3007 8517 3016 8551
rect 2964 8508 3016 8517
rect 3424 8508 3476 8560
rect 2320 8483 2372 8492
rect 2320 8449 2329 8483
rect 2329 8449 2363 8483
rect 2363 8449 2372 8483
rect 2320 8440 2372 8449
rect 1768 8372 1820 8424
rect 2780 8372 2832 8424
rect 5540 8508 5592 8560
rect 6000 8551 6052 8560
rect 6000 8517 6009 8551
rect 6009 8517 6043 8551
rect 6043 8517 6052 8551
rect 6000 8508 6052 8517
rect 13544 8440 13596 8492
rect 1400 8236 1452 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 848 8032 900 8084
rect 4436 8032 4488 8084
rect 7472 8032 7524 8084
rect 3148 7896 3200 7948
rect 4068 7939 4120 7948
rect 4068 7905 4077 7939
rect 4077 7905 4111 7939
rect 4111 7905 4120 7939
rect 4068 7896 4120 7905
rect 4896 7896 4948 7948
rect 1492 7828 1544 7880
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1492 7488 1544 7540
rect 4068 7531 4120 7540
rect 4068 7497 4077 7531
rect 4077 7497 4111 7531
rect 4111 7497 4120 7531
rect 4068 7488 4120 7497
rect 4896 7488 4948 7540
rect 27620 7420 27672 7472
rect 24216 7284 24268 7336
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1584 6987 1636 6996
rect 1584 6953 1593 6987
rect 1593 6953 1627 6987
rect 1627 6953 1636 6987
rect 1584 6944 1636 6953
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 1400 6400 1452 6452
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 27528 5856 27580 5908
rect 24124 5720 24176 5772
rect 24676 5720 24728 5772
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 24676 5355 24728 5364
rect 24676 5321 24685 5355
rect 24685 5321 24719 5355
rect 24719 5321 24728 5355
rect 24676 5312 24728 5321
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 3056 2932 3108 2984
rect 8944 2796 8996 2848
rect 14280 2796 14332 2848
rect 19248 2796 19300 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 7840 2592 7892 2644
rect 8116 2592 8168 2644
rect 12164 2592 12216 2644
rect 21364 2592 21416 2644
rect 24952 2592 25004 2644
rect 5540 2524 5592 2576
rect 7380 2456 7432 2508
rect 19248 2524 19300 2576
rect 7380 2295 7432 2304
rect 7380 2261 7389 2295
rect 7389 2261 7423 2295
rect 7423 2261 7432 2295
rect 7380 2252 7432 2261
rect 14096 2499 14148 2508
rect 14096 2465 14105 2499
rect 14105 2465 14139 2499
rect 14139 2465 14148 2499
rect 14096 2456 14148 2465
rect 18880 2431 18932 2440
rect 18880 2397 18889 2431
rect 18889 2397 18923 2431
rect 18923 2397 18932 2431
rect 18880 2388 18932 2397
rect 16120 2320 16172 2372
rect 20076 2320 20128 2372
rect 9220 2252 9272 2304
rect 24768 2388 24820 2440
rect 22100 2252 22152 2304
rect 22192 2252 22244 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 15844 144 15896 196
rect 11704 76 11756 128
<< metal2 >>
rect 570 27520 626 28000
rect 1766 27554 1822 28000
rect 3054 27554 3110 28000
rect 4342 27554 4398 28000
rect 1688 27526 1822 27554
rect 110 24304 166 24313
rect 110 24239 166 24248
rect 124 24206 152 24239
rect 112 24200 164 24206
rect 112 24142 164 24148
rect 112 23520 164 23526
rect 112 23462 164 23468
rect 20 22976 72 22982
rect 20 22918 72 22924
rect 32 20097 60 22918
rect 124 21185 152 23462
rect 110 21176 166 21185
rect 110 21111 166 21120
rect 18 20088 74 20097
rect 18 20023 74 20032
rect 584 14550 612 27520
rect 1492 23656 1544 23662
rect 1492 23598 1544 23604
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1412 16794 1440 20334
rect 1504 18193 1532 23598
rect 1582 21720 1638 21729
rect 1582 21655 1638 21664
rect 1596 20602 1624 21655
rect 1584 20596 1636 20602
rect 1584 20538 1636 20544
rect 1688 19417 1716 27526
rect 1766 27520 1822 27526
rect 2884 27526 3110 27554
rect 2318 26888 2374 26897
rect 2318 26823 2374 26832
rect 1858 24848 1914 24857
rect 1858 24783 1914 24792
rect 1872 24750 1900 24783
rect 1860 24744 1912 24750
rect 1860 24686 1912 24692
rect 1952 24200 2004 24206
rect 1952 24142 2004 24148
rect 2044 24200 2096 24206
rect 2044 24142 2096 24148
rect 1964 23866 1992 24142
rect 1952 23860 2004 23866
rect 1952 23802 2004 23808
rect 1768 22500 1820 22506
rect 1768 22442 1820 22448
rect 1780 21690 1808 22442
rect 1952 22432 2004 22438
rect 1952 22374 2004 22380
rect 1964 22166 1992 22374
rect 1952 22160 2004 22166
rect 1952 22102 2004 22108
rect 1860 22024 1912 22030
rect 1860 21966 1912 21972
rect 1768 21684 1820 21690
rect 1768 21626 1820 21632
rect 1780 21418 1808 21626
rect 1768 21412 1820 21418
rect 1768 21354 1820 21360
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 1674 19408 1730 19417
rect 1780 19378 1808 19858
rect 1674 19343 1730 19352
rect 1768 19372 1820 19378
rect 1490 18184 1546 18193
rect 1490 18119 1546 18128
rect 1400 16788 1452 16794
rect 1400 16730 1452 16736
rect 664 14952 716 14958
rect 664 14894 716 14900
rect 572 14544 624 14550
rect 572 14486 624 14492
rect 112 9444 164 9450
rect 112 9386 164 9392
rect 124 3505 152 9386
rect 110 3496 166 3505
rect 110 3431 166 3440
rect 676 82 704 14894
rect 1504 14618 1532 18119
rect 1688 17202 1716 19343
rect 1768 19314 1820 19320
rect 1780 19281 1808 19314
rect 1766 19272 1822 19281
rect 1766 19207 1822 19216
rect 1768 18148 1820 18154
rect 1768 18090 1820 18096
rect 1780 17746 1808 18090
rect 1768 17740 1820 17746
rect 1768 17682 1820 17688
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1582 15464 1638 15473
rect 1582 15399 1638 15408
rect 1492 14612 1544 14618
rect 1492 14554 1544 14560
rect 1400 14408 1452 14414
rect 1122 14376 1178 14385
rect 1400 14350 1452 14356
rect 1122 14311 1178 14320
rect 1136 12986 1164 14311
rect 1124 12980 1176 12986
rect 1124 12922 1176 12928
rect 1308 12300 1360 12306
rect 1308 12242 1360 12248
rect 1320 11558 1348 12242
rect 1308 11552 1360 11558
rect 1308 11494 1360 11500
rect 1320 9518 1348 11494
rect 1412 11218 1440 14350
rect 1504 13870 1532 14554
rect 1596 14074 1624 15399
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1492 13864 1544 13870
rect 1872 13814 1900 21966
rect 1964 21060 1992 22102
rect 2056 21554 2084 24142
rect 2228 23656 2280 23662
rect 2228 23598 2280 23604
rect 2240 23497 2268 23598
rect 2226 23488 2282 23497
rect 2226 23423 2282 23432
rect 2332 23186 2360 26823
rect 2320 23180 2372 23186
rect 2320 23122 2372 23128
rect 2780 23180 2832 23186
rect 2780 23122 2832 23128
rect 2320 22976 2372 22982
rect 2320 22918 2372 22924
rect 2044 21548 2096 21554
rect 2044 21490 2096 21496
rect 2044 21072 2096 21078
rect 1964 21032 2044 21060
rect 2044 21014 2096 21020
rect 2056 20262 2084 21014
rect 1952 20256 2004 20262
rect 1952 20198 2004 20204
rect 2044 20256 2096 20262
rect 2044 20198 2096 20204
rect 1964 18698 1992 20198
rect 2136 19712 2188 19718
rect 2136 19654 2188 19660
rect 2148 19242 2176 19654
rect 2136 19236 2188 19242
rect 2136 19178 2188 19184
rect 2148 18902 2176 19178
rect 2136 18896 2188 18902
rect 2136 18838 2188 18844
rect 1952 18692 2004 18698
rect 1952 18634 2004 18640
rect 1964 17746 1992 18634
rect 1952 17740 2004 17746
rect 1952 17682 2004 17688
rect 2228 16652 2280 16658
rect 2228 16594 2280 16600
rect 1952 16040 2004 16046
rect 1952 15982 2004 15988
rect 1964 15638 1992 15982
rect 1952 15632 2004 15638
rect 1952 15574 2004 15580
rect 2136 15428 2188 15434
rect 2136 15370 2188 15376
rect 2148 15026 2176 15370
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 1952 14544 2004 14550
rect 1952 14486 2004 14492
rect 1964 14074 1992 14486
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 1492 13806 1544 13812
rect 1688 13786 1900 13814
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1412 10266 1440 11154
rect 1400 10260 1452 10266
rect 1400 10202 1452 10208
rect 1596 9722 1624 11630
rect 1584 9716 1636 9722
rect 1584 9658 1636 9664
rect 1308 9512 1360 9518
rect 1308 9454 1360 9460
rect 848 8084 900 8090
rect 848 8026 900 8032
rect 860 7993 888 8026
rect 846 7984 902 7993
rect 846 7919 902 7928
rect 1320 1057 1348 9454
rect 1398 9208 1454 9217
rect 1398 9143 1454 9152
rect 1584 9172 1636 9178
rect 1412 8294 1440 9143
rect 1584 9114 1636 9120
rect 1596 9081 1624 9114
rect 1582 9072 1638 9081
rect 1582 9007 1638 9016
rect 1688 8634 1716 13786
rect 1766 12336 1822 12345
rect 1766 12271 1822 12280
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1780 8430 1808 12271
rect 1858 10296 1914 10305
rect 1858 10231 1914 10240
rect 1872 10130 1900 10231
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1400 8288 1452 8294
rect 1400 8230 1452 8236
rect 1412 6866 1440 8230
rect 1490 7984 1546 7993
rect 1490 7919 1546 7928
rect 1504 7886 1532 7919
rect 1492 7880 1544 7886
rect 1492 7822 1544 7828
rect 1504 7546 1532 7822
rect 1492 7540 1544 7546
rect 1492 7482 1544 7488
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1596 6905 1624 6938
rect 1582 6896 1638 6905
rect 1400 6860 1452 6866
rect 1582 6831 1638 6840
rect 1400 6802 1452 6808
rect 1412 6458 1440 6802
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1872 3097 1900 9862
rect 1964 9110 1992 13874
rect 2056 13258 2084 14418
rect 2136 14340 2188 14346
rect 2136 14282 2188 14288
rect 2148 14006 2176 14282
rect 2136 14000 2188 14006
rect 2136 13942 2188 13948
rect 2240 13326 2268 16594
rect 2332 15910 2360 22918
rect 2792 22778 2820 23122
rect 2780 22772 2832 22778
rect 2780 22714 2832 22720
rect 2504 22024 2556 22030
rect 2504 21966 2556 21972
rect 2516 21554 2544 21966
rect 2504 21548 2556 21554
rect 2504 21490 2556 21496
rect 2516 19990 2544 21490
rect 2884 21298 2912 27526
rect 3054 27520 3110 27526
rect 4172 27526 4398 27554
rect 3146 25800 3202 25809
rect 3146 25735 3202 25744
rect 3160 23662 3188 25735
rect 3148 23656 3200 23662
rect 3148 23598 3200 23604
rect 3516 23520 3568 23526
rect 3516 23462 3568 23468
rect 3792 23520 3844 23526
rect 3792 23462 3844 23468
rect 3240 22976 3292 22982
rect 3240 22918 3292 22924
rect 3148 22568 3200 22574
rect 3148 22510 3200 22516
rect 3056 22432 3108 22438
rect 3056 22374 3108 22380
rect 2792 21270 2912 21298
rect 2596 20256 2648 20262
rect 2596 20198 2648 20204
rect 2504 19984 2556 19990
rect 2504 19926 2556 19932
rect 2608 18970 2636 20198
rect 2688 19372 2740 19378
rect 2688 19314 2740 19320
rect 2596 18964 2648 18970
rect 2596 18906 2648 18912
rect 2596 18828 2648 18834
rect 2596 18770 2648 18776
rect 2412 18760 2464 18766
rect 2412 18702 2464 18708
rect 2424 18222 2452 18702
rect 2412 18216 2464 18222
rect 2412 18158 2464 18164
rect 2608 17882 2636 18770
rect 2700 18426 2728 19314
rect 2688 18420 2740 18426
rect 2688 18362 2740 18368
rect 2596 17876 2648 17882
rect 2596 17818 2648 17824
rect 2504 17740 2556 17746
rect 2504 17682 2556 17688
rect 2516 17338 2544 17682
rect 2596 17672 2648 17678
rect 2596 17614 2648 17620
rect 2504 17332 2556 17338
rect 2504 17274 2556 17280
rect 2412 17060 2464 17066
rect 2412 17002 2464 17008
rect 2424 16726 2452 17002
rect 2412 16720 2464 16726
rect 2412 16662 2464 16668
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 2424 16046 2452 16390
rect 2412 16040 2464 16046
rect 2412 15982 2464 15988
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 2320 15564 2372 15570
rect 2320 15506 2372 15512
rect 2332 14890 2360 15506
rect 2424 14958 2452 15982
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 2320 14884 2372 14890
rect 2320 14826 2372 14832
rect 2320 14068 2372 14074
rect 2320 14010 2372 14016
rect 2332 13394 2360 14010
rect 2608 13870 2636 17614
rect 2688 17196 2740 17202
rect 2688 17138 2740 17144
rect 2700 16522 2728 17138
rect 2792 16726 2820 21270
rect 2872 21140 2924 21146
rect 2872 21082 2924 21088
rect 2884 20466 2912 21082
rect 2964 20800 3016 20806
rect 2964 20742 3016 20748
rect 2872 20460 2924 20466
rect 2872 20402 2924 20408
rect 2976 20330 3004 20742
rect 2964 20324 3016 20330
rect 2964 20266 3016 20272
rect 2976 19786 3004 20266
rect 2964 19780 3016 19786
rect 2964 19722 3016 19728
rect 2976 19514 3004 19722
rect 2964 19508 3016 19514
rect 2964 19450 3016 19456
rect 2964 19236 3016 19242
rect 2964 19178 3016 19184
rect 2976 18426 3004 19178
rect 2964 18420 3016 18426
rect 2964 18362 3016 18368
rect 3068 18290 3096 22374
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 3068 17882 3096 18226
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 2780 16720 2832 16726
rect 2780 16662 2832 16668
rect 2688 16516 2740 16522
rect 2688 16458 2740 16464
rect 2700 16250 2728 16458
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 2792 15706 2820 16662
rect 2884 16046 2912 17682
rect 3056 16448 3108 16454
rect 3056 16390 3108 16396
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2792 15162 2820 15642
rect 3068 15609 3096 16390
rect 3054 15600 3110 15609
rect 3054 15535 3110 15544
rect 3160 15502 3188 22510
rect 3252 21078 3280 22918
rect 3528 21078 3556 23462
rect 3608 21888 3660 21894
rect 3608 21830 3660 21836
rect 3620 21418 3648 21830
rect 3608 21412 3660 21418
rect 3608 21354 3660 21360
rect 3240 21072 3292 21078
rect 3240 21014 3292 21020
rect 3516 21072 3568 21078
rect 3516 21014 3568 21020
rect 3332 20460 3384 20466
rect 3332 20402 3384 20408
rect 3240 19984 3292 19990
rect 3240 19926 3292 19932
rect 3252 19514 3280 19926
rect 3344 19854 3372 20402
rect 3620 20058 3648 21354
rect 3700 20324 3752 20330
rect 3700 20266 3752 20272
rect 3608 20052 3660 20058
rect 3608 19994 3660 20000
rect 3332 19848 3384 19854
rect 3332 19790 3384 19796
rect 3516 19848 3568 19854
rect 3516 19790 3568 19796
rect 3240 19508 3292 19514
rect 3240 19450 3292 19456
rect 3240 16244 3292 16250
rect 3240 16186 3292 16192
rect 3252 15502 3280 16186
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 3252 15162 3280 15438
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 3056 14952 3108 14958
rect 3056 14894 3108 14900
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2688 14000 2740 14006
rect 2688 13942 2740 13948
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2412 13456 2464 13462
rect 2412 13398 2464 13404
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2228 13320 2280 13326
rect 2228 13262 2280 13268
rect 2044 13252 2096 13258
rect 2044 13194 2096 13200
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 2056 11898 2084 12038
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 2056 11694 2084 11834
rect 2148 11694 2176 13126
rect 2332 12986 2360 13330
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 2044 11008 2096 11014
rect 2148 10996 2176 11630
rect 2096 10968 2176 10996
rect 2044 10950 2096 10956
rect 2056 10606 2084 10950
rect 2044 10600 2096 10606
rect 2044 10542 2096 10548
rect 1952 9104 2004 9110
rect 1952 9046 2004 9052
rect 1858 3088 1914 3097
rect 1858 3023 1914 3032
rect 2056 2009 2084 10542
rect 2332 10112 2360 12174
rect 2424 11694 2452 13398
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2424 11014 2452 11630
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2516 10674 2544 12786
rect 2608 12782 2636 13806
rect 2700 13734 2728 13942
rect 2884 13814 2912 14758
rect 3068 14618 3096 14894
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 2976 13870 3004 14010
rect 2792 13786 2912 13814
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 3344 13814 3372 19790
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 3436 18834 3464 19654
rect 3424 18828 3476 18834
rect 3424 18770 3476 18776
rect 3528 17610 3556 19790
rect 3608 19712 3660 19718
rect 3608 19654 3660 19660
rect 3620 19378 3648 19654
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 3712 19310 3740 20266
rect 3804 19854 3832 23462
rect 3884 21548 3936 21554
rect 3884 21490 3936 21496
rect 3896 21146 3924 21490
rect 3884 21140 3936 21146
rect 3884 21082 3936 21088
rect 3792 19848 3844 19854
rect 3792 19790 3844 19796
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 3790 19408 3846 19417
rect 3884 19372 3936 19378
rect 3846 19352 3884 19360
rect 3790 19343 3884 19352
rect 3804 19320 3884 19343
rect 3804 19314 3936 19320
rect 3700 19304 3752 19310
rect 3804 19306 3924 19314
rect 3988 19310 4016 19450
rect 3700 19246 3752 19252
rect 3896 19242 3924 19306
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3884 19236 3936 19242
rect 3884 19178 3936 19184
rect 3792 18896 3844 18902
rect 3792 18838 3844 18844
rect 3804 18630 3832 18838
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 3804 18154 3832 18566
rect 3792 18148 3844 18154
rect 3792 18090 3844 18096
rect 3516 17604 3568 17610
rect 3516 17546 3568 17552
rect 3424 17536 3476 17542
rect 3424 17478 3476 17484
rect 3436 17134 3464 17478
rect 3424 17128 3476 17134
rect 3424 17070 3476 17076
rect 3700 17128 3752 17134
rect 3700 17070 3752 17076
rect 3436 16794 3464 17070
rect 3424 16788 3476 16794
rect 3424 16730 3476 16736
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3528 16250 3556 16526
rect 3516 16244 3568 16250
rect 3516 16186 3568 16192
rect 3516 16040 3568 16046
rect 3516 15982 3568 15988
rect 3528 14958 3556 15982
rect 3712 15706 3740 17070
rect 3700 15700 3752 15706
rect 3700 15642 3752 15648
rect 3516 14952 3568 14958
rect 3568 14912 3648 14940
rect 3516 14894 3568 14900
rect 3056 13796 3108 13802
rect 2688 13728 2740 13734
rect 2688 13670 2740 13676
rect 2700 13190 2728 13670
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2516 10130 2544 10610
rect 2700 10130 2728 12922
rect 2412 10124 2464 10130
rect 2332 10084 2412 10112
rect 2412 10066 2464 10072
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2424 9178 2452 10066
rect 2516 9722 2544 10066
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2700 9586 2728 10066
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2332 8498 2360 8978
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2332 8401 2360 8434
rect 2792 8430 2820 13786
rect 3344 13786 3556 13814
rect 3056 13738 3108 13744
rect 3068 13462 3096 13738
rect 3056 13456 3108 13462
rect 3056 13398 3108 13404
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2884 12238 2912 13126
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 3160 12782 3188 12922
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2976 12170 3004 12650
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 2964 12164 3016 12170
rect 2964 12106 3016 12112
rect 2872 11620 2924 11626
rect 2872 11562 2924 11568
rect 2884 11218 2912 11562
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2884 10470 2912 11154
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3160 10674 3188 11086
rect 3332 11076 3384 11082
rect 3332 11018 3384 11024
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2884 8634 2912 10406
rect 3160 10266 3188 10610
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 3344 10130 3372 11018
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2976 8566 3004 8978
rect 2964 8560 3016 8566
rect 2964 8502 3016 8508
rect 2780 8424 2832 8430
rect 2318 8392 2374 8401
rect 2780 8366 2832 8372
rect 2318 8327 2374 8336
rect 3068 2990 3096 9522
rect 3160 7954 3188 9998
rect 3436 8566 3464 12582
rect 3528 9586 3556 13786
rect 3620 13530 3648 14912
rect 3700 14000 3752 14006
rect 3700 13942 3752 13948
rect 3608 13524 3660 13530
rect 3608 13466 3660 13472
rect 3608 12640 3660 12646
rect 3608 12582 3660 12588
rect 3620 9926 3648 12582
rect 3712 12442 3740 13942
rect 3804 13190 3832 18090
rect 3988 17882 4016 19246
rect 4080 18970 4108 19654
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 3976 17876 4028 17882
rect 3976 17818 4028 17824
rect 3884 17196 3936 17202
rect 3884 17138 3936 17144
rect 3896 16726 3924 17138
rect 3884 16720 3936 16726
rect 3884 16662 3936 16668
rect 4172 16402 4200 27526
rect 4342 27520 4398 27526
rect 5630 27520 5686 28000
rect 6918 27554 6974 28000
rect 6656 27526 6974 27554
rect 5644 25226 5672 27520
rect 5632 25220 5684 25226
rect 5632 25162 5684 25168
rect 6552 25220 6604 25226
rect 6552 25162 6604 25168
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6092 24268 6144 24274
rect 6092 24210 6144 24216
rect 6000 24064 6052 24070
rect 6000 24006 6052 24012
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 4804 23724 4856 23730
rect 4804 23666 4856 23672
rect 4620 22092 4672 22098
rect 4620 22034 4672 22040
rect 4632 21690 4660 22034
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4620 21684 4672 21690
rect 4620 21626 4672 21632
rect 4528 20936 4580 20942
rect 4528 20878 4580 20884
rect 4540 20262 4568 20878
rect 4528 20256 4580 20262
rect 4528 20198 4580 20204
rect 4540 18086 4568 20198
rect 4632 20058 4660 21626
rect 4724 20602 4752 21830
rect 4712 20596 4764 20602
rect 4712 20538 4764 20544
rect 4620 20052 4672 20058
rect 4620 19994 4672 20000
rect 4620 19372 4672 19378
rect 4620 19314 4672 19320
rect 4632 18834 4660 19314
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 4632 18426 4660 18770
rect 4724 18698 4752 18770
rect 4712 18692 4764 18698
rect 4712 18634 4764 18640
rect 4620 18420 4672 18426
rect 4620 18362 4672 18368
rect 4632 18222 4660 18362
rect 4620 18216 4672 18222
rect 4620 18158 4672 18164
rect 4528 18080 4580 18086
rect 4528 18022 4580 18028
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4528 17876 4580 17882
rect 4528 17818 4580 17824
rect 4540 17746 4568 17818
rect 4528 17740 4580 17746
rect 4528 17682 4580 17688
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 4264 17066 4292 17274
rect 4436 17196 4488 17202
rect 4540 17184 4568 17682
rect 4488 17156 4568 17184
rect 4436 17138 4488 17144
rect 4252 17060 4304 17066
rect 4252 17002 4304 17008
rect 4448 16658 4476 17138
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 4080 16374 4200 16402
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3896 13814 3924 15846
rect 4080 15026 4108 16374
rect 4448 16250 4476 16594
rect 4436 16244 4488 16250
rect 4436 16186 4488 16192
rect 4252 16176 4304 16182
rect 4252 16118 4304 16124
rect 4264 15570 4292 16118
rect 4448 16046 4476 16186
rect 4436 16040 4488 16046
rect 4436 15982 4488 15988
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4080 14550 4108 14962
rect 4264 14958 4292 15506
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 4068 14544 4120 14550
rect 4068 14486 4120 14492
rect 4264 14482 4292 14894
rect 4448 14618 4476 15982
rect 4436 14612 4488 14618
rect 4436 14554 4488 14560
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 4264 14278 4292 14418
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4068 13864 4120 13870
rect 3896 13786 4016 13814
rect 4264 13814 4292 14214
rect 4068 13806 4120 13812
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3988 12458 4016 13786
rect 4080 13258 4108 13806
rect 4172 13786 4292 13814
rect 4436 13864 4488 13870
rect 4632 13814 4660 18022
rect 4816 17882 4844 23666
rect 4896 23180 4948 23186
rect 4896 23122 4948 23128
rect 4908 22710 4936 23122
rect 4988 22976 5040 22982
rect 4988 22918 5040 22924
rect 5264 22976 5316 22982
rect 6012 22953 6040 24006
rect 6104 23730 6132 24210
rect 6460 24064 6512 24070
rect 6460 24006 6512 24012
rect 6092 23724 6144 23730
rect 6092 23666 6144 23672
rect 6276 23588 6328 23594
rect 6276 23530 6328 23536
rect 6092 23112 6144 23118
rect 6092 23054 6144 23060
rect 5264 22918 5316 22924
rect 5998 22944 6054 22953
rect 4896 22704 4948 22710
rect 4896 22646 4948 22652
rect 4896 21072 4948 21078
rect 4896 21014 4948 21020
rect 4908 20330 4936 21014
rect 5000 20466 5028 22918
rect 5276 22574 5304 22918
rect 5622 22876 5918 22896
rect 5998 22879 6054 22888
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5264 22568 5316 22574
rect 5264 22510 5316 22516
rect 5276 21690 5304 22510
rect 6104 22166 6132 23054
rect 6184 22500 6236 22506
rect 6184 22442 6236 22448
rect 6196 22166 6224 22442
rect 6092 22160 6144 22166
rect 6092 22102 6144 22108
rect 6184 22160 6236 22166
rect 6184 22102 6236 22108
rect 5540 21888 5592 21894
rect 5540 21830 5592 21836
rect 5264 21684 5316 21690
rect 5264 21626 5316 21632
rect 5276 21400 5304 21626
rect 5552 21554 5580 21830
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5356 21412 5408 21418
rect 5276 21372 5356 21400
rect 5356 21354 5408 21360
rect 5368 21146 5396 21354
rect 5356 21140 5408 21146
rect 5356 21082 5408 21088
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 4988 20460 5040 20466
rect 4988 20402 5040 20408
rect 5276 20330 5304 20538
rect 5552 20466 5580 21490
rect 6000 21480 6052 21486
rect 6000 21422 6052 21428
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 4896 20324 4948 20330
rect 4896 20266 4948 20272
rect 5264 20324 5316 20330
rect 5264 20266 5316 20272
rect 4908 19990 4936 20266
rect 5356 20052 5408 20058
rect 5356 19994 5408 20000
rect 4896 19984 4948 19990
rect 4896 19926 4948 19932
rect 4908 19310 4936 19926
rect 5264 19372 5316 19378
rect 5264 19314 5316 19320
rect 4896 19304 4948 19310
rect 4896 19246 4948 19252
rect 5276 19122 5304 19314
rect 5368 19242 5396 19994
rect 5552 19378 5580 20402
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 5356 19236 5408 19242
rect 5356 19178 5408 19184
rect 5540 19236 5592 19242
rect 5540 19178 5592 19184
rect 5552 19122 5580 19178
rect 5276 19094 5580 19122
rect 6012 18884 6040 21422
rect 6104 21146 6132 22102
rect 6196 21690 6224 22102
rect 6184 21684 6236 21690
rect 6184 21626 6236 21632
rect 6092 21140 6144 21146
rect 6092 21082 6144 21088
rect 6184 20256 6236 20262
rect 6184 20198 6236 20204
rect 6092 19168 6144 19174
rect 6196 19156 6224 20198
rect 6288 20074 6316 23530
rect 6368 22432 6420 22438
rect 6368 22374 6420 22380
rect 6380 22030 6408 22374
rect 6368 22024 6420 22030
rect 6368 21966 6420 21972
rect 6380 21554 6408 21966
rect 6368 21548 6420 21554
rect 6368 21490 6420 21496
rect 6288 20046 6408 20074
rect 6276 19916 6328 19922
rect 6276 19858 6328 19864
rect 6288 19514 6316 19858
rect 6276 19508 6328 19514
rect 6276 19450 6328 19456
rect 6144 19128 6224 19156
rect 6092 19110 6144 19116
rect 6196 18970 6224 19128
rect 6276 19168 6328 19174
rect 6276 19110 6328 19116
rect 6184 18964 6236 18970
rect 6184 18906 6236 18912
rect 6012 18856 6132 18884
rect 5448 18828 5500 18834
rect 5448 18770 5500 18776
rect 5080 18760 5132 18766
rect 5080 18702 5132 18708
rect 5092 18222 5120 18702
rect 5460 18222 5488 18770
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 4896 15496 4948 15502
rect 4896 15438 4948 15444
rect 4436 13806 4488 13812
rect 4172 13394 4200 13786
rect 4448 13734 4476 13806
rect 4540 13786 4660 13814
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 4250 13424 4306 13433
rect 4160 13388 4212 13394
rect 4250 13359 4306 13368
rect 4160 13330 4212 13336
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 4172 12646 4200 13330
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3804 12430 4016 12458
rect 4264 12442 4292 13359
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 4252 12436 4304 12442
rect 3712 11694 3740 12378
rect 3700 11688 3752 11694
rect 3700 11630 3752 11636
rect 3804 10742 3832 12430
rect 4252 12378 4304 12384
rect 3976 12368 4028 12374
rect 3976 12310 4028 12316
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3792 10736 3844 10742
rect 3792 10678 3844 10684
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3698 9616 3754 9625
rect 3516 9580 3568 9586
rect 3896 9586 3924 11494
rect 3988 11354 4016 12310
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 4080 11898 4108 12242
rect 4448 12170 4476 12582
rect 4436 12164 4488 12170
rect 4436 12106 4488 12112
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4172 10266 4200 11086
rect 4264 10810 4292 11222
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4252 10532 4304 10538
rect 4252 10474 4304 10480
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 3698 9551 3754 9560
rect 3884 9580 3936 9586
rect 3516 9522 3568 9528
rect 3712 9518 3740 9551
rect 3884 9522 3936 9528
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 3516 9444 3568 9450
rect 3516 9386 3568 9392
rect 3424 8560 3476 8566
rect 3424 8502 3476 8508
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 3056 2984 3108 2990
rect 3056 2926 3108 2932
rect 2042 2000 2098 2009
rect 2042 1935 2098 1944
rect 1306 1048 1362 1057
rect 1306 983 1362 992
rect 1030 82 1086 480
rect 676 54 1086 82
rect 1030 0 1086 54
rect 3146 82 3202 480
rect 3528 82 3556 9386
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3620 8974 3648 9318
rect 3896 9178 3924 9522
rect 4264 9450 4292 10474
rect 4252 9444 4304 9450
rect 4252 9386 4304 9392
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 4448 8090 4476 12106
rect 4540 11898 4568 13786
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4632 12374 4660 13670
rect 4712 13456 4764 13462
rect 4712 13398 4764 13404
rect 4724 12442 4752 13398
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4620 12368 4672 12374
rect 4620 12310 4672 12316
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4908 7954 4936 15438
rect 5000 14958 5028 17274
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 5184 16658 5212 16730
rect 5460 16658 5488 18158
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5552 16998 5580 17478
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5172 16652 5224 16658
rect 5172 16594 5224 16600
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5184 16046 5212 16594
rect 5460 16046 5488 16594
rect 5552 16114 5580 16934
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 5184 15638 5212 15982
rect 5460 15706 5488 15982
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5172 15632 5224 15638
rect 5172 15574 5224 15580
rect 5356 15632 5408 15638
rect 5356 15574 5408 15580
rect 5080 15360 5132 15366
rect 5080 15302 5132 15308
rect 5092 15162 5120 15302
rect 5368 15162 5396 15574
rect 5080 15156 5132 15162
rect 5080 15098 5132 15104
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 4988 14952 5040 14958
rect 4988 14894 5040 14900
rect 5000 14618 5028 14894
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 5172 14476 5224 14482
rect 5172 14418 5224 14424
rect 5184 14074 5212 14418
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5368 13462 5396 15098
rect 5448 15020 5500 15026
rect 5448 14962 5500 14968
rect 5460 14482 5488 14962
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5552 14414 5580 16050
rect 6012 16046 6040 18702
rect 6104 17746 6132 18856
rect 6288 18834 6316 19110
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6092 17740 6144 17746
rect 6092 17682 6144 17688
rect 6104 17338 6132 17682
rect 6092 17332 6144 17338
rect 6092 17274 6144 17280
rect 6196 16658 6224 18022
rect 6288 17814 6316 18770
rect 6276 17808 6328 17814
rect 6276 17750 6328 17756
rect 6380 17202 6408 20046
rect 6472 19990 6500 24006
rect 6564 23474 6592 25162
rect 6656 23866 6684 27526
rect 6918 27520 6974 27526
rect 8114 27554 8170 28000
rect 8114 27526 8248 27554
rect 8114 27520 8170 27526
rect 6920 24268 6972 24274
rect 6920 24210 6972 24216
rect 6828 24132 6880 24138
rect 6828 24074 6880 24080
rect 6644 23860 6696 23866
rect 6644 23802 6696 23808
rect 6644 23656 6696 23662
rect 6644 23598 6696 23604
rect 6656 23474 6684 23598
rect 6564 23446 6684 23474
rect 6460 19984 6512 19990
rect 6460 19926 6512 19932
rect 6460 19848 6512 19854
rect 6460 19790 6512 19796
rect 6472 19446 6500 19790
rect 6460 19440 6512 19446
rect 6460 19382 6512 19388
rect 6552 18828 6604 18834
rect 6552 18770 6604 18776
rect 6564 18426 6592 18770
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6656 18222 6684 23446
rect 6736 22976 6788 22982
rect 6736 22918 6788 22924
rect 6748 22438 6776 22918
rect 6736 22432 6788 22438
rect 6736 22374 6788 22380
rect 6840 21962 6868 24074
rect 6932 23594 6960 24210
rect 8220 23798 8248 27526
rect 9402 27520 9458 28000
rect 10690 27554 10746 28000
rect 11978 27554 12034 28000
rect 10690 27526 10916 27554
rect 10690 27520 10746 27526
rect 9416 25226 9444 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 9404 25220 9456 25226
rect 9404 25162 9456 25168
rect 8668 24676 8720 24682
rect 8668 24618 8720 24624
rect 8208 23792 8260 23798
rect 8208 23734 8260 23740
rect 6920 23588 6972 23594
rect 6920 23530 6972 23536
rect 7748 23520 7800 23526
rect 7748 23462 7800 23468
rect 7564 22432 7616 22438
rect 7564 22374 7616 22380
rect 6828 21956 6880 21962
rect 6828 21898 6880 21904
rect 6840 21468 6868 21898
rect 6920 21480 6972 21486
rect 6840 21440 6920 21468
rect 6840 21146 6868 21440
rect 6920 21422 6972 21428
rect 7472 21412 7524 21418
rect 7472 21354 7524 21360
rect 6828 21140 6880 21146
rect 6828 21082 6880 21088
rect 7484 20942 7512 21354
rect 7472 20936 7524 20942
rect 7472 20878 7524 20884
rect 7484 20058 7512 20878
rect 7472 20052 7524 20058
rect 7472 19994 7524 20000
rect 7576 19990 7604 22374
rect 7760 22234 7788 23462
rect 8024 23180 8076 23186
rect 8024 23122 8076 23128
rect 8036 22438 8064 23122
rect 7840 22432 7892 22438
rect 7840 22374 7892 22380
rect 8024 22432 8076 22438
rect 8024 22374 8076 22380
rect 7748 22228 7800 22234
rect 7748 22170 7800 22176
rect 7748 21140 7800 21146
rect 7748 21082 7800 21088
rect 7760 20330 7788 21082
rect 7748 20324 7800 20330
rect 7748 20266 7800 20272
rect 7760 20058 7788 20266
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 6736 19984 6788 19990
rect 6736 19926 6788 19932
rect 7564 19984 7616 19990
rect 7564 19926 7616 19932
rect 6644 18216 6696 18222
rect 6644 18158 6696 18164
rect 6748 17746 6776 19926
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 6828 18760 6880 18766
rect 6828 18702 6880 18708
rect 6736 17740 6788 17746
rect 6736 17682 6788 17688
rect 6748 17202 6776 17682
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6748 16794 6776 17138
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 6104 16114 6132 16526
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6000 16040 6052 16046
rect 6000 15982 6052 15988
rect 6092 15972 6144 15978
rect 6092 15914 6144 15920
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5356 13456 5408 13462
rect 5078 13424 5134 13433
rect 5356 13398 5408 13404
rect 5078 13359 5134 13368
rect 5092 12918 5120 13359
rect 5080 12912 5132 12918
rect 5080 12854 5132 12860
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 5000 11830 5028 12582
rect 5092 12442 5120 12854
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 4988 11824 5040 11830
rect 4988 11766 5040 11772
rect 5000 11626 5028 11766
rect 4988 11620 5040 11626
rect 5368 11608 5396 12854
rect 5460 11762 5488 13806
rect 5552 13530 5580 14350
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 6012 13394 6040 15846
rect 6104 15502 6132 15914
rect 6196 15910 6224 16594
rect 6644 15972 6696 15978
rect 6644 15914 6696 15920
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 6656 15638 6684 15914
rect 6644 15632 6696 15638
rect 6644 15574 6696 15580
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6104 14618 6132 15438
rect 6656 15094 6684 15574
rect 6840 15201 6868 18702
rect 7196 18080 7248 18086
rect 7196 18022 7248 18028
rect 6920 17604 6972 17610
rect 6920 17546 6972 17552
rect 6826 15192 6882 15201
rect 6826 15127 6882 15136
rect 6932 15094 6960 17546
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6644 15088 6696 15094
rect 6644 15030 6696 15036
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 6092 14612 6144 14618
rect 6092 14554 6144 14560
rect 6184 14476 6236 14482
rect 6184 14418 6236 14424
rect 6196 14074 6224 14418
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 6092 13456 6144 13462
rect 6092 13398 6144 13404
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5552 12696 5580 13262
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6104 12986 6132 13398
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 5816 12708 5868 12714
rect 5552 12668 5816 12696
rect 5816 12650 5868 12656
rect 5828 12442 5856 12650
rect 6104 12646 6132 12922
rect 6380 12850 6408 13126
rect 6656 12986 6684 15030
rect 7024 14822 7052 15302
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 7116 13814 7144 17274
rect 7208 15026 7236 18022
rect 7392 17649 7420 19246
rect 7576 18970 7604 19926
rect 7564 18964 7616 18970
rect 7564 18906 7616 18912
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7668 18222 7696 18566
rect 7760 18426 7788 19994
rect 7748 18420 7800 18426
rect 7748 18362 7800 18368
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 7472 17672 7524 17678
rect 7378 17640 7434 17649
rect 7472 17614 7524 17620
rect 7378 17575 7434 17584
rect 7484 16794 7512 17614
rect 7668 17202 7696 18158
rect 7760 18154 7788 18362
rect 7852 18329 7880 22374
rect 7932 22228 7984 22234
rect 7932 22170 7984 22176
rect 7944 21350 7972 22170
rect 7932 21344 7984 21350
rect 7932 21286 7984 21292
rect 7944 21078 7972 21286
rect 7932 21072 7984 21078
rect 7932 21014 7984 21020
rect 7944 20262 7972 21014
rect 8036 20602 8064 22374
rect 8220 21010 8248 23734
rect 8484 23656 8536 23662
rect 8484 23598 8536 23604
rect 8392 23520 8444 23526
rect 8392 23462 8444 23468
rect 8404 21622 8432 23462
rect 8496 22710 8524 23598
rect 8680 23322 8708 24618
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10600 24064 10652 24070
rect 10600 24006 10652 24012
rect 10612 23662 10640 24006
rect 10600 23656 10652 23662
rect 10652 23616 10732 23644
rect 10600 23598 10652 23604
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 8668 23316 8720 23322
rect 8668 23258 8720 23264
rect 8576 22976 8628 22982
rect 8576 22918 8628 22924
rect 8484 22704 8536 22710
rect 8484 22646 8536 22652
rect 8392 21616 8444 21622
rect 8392 21558 8444 21564
rect 8404 21146 8432 21558
rect 8392 21140 8444 21146
rect 8392 21082 8444 21088
rect 8116 21004 8168 21010
rect 8116 20946 8168 20952
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 8024 20596 8076 20602
rect 8024 20538 8076 20544
rect 7932 20256 7984 20262
rect 7932 20198 7984 20204
rect 7944 20058 7972 20198
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 7944 18834 7972 19994
rect 8036 18873 8064 20538
rect 8022 18864 8078 18873
rect 7932 18828 7984 18834
rect 8022 18799 8078 18808
rect 7932 18770 7984 18776
rect 8128 18766 8156 20946
rect 8496 20754 8524 22646
rect 8588 22506 8616 22918
rect 8680 22642 8708 23258
rect 10416 23248 10468 23254
rect 10416 23190 10468 23196
rect 10428 23089 10456 23190
rect 10414 23080 10470 23089
rect 9496 23044 9548 23050
rect 10414 23015 10470 23024
rect 9496 22986 9548 22992
rect 8668 22636 8720 22642
rect 8668 22578 8720 22584
rect 8576 22500 8628 22506
rect 8576 22442 8628 22448
rect 8944 22500 8996 22506
rect 8944 22442 8996 22448
rect 8588 21418 8616 22442
rect 8760 22024 8812 22030
rect 8760 21966 8812 21972
rect 8772 21554 8800 21966
rect 8956 21554 8984 22442
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 8760 21548 8812 21554
rect 8760 21490 8812 21496
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 8576 21412 8628 21418
rect 8576 21354 8628 21360
rect 8588 20806 8616 21354
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8404 20726 8524 20754
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 8220 18902 8248 19110
rect 8208 18896 8260 18902
rect 8208 18838 8260 18844
rect 8116 18760 8168 18766
rect 8116 18702 8168 18708
rect 7838 18320 7894 18329
rect 7838 18255 7894 18264
rect 7748 18148 7800 18154
rect 7748 18090 7800 18096
rect 7760 17814 7788 18090
rect 8128 17882 8156 18702
rect 8220 17882 8248 18838
rect 8116 17876 8168 17882
rect 8116 17818 8168 17824
rect 8208 17876 8260 17882
rect 8208 17818 8260 17824
rect 7748 17808 7800 17814
rect 7748 17750 7800 17756
rect 7760 17338 7788 17750
rect 8220 17338 8248 17818
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 7300 15706 7328 16050
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7208 14618 7236 14962
rect 7472 14884 7524 14890
rect 7472 14826 7524 14832
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 7116 13786 7236 13814
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 5816 12436 5868 12442
rect 5816 12378 5868 12384
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5552 11762 5580 12242
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5448 11620 5500 11626
rect 5368 11580 5448 11608
rect 4988 11562 5040 11568
rect 5448 11562 5500 11568
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5276 10538 5304 11086
rect 5356 11076 5408 11082
rect 5356 11018 5408 11024
rect 5368 10538 5396 11018
rect 5460 10996 5488 11562
rect 5552 11354 5580 11698
rect 5908 11620 5960 11626
rect 5908 11562 5960 11568
rect 5920 11354 5948 11562
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5908 11348 5960 11354
rect 5908 11290 5960 11296
rect 6012 11218 6040 12174
rect 6104 11286 6132 12582
rect 6276 12368 6328 12374
rect 6276 12310 6328 12316
rect 6288 11898 6316 12310
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6288 11286 6316 11834
rect 6092 11280 6144 11286
rect 6092 11222 6144 11228
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 5540 11008 5592 11014
rect 5460 10968 5540 10996
rect 5540 10950 5592 10956
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 5092 9654 5120 9998
rect 5276 9926 5304 10474
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5356 10192 5408 10198
rect 5460 10180 5488 10406
rect 5408 10152 5488 10180
rect 5356 10134 5408 10140
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5184 9110 5212 9318
rect 5276 9110 5304 9862
rect 5368 9450 5396 10134
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5172 9104 5224 9110
rect 5172 9046 5224 9052
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 5184 8634 5212 9046
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5552 8566 5580 10950
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6012 10266 6040 11154
rect 6104 10470 6132 11222
rect 6380 10674 6408 12786
rect 7024 12714 7052 13126
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6288 9722 6316 10134
rect 6380 9994 6408 10610
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6564 9722 6592 9862
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6564 9382 6592 9658
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6656 9178 6684 12582
rect 7012 12300 7064 12306
rect 7116 12288 7144 13126
rect 7208 12442 7236 13786
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7064 12260 7144 12288
rect 7012 12242 7064 12248
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6932 11694 6960 12038
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6748 9654 6776 11494
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6840 10674 6868 11290
rect 7024 11150 7052 12242
rect 7484 12073 7512 14826
rect 7470 12064 7526 12073
rect 7470 11999 7526 12008
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 7484 9994 7512 11494
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6012 8566 6040 8910
rect 7024 8838 7052 9522
rect 7208 9110 7236 9522
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 7024 8634 7052 8774
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 7484 8090 7512 9930
rect 7576 8906 7604 10474
rect 7668 9178 7696 17002
rect 7760 16114 7788 17274
rect 8220 16998 8248 17274
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 7932 16652 7984 16658
rect 7932 16594 7984 16600
rect 7944 16250 7972 16594
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8312 16250 8340 16390
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 7760 15978 7788 16050
rect 7748 15972 7800 15978
rect 7748 15914 7800 15920
rect 7944 15706 7972 16186
rect 8312 15910 8340 16186
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7944 15162 7972 15642
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 8128 15026 8156 15438
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 8128 14414 8156 14962
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 7852 12442 7880 13262
rect 7944 13190 7972 13806
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 7852 11354 7880 12378
rect 7932 11620 7984 11626
rect 7984 11580 8064 11608
rect 7932 11562 7984 11568
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 8036 11218 8064 11580
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 7852 10810 7880 11154
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 8036 10538 8064 11154
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7760 10198 7788 10406
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7852 9382 7880 9998
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7576 8634 7604 8842
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4080 7546 4108 7890
rect 4908 7546 4936 7890
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5446 5400 5502 5409
rect 5622 5392 5918 5412
rect 5446 5335 5502 5344
rect 5460 5137 5488 5335
rect 5446 5128 5502 5137
rect 5446 5063 5502 5072
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 7852 2650 7880 9318
rect 8128 2650 8156 14214
rect 8404 13814 8432 20726
rect 8680 20466 8708 21286
rect 9312 21004 9364 21010
rect 9312 20946 9364 20952
rect 8760 20528 8812 20534
rect 8760 20470 8812 20476
rect 8668 20460 8720 20466
rect 8668 20402 8720 20408
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8588 17066 8616 19110
rect 8576 17060 8628 17066
rect 8576 17002 8628 17008
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 8496 15978 8524 16390
rect 8484 15972 8536 15978
rect 8484 15914 8536 15920
rect 8312 13802 8432 13814
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 8300 13796 8432 13802
rect 8352 13786 8432 13796
rect 8300 13738 8352 13744
rect 8220 12850 8248 13738
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 8312 12986 8340 13398
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 8312 12714 8340 12922
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8220 11014 8248 12242
rect 8312 11830 8340 12650
rect 8392 12300 8444 12306
rect 8392 12242 8444 12248
rect 8300 11824 8352 11830
rect 8300 11766 8352 11772
rect 8404 11558 8432 12242
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8220 10130 8248 10950
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8496 9586 8524 15914
rect 8576 14884 8628 14890
rect 8576 14826 8628 14832
rect 8588 14550 8616 14826
rect 8576 14544 8628 14550
rect 8576 14486 8628 14492
rect 8588 14074 8616 14486
rect 8576 14068 8628 14074
rect 8576 14010 8628 14016
rect 8576 13796 8628 13802
rect 8576 13738 8628 13744
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8588 5137 8616 13738
rect 8680 11529 8708 20402
rect 8772 19990 8800 20470
rect 9220 20460 9272 20466
rect 9220 20402 9272 20408
rect 9128 20256 9180 20262
rect 9128 20198 9180 20204
rect 9140 20058 9168 20198
rect 9128 20052 9180 20058
rect 9128 19994 9180 20000
rect 8760 19984 8812 19990
rect 8760 19926 8812 19932
rect 9232 19378 9260 20402
rect 9324 20262 9352 20946
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 9220 19372 9272 19378
rect 9220 19314 9272 19320
rect 9036 19236 9088 19242
rect 9036 19178 9088 19184
rect 9048 18358 9076 19178
rect 9232 18970 9260 19314
rect 9324 19281 9352 20198
rect 9310 19272 9366 19281
rect 9310 19207 9366 19216
rect 9220 18964 9272 18970
rect 9220 18906 9272 18912
rect 9128 18692 9180 18698
rect 9128 18634 9180 18640
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 8942 18184 8998 18193
rect 8942 18119 8998 18128
rect 8956 16697 8984 18119
rect 9140 17270 9168 18634
rect 9416 17338 9444 21830
rect 9508 20330 9536 22986
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 9588 22092 9640 22098
rect 9588 22034 9640 22040
rect 9600 21350 9628 22034
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 10060 21418 10088 21830
rect 9772 21412 9824 21418
rect 9772 21354 9824 21360
rect 10048 21412 10100 21418
rect 10048 21354 10100 21360
rect 10140 21412 10192 21418
rect 10140 21354 10192 21360
rect 9588 21344 9640 21350
rect 9588 21286 9640 21292
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9496 20324 9548 20330
rect 9496 20266 9548 20272
rect 9508 19990 9536 20266
rect 9600 20262 9628 20742
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 9496 19984 9548 19990
rect 9496 19926 9548 19932
rect 9588 19916 9640 19922
rect 9588 19858 9640 19864
rect 9600 19174 9628 19858
rect 9588 19168 9640 19174
rect 9588 19110 9640 19116
rect 9692 18970 9720 20742
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9692 18426 9720 18906
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9784 18306 9812 21354
rect 10152 21078 10180 21354
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10140 21072 10192 21078
rect 10140 21014 10192 21020
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10232 19916 10284 19922
rect 10232 19858 10284 19864
rect 10244 19514 10272 19858
rect 10704 19514 10732 23616
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 10796 19922 10824 21830
rect 10784 19916 10836 19922
rect 10784 19858 10836 19864
rect 10232 19508 10284 19514
rect 10232 19450 10284 19456
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9876 18902 9904 19110
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 9864 18896 9916 18902
rect 9864 18838 9916 18844
rect 9692 18278 9812 18306
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 8942 16688 8998 16697
rect 8942 16623 8998 16632
rect 9312 15972 9364 15978
rect 9312 15914 9364 15920
rect 9324 15638 9352 15914
rect 9312 15632 9364 15638
rect 9312 15574 9364 15580
rect 9324 15473 9352 15574
rect 9310 15464 9366 15473
rect 9310 15399 9366 15408
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9036 14000 9088 14006
rect 9036 13942 9088 13948
rect 9048 13326 9076 13942
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 9048 12442 9076 12786
rect 9140 12782 9168 13670
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8772 11762 8800 12174
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8666 11520 8722 11529
rect 8666 11455 8722 11464
rect 8680 7857 8708 11455
rect 8772 11354 8800 11698
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 9232 10810 9260 11562
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 9324 10266 9352 14010
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9416 11286 9444 12174
rect 9404 11280 9456 11286
rect 9456 11240 9628 11268
rect 9404 11222 9456 11228
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9416 10470 9444 11086
rect 9496 11076 9548 11082
rect 9496 11018 9548 11024
rect 9508 10810 9536 11018
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8864 9722 8892 10066
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 9416 9586 9444 10406
rect 9600 10130 9628 11240
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 8666 7848 8722 7857
rect 8666 7783 8722 7792
rect 8574 5128 8630 5137
rect 8574 5063 8630 5072
rect 9692 4154 9720 18278
rect 9876 18154 9904 18838
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 9864 18148 9916 18154
rect 9864 18090 9916 18096
rect 9968 17882 9996 18226
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 9956 17876 10008 17882
rect 9956 17818 10008 17824
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 10600 17740 10652 17746
rect 10600 17682 10652 17688
rect 10152 16998 10180 17682
rect 10612 17270 10640 17682
rect 10600 17264 10652 17270
rect 10600 17206 10652 17212
rect 10612 17134 10640 17206
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9784 15910 9812 16526
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 9784 15706 9812 15846
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 10060 15162 10088 15506
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 10152 13530 10180 16934
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10704 15638 10732 19450
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10796 18834 10824 19314
rect 10888 18873 10916 27526
rect 11624 27526 12034 27554
rect 11336 24608 11388 24614
rect 11336 24550 11388 24556
rect 11348 24274 11376 24550
rect 11624 24410 11652 27526
rect 11978 27520 12034 27526
rect 13266 27520 13322 28000
rect 14554 27520 14610 28000
rect 15750 27520 15806 28000
rect 17038 27554 17094 28000
rect 16684 27526 17094 27554
rect 12164 25356 12216 25362
rect 12164 25298 12216 25304
rect 12716 25356 12768 25362
rect 12716 25298 12768 25304
rect 12176 24614 12204 25298
rect 12440 25152 12492 25158
rect 12440 25094 12492 25100
rect 12532 25152 12584 25158
rect 12532 25094 12584 25100
rect 12256 24676 12308 24682
rect 12256 24618 12308 24624
rect 12164 24608 12216 24614
rect 12164 24550 12216 24556
rect 11612 24404 11664 24410
rect 11612 24346 11664 24352
rect 11336 24268 11388 24274
rect 11336 24210 11388 24216
rect 11348 23866 11376 24210
rect 11336 23860 11388 23866
rect 11336 23802 11388 23808
rect 10968 23656 11020 23662
rect 10968 23598 11020 23604
rect 10980 23526 11008 23598
rect 11060 23588 11112 23594
rect 11060 23530 11112 23536
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 11072 21010 11100 23530
rect 11336 23520 11388 23526
rect 11336 23462 11388 23468
rect 11348 22574 11376 23462
rect 11704 23112 11756 23118
rect 11704 23054 11756 23060
rect 11716 22778 11744 23054
rect 12072 23044 12124 23050
rect 12072 22986 12124 22992
rect 11704 22772 11756 22778
rect 11704 22714 11756 22720
rect 11336 22568 11388 22574
rect 11336 22510 11388 22516
rect 11152 22432 11204 22438
rect 11152 22374 11204 22380
rect 11164 22030 11192 22374
rect 11244 22160 11296 22166
rect 11244 22102 11296 22108
rect 11152 22024 11204 22030
rect 11152 21966 11204 21972
rect 11164 21690 11192 21966
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 11256 21350 11284 22102
rect 11348 21962 11376 22510
rect 12084 21962 12112 22986
rect 12176 22710 12204 24550
rect 12164 22704 12216 22710
rect 12164 22646 12216 22652
rect 11336 21956 11388 21962
rect 11336 21898 11388 21904
rect 12072 21956 12124 21962
rect 12072 21898 12124 21904
rect 12084 21622 12112 21898
rect 12072 21616 12124 21622
rect 12072 21558 12124 21564
rect 11244 21344 11296 21350
rect 11244 21286 11296 21292
rect 12164 21344 12216 21350
rect 12164 21286 12216 21292
rect 11256 21078 11284 21286
rect 12176 21146 12204 21286
rect 12164 21140 12216 21146
rect 12164 21082 12216 21088
rect 11244 21072 11296 21078
rect 11244 21014 11296 21020
rect 11060 21004 11112 21010
rect 11060 20946 11112 20952
rect 11072 20058 11100 20946
rect 11256 20602 11284 21014
rect 11244 20596 11296 20602
rect 11244 20538 11296 20544
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11624 19378 11652 19790
rect 11612 19372 11664 19378
rect 11612 19314 11664 19320
rect 11428 19236 11480 19242
rect 11428 19178 11480 19184
rect 10874 18864 10930 18873
rect 10784 18828 10836 18834
rect 10874 18799 10930 18808
rect 10784 18770 10836 18776
rect 10796 18737 10824 18770
rect 10968 18760 11020 18766
rect 10782 18728 10838 18737
rect 10968 18702 11020 18708
rect 10782 18663 10838 18672
rect 10980 18086 11008 18702
rect 11440 18698 11468 19178
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11716 18970 11744 19110
rect 11704 18964 11756 18970
rect 11704 18906 11756 18912
rect 11428 18692 11480 18698
rect 11428 18634 11480 18640
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 10980 17814 11008 18022
rect 11440 17882 11468 18634
rect 11716 18426 11744 18906
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11612 18352 11664 18358
rect 11518 18320 11574 18329
rect 11612 18294 11664 18300
rect 11518 18255 11574 18264
rect 11532 18222 11560 18255
rect 11520 18216 11572 18222
rect 11520 18158 11572 18164
rect 11624 17882 11652 18294
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11612 17876 11664 17882
rect 11612 17818 11664 17824
rect 10968 17808 11020 17814
rect 10968 17750 11020 17756
rect 11440 17270 11468 17818
rect 11624 17678 11652 17818
rect 11612 17672 11664 17678
rect 11612 17614 11664 17620
rect 10784 17264 10836 17270
rect 10784 17206 10836 17212
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 10796 16028 10824 17206
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 11072 16794 11100 16934
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 11716 16726 11744 18362
rect 11888 17808 11940 17814
rect 11888 17750 11940 17756
rect 11900 16998 11928 17750
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12176 17202 12204 17614
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11704 16720 11756 16726
rect 11704 16662 11756 16668
rect 11716 16250 11744 16662
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 10876 16040 10928 16046
rect 10796 16000 10876 16028
rect 10796 15706 10824 16000
rect 10876 15982 10928 15988
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10704 15162 10732 15574
rect 11348 15502 11376 16050
rect 11716 15706 11744 16186
rect 11900 15706 11928 16934
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 12268 15502 12296 24618
rect 12452 24274 12480 25094
rect 12440 24268 12492 24274
rect 12440 24210 12492 24216
rect 12544 23730 12572 25094
rect 12728 24954 12756 25298
rect 13280 24954 13308 27520
rect 13544 25220 13596 25226
rect 13544 25162 13596 25168
rect 12716 24948 12768 24954
rect 12716 24890 12768 24896
rect 13268 24948 13320 24954
rect 13268 24890 13320 24896
rect 13452 24268 13504 24274
rect 13452 24210 13504 24216
rect 13464 23866 13492 24210
rect 13556 24177 13584 25162
rect 14096 24744 14148 24750
rect 14096 24686 14148 24692
rect 13542 24168 13598 24177
rect 13542 24103 13598 24112
rect 13452 23860 13504 23866
rect 13452 23802 13504 23808
rect 12532 23724 12584 23730
rect 12532 23666 12584 23672
rect 12808 23724 12860 23730
rect 12808 23666 12860 23672
rect 12544 23322 12572 23666
rect 12716 23520 12768 23526
rect 12716 23462 12768 23468
rect 12532 23316 12584 23322
rect 12532 23258 12584 23264
rect 12728 23254 12756 23462
rect 12716 23248 12768 23254
rect 12716 23190 12768 23196
rect 12532 22976 12584 22982
rect 12532 22918 12584 22924
rect 12544 22506 12572 22918
rect 12532 22500 12584 22506
rect 12532 22442 12584 22448
rect 12624 22500 12676 22506
rect 12624 22442 12676 22448
rect 12636 22234 12664 22442
rect 12728 22438 12756 23190
rect 12820 22982 12848 23666
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 13268 22704 13320 22710
rect 13268 22646 13320 22652
rect 12716 22432 12768 22438
rect 12716 22374 12768 22380
rect 12624 22228 12676 22234
rect 12624 22170 12676 22176
rect 12440 21684 12492 21690
rect 12440 21626 12492 21632
rect 12348 19440 12400 19446
rect 12348 19382 12400 19388
rect 12360 18630 12388 19382
rect 12348 18624 12400 18630
rect 12348 18566 12400 18572
rect 12360 17066 12388 18566
rect 12348 17060 12400 17066
rect 12348 17002 12400 17008
rect 12360 16726 12388 17002
rect 12348 16720 12400 16726
rect 12348 16662 12400 16668
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14618 10732 15098
rect 11164 15094 11192 15302
rect 11348 15162 11376 15438
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 11244 14884 11296 14890
rect 11244 14826 11296 14832
rect 11520 14884 11572 14890
rect 11520 14826 11572 14832
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10244 14074 10272 14418
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10704 13841 10732 14418
rect 11256 14278 11284 14826
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11256 14074 11284 14214
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11532 13938 11560 14826
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 11992 14618 12020 14758
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11992 14006 12020 14554
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 11980 14000 12032 14006
rect 11980 13942 12032 13948
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 11520 13932 11572 13938
rect 11520 13874 11572 13880
rect 10690 13832 10746 13841
rect 10690 13767 10746 13776
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9876 13297 9904 13330
rect 9862 13288 9918 13297
rect 9862 13223 9918 13232
rect 10704 13190 10732 13767
rect 10796 13530 10824 13874
rect 11992 13802 12020 13942
rect 11980 13796 12032 13802
rect 11980 13738 12032 13744
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11900 13530 11928 13670
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11992 13462 12020 13738
rect 12268 13530 12296 14350
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 11980 13456 12032 13462
rect 11980 13398 12032 13404
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10428 12782 10456 13126
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 9784 12306 9812 12718
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10796 12442 10824 13330
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 10980 12850 11008 13262
rect 11704 13252 11756 13258
rect 11704 13194 11756 13200
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 10966 12608 11022 12617
rect 10966 12543 11022 12552
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9784 11626 9812 12242
rect 10876 11688 10928 11694
rect 10796 11648 10876 11676
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9876 11286 9904 11494
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 9876 10810 9904 11222
rect 10796 11014 10824 11648
rect 10876 11630 10928 11636
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10704 10266 10732 10542
rect 10796 10538 10824 10950
rect 10784 10532 10836 10538
rect 10784 10474 10836 10480
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10336 9722 10364 10066
rect 10796 9994 10824 10474
rect 10784 9988 10836 9994
rect 10784 9930 10836 9936
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10980 7993 11008 12543
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11440 11218 11468 12378
rect 11716 12306 11744 13194
rect 11992 12918 12020 13398
rect 11980 12912 12032 12918
rect 11980 12854 12032 12860
rect 12452 12617 12480 21626
rect 12532 20800 12584 20806
rect 12532 20742 12584 20748
rect 12624 20800 12676 20806
rect 12728 20788 12756 22374
rect 13280 22030 13308 22646
rect 13452 22160 13504 22166
rect 13452 22102 13504 22108
rect 12992 22024 13044 22030
rect 12992 21966 13044 21972
rect 13268 22024 13320 22030
rect 13268 21966 13320 21972
rect 13004 21418 13032 21966
rect 13280 21554 13308 21966
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 12992 21412 13044 21418
rect 12992 21354 13044 21360
rect 12808 20936 12860 20942
rect 12808 20878 12860 20884
rect 12676 20760 12756 20788
rect 12624 20742 12676 20748
rect 12544 20466 12572 20742
rect 12532 20460 12584 20466
rect 12532 20402 12584 20408
rect 12544 20369 12572 20402
rect 12530 20360 12586 20369
rect 12636 20330 12664 20742
rect 12530 20295 12586 20304
rect 12624 20324 12676 20330
rect 12624 20266 12676 20272
rect 12820 20058 12848 20878
rect 13004 20534 13032 21354
rect 13464 21350 13492 22102
rect 13556 21690 13584 24103
rect 13820 23656 13872 23662
rect 13820 23598 13872 23604
rect 13728 23180 13780 23186
rect 13728 23122 13780 23128
rect 13740 22778 13768 23122
rect 13728 22772 13780 22778
rect 13728 22714 13780 22720
rect 13544 21684 13596 21690
rect 13544 21626 13596 21632
rect 13544 21480 13596 21486
rect 13544 21422 13596 21428
rect 13452 21344 13504 21350
rect 13452 21286 13504 21292
rect 12992 20528 13044 20534
rect 12992 20470 13044 20476
rect 12808 20052 12860 20058
rect 12808 19994 12860 20000
rect 13464 19922 13492 21286
rect 13556 21078 13584 21422
rect 13544 21072 13596 21078
rect 13544 21014 13596 21020
rect 13556 20262 13584 21014
rect 13740 20602 13768 22714
rect 13832 21894 13860 23598
rect 14108 23497 14136 24686
rect 14568 24410 14596 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15200 24744 15252 24750
rect 15200 24686 15252 24692
rect 14556 24404 14608 24410
rect 14556 24346 14608 24352
rect 15212 24177 15240 24686
rect 15384 24676 15436 24682
rect 15384 24618 15436 24624
rect 15198 24168 15254 24177
rect 15198 24103 15254 24112
rect 14188 24064 14240 24070
rect 14188 24006 14240 24012
rect 14200 23662 14228 24006
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14648 23724 14700 23730
rect 14648 23666 14700 23672
rect 14188 23656 14240 23662
rect 14188 23598 14240 23604
rect 14094 23488 14150 23497
rect 14094 23423 14150 23432
rect 14200 23186 14228 23598
rect 14188 23180 14240 23186
rect 14188 23122 14240 23128
rect 13912 22636 13964 22642
rect 13912 22578 13964 22584
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13728 20596 13780 20602
rect 13728 20538 13780 20544
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 13556 19990 13584 20198
rect 13544 19984 13596 19990
rect 13544 19926 13596 19932
rect 13452 19916 13504 19922
rect 13452 19858 13504 19864
rect 13556 19861 13584 19926
rect 13636 19916 13688 19922
rect 13636 19858 13688 19864
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13372 19378 13400 19790
rect 13648 19514 13676 19858
rect 13636 19508 13688 19514
rect 13636 19450 13688 19456
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 12532 19236 12584 19242
rect 12532 19178 12584 19184
rect 12624 19236 12676 19242
rect 12624 19178 12676 19184
rect 12544 18630 12572 19178
rect 12636 18902 12664 19178
rect 13648 19145 13676 19450
rect 13924 19446 13952 22578
rect 14200 22438 14228 23122
rect 14370 22944 14426 22953
rect 14370 22879 14426 22888
rect 14384 22642 14412 22879
rect 14372 22636 14424 22642
rect 14372 22578 14424 22584
rect 14188 22432 14240 22438
rect 14188 22374 14240 22380
rect 14004 20460 14056 20466
rect 14004 20402 14056 20408
rect 13912 19440 13964 19446
rect 13912 19382 13964 19388
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13740 19174 13768 19246
rect 13728 19168 13780 19174
rect 13634 19136 13690 19145
rect 13728 19110 13780 19116
rect 13634 19071 13690 19080
rect 12624 18896 12676 18902
rect 12624 18838 12676 18844
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12636 18154 12664 18838
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 12624 18148 12676 18154
rect 12624 18090 12676 18096
rect 12912 17542 12940 18226
rect 13004 17785 13032 18566
rect 13556 18086 13584 18702
rect 13636 18352 13688 18358
rect 13636 18294 13688 18300
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13556 17921 13584 18022
rect 13542 17912 13598 17921
rect 13542 17847 13598 17856
rect 12990 17776 13046 17785
rect 12990 17711 13046 17720
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 12900 17536 12952 17542
rect 12900 17478 12952 17484
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12820 16794 12848 16934
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12544 15910 12572 16390
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 12636 15366 12664 15982
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12532 14340 12584 14346
rect 12532 14282 12584 14288
rect 12544 13938 12572 14282
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12544 13530 12572 13874
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12636 12646 12664 15302
rect 12912 15162 12940 17478
rect 13556 16998 13584 17682
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 13556 16182 13584 16934
rect 13648 16658 13676 18294
rect 13740 17746 13768 19110
rect 13820 18896 13872 18902
rect 13820 18838 13872 18844
rect 13832 18426 13860 18838
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13924 18358 13952 19382
rect 13912 18352 13964 18358
rect 13912 18294 13964 18300
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 14016 17542 14044 20402
rect 14096 20256 14148 20262
rect 14096 20198 14148 20204
rect 14108 20058 14136 20198
rect 14096 20052 14148 20058
rect 14096 19994 14148 20000
rect 14200 19922 14228 22374
rect 14384 22234 14412 22578
rect 14464 22500 14516 22506
rect 14464 22442 14516 22448
rect 14372 22228 14424 22234
rect 14372 22170 14424 22176
rect 14476 22166 14504 22442
rect 14464 22160 14516 22166
rect 14464 22102 14516 22108
rect 14660 21554 14688 23666
rect 15396 23118 15424 24618
rect 15764 24274 15792 27520
rect 15752 24268 15804 24274
rect 15752 24210 15804 24216
rect 15764 23866 15792 24210
rect 15936 24132 15988 24138
rect 15936 24074 15988 24080
rect 15752 23860 15804 23866
rect 15752 23802 15804 23808
rect 15948 23730 15976 24074
rect 16212 24064 16264 24070
rect 16212 24006 16264 24012
rect 16304 24064 16356 24070
rect 16304 24006 16356 24012
rect 15936 23724 15988 23730
rect 15936 23666 15988 23672
rect 16120 23724 16172 23730
rect 16120 23666 16172 23672
rect 15752 23520 15804 23526
rect 15752 23462 15804 23468
rect 15476 23248 15528 23254
rect 15476 23190 15528 23196
rect 14832 23112 14884 23118
rect 14832 23054 14884 23060
rect 15384 23112 15436 23118
rect 15384 23054 15436 23060
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 14660 21146 14688 21490
rect 14648 21140 14700 21146
rect 14648 21082 14700 21088
rect 14844 21010 14872 23054
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15396 22234 15424 23054
rect 15488 22506 15516 23190
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15672 22642 15700 23054
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 15476 22500 15528 22506
rect 15476 22442 15528 22448
rect 15384 22228 15436 22234
rect 15384 22170 15436 22176
rect 15292 22160 15344 22166
rect 15292 22102 15344 22108
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15304 21146 15332 22102
rect 15488 21690 15516 22442
rect 15476 21684 15528 21690
rect 15476 21626 15528 21632
rect 15384 21344 15436 21350
rect 15384 21286 15436 21292
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15396 21078 15424 21286
rect 15384 21072 15436 21078
rect 15384 21014 15436 21020
rect 14832 21004 14884 21010
rect 14832 20946 14884 20952
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 14384 20398 14412 20742
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 14200 18630 14228 19858
rect 14384 19378 14412 20334
rect 14844 20058 14872 20946
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15396 20262 15424 21014
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15396 20058 15424 20198
rect 14832 20052 14884 20058
rect 14832 19994 14884 20000
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14740 19712 14792 19718
rect 14740 19654 14792 19660
rect 14752 19378 14780 19654
rect 14372 19372 14424 19378
rect 14740 19372 14792 19378
rect 14424 19320 14504 19334
rect 14372 19314 14504 19320
rect 14740 19314 14792 19320
rect 14384 19310 14504 19314
rect 14384 19306 14516 19310
rect 14464 19304 14516 19306
rect 14464 19246 14516 19252
rect 14554 19136 14610 19145
rect 14554 19071 14610 19080
rect 14568 18698 14596 19071
rect 14844 18970 14872 19790
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15396 19514 15424 19994
rect 15384 19508 15436 19514
rect 15384 19450 15436 19456
rect 14832 18964 14884 18970
rect 14832 18906 14884 18912
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14188 18624 14240 18630
rect 14188 18566 14240 18572
rect 14096 17740 14148 17746
rect 14200 17728 14228 18566
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14648 18216 14700 18222
rect 14648 18158 14700 18164
rect 14556 18148 14608 18154
rect 14556 18090 14608 18096
rect 14148 17700 14228 17728
rect 14096 17682 14148 17688
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 14108 16998 14136 17682
rect 14568 17066 14596 18090
rect 14660 17610 14688 18158
rect 15488 17746 15516 18702
rect 15568 18080 15620 18086
rect 15568 18022 15620 18028
rect 15476 17740 15528 17746
rect 15476 17682 15528 17688
rect 14648 17604 14700 17610
rect 14648 17546 14700 17552
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14740 17128 14792 17134
rect 14740 17070 14792 17076
rect 14556 17060 14608 17066
rect 14556 17002 14608 17008
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13544 16176 13596 16182
rect 13544 16118 13596 16124
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 13004 15706 13032 15982
rect 13648 15978 13676 16594
rect 14108 16522 14136 16934
rect 14752 16726 14780 17070
rect 14740 16720 14792 16726
rect 14740 16662 14792 16668
rect 14096 16516 14148 16522
rect 14096 16458 14148 16464
rect 14108 16250 14136 16458
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14096 16244 14148 16250
rect 14096 16186 14148 16192
rect 15580 16114 15608 18022
rect 15672 16590 15700 22578
rect 15764 22166 15792 23462
rect 16132 23118 16160 23666
rect 16224 23254 16252 24006
rect 16316 23322 16344 24006
rect 16304 23316 16356 23322
rect 16304 23258 16356 23264
rect 16212 23248 16264 23254
rect 16212 23190 16264 23196
rect 16120 23112 16172 23118
rect 16040 23072 16120 23100
rect 15752 22160 15804 22166
rect 15752 22102 15804 22108
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 15948 21690 15976 21966
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 15752 20256 15804 20262
rect 15752 20198 15804 20204
rect 15764 19786 15792 20198
rect 15752 19780 15804 19786
rect 15752 19722 15804 19728
rect 15764 18902 15792 19722
rect 15752 18896 15804 18902
rect 15752 18838 15804 18844
rect 15764 18086 15792 18838
rect 16040 18766 16068 23072
rect 16120 23054 16172 23060
rect 16316 22710 16344 23258
rect 16304 22704 16356 22710
rect 16304 22646 16356 22652
rect 16212 22636 16264 22642
rect 16212 22578 16264 22584
rect 16224 22166 16252 22578
rect 16212 22160 16264 22166
rect 16212 22102 16264 22108
rect 16224 20534 16252 22102
rect 16488 21888 16540 21894
rect 16488 21830 16540 21836
rect 16500 21486 16528 21830
rect 16580 21616 16632 21622
rect 16580 21558 16632 21564
rect 16488 21480 16540 21486
rect 16488 21422 16540 21428
rect 16212 20528 16264 20534
rect 16132 20488 16212 20516
rect 16132 19378 16160 20488
rect 16212 20470 16264 20476
rect 16212 19712 16264 19718
rect 16212 19654 16264 19660
rect 16224 19514 16252 19654
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 16120 19236 16172 19242
rect 16224 19224 16252 19450
rect 16172 19196 16252 19224
rect 16120 19178 16172 19184
rect 16028 18760 16080 18766
rect 16028 18702 16080 18708
rect 16040 18290 16068 18702
rect 16500 18408 16528 21422
rect 16592 21146 16620 21558
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 16592 20466 16620 21082
rect 16580 20460 16632 20466
rect 16580 20402 16632 20408
rect 16684 18698 16712 27526
rect 17038 27520 17094 27526
rect 18326 27554 18382 28000
rect 19614 27554 19670 28000
rect 18326 27526 18644 27554
rect 18326 27520 18382 27526
rect 18616 24274 18644 27526
rect 19352 27526 19670 27554
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 18604 24268 18656 24274
rect 18604 24210 18656 24216
rect 16960 23594 16988 24210
rect 17316 23860 17368 23866
rect 17316 23802 17368 23808
rect 16948 23588 17000 23594
rect 16948 23530 17000 23536
rect 17328 23254 17356 23802
rect 18616 23798 18644 24210
rect 18880 24064 18932 24070
rect 18880 24006 18932 24012
rect 18604 23792 18656 23798
rect 18604 23734 18656 23740
rect 17776 23656 17828 23662
rect 17776 23598 17828 23604
rect 16948 23248 17000 23254
rect 16948 23190 17000 23196
rect 17040 23248 17092 23254
rect 17040 23190 17092 23196
rect 17316 23248 17368 23254
rect 17316 23190 17368 23196
rect 16960 22778 16988 23190
rect 16948 22772 17000 22778
rect 16948 22714 17000 22720
rect 17052 22642 17080 23190
rect 17788 23089 17816 23598
rect 18892 23322 18920 24006
rect 19352 23866 19380 27526
rect 19614 27520 19670 27526
rect 20902 27520 20958 28000
rect 22098 27520 22154 28000
rect 23386 27520 23442 28000
rect 24674 27520 24730 28000
rect 24952 27532 25004 27538
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20352 24064 20404 24070
rect 20352 24006 20404 24012
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 19340 23656 19392 23662
rect 19340 23598 19392 23604
rect 18880 23316 18932 23322
rect 18880 23258 18932 23264
rect 18236 23248 18288 23254
rect 18236 23190 18288 23196
rect 17774 23080 17830 23089
rect 17774 23015 17830 23024
rect 18248 22778 18276 23190
rect 18328 22976 18380 22982
rect 18328 22918 18380 22924
rect 18236 22772 18288 22778
rect 18236 22714 18288 22720
rect 17040 22636 17092 22642
rect 17040 22578 17092 22584
rect 18340 22166 18368 22918
rect 18892 22710 18920 23258
rect 18880 22704 18932 22710
rect 18880 22646 18932 22652
rect 18972 22704 19024 22710
rect 18972 22646 19024 22652
rect 18328 22160 18380 22166
rect 18328 22102 18380 22108
rect 18420 22160 18472 22166
rect 18420 22102 18472 22108
rect 18052 21888 18104 21894
rect 18052 21830 18104 21836
rect 18064 21554 18092 21830
rect 18340 21690 18368 22102
rect 18432 21690 18460 22102
rect 18984 22030 19012 22646
rect 18972 22024 19024 22030
rect 18972 21966 19024 21972
rect 18328 21684 18380 21690
rect 18328 21626 18380 21632
rect 18420 21684 18472 21690
rect 18420 21626 18472 21632
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 17132 21412 17184 21418
rect 17132 21354 17184 21360
rect 16764 21004 16816 21010
rect 16764 20946 16816 20952
rect 17144 20992 17172 21354
rect 17776 21344 17828 21350
rect 17776 21286 17828 21292
rect 17224 21004 17276 21010
rect 17144 20964 17224 20992
rect 16776 20602 16804 20946
rect 17144 20602 17172 20964
rect 17224 20946 17276 20952
rect 16764 20596 16816 20602
rect 16764 20538 16816 20544
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 17144 19854 17172 20538
rect 17788 20262 17816 21286
rect 18432 21146 18460 21626
rect 18420 21140 18472 21146
rect 18420 21082 18472 21088
rect 17868 20936 17920 20942
rect 17868 20878 17920 20884
rect 18696 20936 18748 20942
rect 18696 20878 18748 20884
rect 17880 20466 17908 20878
rect 17868 20460 17920 20466
rect 17868 20402 17920 20408
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17788 20058 17816 20198
rect 17880 20058 17908 20402
rect 17776 20052 17828 20058
rect 17776 19994 17828 20000
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17592 19916 17644 19922
rect 17592 19858 17644 19864
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 17144 19514 17172 19790
rect 17132 19508 17184 19514
rect 17132 19450 17184 19456
rect 17604 19446 17632 19858
rect 17592 19440 17644 19446
rect 17592 19382 17644 19388
rect 17788 19310 17816 19994
rect 18708 19990 18736 20878
rect 18696 19984 18748 19990
rect 18696 19926 18748 19932
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17776 19304 17828 19310
rect 17776 19246 17828 19252
rect 16764 19236 16816 19242
rect 16764 19178 16816 19184
rect 16672 18692 16724 18698
rect 16672 18634 16724 18640
rect 16500 18380 16620 18408
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 16488 18284 16540 18290
rect 16488 18226 16540 18232
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 16224 17882 16252 18022
rect 16500 17882 16528 18226
rect 16212 17876 16264 17882
rect 16212 17818 16264 17824
rect 16488 17876 16540 17882
rect 16488 17818 16540 17824
rect 16028 17808 16080 17814
rect 16028 17750 16080 17756
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 15856 16726 15884 16934
rect 15844 16720 15896 16726
rect 15844 16662 15896 16668
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 15672 16182 15700 16526
rect 15856 16250 15884 16662
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15660 16176 15712 16182
rect 15660 16118 15712 16124
rect 15752 16176 15804 16182
rect 15752 16118 15804 16124
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15028 15978 15056 16050
rect 13636 15972 13688 15978
rect 13636 15914 13688 15920
rect 15016 15972 15068 15978
rect 15016 15914 15068 15920
rect 14832 15904 14884 15910
rect 14832 15846 14884 15852
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 14188 15632 14240 15638
rect 14188 15574 14240 15580
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 13188 15026 13216 15438
rect 13728 15360 13780 15366
rect 13728 15302 13780 15308
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 13176 15020 13228 15026
rect 13228 14980 13308 15008
rect 13176 14962 13228 14968
rect 12912 14550 12940 14962
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 12900 14544 12952 14550
rect 12900 14486 12952 14492
rect 12714 13832 12770 13841
rect 12714 13767 12770 13776
rect 12728 13734 12756 13767
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 13188 13530 13216 14826
rect 13280 14278 13308 14980
rect 13452 14612 13504 14618
rect 13452 14554 13504 14560
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13280 13938 13308 14214
rect 13464 14074 13492 14554
rect 13636 14408 13688 14414
rect 13740 14396 13768 15302
rect 13924 14822 13952 15438
rect 14002 15192 14058 15201
rect 14002 15127 14058 15136
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13688 14368 13768 14396
rect 13636 14350 13688 14356
rect 13740 14074 13768 14368
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13740 13814 13768 14010
rect 13924 13938 13952 14758
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 14016 13870 14044 15127
rect 14200 15094 14228 15574
rect 14844 15366 14872 15846
rect 15384 15632 15436 15638
rect 15304 15592 15384 15620
rect 14832 15360 14884 15366
rect 14832 15302 14884 15308
rect 14188 15088 14240 15094
rect 14188 15030 14240 15036
rect 14200 14006 14228 15030
rect 14188 14000 14240 14006
rect 14188 13942 14240 13948
rect 13556 13786 13768 13814
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13452 13456 13504 13462
rect 13452 13398 13504 13404
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12624 12640 12676 12646
rect 12438 12608 12494 12617
rect 12624 12582 12676 12588
rect 12438 12543 12494 12552
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11716 11898 11744 12242
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11808 11694 11836 12242
rect 12636 12170 12664 12582
rect 12728 12374 12756 13262
rect 13464 12646 13492 13398
rect 13556 12918 13584 13786
rect 14740 13456 14792 13462
rect 14740 13398 14792 13404
rect 14752 13297 14780 13398
rect 14738 13288 14794 13297
rect 14738 13223 14794 13232
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13544 12912 13596 12918
rect 13544 12854 13596 12860
rect 13924 12714 13952 13126
rect 14752 12986 14780 13223
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 14016 12714 14044 12922
rect 13912 12708 13964 12714
rect 13912 12650 13964 12656
rect 14004 12708 14056 12714
rect 14004 12650 14056 12656
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 12716 12368 12768 12374
rect 12716 12310 12768 12316
rect 12624 12164 12676 12170
rect 12624 12106 12676 12112
rect 12636 11830 12664 12106
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 12624 11824 12676 11830
rect 12624 11766 12676 11772
rect 13096 11762 13124 12038
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 13464 11626 13492 12582
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13740 11830 13768 12174
rect 13832 11898 13860 12310
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13452 11620 13504 11626
rect 13452 11562 13504 11568
rect 13464 11354 13492 11562
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 11428 11212 11480 11218
rect 11428 11154 11480 11160
rect 11440 10810 11468 11154
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11058 10704 11114 10713
rect 11058 10639 11114 10648
rect 11072 10606 11100 10639
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 12268 10198 12296 10950
rect 13464 10810 13492 11290
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 13004 10470 13032 10542
rect 13556 10470 13584 11086
rect 13648 10538 13676 11494
rect 13636 10532 13688 10538
rect 13636 10474 13688 10480
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 12256 10192 12308 10198
rect 12256 10134 12308 10140
rect 12716 10192 12768 10198
rect 12716 10134 12768 10140
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 12176 9382 12204 9998
rect 12728 9722 12756 10134
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12820 9586 12848 10406
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 10966 7984 11022 7993
rect 10966 7919 11022 7928
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 9692 4126 9812 4154
rect 8944 2848 8996 2854
rect 8944 2790 8996 2796
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 5540 2576 5592 2582
rect 8956 2553 8984 2790
rect 5540 2518 5592 2524
rect 8942 2544 8998 2553
rect 3146 54 3556 82
rect 5262 82 5318 480
rect 5552 82 5580 2518
rect 7380 2508 7432 2514
rect 8942 2479 8998 2488
rect 7380 2450 7432 2456
rect 7392 2310 7420 2450
rect 7380 2304 7432 2310
rect 7380 2246 7432 2252
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5262 54 5580 82
rect 7392 82 7420 2246
rect 7470 82 7526 480
rect 7392 54 7526 82
rect 9232 82 9260 2246
rect 9784 1873 9812 4126
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 12176 2650 12204 9318
rect 13004 9081 13032 10406
rect 13556 10198 13584 10406
rect 13740 10198 13768 11766
rect 13832 11354 13860 11834
rect 13924 11762 13952 12650
rect 14648 12300 14700 12306
rect 14648 12242 14700 12248
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 14108 11082 14136 12174
rect 14660 12073 14688 12242
rect 14646 12064 14702 12073
rect 14646 11999 14702 12008
rect 14660 11898 14688 11999
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14096 11076 14148 11082
rect 14096 11018 14148 11024
rect 14108 10742 14136 11018
rect 14752 10742 14780 11630
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 13924 10266 13952 10610
rect 14844 10266 14872 15302
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15108 15088 15160 15094
rect 15108 15030 15160 15036
rect 14924 14952 14976 14958
rect 14922 14920 14924 14929
rect 14976 14920 14978 14929
rect 14922 14855 14978 14864
rect 14936 14822 14964 14855
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 15120 14550 15148 15030
rect 15304 14822 15332 15592
rect 15384 15574 15436 15580
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15304 14550 15332 14758
rect 15396 14618 15424 15438
rect 15764 15178 15792 16118
rect 15948 16046 15976 17478
rect 16040 17066 16068 17750
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16316 17338 16344 17614
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 16028 17060 16080 17066
rect 16028 17002 16080 17008
rect 15936 16040 15988 16046
rect 15936 15982 15988 15988
rect 16488 16040 16540 16046
rect 16488 15982 16540 15988
rect 15844 15428 15896 15434
rect 15844 15370 15896 15376
rect 15580 15162 15792 15178
rect 15568 15156 15792 15162
rect 15620 15150 15792 15156
rect 15568 15098 15620 15104
rect 15580 15026 15608 15098
rect 15752 15088 15804 15094
rect 15752 15030 15804 15036
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15384 14612 15436 14618
rect 15384 14554 15436 14560
rect 15108 14544 15160 14550
rect 15108 14486 15160 14492
rect 15292 14544 15344 14550
rect 15292 14486 15344 14492
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 15304 13802 15332 13942
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14936 13297 14964 13330
rect 14922 13288 14978 13297
rect 14922 13223 14978 13232
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15304 11694 15332 13466
rect 15396 13326 15424 13670
rect 15384 13320 15436 13326
rect 15580 13297 15608 14350
rect 15384 13262 15436 13268
rect 15566 13288 15622 13297
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15304 11354 15332 11630
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15396 10810 15424 13262
rect 15566 13223 15622 13232
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15382 10568 15438 10577
rect 15580 10538 15608 11834
rect 15382 10503 15438 10512
rect 15476 10532 15528 10538
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 13544 10192 13596 10198
rect 13544 10134 13596 10140
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13820 10192 13872 10198
rect 13820 10134 13872 10140
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13372 9178 13400 9522
rect 13464 9450 13492 9658
rect 13452 9444 13504 9450
rect 13452 9386 13504 9392
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 12990 9072 13046 9081
rect 12990 9007 13046 9016
rect 13556 8498 13584 9658
rect 13832 9586 13860 10134
rect 15396 10130 15424 10503
rect 15476 10474 15528 10480
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15488 10266 15516 10474
rect 15476 10260 15528 10266
rect 15476 10202 15528 10208
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 14200 9722 14228 10066
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 15396 9450 15424 10066
rect 15384 9444 15436 9450
rect 15384 9386 15436 9392
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 15672 8401 15700 14962
rect 15764 14006 15792 15030
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15764 13326 15792 13942
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15764 10266 15792 11154
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15658 8392 15714 8401
rect 15658 8327 15714 8336
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14094 5128 14150 5137
rect 14094 5063 14150 5072
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 14108 2514 14136 5063
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14280 2848 14332 2854
rect 14280 2790 14332 2796
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 9770 1864 9826 1873
rect 9770 1799 9826 1808
rect 9586 82 9642 480
rect 9232 54 9642 82
rect 3146 0 3202 54
rect 5262 0 5318 54
rect 7470 0 7526 54
rect 9586 0 9642 54
rect 11702 128 11758 480
rect 11702 76 11704 128
rect 11756 76 11758 128
rect 11702 0 11758 76
rect 13910 82 13966 480
rect 14292 82 14320 2790
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15856 202 15884 15370
rect 16500 15366 16528 15982
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16212 14884 16264 14890
rect 16212 14826 16264 14832
rect 16028 14544 16080 14550
rect 16028 14486 16080 14492
rect 16040 13734 16068 14486
rect 16120 14340 16172 14346
rect 16120 14282 16172 14288
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 16040 13462 16068 13670
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 15936 13252 15988 13258
rect 15936 13194 15988 13200
rect 15948 12102 15976 13194
rect 16132 12918 16160 14282
rect 16120 12912 16172 12918
rect 16120 12854 16172 12860
rect 16224 12714 16252 14826
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 16304 13728 16356 13734
rect 16304 13670 16356 13676
rect 16212 12708 16264 12714
rect 16212 12650 16264 12656
rect 16316 12442 16344 13670
rect 16408 13190 16436 14418
rect 16500 13734 16528 15302
rect 16592 14482 16620 18380
rect 16776 18290 16804 19178
rect 17880 19174 17908 19790
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18512 19440 18564 19446
rect 18512 19382 18564 19388
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 17880 18834 17908 19110
rect 18064 18970 18092 19246
rect 18420 19236 18472 19242
rect 18420 19178 18472 19184
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 17868 18828 17920 18834
rect 17868 18770 17920 18776
rect 17880 18426 17908 18770
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 16672 17264 16724 17270
rect 16672 17206 16724 17212
rect 16684 15162 16712 17206
rect 16776 17134 16804 18226
rect 17236 17882 17264 18362
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17040 17740 17092 17746
rect 17040 17682 17092 17688
rect 17052 17649 17080 17682
rect 17038 17640 17094 17649
rect 17038 17575 17094 17584
rect 17052 17338 17080 17575
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16776 16794 16804 17070
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16764 15972 16816 15978
rect 16764 15914 16816 15920
rect 16672 15156 16724 15162
rect 16672 15098 16724 15104
rect 16684 14958 16712 15098
rect 16672 14952 16724 14958
rect 16672 14894 16724 14900
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16488 13728 16540 13734
rect 16488 13670 16540 13676
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 16488 12368 16540 12374
rect 16488 12310 16540 12316
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 15948 9722 15976 12038
rect 16500 11898 16528 12310
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16396 11620 16448 11626
rect 16396 11562 16448 11568
rect 16408 11286 16436 11562
rect 16396 11280 16448 11286
rect 16396 11222 16448 11228
rect 16408 10674 16436 11222
rect 16776 11218 16804 15914
rect 16868 15570 16896 16934
rect 17328 16658 17356 17138
rect 17880 16658 17908 18362
rect 17972 18086 18000 18702
rect 18432 18426 18460 19178
rect 18420 18420 18472 18426
rect 18420 18362 18472 18368
rect 18432 18154 18460 18362
rect 18420 18148 18472 18154
rect 18420 18090 18472 18096
rect 17960 18080 18012 18086
rect 17960 18022 18012 18028
rect 17316 16652 17368 16658
rect 17868 16652 17920 16658
rect 17316 16594 17368 16600
rect 17788 16612 17868 16640
rect 17132 15972 17184 15978
rect 17132 15914 17184 15920
rect 17144 15570 17172 15914
rect 17328 15706 17356 16594
rect 17788 16250 17816 16612
rect 17868 16594 17920 16600
rect 17868 16448 17920 16454
rect 17868 16390 17920 16396
rect 17776 16244 17828 16250
rect 17776 16186 17828 16192
rect 17880 16046 17908 16390
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 17132 15564 17184 15570
rect 17132 15506 17184 15512
rect 16868 15162 16896 15506
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 17144 14074 17172 14418
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 17696 13814 17724 15642
rect 17776 15564 17828 15570
rect 17776 15506 17828 15512
rect 17788 15162 17816 15506
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17880 14550 17908 15982
rect 17868 14544 17920 14550
rect 17868 14486 17920 14492
rect 17972 14385 18000 18022
rect 18432 17882 18460 18090
rect 18420 17876 18472 17882
rect 18420 17818 18472 17824
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 18156 17338 18184 17614
rect 18432 17338 18460 17818
rect 18144 17332 18196 17338
rect 18144 17274 18196 17280
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18052 17264 18104 17270
rect 18052 17206 18104 17212
rect 18064 17066 18092 17206
rect 18052 17060 18104 17066
rect 18052 17002 18104 17008
rect 18064 16250 18092 17002
rect 18156 16726 18184 17274
rect 18524 17066 18552 19382
rect 18616 18737 18644 19654
rect 18880 19508 18932 19514
rect 18880 19450 18932 19456
rect 18696 18760 18748 18766
rect 18602 18728 18658 18737
rect 18696 18702 18748 18708
rect 18602 18663 18658 18672
rect 18708 18290 18736 18702
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18512 17060 18564 17066
rect 18512 17002 18564 17008
rect 18524 16794 18552 17002
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18144 16720 18196 16726
rect 18144 16662 18196 16668
rect 18892 16658 18920 19450
rect 18984 18748 19012 21966
rect 19064 21140 19116 21146
rect 19064 21082 19116 21088
rect 19076 20330 19104 21082
rect 19064 20324 19116 20330
rect 19064 20266 19116 20272
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19168 19514 19196 19858
rect 19156 19508 19208 19514
rect 19156 19450 19208 19456
rect 19260 18970 19288 19994
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19156 18896 19208 18902
rect 19156 18838 19208 18844
rect 19064 18760 19116 18766
rect 18984 18720 19064 18748
rect 19064 18702 19116 18708
rect 19076 18358 19104 18702
rect 19064 18352 19116 18358
rect 19064 18294 19116 18300
rect 18972 17604 19024 17610
rect 18972 17546 19024 17552
rect 18984 16794 19012 17546
rect 19076 17270 19104 18294
rect 19168 17882 19196 18838
rect 19248 18760 19300 18766
rect 19352 18737 19380 23598
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 20364 22642 20392 24006
rect 20916 23866 20944 27520
rect 21454 25392 21510 25401
rect 21454 25327 21510 25336
rect 21468 24274 21496 25327
rect 21456 24268 21508 24274
rect 21456 24210 21508 24216
rect 21468 23866 21496 24210
rect 20904 23860 20956 23866
rect 20904 23802 20956 23808
rect 21456 23860 21508 23866
rect 21456 23802 21508 23808
rect 20904 23520 20956 23526
rect 20956 23480 21036 23508
rect 20904 23462 20956 23468
rect 21008 23118 21036 23480
rect 22112 23474 22140 27520
rect 22558 24168 22614 24177
rect 22558 24103 22614 24112
rect 21928 23446 22140 23474
rect 21364 23248 21416 23254
rect 21364 23190 21416 23196
rect 20996 23112 21048 23118
rect 20996 23054 21048 23060
rect 21272 23112 21324 23118
rect 21272 23054 21324 23060
rect 21008 22778 21036 23054
rect 21088 22976 21140 22982
rect 21088 22918 21140 22924
rect 20996 22772 21048 22778
rect 20996 22714 21048 22720
rect 20352 22636 20404 22642
rect 20352 22578 20404 22584
rect 19984 22500 20036 22506
rect 19984 22442 20036 22448
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19892 21956 19944 21962
rect 19892 21898 19944 21904
rect 19904 21554 19932 21898
rect 19892 21548 19944 21554
rect 19892 21490 19944 21496
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19536 21146 19564 21286
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19996 21146 20024 22442
rect 20364 22234 20392 22578
rect 20352 22228 20404 22234
rect 20352 22170 20404 22176
rect 20996 22160 21048 22166
rect 20996 22102 21048 22108
rect 21008 21690 21036 22102
rect 21100 22030 21128 22918
rect 21284 22642 21312 23054
rect 21376 22710 21404 23190
rect 21364 22704 21416 22710
rect 21364 22646 21416 22652
rect 21272 22636 21324 22642
rect 21272 22578 21324 22584
rect 21284 22030 21312 22578
rect 21088 22024 21140 22030
rect 21088 21966 21140 21972
rect 21272 22024 21324 22030
rect 21272 21966 21324 21972
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 20536 21412 20588 21418
rect 20536 21354 20588 21360
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 19524 21140 19576 21146
rect 19984 21140 20036 21146
rect 19524 21082 19576 21088
rect 19904 21100 19984 21128
rect 19904 20602 19932 21100
rect 19984 21082 20036 21088
rect 19984 20936 20036 20942
rect 19984 20878 20036 20884
rect 19892 20596 19944 20602
rect 19892 20538 19944 20544
rect 19904 20312 19932 20538
rect 19996 20466 20024 20878
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 19984 20324 20036 20330
rect 19904 20284 19984 20312
rect 19984 20266 20036 20272
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 20272 20058 20300 20402
rect 20260 20052 20312 20058
rect 20260 19994 20312 20000
rect 20272 19378 20300 19994
rect 20260 19372 20312 19378
rect 20260 19314 20312 19320
rect 19984 19236 20036 19242
rect 19984 19178 20036 19184
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19248 18702 19300 18708
rect 19338 18728 19394 18737
rect 19260 17921 19288 18702
rect 19338 18663 19394 18672
rect 19246 17912 19302 17921
rect 19156 17876 19208 17882
rect 19246 17847 19302 17856
rect 19156 17818 19208 17824
rect 19064 17264 19116 17270
rect 19064 17206 19116 17212
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 18880 16652 18932 16658
rect 18880 16594 18932 16600
rect 18892 16250 18920 16594
rect 18052 16244 18104 16250
rect 18880 16244 18932 16250
rect 18052 16186 18104 16192
rect 18800 16204 18880 16232
rect 18064 15960 18092 16186
rect 18144 15972 18196 15978
rect 18064 15932 18144 15960
rect 18144 15914 18196 15920
rect 18156 15638 18184 15914
rect 18144 15632 18196 15638
rect 18144 15574 18196 15580
rect 18156 15162 18184 15574
rect 18512 15360 18564 15366
rect 18512 15302 18564 15308
rect 18144 15156 18196 15162
rect 18196 15116 18276 15144
rect 18144 15098 18196 15104
rect 17958 14376 18014 14385
rect 17958 14311 18014 14320
rect 18052 13864 18104 13870
rect 17696 13786 17816 13814
rect 18052 13806 18104 13812
rect 17132 13388 17184 13394
rect 17132 13330 17184 13336
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17144 12986 17172 13330
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17512 12646 17540 13330
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 16868 11898 16896 12174
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16960 11830 16988 12106
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 16764 11212 16816 11218
rect 16764 11154 16816 11160
rect 16672 11008 16724 11014
rect 16672 10950 16724 10956
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 16684 10198 16712 10950
rect 16672 10192 16724 10198
rect 16672 10134 16724 10140
rect 16684 9722 16712 10134
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 15936 9716 15988 9722
rect 15936 9658 15988 9664
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16776 9382 16804 9998
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16868 5273 16896 11630
rect 16960 10062 16988 11766
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17604 10266 17632 11154
rect 17788 10810 17816 13786
rect 18064 13462 18092 13806
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 17972 11218 18000 12582
rect 18156 12306 18184 13670
rect 18248 13530 18276 15116
rect 18524 15026 18552 15302
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18616 14890 18644 14962
rect 18604 14884 18656 14890
rect 18604 14826 18656 14832
rect 18616 14618 18644 14826
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18432 13870 18460 14214
rect 18420 13864 18472 13870
rect 18420 13806 18472 13812
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18432 13326 18460 13806
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 18144 12300 18196 12306
rect 18144 12242 18196 12248
rect 18156 11898 18184 12242
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17776 10804 17828 10810
rect 17776 10746 17828 10752
rect 17788 10713 17816 10746
rect 17972 10742 18000 11154
rect 17960 10736 18012 10742
rect 17774 10704 17830 10713
rect 17960 10678 18012 10684
rect 17774 10639 17830 10648
rect 17788 10606 17816 10639
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 17960 10532 18012 10538
rect 17960 10474 18012 10480
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16854 5264 16910 5273
rect 16854 5199 16910 5208
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 15844 196 15896 202
rect 15844 138 15896 144
rect 13910 54 14320 82
rect 16026 82 16082 480
rect 16132 82 16160 2314
rect 16026 54 16160 82
rect 17972 82 18000 10474
rect 18156 10266 18184 10542
rect 18340 10470 18368 12718
rect 18524 11762 18552 14214
rect 18800 14074 18828 16204
rect 18880 16186 18932 16192
rect 18880 15904 18932 15910
rect 18880 15846 18932 15852
rect 18892 14550 18920 15846
rect 19064 15428 19116 15434
rect 19064 15370 19116 15376
rect 18880 14544 18932 14550
rect 18880 14486 18932 14492
rect 18892 14074 18920 14486
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 18696 13456 18748 13462
rect 19076 13433 19104 15370
rect 19156 14884 19208 14890
rect 19156 14826 19208 14832
rect 19168 14414 19196 14826
rect 19156 14408 19208 14414
rect 19156 14350 19208 14356
rect 19168 13802 19196 14350
rect 19352 14278 19380 18663
rect 19996 18630 20024 19178
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19996 18426 20024 18566
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19444 17338 19472 17478
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19982 16688 20038 16697
rect 19708 16652 19760 16658
rect 20088 16674 20116 19110
rect 20168 18896 20220 18902
rect 20168 18838 20220 18844
rect 20038 16646 20116 16674
rect 19982 16623 20038 16632
rect 19708 16594 19760 16600
rect 19720 16454 19748 16594
rect 19708 16448 19760 16454
rect 19708 16390 19760 16396
rect 19720 16250 19748 16390
rect 19708 16244 19760 16250
rect 19708 16186 19760 16192
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19536 14618 19564 14758
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19996 13814 20024 16623
rect 20076 15700 20128 15706
rect 20076 15642 20128 15648
rect 20088 14890 20116 15642
rect 20180 15570 20208 18838
rect 20272 18290 20300 19314
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 20168 15564 20220 15570
rect 20220 15524 20300 15552
rect 20168 15506 20220 15512
rect 20168 15360 20220 15366
rect 20168 15302 20220 15308
rect 20076 14884 20128 14890
rect 20076 14826 20128 14832
rect 20088 14550 20116 14826
rect 20180 14550 20208 15302
rect 20076 14544 20128 14550
rect 20076 14486 20128 14492
rect 20168 14544 20220 14550
rect 20168 14486 20220 14492
rect 20272 14482 20300 15524
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 19156 13796 19208 13802
rect 19996 13786 20208 13814
rect 19156 13738 19208 13744
rect 18696 13398 18748 13404
rect 19062 13424 19118 13433
rect 18708 12646 18736 13398
rect 19062 13359 19118 13368
rect 19168 13190 19196 13738
rect 19432 13728 19484 13734
rect 19432 13670 19484 13676
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19156 13184 19208 13190
rect 19156 13126 19208 13132
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18708 12374 18736 12582
rect 18696 12368 18748 12374
rect 18696 12310 18748 12316
rect 18708 11898 18736 12310
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18512 11756 18564 11762
rect 18512 11698 18564 11704
rect 18512 11620 18564 11626
rect 18512 11562 18564 11568
rect 18604 11620 18656 11626
rect 18604 11562 18656 11568
rect 18524 11354 18552 11562
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 18616 11286 18644 11562
rect 18604 11280 18656 11286
rect 18604 11222 18656 11228
rect 19076 11218 19104 12038
rect 19168 11762 19196 13126
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19260 11898 19288 12038
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 19156 11756 19208 11762
rect 19156 11698 19208 11704
rect 19260 11626 19288 11834
rect 19248 11620 19300 11626
rect 19248 11562 19300 11568
rect 19352 11218 19380 13262
rect 19444 12986 19472 13670
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19996 13394 20024 13670
rect 19524 13388 19576 13394
rect 19524 13330 19576 13336
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19536 12442 19564 13330
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19524 12436 19576 12442
rect 19524 12378 19576 12384
rect 20088 12102 20116 12718
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19064 11212 19116 11218
rect 19064 11154 19116 11160
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19076 10810 19104 11154
rect 19352 10810 19380 11154
rect 19536 10810 19564 11290
rect 20088 11286 20116 12038
rect 20076 11280 20128 11286
rect 20076 11222 20128 11228
rect 19064 10804 19116 10810
rect 19064 10746 19116 10752
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19352 10606 19380 10746
rect 19340 10600 19392 10606
rect 19340 10542 19392 10548
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 19444 9654 19472 10542
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19246 9072 19302 9081
rect 19246 9007 19302 9016
rect 19260 2854 19288 9007
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 19260 2582 19288 2790
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19248 2576 19300 2582
rect 18878 2544 18934 2553
rect 19248 2518 19300 2524
rect 18878 2479 18934 2488
rect 18892 2446 18920 2479
rect 18880 2440 18932 2446
rect 20180 2417 20208 13786
rect 20258 12200 20314 12209
rect 20258 12135 20314 12144
rect 20272 10810 20300 12135
rect 20260 10804 20312 10810
rect 20260 10746 20312 10752
rect 20364 9625 20392 16934
rect 20456 16114 20484 21286
rect 20548 19378 20576 21354
rect 21008 20602 21036 21626
rect 21100 21146 21128 21966
rect 21088 21140 21140 21146
rect 21088 21082 21140 21088
rect 20996 20596 21048 20602
rect 20996 20538 21048 20544
rect 21270 20360 21326 20369
rect 21270 20295 21326 20304
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20548 18902 20576 19314
rect 20824 19174 20852 19858
rect 21284 19378 21312 20295
rect 21376 19446 21404 22646
rect 21928 21690 21956 23446
rect 22572 23186 22600 24103
rect 23400 23594 23428 27520
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24688 23866 24716 27520
rect 25962 27532 26018 28000
rect 25962 27520 25964 27532
rect 24952 27474 25004 27480
rect 26016 27520 26018 27532
rect 27250 27520 27306 28000
rect 25964 27474 26016 27480
rect 24676 23860 24728 23866
rect 24676 23802 24728 23808
rect 23388 23588 23440 23594
rect 23388 23530 23440 23536
rect 22744 23520 22796 23526
rect 22744 23462 22796 23468
rect 22560 23180 22612 23186
rect 22560 23122 22612 23128
rect 22572 22778 22600 23122
rect 22560 22772 22612 22778
rect 22560 22714 22612 22720
rect 21916 21684 21968 21690
rect 21916 21626 21968 21632
rect 21928 21486 21956 21626
rect 21916 21480 21968 21486
rect 21916 21422 21968 21428
rect 21640 20596 21692 20602
rect 21640 20538 21692 20544
rect 21652 20330 21680 20538
rect 21548 20324 21600 20330
rect 21548 20266 21600 20272
rect 21640 20324 21692 20330
rect 21640 20266 21692 20272
rect 21560 20058 21588 20266
rect 21548 20052 21600 20058
rect 21548 19994 21600 20000
rect 21364 19440 21416 19446
rect 21364 19382 21416 19388
rect 21272 19372 21324 19378
rect 21272 19314 21324 19320
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 20536 18896 20588 18902
rect 20536 18838 20588 18844
rect 21376 18154 21404 19382
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 21916 19168 21968 19174
rect 21916 19110 21968 19116
rect 21822 18864 21878 18873
rect 21822 18799 21878 18808
rect 21732 18692 21784 18698
rect 21732 18634 21784 18640
rect 20536 18148 20588 18154
rect 20536 18090 20588 18096
rect 21364 18148 21416 18154
rect 21364 18090 21416 18096
rect 20548 17882 20576 18090
rect 20536 17876 20588 17882
rect 20536 17818 20588 17824
rect 20548 17338 20576 17818
rect 20628 17740 20680 17746
rect 20628 17682 20680 17688
rect 21364 17740 21416 17746
rect 21364 17682 21416 17688
rect 20640 17338 20668 17682
rect 20536 17332 20588 17338
rect 20536 17274 20588 17280
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 21376 17241 21404 17682
rect 21362 17232 21418 17241
rect 21362 17167 21418 17176
rect 21376 17134 21404 17167
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 21272 16652 21324 16658
rect 21272 16594 21324 16600
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20456 15706 20484 16050
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20640 15094 20668 16050
rect 21284 15910 21312 16594
rect 21744 16046 21772 18634
rect 21836 16658 21864 18799
rect 21928 17785 21956 19110
rect 21914 17776 21970 17785
rect 21914 17711 21970 17720
rect 21824 16652 21876 16658
rect 21824 16594 21876 16600
rect 21836 16250 21864 16594
rect 21916 16448 21968 16454
rect 21916 16390 21968 16396
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 21732 16040 21784 16046
rect 21732 15982 21784 15988
rect 21364 15972 21416 15978
rect 21364 15914 21416 15920
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21088 15632 21140 15638
rect 21088 15574 21140 15580
rect 21180 15632 21232 15638
rect 21284 15609 21312 15846
rect 21180 15574 21232 15580
rect 21270 15600 21326 15609
rect 21100 15162 21128 15574
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 20628 15088 20680 15094
rect 20628 15030 20680 15036
rect 20640 13462 20668 15030
rect 21100 14890 21128 15098
rect 21192 15026 21220 15574
rect 21270 15535 21326 15544
rect 21376 15162 21404 15914
rect 21364 15156 21416 15162
rect 21364 15098 21416 15104
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 21376 14890 21404 15098
rect 21088 14884 21140 14890
rect 21088 14826 21140 14832
rect 21364 14884 21416 14890
rect 21364 14826 21416 14832
rect 21640 14816 21692 14822
rect 21640 14758 21692 14764
rect 20996 14476 21048 14482
rect 20996 14418 21048 14424
rect 21008 14074 21036 14418
rect 21548 14272 21600 14278
rect 21548 14214 21600 14220
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 21560 14006 21588 14214
rect 21548 14000 21600 14006
rect 21548 13942 21600 13948
rect 20812 13932 20864 13938
rect 20812 13874 20864 13880
rect 20628 13456 20680 13462
rect 20628 13398 20680 13404
rect 20640 12442 20668 13398
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 20824 10538 20852 13874
rect 21560 13870 21588 13942
rect 21548 13864 21600 13870
rect 21548 13806 21600 13812
rect 21180 13796 21232 13802
rect 21180 13738 21232 13744
rect 21192 13326 21220 13738
rect 21272 13456 21324 13462
rect 21272 13398 21324 13404
rect 21456 13456 21508 13462
rect 21456 13398 21508 13404
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 21192 12918 21220 13262
rect 21284 12986 21312 13398
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21180 12912 21232 12918
rect 21180 12854 21232 12860
rect 21088 12368 21140 12374
rect 21088 12310 21140 12316
rect 21100 11898 21128 12310
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 21100 11626 21128 11834
rect 21088 11620 21140 11626
rect 21088 11562 21140 11568
rect 21376 11558 21404 12174
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 20916 11354 20944 11494
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 20812 10532 20864 10538
rect 20812 10474 20864 10480
rect 20916 10470 20944 11154
rect 20904 10464 20956 10470
rect 20904 10406 20956 10412
rect 20350 9616 20406 9625
rect 20350 9551 20406 9560
rect 20916 9081 20944 10406
rect 20902 9072 20958 9081
rect 20902 9007 20958 9016
rect 21376 2650 21404 11494
rect 21468 9450 21496 13398
rect 21652 13297 21680 14758
rect 21744 14482 21772 15982
rect 21928 15706 21956 16390
rect 21916 15700 21968 15706
rect 21916 15642 21968 15648
rect 21928 15026 21956 15642
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 22020 15026 22048 15438
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 21732 14476 21784 14482
rect 21732 14418 21784 14424
rect 21730 14376 21786 14385
rect 21730 14311 21786 14320
rect 21744 14278 21772 14311
rect 21732 14272 21784 14278
rect 21732 14214 21784 14220
rect 21744 13802 21772 14214
rect 22020 13814 22048 14962
rect 22112 14929 22140 19246
rect 22652 16992 22704 16998
rect 22652 16934 22704 16940
rect 22664 15434 22692 16934
rect 22652 15428 22704 15434
rect 22652 15370 22704 15376
rect 22664 15162 22692 15370
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22098 14920 22154 14929
rect 22098 14855 22154 14864
rect 22112 14657 22140 14855
rect 22098 14648 22154 14657
rect 22098 14583 22154 14592
rect 22100 14476 22152 14482
rect 22100 14418 22152 14424
rect 21732 13796 21784 13802
rect 21732 13738 21784 13744
rect 21928 13786 22048 13814
rect 21638 13288 21694 13297
rect 21638 13223 21694 13232
rect 21928 12714 21956 13786
rect 22112 13734 22140 14418
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22112 13462 22140 13670
rect 22100 13456 22152 13462
rect 22100 13398 22152 13404
rect 22008 12912 22060 12918
rect 22008 12854 22060 12860
rect 21916 12708 21968 12714
rect 21916 12650 21968 12656
rect 21928 12102 21956 12650
rect 21916 12096 21968 12102
rect 21916 12038 21968 12044
rect 21928 11762 21956 12038
rect 22020 11898 22048 12854
rect 22756 12170 22784 23462
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24030 18728 24086 18737
rect 24030 18663 24086 18672
rect 23664 16244 23716 16250
rect 23664 16186 23716 16192
rect 23676 15570 23704 16186
rect 23664 15564 23716 15570
rect 23664 15506 23716 15512
rect 22928 14476 22980 14482
rect 22928 14418 22980 14424
rect 22940 13938 22968 14418
rect 22928 13932 22980 13938
rect 22928 13874 22980 13880
rect 22744 12164 22796 12170
rect 22744 12106 22796 12112
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 21916 11756 21968 11762
rect 21916 11698 21968 11704
rect 22020 11694 22048 11834
rect 22008 11688 22060 11694
rect 22008 11630 22060 11636
rect 21916 11552 21968 11558
rect 21916 11494 21968 11500
rect 21928 11218 21956 11494
rect 21916 11212 21968 11218
rect 21916 11154 21968 11160
rect 24044 10606 24072 18663
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24766 17368 24822 17377
rect 24766 17303 24822 17312
rect 24780 16794 24808 17303
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 24676 16652 24728 16658
rect 24676 16594 24728 16600
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24688 16250 24716 16594
rect 24676 16244 24728 16250
rect 24676 16186 24728 16192
rect 24124 16040 24176 16046
rect 24124 15982 24176 15988
rect 24766 16008 24822 16017
rect 24136 15473 24164 15982
rect 24766 15943 24822 15952
rect 24780 15706 24808 15943
rect 24768 15700 24820 15706
rect 24768 15642 24820 15648
rect 24216 15564 24268 15570
rect 24216 15506 24268 15512
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24122 15464 24178 15473
rect 24122 15399 24178 15408
rect 24124 14476 24176 14482
rect 24124 14418 24176 14424
rect 24136 13734 24164 14418
rect 24124 13728 24176 13734
rect 24124 13670 24176 13676
rect 24136 12617 24164 13670
rect 24122 12608 24178 12617
rect 24122 12543 24178 12552
rect 24228 11370 24256 15506
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24688 15162 24716 15506
rect 24964 15162 24992 27474
rect 25976 27443 26004 27474
rect 27264 23866 27292 27520
rect 27618 27296 27674 27305
rect 27618 27231 27674 27240
rect 27632 25362 27660 27231
rect 27620 25356 27672 25362
rect 27620 25298 27672 25304
rect 27252 23860 27304 23866
rect 27252 23802 27304 23808
rect 25134 22672 25190 22681
rect 25134 22607 25190 22616
rect 25148 21690 25176 22607
rect 25136 21684 25188 21690
rect 25136 21626 25188 21632
rect 25148 21486 25176 21626
rect 25136 21480 25188 21486
rect 25136 21422 25188 21428
rect 25502 21312 25558 21321
rect 25502 21247 25558 21256
rect 25134 20088 25190 20097
rect 25134 20023 25190 20032
rect 25148 19514 25176 20023
rect 25516 19922 25544 21247
rect 25504 19916 25556 19922
rect 25504 19858 25556 19864
rect 25516 19514 25544 19858
rect 25136 19508 25188 19514
rect 25136 19450 25188 19456
rect 25504 19508 25556 19514
rect 25504 19450 25556 19456
rect 25148 19310 25176 19450
rect 25136 19304 25188 19310
rect 25136 19246 25188 19252
rect 25134 18728 25190 18737
rect 25134 18663 25190 18672
rect 25148 17338 25176 18663
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 25148 17134 25176 17274
rect 25136 17128 25188 17134
rect 25136 17070 25188 17076
rect 24676 15156 24728 15162
rect 24676 15098 24728 15104
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 24964 14958 24992 15098
rect 24952 14952 25004 14958
rect 24952 14894 25004 14900
rect 25410 14784 25466 14793
rect 25410 14719 25466 14728
rect 25424 14618 25452 14719
rect 25412 14612 25464 14618
rect 25412 14554 25464 14560
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 26424 12640 26476 12646
rect 26424 12582 26476 12588
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24136 11342 24256 11370
rect 24032 10600 24084 10606
rect 24032 10542 24084 10548
rect 21730 9616 21786 9625
rect 21730 9551 21786 9560
rect 21456 9444 21508 9450
rect 21456 9386 21508 9392
rect 21364 2644 21416 2650
rect 21364 2586 21416 2592
rect 18880 2382 18932 2388
rect 20166 2408 20222 2417
rect 20076 2372 20128 2378
rect 20166 2343 20222 2352
rect 20076 2314 20128 2320
rect 18234 82 18290 480
rect 17972 54 18290 82
rect 20088 82 20116 2314
rect 21468 1193 21496 9386
rect 21744 9042 21772 9551
rect 21732 9036 21784 9042
rect 21732 8978 21784 8984
rect 24136 5778 24164 11342
rect 24216 11212 24268 11218
rect 24216 11154 24268 11160
rect 24228 10810 24256 11154
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24766 10840 24822 10849
rect 24216 10804 24268 10810
rect 24766 10775 24822 10784
rect 24216 10746 24268 10752
rect 24780 10742 24808 10775
rect 24768 10736 24820 10742
rect 24768 10678 24820 10684
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 25136 9376 25188 9382
rect 24766 9344 24822 9353
rect 25136 9318 25188 9324
rect 24766 9279 24822 9288
rect 24780 9178 24808 9279
rect 24768 9172 24820 9178
rect 24768 9114 24820 9120
rect 25148 9081 25176 9318
rect 25134 9072 25190 9081
rect 24676 9036 24728 9042
rect 25134 9007 25190 9016
rect 24676 8978 24728 8984
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24688 8634 24716 8978
rect 24676 8628 24728 8634
rect 24676 8570 24728 8576
rect 24214 7848 24270 7857
rect 24214 7783 24270 7792
rect 24228 7342 24256 7783
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24216 7336 24268 7342
rect 24216 7278 24268 7284
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24124 5772 24176 5778
rect 24124 5714 24176 5720
rect 24676 5772 24728 5778
rect 24676 5714 24728 5720
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 5370 24716 5714
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24950 2816 25006 2825
rect 24950 2751 25006 2760
rect 24964 2650 24992 2751
rect 24952 2644 25004 2650
rect 24952 2586 25004 2592
rect 24768 2440 24820 2446
rect 24768 2382 24820 2388
rect 22100 2304 22152 2310
rect 22100 2246 22152 2252
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 21454 1184 21510 1193
rect 21454 1119 21510 1128
rect 20350 82 20406 480
rect 20088 54 20406 82
rect 22112 82 22140 2246
rect 22204 1873 22232 2246
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 22190 1864 22246 1873
rect 22190 1799 22246 1808
rect 22466 82 22522 480
rect 22112 54 22522 82
rect 13910 0 13966 54
rect 16026 0 16082 54
rect 18234 0 18290 54
rect 20350 0 20406 54
rect 22466 0 22522 54
rect 24674 82 24730 480
rect 24780 82 24808 2382
rect 24674 54 24808 82
rect 26436 82 26464 12582
rect 27712 11008 27764 11014
rect 27712 10950 27764 10956
rect 27620 7472 27672 7478
rect 27620 7414 27672 7420
rect 27632 7313 27660 7414
rect 27618 7304 27674 7313
rect 27618 7239 27674 7248
rect 27618 5944 27674 5953
rect 27540 5914 27618 5930
rect 27528 5908 27618 5914
rect 27580 5902 27618 5908
rect 27618 5879 27674 5888
rect 27528 5850 27580 5856
rect 27724 4593 27752 10950
rect 27710 4584 27766 4593
rect 27710 4519 27766 4528
rect 26790 82 26846 480
rect 26436 54 26846 82
rect 24674 0 24730 54
rect 26790 0 26846 54
<< via2 >>
rect 110 24248 166 24304
rect 110 21120 166 21176
rect 18 20032 74 20088
rect 1582 21664 1638 21720
rect 2318 26832 2374 26888
rect 1858 24792 1914 24848
rect 1674 19352 1730 19408
rect 1490 18128 1546 18184
rect 110 3440 166 3496
rect 1766 19216 1822 19272
rect 1582 15408 1638 15464
rect 1122 14320 1178 14376
rect 2226 23432 2282 23488
rect 846 7928 902 7984
rect 1398 9152 1454 9208
rect 1582 9016 1638 9072
rect 1766 12280 1822 12336
rect 1858 10240 1914 10296
rect 1490 7928 1546 7984
rect 1582 6840 1638 6896
rect 3146 25744 3202 25800
rect 3054 15544 3110 15600
rect 1858 3032 1914 3088
rect 3790 19352 3846 19408
rect 2318 8336 2374 8392
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5998 22888 6054 22944
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 4250 13368 4306 13424
rect 3698 9560 3754 9616
rect 2042 1944 2098 2000
rect 1306 992 1362 1048
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5078 13368 5134 13424
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 6826 15136 6882 15192
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 7378 17584 7434 17640
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 8022 18808 8078 18864
rect 10414 23024 10470 23080
rect 7838 18264 7894 18320
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 7470 12008 7526 12064
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5446 5344 5502 5400
rect 5446 5072 5502 5128
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 9310 19216 9366 19272
rect 8942 18128 8998 18184
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 8942 16632 8998 16688
rect 9310 15408 9366 15464
rect 8666 11464 8722 11520
rect 8666 7792 8722 7848
rect 8574 5072 8630 5128
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10874 18808 10930 18864
rect 10782 18672 10838 18728
rect 11518 18264 11574 18320
rect 13542 24112 13598 24168
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10690 13776 10746 13832
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 9862 13232 9918 13288
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10966 12552 11022 12608
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 12530 20304 12586 20360
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 15198 24112 15254 24168
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14094 23432 14150 23488
rect 14370 22888 14426 22944
rect 13634 19080 13690 19136
rect 13542 17856 13598 17912
rect 12990 17720 13046 17776
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14554 19080 14610 19136
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 17774 23024 17830 23080
rect 12714 13776 12770 13832
rect 14002 15136 14058 15192
rect 12438 12552 12494 12608
rect 14738 13232 14794 13288
rect 11058 10648 11114 10704
rect 10966 7928 11022 7984
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 8942 2488 8998 2544
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 14646 12008 14702 12064
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14922 14900 14924 14920
rect 14924 14900 14976 14920
rect 14976 14900 14978 14920
rect 14922 14864 14978 14900
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14922 13232 14978 13288
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15566 13232 15622 13288
rect 15382 10512 15438 10568
rect 12990 9016 13046 9072
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15658 8336 15714 8392
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14094 5072 14150 5128
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 9770 1808 9826 1864
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 17038 17584 17094 17640
rect 18602 18672 18658 18728
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 21454 25336 21510 25392
rect 22558 24112 22614 24168
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19338 18672 19394 18728
rect 19246 17856 19302 17912
rect 17958 14320 18014 14376
rect 17774 10648 17830 10704
rect 16854 5208 16910 5264
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19982 16632 20038 16688
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19062 13368 19118 13424
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19246 9016 19302 9072
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 18878 2488 18934 2544
rect 20258 12144 20314 12200
rect 21270 20304 21326 20360
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 21822 18808 21878 18864
rect 21362 17176 21418 17232
rect 21914 17720 21970 17776
rect 21270 15544 21326 15600
rect 20350 9560 20406 9616
rect 20902 9016 20958 9072
rect 21730 14320 21786 14376
rect 22098 14864 22154 14920
rect 22098 14592 22154 14648
rect 21638 13232 21694 13288
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24030 18672 24086 18728
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24766 17312 24822 17368
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24766 15952 24822 16008
rect 24122 15408 24178 15464
rect 24122 12552 24178 12608
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 27618 27240 27674 27296
rect 25134 22616 25190 22672
rect 25502 21256 25558 21312
rect 25134 20032 25190 20088
rect 25134 18672 25190 18728
rect 25410 14728 25466 14784
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 21730 9560 21786 9616
rect 20166 2352 20222 2408
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24766 10784 24822 10840
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24766 9288 24822 9344
rect 25134 9016 25190 9072
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24214 7792 24270 7848
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24950 2760 25006 2816
rect 21454 1128 21510 1184
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 22190 1808 22246 1864
rect 27618 7248 27674 7304
rect 27618 5888 27674 5944
rect 27710 4528 27766 4584
<< metal3 >>
rect 0 27344 480 27464
rect 62 26890 122 27344
rect 27520 27296 28000 27328
rect 27520 27240 27618 27296
rect 27674 27240 28000 27296
rect 27520 27208 28000 27240
rect 2313 26890 2379 26893
rect 62 26888 2379 26890
rect 62 26832 2318 26888
rect 2374 26832 2379 26888
rect 62 26830 2379 26832
rect 2313 26827 2379 26830
rect 0 26256 480 26376
rect 62 25802 122 26256
rect 27520 25848 28000 25968
rect 3141 25802 3207 25805
rect 62 25800 3207 25802
rect 62 25744 3146 25800
rect 3202 25744 3207 25800
rect 62 25742 3207 25744
rect 3141 25739 3207 25742
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25304 480 25424
rect 21449 25394 21515 25397
rect 27662 25394 27722 25848
rect 21449 25392 27722 25394
rect 21449 25336 21454 25392
rect 21510 25336 27722 25392
rect 21449 25334 27722 25336
rect 21449 25331 21515 25334
rect 62 24850 122 25304
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 1853 24850 1919 24853
rect 62 24848 1919 24850
rect 62 24792 1858 24848
rect 1914 24792 1919 24848
rect 62 24790 1919 24792
rect 1853 24787 1919 24790
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 27520 24488 28000 24608
rect 19610 24447 19930 24448
rect 0 24304 480 24336
rect 0 24248 110 24304
rect 166 24248 480 24304
rect 0 24216 480 24248
rect 13537 24170 13603 24173
rect 15193 24170 15259 24173
rect 13537 24168 15259 24170
rect 13537 24112 13542 24168
rect 13598 24112 15198 24168
rect 15254 24112 15259 24168
rect 13537 24110 15259 24112
rect 13537 24107 13603 24110
rect 15193 24107 15259 24110
rect 22553 24170 22619 24173
rect 27662 24170 27722 24488
rect 22553 24168 27722 24170
rect 22553 24112 22558 24168
rect 22614 24112 27722 24168
rect 22553 24110 27722 24112
rect 22553 24107 22619 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 2221 23490 2287 23493
rect 62 23488 2287 23490
rect 62 23432 2226 23488
rect 2282 23432 2287 23488
rect 62 23430 2287 23432
rect 62 23248 122 23430
rect 2221 23427 2287 23430
rect 14089 23490 14155 23493
rect 14590 23490 14596 23492
rect 14089 23488 14596 23490
rect 14089 23432 14094 23488
rect 14150 23432 14596 23488
rect 14089 23430 14596 23432
rect 14089 23427 14155 23430
rect 14590 23428 14596 23430
rect 14660 23428 14666 23492
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 0 23128 480 23248
rect 27520 23128 28000 23248
rect 10409 23082 10475 23085
rect 17769 23082 17835 23085
rect 10409 23080 17835 23082
rect 10409 23024 10414 23080
rect 10470 23024 17774 23080
rect 17830 23024 17835 23080
rect 10409 23022 17835 23024
rect 10409 23019 10475 23022
rect 17769 23019 17835 23022
rect 5993 22946 6059 22949
rect 14365 22946 14431 22949
rect 5993 22944 14431 22946
rect 5993 22888 5998 22944
rect 6054 22888 14370 22944
rect 14426 22888 14431 22944
rect 5993 22886 14431 22888
rect 5993 22883 6059 22886
rect 14365 22883 14431 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 25129 22674 25195 22677
rect 27662 22674 27722 23128
rect 25129 22672 27722 22674
rect 25129 22616 25134 22672
rect 25190 22616 27722 22672
rect 25129 22614 27722 22616
rect 25129 22611 25195 22614
rect 10277 22336 10597 22337
rect 0 22176 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 62 21722 122 22176
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 27520 21768 28000 21888
rect 24277 21727 24597 21728
rect 1577 21722 1643 21725
rect 62 21720 1643 21722
rect 62 21664 1582 21720
rect 1638 21664 1643 21720
rect 62 21662 1643 21664
rect 1577 21659 1643 21662
rect 25497 21314 25563 21317
rect 27662 21314 27722 21768
rect 25497 21312 27722 21314
rect 25497 21256 25502 21312
rect 25558 21256 27722 21312
rect 25497 21254 27722 21256
rect 25497 21251 25563 21254
rect 10277 21248 10597 21249
rect 0 21176 480 21208
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 0 21120 110 21176
rect 166 21120 480 21176
rect 0 21088 480 21120
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 27520 20544 28000 20664
rect 12525 20362 12591 20365
rect 21265 20362 21331 20365
rect 12525 20360 21331 20362
rect 12525 20304 12530 20360
rect 12586 20304 21270 20360
rect 21326 20304 21331 20360
rect 12525 20302 21331 20304
rect 12525 20299 12591 20302
rect 21265 20299 21331 20302
rect 10277 20160 10597 20161
rect 0 20088 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 0 20032 18 20088
rect 74 20032 480 20088
rect 0 20000 480 20032
rect 25129 20090 25195 20093
rect 27662 20090 27722 20544
rect 25129 20088 27722 20090
rect 25129 20032 25134 20088
rect 25190 20032 27722 20088
rect 25129 20030 27722 20032
rect 25129 20027 25195 20030
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 1669 19410 1735 19413
rect 3785 19410 3851 19413
rect 1669 19408 3851 19410
rect 1669 19352 1674 19408
rect 1730 19352 3790 19408
rect 3846 19352 3851 19408
rect 1669 19350 3851 19352
rect 1669 19347 1735 19350
rect 3785 19347 3851 19350
rect 1761 19274 1827 19277
rect 9305 19274 9371 19277
rect 1761 19272 9371 19274
rect 1761 19216 1766 19272
rect 1822 19216 9310 19272
rect 9366 19216 9371 19272
rect 1761 19214 9371 19216
rect 1761 19211 1827 19214
rect 9305 19211 9371 19214
rect 27520 19184 28000 19304
rect 0 19140 480 19168
rect 0 19076 60 19140
rect 124 19076 480 19140
rect 0 19048 480 19076
rect 13629 19138 13695 19141
rect 14549 19138 14615 19141
rect 13629 19136 14615 19138
rect 13629 19080 13634 19136
rect 13690 19080 14554 19136
rect 14610 19080 14615 19136
rect 13629 19078 14615 19080
rect 13629 19075 13695 19078
rect 14549 19075 14615 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 54 18804 60 18868
rect 124 18866 130 18868
rect 8017 18866 8083 18869
rect 124 18864 8083 18866
rect 124 18808 8022 18864
rect 8078 18808 8083 18864
rect 124 18806 8083 18808
rect 124 18804 130 18806
rect 8017 18803 8083 18806
rect 10869 18866 10935 18869
rect 21817 18866 21883 18869
rect 10869 18864 21883 18866
rect 10869 18808 10874 18864
rect 10930 18808 21822 18864
rect 21878 18808 21883 18864
rect 10869 18806 21883 18808
rect 10869 18803 10935 18806
rect 21817 18803 21883 18806
rect 10777 18730 10843 18733
rect 18597 18730 18663 18733
rect 10777 18728 18663 18730
rect 10777 18672 10782 18728
rect 10838 18672 18602 18728
rect 18658 18672 18663 18728
rect 10777 18670 18663 18672
rect 10777 18667 10843 18670
rect 18597 18667 18663 18670
rect 19333 18730 19399 18733
rect 24025 18730 24091 18733
rect 19333 18728 24091 18730
rect 19333 18672 19338 18728
rect 19394 18672 24030 18728
rect 24086 18672 24091 18728
rect 19333 18670 24091 18672
rect 19333 18667 19399 18670
rect 24025 18667 24091 18670
rect 25129 18730 25195 18733
rect 27662 18730 27722 19184
rect 25129 18728 27722 18730
rect 25129 18672 25134 18728
rect 25190 18672 27722 18728
rect 25129 18670 27722 18672
rect 25129 18667 25195 18670
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 7833 18322 7899 18325
rect 11513 18322 11579 18325
rect 62 18320 11579 18322
rect 62 18264 7838 18320
rect 7894 18264 11518 18320
rect 11574 18264 11579 18320
rect 62 18262 11579 18264
rect 62 18080 122 18262
rect 7833 18259 7899 18262
rect 11513 18259 11579 18262
rect 1485 18186 1551 18189
rect 8937 18186 9003 18189
rect 1485 18184 9003 18186
rect 1485 18128 1490 18184
rect 1546 18128 8942 18184
rect 8998 18128 9003 18184
rect 1485 18126 9003 18128
rect 1485 18123 1551 18126
rect 8937 18123 9003 18126
rect 0 17960 480 18080
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 13537 17914 13603 17917
rect 19241 17914 19307 17917
rect 13537 17912 19307 17914
rect 13537 17856 13542 17912
rect 13598 17856 19246 17912
rect 19302 17856 19307 17912
rect 13537 17854 19307 17856
rect 13537 17851 13603 17854
rect 19241 17851 19307 17854
rect 27520 17824 28000 17944
rect 12985 17778 13051 17781
rect 21909 17778 21975 17781
rect 12985 17776 21975 17778
rect 12985 17720 12990 17776
rect 13046 17720 21914 17776
rect 21970 17720 21975 17776
rect 12985 17718 21975 17720
rect 12985 17715 13051 17718
rect 21909 17715 21975 17718
rect 7373 17642 7439 17645
rect 17033 17642 17099 17645
rect 7373 17640 17099 17642
rect 7373 17584 7378 17640
rect 7434 17584 17038 17640
rect 17094 17584 17099 17640
rect 7373 17582 17099 17584
rect 7373 17579 7439 17582
rect 17033 17579 17099 17582
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 54 17308 60 17372
rect 124 17370 130 17372
rect 24761 17370 24827 17373
rect 27662 17370 27722 17824
rect 124 17310 674 17370
rect 124 17308 130 17310
rect 614 17234 674 17310
rect 24761 17368 27722 17370
rect 24761 17312 24766 17368
rect 24822 17312 27722 17368
rect 24761 17310 27722 17312
rect 24761 17307 24827 17310
rect 21357 17234 21423 17237
rect 614 17232 21423 17234
rect 614 17176 21362 17232
rect 21418 17176 21423 17232
rect 614 17174 21423 17176
rect 21357 17171 21423 17174
rect 0 17100 480 17128
rect 0 17036 60 17100
rect 124 17036 480 17100
rect 0 17008 480 17036
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 8937 16690 9003 16693
rect 19977 16690 20043 16693
rect 8937 16688 20043 16690
rect 8937 16632 8942 16688
rect 8998 16632 19982 16688
rect 20038 16632 20043 16688
rect 8937 16630 20043 16632
rect 8937 16627 9003 16630
rect 19977 16627 20043 16630
rect 27520 16464 28000 16584
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 0 15920 480 16040
rect 24761 16010 24827 16013
rect 27662 16010 27722 16464
rect 24761 16008 27722 16010
rect 24761 15952 24766 16008
rect 24822 15952 27722 16008
rect 24761 15950 27722 15952
rect 24761 15947 24827 15950
rect 62 15466 122 15920
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 3049 15602 3115 15605
rect 21265 15602 21331 15605
rect 3049 15600 21331 15602
rect 3049 15544 3054 15600
rect 3110 15544 21270 15600
rect 21326 15544 21331 15600
rect 3049 15542 21331 15544
rect 3049 15539 3115 15542
rect 21265 15539 21331 15542
rect 1577 15466 1643 15469
rect 62 15464 1643 15466
rect 62 15408 1582 15464
rect 1638 15408 1643 15464
rect 62 15406 1643 15408
rect 1577 15403 1643 15406
rect 9305 15466 9371 15469
rect 24117 15466 24183 15469
rect 9305 15464 24183 15466
rect 9305 15408 9310 15464
rect 9366 15408 24122 15464
rect 24178 15408 24183 15464
rect 9305 15406 24183 15408
rect 9305 15403 9371 15406
rect 24117 15403 24183 15406
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 6821 15194 6887 15197
rect 13997 15194 14063 15197
rect 6821 15192 14063 15194
rect 6821 15136 6826 15192
rect 6882 15136 14002 15192
rect 14058 15136 14063 15192
rect 6821 15134 14063 15136
rect 6821 15131 6887 15134
rect 13997 15131 14063 15134
rect 27520 15104 28000 15224
rect 0 14832 480 14952
rect 14917 14922 14983 14925
rect 22093 14922 22159 14925
rect 14917 14920 22159 14922
rect 14917 14864 14922 14920
rect 14978 14864 22098 14920
rect 22154 14864 22159 14920
rect 14917 14862 22159 14864
rect 14917 14859 14983 14862
rect 22093 14859 22159 14862
rect 62 14378 122 14832
rect 25405 14786 25471 14789
rect 27662 14786 27722 15104
rect 25405 14784 27722 14786
rect 25405 14728 25410 14784
rect 25466 14728 27722 14784
rect 25405 14726 27722 14728
rect 25405 14723 25471 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 22093 14650 22159 14653
rect 22093 14648 27722 14650
rect 22093 14592 22098 14648
rect 22154 14592 27722 14648
rect 22093 14590 27722 14592
rect 22093 14587 22159 14590
rect 1117 14378 1183 14381
rect 62 14376 1183 14378
rect 62 14320 1122 14376
rect 1178 14320 1183 14376
rect 62 14318 1183 14320
rect 1117 14315 1183 14318
rect 17953 14378 18019 14381
rect 21725 14378 21791 14381
rect 17953 14376 21791 14378
rect 17953 14320 17958 14376
rect 18014 14320 21730 14376
rect 21786 14320 21791 14376
rect 17953 14318 21791 14320
rect 17953 14315 18019 14318
rect 21725 14315 21791 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 27662 14000 27722 14590
rect 0 13880 480 14000
rect 27520 13880 28000 14000
rect 62 13426 122 13880
rect 10685 13834 10751 13837
rect 12709 13834 12775 13837
rect 10685 13832 12775 13834
rect 10685 13776 10690 13832
rect 10746 13776 12714 13832
rect 12770 13776 12775 13832
rect 10685 13774 12775 13776
rect 10685 13771 10751 13774
rect 12709 13771 12775 13774
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 4245 13426 4311 13429
rect 62 13424 4311 13426
rect 62 13368 4250 13424
rect 4306 13368 4311 13424
rect 62 13366 4311 13368
rect 4245 13363 4311 13366
rect 5073 13426 5139 13429
rect 19057 13426 19123 13429
rect 5073 13424 19123 13426
rect 5073 13368 5078 13424
rect 5134 13368 19062 13424
rect 19118 13368 19123 13424
rect 5073 13366 19123 13368
rect 5073 13363 5139 13366
rect 19057 13363 19123 13366
rect 9857 13290 9923 13293
rect 14733 13290 14799 13293
rect 9857 13288 14799 13290
rect 9857 13232 9862 13288
rect 9918 13232 14738 13288
rect 14794 13232 14799 13288
rect 9857 13230 14799 13232
rect 9857 13227 9923 13230
rect 14733 13227 14799 13230
rect 14917 13290 14983 13293
rect 15561 13290 15627 13293
rect 21633 13290 21699 13293
rect 14917 13288 21699 13290
rect 14917 13232 14922 13288
rect 14978 13232 15566 13288
rect 15622 13232 21638 13288
rect 21694 13232 21699 13288
rect 14917 13230 21699 13232
rect 14917 13227 14983 13230
rect 15561 13227 15627 13230
rect 21633 13227 21699 13230
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 0 12792 480 12912
rect 62 12338 122 12792
rect 10961 12610 11027 12613
rect 12433 12610 12499 12613
rect 18638 12610 18644 12612
rect 10961 12608 18644 12610
rect 10961 12552 10966 12608
rect 11022 12552 12438 12608
rect 12494 12552 18644 12608
rect 10961 12550 18644 12552
rect 10961 12547 11027 12550
rect 12433 12547 12499 12550
rect 18638 12548 18644 12550
rect 18708 12548 18714 12612
rect 23422 12548 23428 12612
rect 23492 12610 23498 12612
rect 24117 12610 24183 12613
rect 23492 12608 24183 12610
rect 23492 12552 24122 12608
rect 24178 12552 24183 12608
rect 23492 12550 24183 12552
rect 23492 12548 23498 12550
rect 24117 12547 24183 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 27520 12520 28000 12640
rect 19610 12479 19930 12480
rect 1761 12338 1827 12341
rect 62 12336 1827 12338
rect 62 12280 1766 12336
rect 1822 12280 1827 12336
rect 62 12278 1827 12280
rect 1761 12275 1827 12278
rect 20253 12202 20319 12205
rect 27662 12202 27722 12520
rect 20253 12200 27722 12202
rect 20253 12144 20258 12200
rect 20314 12144 27722 12200
rect 20253 12142 27722 12144
rect 20253 12139 20319 12142
rect 7465 12066 7531 12069
rect 14641 12066 14707 12069
rect 7465 12064 14707 12066
rect 7465 12008 7470 12064
rect 7526 12008 14646 12064
rect 14702 12008 14707 12064
rect 7465 12006 14707 12008
rect 7465 12003 7531 12006
rect 14641 12003 14707 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 0 11796 480 11824
rect 0 11732 60 11796
rect 124 11732 480 11796
rect 0 11704 480 11732
rect 54 11460 60 11524
rect 124 11522 130 11524
rect 8661 11522 8727 11525
rect 124 11520 8727 11522
rect 124 11464 8666 11520
rect 8722 11464 8727 11520
rect 124 11462 8727 11464
rect 124 11460 130 11462
rect 8661 11459 8727 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 27520 11160 28000 11280
rect 5610 10912 5930 10913
rect 0 10752 480 10872
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 24761 10842 24827 10845
rect 27662 10842 27722 11160
rect 24761 10840 27722 10842
rect 24761 10784 24766 10840
rect 24822 10784 27722 10840
rect 24761 10782 27722 10784
rect 24761 10779 24827 10782
rect 62 10298 122 10752
rect 11053 10706 11119 10709
rect 17769 10706 17835 10709
rect 11053 10704 17835 10706
rect 11053 10648 11058 10704
rect 11114 10648 17774 10704
rect 17830 10648 17835 10704
rect 11053 10646 17835 10648
rect 11053 10643 11119 10646
rect 17769 10643 17835 10646
rect 14590 10508 14596 10572
rect 14660 10570 14666 10572
rect 15377 10570 15443 10573
rect 14660 10568 15443 10570
rect 14660 10512 15382 10568
rect 15438 10512 15443 10568
rect 14660 10510 15443 10512
rect 14660 10508 14666 10510
rect 15377 10507 15443 10510
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 1853 10298 1919 10301
rect 62 10296 1919 10298
rect 62 10240 1858 10296
rect 1914 10240 1919 10296
rect 62 10238 1919 10240
rect 1853 10235 1919 10238
rect 5610 9824 5930 9825
rect 0 9664 480 9784
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 27520 9800 28000 9920
rect 24277 9759 24597 9760
rect 62 9210 122 9664
rect 3693 9618 3759 9621
rect 20345 9618 20411 9621
rect 21725 9618 21791 9621
rect 3693 9616 21791 9618
rect 3693 9560 3698 9616
rect 3754 9560 20350 9616
rect 20406 9560 21730 9616
rect 21786 9560 21791 9616
rect 3693 9558 21791 9560
rect 3693 9555 3759 9558
rect 20345 9555 20411 9558
rect 21725 9555 21791 9558
rect 24761 9346 24827 9349
rect 27662 9346 27722 9800
rect 24761 9344 27722 9346
rect 24761 9288 24766 9344
rect 24822 9288 27722 9344
rect 24761 9286 27722 9288
rect 24761 9283 24827 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 1393 9210 1459 9213
rect 62 9208 1459 9210
rect 62 9152 1398 9208
rect 1454 9152 1459 9208
rect 62 9150 1459 9152
rect 1393 9147 1459 9150
rect 54 9012 60 9076
rect 124 9074 130 9076
rect 1577 9074 1643 9077
rect 124 9072 1643 9074
rect 124 9016 1582 9072
rect 1638 9016 1643 9072
rect 124 9014 1643 9016
rect 124 9012 130 9014
rect 1577 9011 1643 9014
rect 12985 9074 13051 9077
rect 19241 9074 19307 9077
rect 20897 9074 20963 9077
rect 12985 9072 20963 9074
rect 12985 9016 12990 9072
rect 13046 9016 19246 9072
rect 19302 9016 20902 9072
rect 20958 9016 20963 9072
rect 12985 9014 20963 9016
rect 12985 9011 13051 9014
rect 19241 9011 19307 9014
rect 20897 9011 20963 9014
rect 25129 9074 25195 9077
rect 25129 9072 27722 9074
rect 25129 9016 25134 9072
rect 25190 9016 27722 9072
rect 25129 9014 27722 9016
rect 25129 9011 25195 9014
rect 0 8804 480 8832
rect 0 8740 60 8804
rect 124 8740 480 8804
rect 0 8712 480 8740
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 27662 8560 27722 9014
rect 27520 8440 28000 8560
rect 2313 8394 2379 8397
rect 15653 8394 15719 8397
rect 2313 8392 15719 8394
rect 2313 8336 2318 8392
rect 2374 8336 15658 8392
rect 15714 8336 15719 8392
rect 2313 8334 15719 8336
rect 2313 8331 2379 8334
rect 15653 8331 15719 8334
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 54 7924 60 7988
rect 124 7986 130 7988
rect 841 7986 907 7989
rect 124 7984 907 7986
rect 124 7928 846 7984
rect 902 7928 907 7984
rect 124 7926 907 7928
rect 124 7924 130 7926
rect 841 7923 907 7926
rect 1485 7986 1551 7989
rect 10961 7986 11027 7989
rect 1485 7984 11027 7986
rect 1485 7928 1490 7984
rect 1546 7928 10966 7984
rect 11022 7928 11027 7984
rect 1485 7926 11027 7928
rect 1485 7923 1551 7926
rect 10961 7923 11027 7926
rect 8661 7850 8727 7853
rect 24209 7850 24275 7853
rect 8661 7848 24275 7850
rect 8661 7792 8666 7848
rect 8722 7792 24214 7848
rect 24270 7792 24275 7848
rect 8661 7790 24275 7792
rect 8661 7787 8727 7790
rect 24209 7787 24275 7790
rect 0 7716 480 7744
rect 0 7652 60 7716
rect 124 7652 480 7716
rect 0 7624 480 7652
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 27520 7304 28000 7336
rect 27520 7248 27618 7304
rect 27674 7248 28000 7304
rect 27520 7216 28000 7248
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 54 6836 60 6900
rect 124 6898 130 6900
rect 1577 6898 1643 6901
rect 124 6896 1643 6898
rect 124 6840 1582 6896
rect 1638 6840 1643 6896
rect 124 6838 1643 6840
rect 124 6836 130 6838
rect 1577 6835 1643 6838
rect 0 6628 480 6656
rect 0 6564 60 6628
rect 124 6564 480 6628
rect 0 6536 480 6564
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 27520 5944 28000 5976
rect 27520 5888 27618 5944
rect 27674 5888 28000 5944
rect 27520 5856 28000 5888
rect 0 5584 480 5704
rect 62 5402 122 5584
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 5441 5402 5507 5405
rect 62 5400 5507 5402
rect 62 5344 5446 5400
rect 5502 5344 5507 5400
rect 62 5342 5507 5344
rect 5441 5339 5507 5342
rect 16849 5266 16915 5269
rect 62 5264 16915 5266
rect 62 5208 16854 5264
rect 16910 5208 16915 5264
rect 62 5206 16915 5208
rect 62 4616 122 5206
rect 16849 5203 16915 5206
rect 5441 5130 5507 5133
rect 8569 5130 8635 5133
rect 14089 5130 14155 5133
rect 5441 5128 14155 5130
rect 5441 5072 5446 5128
rect 5502 5072 8574 5128
rect 8630 5072 14094 5128
rect 14150 5072 14155 5128
rect 5441 5070 14155 5072
rect 5441 5067 5507 5070
rect 8569 5067 8635 5070
rect 14089 5067 14155 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 0 4496 480 4616
rect 27520 4584 28000 4616
rect 27520 4528 27710 4584
rect 27766 4528 28000 4584
rect 27520 4496 28000 4528
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 0 3496 480 3528
rect 0 3440 110 3496
rect 166 3440 480 3496
rect 0 3408 480 3440
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 27520 3136 28000 3256
rect 1853 3090 1919 3093
rect 62 3088 1919 3090
rect 62 3032 1858 3088
rect 1914 3032 1919 3088
rect 62 3030 1919 3032
rect 62 2576 122 3030
rect 1853 3027 1919 3030
rect 24945 2818 25011 2821
rect 27662 2818 27722 3136
rect 24945 2816 27722 2818
rect 24945 2760 24950 2816
rect 25006 2760 27722 2816
rect 24945 2758 27722 2760
rect 24945 2755 25011 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 0 2456 480 2576
rect 8937 2546 9003 2549
rect 18873 2546 18939 2549
rect 8937 2544 18939 2546
rect 8937 2488 8942 2544
rect 8998 2488 18878 2544
rect 18934 2488 18939 2544
rect 8937 2486 18939 2488
rect 8937 2483 9003 2486
rect 18873 2483 18939 2486
rect 20161 2410 20227 2413
rect 27654 2410 27660 2412
rect 20161 2408 27660 2410
rect 20161 2352 20166 2408
rect 20222 2352 27660 2408
rect 20161 2350 27660 2352
rect 20161 2347 20227 2350
rect 27654 2348 27660 2350
rect 27724 2348 27730 2412
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 2037 2002 2103 2005
rect 62 2000 2103 2002
rect 62 1944 2042 2000
rect 2098 1944 2103 2000
rect 62 1942 2103 1944
rect 62 1488 122 1942
rect 2037 1939 2103 1942
rect 9765 1866 9831 1869
rect 22185 1866 22251 1869
rect 9765 1864 22251 1866
rect 9765 1808 9770 1864
rect 9826 1808 22190 1864
rect 22246 1808 22251 1864
rect 9765 1806 22251 1808
rect 9765 1803 9831 1806
rect 22185 1803 22251 1806
rect 27520 1868 28000 1896
rect 27520 1804 27660 1868
rect 27724 1804 28000 1868
rect 27520 1776 28000 1804
rect 0 1368 480 1488
rect 21449 1186 21515 1189
rect 21449 1184 27722 1186
rect 21449 1128 21454 1184
rect 21510 1128 27722 1184
rect 21449 1126 27722 1128
rect 21449 1123 21515 1126
rect 1301 1050 1367 1053
rect 62 1048 1367 1050
rect 62 992 1306 1048
rect 1362 992 1367 1048
rect 62 990 1367 992
rect 62 536 122 990
rect 1301 987 1367 990
rect 27662 672 27722 1126
rect 27520 552 28000 672
rect 0 416 480 536
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 14596 23428 14660 23492
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 60 19076 124 19140
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 60 18804 124 18868
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 60 17308 124 17372
rect 60 17036 124 17100
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 18644 12548 18708 12612
rect 23428 12548 23492 12612
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 60 11732 124 11796
rect 60 11460 124 11524
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 14596 10508 14660 10572
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 60 9012 124 9076
rect 60 8740 124 8804
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 60 7924 124 7988
rect 60 7652 124 7716
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 60 6836 124 6900
rect 60 6564 124 6628
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 27660 2348 27724 2412
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 27660 1804 27724 1868
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 59 19140 125 19141
rect 59 19076 60 19140
rect 124 19076 125 19140
rect 59 19075 125 19076
rect 62 18869 122 19075
rect 59 18868 125 18869
rect 59 18804 60 18868
rect 124 18804 125 18868
rect 59 18803 125 18804
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 59 17372 125 17373
rect 59 17308 60 17372
rect 124 17308 125 17372
rect 59 17307 125 17308
rect 62 17101 122 17307
rect 59 17100 125 17101
rect 59 17036 60 17100
rect 124 17036 125 17100
rect 59 17035 125 17036
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 59 11796 125 11797
rect 59 11732 60 11796
rect 124 11732 125 11796
rect 59 11731 125 11732
rect 62 11525 122 11731
rect 59 11524 125 11525
rect 59 11460 60 11524
rect 124 11460 125 11524
rect 59 11459 125 11460
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 59 9076 125 9077
rect 59 9012 60 9076
rect 124 9012 125 9076
rect 59 9011 125 9012
rect 62 8805 122 9011
rect 59 8804 125 8805
rect 59 8740 60 8804
rect 124 8740 125 8804
rect 59 8739 125 8740
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 59 7988 125 7989
rect 59 7924 60 7988
rect 124 7924 125 7988
rect 59 7923 125 7924
rect 62 7717 122 7923
rect 59 7716 125 7717
rect 59 7652 60 7716
rect 124 7652 125 7716
rect 59 7651 125 7652
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 59 6900 125 6901
rect 59 6836 60 6900
rect 124 6836 125 6900
rect 59 6835 125 6836
rect 62 6629 122 6835
rect 59 6628 125 6629
rect 59 6564 60 6628
rect 124 6564 125 6628
rect 59 6563 125 6564
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14595 23492 14661 23493
rect 14595 23428 14596 23492
rect 14660 23428 14661 23492
rect 14595 23427 14661 23428
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 14598 10573 14658 23427
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14595 10572 14661 10573
rect 14595 10508 14596 10572
rect 14660 10508 14661 10572
rect 14595 10507 14661 10508
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 27659 2412 27725 2413
rect 27659 2348 27660 2412
rect 27724 2348 27725 2412
rect 27659 2347 27725 2348
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 27662 1869 27722 2347
rect 27659 1868 27725 1869
rect 27659 1804 27660 1868
rect 27724 1804 27725 1868
rect 27659 1803 27725 1804
<< via4 >>
rect 18558 12612 18794 12698
rect 18558 12548 18644 12612
rect 18644 12548 18708 12612
rect 18708 12548 18794 12612
rect 18558 12462 18794 12548
rect 23342 12612 23578 12698
rect 23342 12548 23428 12612
rect 23428 12548 23492 12612
rect 23492 12548 23578 12612
rect 23342 12462 23578 12548
<< metal5 >>
rect 18516 12698 23620 12740
rect 18516 12462 18558 12698
rect 18794 12462 23342 12698
rect 23578 12462 23620 12698
rect 18516 12420 23620 12462
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_2.tap_buf4_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3864 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_33 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_37
timestamp 1586364061
transform 1 0 4508 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_49
timestamp 1586364061
transform 1 0 5612 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_66
timestamp 1586364061
transform 1 0 7176 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_70
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_77
timestamp 1586364061
transform 1 0 8188 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_81
timestamp 1586364061
transform 1 0 8556 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_112 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _194_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 18860 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_191
timestamp 1586364061
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_195
timestamp 1586364061
transform 1 0 19044 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_0_207 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20148 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_215
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_221
timestamp 1586364061
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_225
timestamp 1586364061
transform 1 0 21804 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_0_238
timestamp 1586364061
transform 1 0 23000 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_233
timestamp 1586364061
transform 1 0 22540 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22724 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _190_
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_259
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_263
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 24564 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_253
timestamp 1586364061
transform 1 0 24380 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_19
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_31
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_43
timestamp 1586364061
transform 1 0 5060 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_55
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 590 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_buf_2  _186_
timestamp 1586364061
transform 1 0 24564 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_259
timestamp 1586364061
transform 1 0 24932 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_271
timestamp 1586364061
transform 1 0 26036 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_buf_2  _191_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_19
timestamp 1586364061
transform 1 0 2852 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_19
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 5060 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_42
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_45
timestamp 1586364061
transform 1 0 5244 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 774 592
use scs8hd_buf_2  _185_
timestamp 1586364061
transform 1 0 24564 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 25116 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_253
timestamp 1586364061
transform 1 0 24380 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_259
timestamp 1586364061
transform 1 0 24932 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_263
timestamp 1586364061
transform 1 0 25300 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_275
timestamp 1586364061
transform 1 0 26404 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _187_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_1  _068_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_19
timestamp 1586364061
transform 1 0 2852 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_35
timestamp 1586364061
transform 1 0 4324 0 -1 8160
box -38 -48 774 592
use scs8hd_buf_1  _151_
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_46
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_58
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_70
timestamp 1586364061
transform 1 0 7544 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_82
timestamp 1586364061
transform 1 0 8648 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_90
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_202
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_6
timestamp 1586364061
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_10
timestamp 1586364061
transform 1 0 2024 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_14
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 590 592
use scs8hd_buf_1  _079_
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 314 592
use scs8hd_buf_1  _166_
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_25
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_29
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5612 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_36
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_47
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 7544 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_55
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 590 592
use scs8hd_decap_8  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 774 592
use scs8hd_decap_12  FILLER_11_72
timestamp 1586364061
transform 1 0 7728 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_84
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_96
timestamp 1586364061
transform 1 0 9936 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_108
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_11_120
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 24564 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_253
timestamp 1586364061
transform 1 0 24380 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_buf_2  _184_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__067__C
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_13
timestamp 1586364061
transform 1 0 2300 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_16
timestamp 1586364061
transform 1 0 2576 0 -1 9248
box -38 -48 406 592
use scs8hd_buf_1  _092_
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4968 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_6  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_8  FILLER_12_51
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 774 592
use scs8hd_buf_1  _107_
timestamp 1586364061
transform 1 0 7544 0 -1 9248
box -38 -48 314 592
use scs8hd_conb_1  _181_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_62
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_66
timestamp 1586364061
transform 1 0 7176 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_73
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_12_85
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_91
timestamp 1586364061
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_134
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_146
timestamp 1586364061
transform 1 0 14536 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_152
timestamp 1586364061
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_buf_2  _199_
timestamp 1586364061
transform 1 0 24564 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_259
timestamp 1586364061
transform 1 0 24932 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_271
timestamp 1586364061
transform 1 0 26036 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_6
timestamp 1586364061
transform 1 0 1656 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 1840 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_buf_1  _077_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_16
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_10
timestamp 1586364061
transform 1 0 2024 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_or3_4  _067_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_26
timestamp 1586364061
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_20
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__B
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_30
timestamp 1586364061
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_45
timestamp 1586364061
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_49
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_52
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_69
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6624 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_buf_1  _069_
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 314 592
use scs8hd_conb_1  _180_
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_75
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_82
timestamp 1586364061
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_6  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_6  FILLER_13_93
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_conb_1  _179_
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_103
timestamp 1586364061
transform 1 0 10580 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_99
timestamp 1586364061
transform 1 0 10212 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_99
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_1  _101_
timestamp 1586364061
transform 1 0 10304 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_102
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_119
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_3  FILLER_13_127
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_138
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_134
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_141
timestamp 1586364061
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_8  FILLER_13_145
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_157
timestamp 1586364061
transform 1 0 15548 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_160
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_156
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_153
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_167
timestamp 1586364061
transform 1 0 16468 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_161
timestamp 1586364061
transform 1 0 15916 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_168
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_164
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_177
timestamp 1586364061
transform 1 0 17388 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_176
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_172
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 17572 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_182
timestamp 1586364061
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_14_181
timestamp 1586364061
transform 1 0 17756 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_186
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_198
timestamp 1586364061
transform 1 0 19320 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_210
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_253
timestamp 1586364061
transform 1 0 24380 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_258
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_262
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_274
timestamp 1586364061
transform 1 0 26312 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_8  _065_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_20
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_35
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8832 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_73
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_77
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_81
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_87
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _154_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_91
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_95
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_99
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_126
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_130
timestamp 1586364061
transform 1 0 13064 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_151
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_164
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_168
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_204
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_214
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_229
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_241
timestamp 1586364061
transform 1 0 23276 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 774 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 24564 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 24380 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_259
timestamp 1586364061
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_263
timestamp 1586364061
transform 1 0 25300 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_275
timestamp 1586364061
transform 1 0 26404 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _089_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _171_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_12
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_41
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_46
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_50
timestamp 1586364061
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_62
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_66
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_79
timestamp 1586364061
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_83
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_87
timestamp 1586364061
transform 1 0 9108 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_107
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11316 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_16_122
timestamp 1586364061
transform 1 0 12328 0 -1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_128
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15732 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_158
timestamp 1586364061
transform 1 0 15640 0 -1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _155_
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_170
timestamp 1586364061
transform 1 0 16744 0 -1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_187
timestamp 1586364061
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_191
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_204
timestamp 1586364061
transform 1 0 19872 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_212
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_218
timestamp 1586364061
transform 1 0 21160 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_230
timestamp 1586364061
transform 1 0 22264 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_242
timestamp 1586364061
transform 1 0 23368 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _188_
timestamp 1586364061
transform 1 0 24564 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_254
timestamp 1586364061
transform 1 0 24472 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_259
timestamp 1586364061
transform 1 0 24932 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_271
timestamp 1586364061
transform 1 0 26036 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_or3_4  _085_
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _170_
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__C
timestamp 1586364061
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_19
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_23
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _168_
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_36
timestamp 1586364061
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_40
timestamp 1586364061
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _172_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_77
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 406 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_94
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_102
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_137
timestamp 1586364061
transform 1 0 13708 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_141
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14996 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_145
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_149
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_164
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_168
timestamp 1586364061
transform 1 0 16560 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_201
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_214
timestamp 1586364061
transform 1 0 20792 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21528 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21988 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_218
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_225
timestamp 1586364061
transform 1 0 21804 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_229
timestamp 1586364061
transform 1 0 22172 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_241
timestamp 1586364061
transform 1 0 23276 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_inv_8  _066_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 2576 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_12
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 406 592
use scs8hd_buf_1  _083_
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 314 592
use scs8hd_buf_2  _198_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__078__C
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_18
timestamp 1586364061
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 4968 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_36
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_40
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_53
timestamp 1586364061
transform 1 0 5980 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_1  _105_
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_57
timestamp 1586364061
transform 1 0 6348 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_61
timestamp 1586364061
transform 1 0 6716 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_67
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 590 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use scs8hd_nor2_4  _084_
timestamp 1586364061
transform 1 0 9752 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_103
timestamp 1586364061
transform 1 0 10580 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_107
timestamp 1586364061
transform 1 0 10948 0 -1 12512
box -38 -48 406 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_6  FILLER_18_120
timestamp 1586364061
transform 1 0 12144 0 -1 12512
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_128
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_132
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 406 592
use scs8hd_buf_1  _128_
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_157
timestamp 1586364061
transform 1 0 15548 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_18_161
timestamp 1586364061
transform 1 0 15916 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_174
timestamp 1586364061
transform 1 0 17112 0 -1 12512
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18216 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_197
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_201
timestamp 1586364061
transform 1 0 19596 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_205
timestamp 1586364061
transform 1 0 19964 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_208
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_224
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_228
timestamp 1586364061
transform 1 0 22080 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_240
timestamp 1586364061
transform 1 0 23184 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_252
timestamp 1586364061
transform 1 0 24288 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_264
timestamp 1586364061
transform 1 0 25392 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_272
timestamp 1586364061
transform 1 0 26128 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 2668 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use scs8hd_inv_8  _081_
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_19
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__C
timestamp 1586364061
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_34
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_19_28
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__165__C
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_or2_4  _071_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 682 592
use scs8hd_or3_4  _078_
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_43
timestamp 1586364061
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_39
timestamp 1586364061
transform 1 0 4692 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__C
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_47
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_52
timestamp 1586364061
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 5520 0 -1 13600
box -38 -48 1050 592
use scs8hd_nor2_4  _167_
timestamp 1586364061
transform 1 0 5060 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_59
timestamp 1586364061
transform 1 0 6532 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_56
timestamp 1586364061
transform 1 0 6256 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6072 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_71
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_64
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_96
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_92
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 9936 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_103
timestamp 1586364061
transform 1 0 10580 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_99
timestamp 1586364061
transform 1 0 10212 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 10396 0 -1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 10948 0 -1 13600
box -38 -48 1050 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_109
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_113
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_121
timestamp 1586364061
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_117
timestamp 1586364061
transform 1 0 11868 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_122
timestamp 1586364061
transform 1 0 12328 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_buf_1  _099_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_130
timestamp 1586364061
transform 1 0 13064 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_126
timestamp 1586364061
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_134
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12696 0 -1 13600
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_152
timestamp 1586364061
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 17020 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_165
timestamp 1586364061
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_169
timestamp 1586364061
transform 1 0 16652 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_186
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_182
timestamp 1586364061
transform 1 0 17848 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_189
timestamp 1586364061
transform 1 0 18492 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 18768 0 -1 13600
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18308 0 1 12512
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_20_203
timestamp 1586364061
transform 1 0 19780 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_202
timestamp 1586364061
transform 1 0 19688 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_198
timestamp 1586364061
transform 1 0 19320 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19872 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19504 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_213
timestamp 1586364061
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_20_207
timestamp 1586364061
transform 1 0 20148 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 20056 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21804 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21620 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21252 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_217
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_221
timestamp 1586364061
transform 1 0 21436 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_234
timestamp 1586364061
transform 1 0 22632 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_242
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_236
timestamp 1586364061
transform 1 0 22816 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_248
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_253
timestamp 1586364061
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_258
timestamp 1586364061
transform 1 0 24840 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_262
timestamp 1586364061
transform 1 0 25208 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_260
timestamp 1586364061
transform 1 0 25024 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_274
timestamp 1586364061
transform 1 0 26312 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_272
timestamp 1586364061
transform 1 0 26128 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_or3_4  _091_
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 866 592
use scs8hd_buf_2  _195_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 2024 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_12
timestamp 1586364061
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use scs8hd_or3_4  _082_
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_25
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_29
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use scs8hd_buf_1  _086_
timestamp 1586364061
transform 1 0 5704 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_42
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_46
timestamp 1586364061
transform 1 0 5336 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _090_
timestamp 1586364061
transform 1 0 7452 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 7268 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_66
timestamp 1586364061
transform 1 0 7176 0 1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _087_
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_78
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_82
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_99
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_buf_1  _075_
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_132
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_136
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15088 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_143
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 314 592
use scs8hd_conb_1  _176_
timestamp 1586364061
transform 1 0 16652 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 16468 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_161
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_165
timestamp 1586364061
transform 1 0 16284 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_172
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_176
timestamp 1586364061
transform 1 0 17296 0 1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_180
timestamp 1586364061
transform 1 0 17664 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_210
timestamp 1586364061
transform 1 0 20424 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_214
timestamp 1586364061
transform 1 0 20792 0 1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22172 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_217
timestamp 1586364061
transform 1 0 21068 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_227
timestamp 1586364061
transform 1 0 21988 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_231
timestamp 1586364061
transform 1 0 22356 0 1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_239
timestamp 1586364061
transform 1 0 23092 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_243
timestamp 1586364061
transform 1 0 23460 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 24564 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_253
timestamp 1586364061
transform 1 0 24380 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_or3_4  _088_
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 314 592
use scs8hd_inv_8  _094_
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 3496 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_19
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_28
timestamp 1586364061
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use scs8hd_inv_8  _072_
timestamp 1586364061
transform 1 0 5612 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__D
timestamp 1586364061
transform 1 0 5428 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_41
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_45
timestamp 1586364061
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_58
timestamp 1586364061
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_62
timestamp 1586364061
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_66
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_70
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_81
timestamp 1586364061
transform 1 0 8556 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_85
timestamp 1586364061
transform 1 0 8924 0 -1 14688
box -38 -48 590 592
use scs8hd_nor2_4  _076_
timestamp 1586364061
transform 1 0 10120 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_91
timestamp 1586364061
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_97
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_107
timestamp 1586364061
transform 1 0 10948 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 11684 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_111
timestamp 1586364061
transform 1 0 11316 0 -1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_126
timestamp 1586364061
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_130
timestamp 1586364061
transform 1 0 13064 0 -1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_143
timestamp 1586364061
transform 1 0 14260 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 17112 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_165
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_173
timestamp 1586364061
transform 1 0 17020 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 18124 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18492 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_183
timestamp 1586364061
transform 1 0 17940 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_187
timestamp 1586364061
transform 1 0 18308 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19964 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20332 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_200
timestamp 1586364061
transform 1 0 19504 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_204
timestamp 1586364061
transform 1 0 19872 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_207
timestamp 1586364061
transform 1 0 20148 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_211
timestamp 1586364061
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21896 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 21344 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_218
timestamp 1586364061
transform 1 0 21160 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_222
timestamp 1586364061
transform 1 0 21528 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_229
timestamp 1586364061
transform 1 0 22172 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22908 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_240
timestamp 1586364061
transform 1 0 23184 0 -1 14688
box -38 -48 1142 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 24564 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  FILLER_22_252
timestamp 1586364061
transform 1 0 24288 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_259
timestamp 1586364061
transform 1 0 24932 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_271
timestamp 1586364061
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_inv_8  _117_
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_12
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_16
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use scs8hd_or3_4  _165_
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_20
timestamp 1586364061
transform 1 0 2944 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_35
timestamp 1586364061
transform 1 0 4324 0 1 14688
box -38 -48 222 592
use scs8hd_or4_4  _127_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5060 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_52
timestamp 1586364061
transform 1 0 5888 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6072 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 6440 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_56
timestamp 1586364061
transform 1 0 6256 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_60
timestamp 1586364061
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use scs8hd_inv_8  _148_
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_77
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_81
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 9936 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 10304 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_94
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_102
timestamp 1586364061
transform 1 0 10488 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_136
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_140
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_151
timestamp 1586364061
transform 1 0 14996 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_164
timestamp 1586364061
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_168
timestamp 1586364061
transform 1 0 16560 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 18216 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19964 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_201
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_214
timestamp 1586364061
transform 1 0 20792 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_218
timestamp 1586364061
transform 1 0 21160 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_231
timestamp 1586364061
transform 1 0 22356 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22540 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_235
timestamp 1586364061
transform 1 0 22724 0 1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_23_243
timestamp 1586364061
transform 1 0 23460 0 1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_249
timestamp 1586364061
transform 1 0 24012 0 1 14688
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 24564 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24932 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_253
timestamp 1586364061
transform 1 0 24380 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_261
timestamp 1586364061
transform 1 0 25116 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_23_273
timestamp 1586364061
transform 1 0 26220 0 1 14688
box -38 -48 406 592
use scs8hd_or3_4  _149_
timestamp 1586364061
transform 1 0 2024 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__073__C
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_8
timestamp 1586364061
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use scs8hd_or3_4  _150_
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__119__C
timestamp 1586364061
transform 1 0 3036 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__C
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_19
timestamp 1586364061
transform 1 0 2852 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 5060 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 5796 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_41
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_45
timestamp 1586364061
transform 1 0 5244 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_49
timestamp 1586364061
transform 1 0 5612 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_53
timestamp 1586364061
transform 1 0 5980 0 -1 15776
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6072 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_65
timestamp 1586364061
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_69
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 774 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_107
timestamp 1586364061
transform 1 0 10948 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 11316 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 12512 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_122
timestamp 1586364061
transform 1 0 12328 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_126
timestamp 1586364061
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_130
timestamp 1586364061
transform 1 0 13064 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_151
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_2  _192_
timestamp 1586364061
transform 1 0 16836 0 -1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 17388 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_168
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_175
timestamp 1586364061
transform 1 0 17204 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18032 0 -1 15776
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_24_179
timestamp 1586364061
transform 1 0 17572 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_183
timestamp 1586364061
transform 1 0 17940 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_195
timestamp 1586364061
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_199
timestamp 1586364061
transform 1 0 19412 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_210
timestamp 1586364061
transform 1 0 20424 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_224
timestamp 1586364061
transform 1 0 21712 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_228
timestamp 1586364061
transform 1 0 22080 0 -1 15776
box -38 -48 406 592
use scs8hd_conb_1  _175_
timestamp 1586364061
transform 1 0 22448 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_235
timestamp 1586364061
transform 1 0 22724 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_247
timestamp 1586364061
transform 1 0 23828 0 -1 15776
box -38 -48 774 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 24564 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_259
timestamp 1586364061
transform 1 0 24932 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_271
timestamp 1586364061
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_nand3_4  _073_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 1 15776
box -38 -48 1326 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 3496 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_20
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_24
timestamp 1586364061
transform 1 0 3312 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_28
timestamp 1586364061
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_32
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_nor4_4  _164_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__D
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_73
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_77
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_90
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_96
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_100
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _138_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_119
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_138
timestamp 1586364061
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_142
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_146
timestamp 1586364061
transform 1 0 14536 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_158
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_162
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_195
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20056 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_199
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_203
timestamp 1586364061
transform 1 0 19780 0 1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21804 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22264 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_217
timestamp 1586364061
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_221
timestamp 1586364061
transform 1 0 21436 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_228
timestamp 1586364061
transform 1 0 22080 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22632 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_248
timestamp 1586364061
transform 1 0 23920 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 24564 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_252
timestamp 1586364061
transform 1 0 24288 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_6
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_10
timestamp 1586364061
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__D
timestamp 1586364061
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 2024 0 1 16864
box -38 -48 222 592
use scs8hd_or4_4  _119_
timestamp 1586364061
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_8  _070_
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_25
timestamp 1586364061
transform 1 0 3404 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_21
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__D
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__C
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_or4_4  _135_
timestamp 1586364061
transform 1 0 3772 0 1 16864
box -38 -48 866 592
use scs8hd_or2_4  _118_
timestamp 1586364061
transform 1 0 5336 0 1 16864
box -38 -48 682 592
use scs8hd_nor4_4  _163_
timestamp 1586364061
transform 1 0 4600 0 -1 16864
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__C
timestamp 1586364061
transform 1 0 4416 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_38
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_42
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_59
timestamp 1586364061
transform 1 0 6532 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_55
timestamp 1586364061
transform 1 0 6164 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 6348 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_71
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_65
timestamp 1586364061
transform 1 0 7084 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 6900 0 -1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 6900 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_76
timestamp 1586364061
transform 1 0 8096 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_72
timestamp 1586364061
transform 1 0 7728 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_89
timestamp 1586364061
transform 1 0 9292 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_86
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_26_82
timestamp 1586364061
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 16864
box -38 -48 866 592
use scs8hd_inv_8  _147_
timestamp 1586364061
transform 1 0 7820 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_97
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_93
timestamp 1586364061
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_97
timestamp 1586364061
transform 1 0 10028 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_101
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 10120 0 -1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11684 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_109
timestamp 1586364061
transform 1 0 11132 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_128
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_132
timestamp 1586364061
transform 1 0 13248 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_138
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_142
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 14720 0 1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14720 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_150
timestamp 1586364061
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_163
timestamp 1586364061
transform 1 0 16100 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_168
timestamp 1586364061
transform 1 0 16560 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_164
timestamp 1586364061
transform 1 0 16192 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16468 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_170
timestamp 1586364061
transform 1 0 16744 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_26_172
timestamp 1586364061
transform 1 0 16928 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 17296 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_3  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_185
timestamp 1586364061
transform 1 0 18124 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_189
timestamp 1586364061
transform 1 0 18492 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18676 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 18860 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19872 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19320 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_200
timestamp 1586364061
transform 1 0 19504 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_207
timestamp 1586364061
transform 1 0 20148 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_211
timestamp 1586364061
transform 1 0 20516 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_222
timestamp 1586364061
transform 1 0 21528 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_218
timestamp 1586364061
transform 1 0 21160 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_218
timestamp 1586364061
transform 1 0 21160 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 314 592
use scs8hd_buf_1  _120_
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21712 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21896 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_226
timestamp 1586364061
transform 1 0 21896 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_229
timestamp 1586364061
transform 1 0 22172 0 -1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_241
timestamp 1586364061
transform 1 0 23276 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_27_238
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 590 592
use scs8hd_decap_8  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 774 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 24564 0 -1 16864
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_253
timestamp 1586364061
transform 1 0 24380 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_259
timestamp 1586364061
transform 1 0 24932 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_253
timestamp 1586364061
transform 1 0 24380 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_258
timestamp 1586364061
transform 1 0 24840 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_262
timestamp 1586364061
transform 1 0 25208 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_271
timestamp 1586364061
transform 1 0 26036 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_27_274
timestamp 1586364061
transform 1 0 26312 0 1 16864
box -38 -48 314 592
use scs8hd_nor3_4  _160_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1472 0 -1 17952
box -38 -48 1234 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_17
timestamp 1586364061
transform 1 0 2668 0 -1 17952
box -38 -48 222 592
use scs8hd_or3_4  _109_
timestamp 1586364061
transform 1 0 4324 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 2852 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_21
timestamp 1586364061
transform 1 0 3036 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 5888 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 5336 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__C
timestamp 1586364061
transform 1 0 5704 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_48
timestamp 1586364061
transform 1 0 5520 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 6900 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_61
timestamp 1586364061
transform 1 0 6716 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_65
timestamp 1586364061
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 10212 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_97
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11776 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_108
timestamp 1586364061
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_112
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_125
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_135
timestamp 1586364061
transform 1 0 13524 0 -1 17952
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_149
timestamp 1586364061
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 17020 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_165
timestamp 1586364061
transform 1 0 16284 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_169
timestamp 1586364061
transform 1 0 16652 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_8  FILLER_28_176
timestamp 1586364061
transform 1 0 17296 0 -1 17952
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18124 0 -1 17952
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_28_184
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_196
timestamp 1586364061
transform 1 0 19136 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19320 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_200
timestamp 1586364061
transform 1 0 19504 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_208
timestamp 1586364061
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_212
timestamp 1586364061
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_218
timestamp 1586364061
transform 1 0 21160 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_230
timestamp 1586364061
transform 1 0 22264 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_242
timestamp 1586364061
transform 1 0 23368 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_254
timestamp 1586364061
transform 1 0 24472 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_266
timestamp 1586364061
transform 1 0 25576 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_274
timestamp 1586364061
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_nor3_4  _159_
timestamp 1586364061
transform 1 0 1564 0 1 17952
box -38 -48 1234 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 3496 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_18
timestamp 1586364061
transform 1 0 2760 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_22
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_28
timestamp 1586364061
transform 1 0 3680 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_32
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use scs8hd_nor3_4  _161_
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_49
timestamp 1586364061
transform 1 0 5612 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__C
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_65
timestamp 1586364061
transform 1 0 7084 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_69
timestamp 1586364061
transform 1 0 7452 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_84
timestamp 1586364061
transform 1 0 8832 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_88
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10948 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_101
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_105
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_112
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_116
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_120
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_140
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14444 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_144
timestamp 1586364061
transform 1 0 14352 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_158
timestamp 1586364061
transform 1 0 15640 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_162
timestamp 1586364061
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 18676 0 1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 18492 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_188
timestamp 1586364061
transform 1 0 18400 0 1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20424 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_202
timestamp 1586364061
transform 1 0 19688 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_206
timestamp 1586364061
transform 1 0 20056 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_219
timestamp 1586364061
transform 1 0 21252 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_231
timestamp 1586364061
transform 1 0 22356 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_243
timestamp 1586364061
transform 1 0 23460 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 1050 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_17
timestamp 1586364061
transform 1 0 2668 0 -1 19040
box -38 -48 222 592
use scs8hd_nor3_4  _162_
timestamp 1586364061
transform 1 0 4324 0 -1 19040
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__159__C
timestamp 1586364061
transform 1 0 2852 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_21
timestamp 1586364061
transform 1 0 3036 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_25
timestamp 1586364061
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_29
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__162__C
timestamp 1586364061
transform 1 0 5704 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_48
timestamp 1586364061
transform 1 0 5520 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_52
timestamp 1586364061
transform 1 0 5888 0 -1 19040
box -38 -48 222 592
use scs8hd_or2_4  _074_
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_63
timestamp 1586364061
transform 1 0 6900 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_67
timestamp 1586364061
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_71
timestamp 1586364061
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_88
timestamp 1586364061
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_106
timestamp 1586364061
transform 1 0 10856 0 -1 19040
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 11316 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12512 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_110
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_122
timestamp 1586364061
transform 1 0 12328 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_126
timestamp 1586364061
transform 1 0 12696 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_139
timestamp 1586364061
transform 1 0 13892 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_143
timestamp 1586364061
transform 1 0 14260 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_147
timestamp 1586364061
transform 1 0 14628 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_3  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 17388 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_174
timestamp 1586364061
transform 1 0 17112 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18952 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18400 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18768 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_186
timestamp 1586364061
transform 1 0 18216 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19964 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_203
timestamp 1586364061
transform 1 0 19780 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_207
timestamp 1586364061
transform 1 0 20148 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_213
timestamp 1586364061
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use scs8hd_conb_1  _174_
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_218
timestamp 1586364061
transform 1 0 21160 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_230
timestamp 1586364061
transform 1 0 22264 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_242
timestamp 1586364061
transform 1 0 23368 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_254
timestamp 1586364061
transform 1 0 24472 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_266
timestamp 1586364061
transform 1 0 25576 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_274
timestamp 1586364061
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2024 0 1 19040
box -38 -48 1050 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 314 592
use scs8hd_or2_4  _095_
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_21
timestamp 1586364061
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_25
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_36
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_40
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_or2_4  _096_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_69
timestamp 1586364061
transform 1 0 7452 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8280 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 9292 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8096 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_73
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_87
timestamp 1586364061
transform 1 0 9108 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_91
timestamp 1586364061
transform 1 0 9476 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_104
timestamp 1586364061
transform 1 0 10672 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_108
timestamp 1586364061
transform 1 0 11040 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_112
timestamp 1586364061
transform 1 0 11408 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_116
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_132
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_136
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_149
timestamp 1586364061
transform 1 0 14812 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_153
timestamp 1586364061
transform 1 0 15180 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_156
timestamp 1586364061
transform 1 0 15456 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_166
timestamp 1586364061
transform 1 0 16376 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_170
timestamp 1586364061
transform 1 0 16744 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_195
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 19596 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_199
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_212
timestamp 1586364061
transform 1 0 20608 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21804 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_217
timestamp 1586364061
transform 1 0 21068 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_223
timestamp 1586364061
transform 1 0 21620 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_227
timestamp 1586364061
transform 1 0 21988 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_239
timestamp 1586364061
transform 1 0 23092 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_243
timestamp 1586364061
transform 1 0 23460 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_253
timestamp 1586364061
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_258
timestamp 1586364061
transform 1 0 24840 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_262
timestamp 1586364061
transform 1 0 25208 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_266
timestamp 1586364061
transform 1 0 25576 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_274
timestamp 1586364061
transform 1 0 26312 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_6
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_12
timestamp 1586364061
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4692 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5888 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4508 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_36
timestamp 1586364061
transform 1 0 4416 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_50
timestamp 1586364061
transform 1 0 5704 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_8  _143_
timestamp 1586364061
transform 1 0 6440 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_54
timestamp 1586364061
transform 1 0 6072 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_67
timestamp 1586364061
transform 1 0 7268 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_71
timestamp 1586364061
transform 1 0 7636 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 590 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_102
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 11592 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11040 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_110
timestamp 1586364061
transform 1 0 11224 0 -1 20128
box -38 -48 406 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 13616 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_125
timestamp 1586364061
transform 1 0 12604 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_135
timestamp 1586364061
transform 1 0 13524 0 -1 20128
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_149
timestamp 1586364061
transform 1 0 14812 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_165
timestamp 1586364061
transform 1 0 16284 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_169
timestamp 1586364061
transform 1 0 16652 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_177
timestamp 1586364061
transform 1 0 17388 0 -1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 17572 0 -1 20128
box -38 -48 866 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 19136 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18952 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_188
timestamp 1586364061
transform 1 0 18400 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_192
timestamp 1586364061
transform 1 0 18768 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_205
timestamp 1586364061
transform 1 0 19964 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_209
timestamp 1586364061
transform 1 0 20332 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_213
timestamp 1586364061
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21436 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_218
timestamp 1586364061
transform 1 0 21160 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_223
timestamp 1586364061
transform 1 0 21620 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_235
timestamp 1586364061
transform 1 0 22724 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_247
timestamp 1586364061
transform 1 0 23828 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_258
timestamp 1586364061
transform 1 0 24840 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_270
timestamp 1586364061
transform 1 0 25944 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_274
timestamp 1586364061
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1656 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_17
timestamp 1586364061
transform 1 0 2668 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_11
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__C
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_25
timestamp 1586364061
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_21
timestamp 1586364061
transform 1 0 3036 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_29
timestamp 1586364061
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_35
timestamp 1586364061
transform 1 0 4324 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_31
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 3772 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4140 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2760 0 1 20128
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4876 0 -1 21216
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5060 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4876 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_52
timestamp 1586364061
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_40
timestamp 1586364061
transform 1 0 4784 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_52
timestamp 1586364061
transform 1 0 5888 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_33_60
timestamp 1586364061
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_56
timestamp 1586364061
transform 1 0 6256 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 6808 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_64
timestamp 1586364061
transform 1 0 6992 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_69
timestamp 1586364061
transform 1 0 7452 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_65
timestamp 1586364061
transform 1 0 7084 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7452 0 -1 21216
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_84
timestamp 1586364061
transform 1 0 8832 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_88
timestamp 1586364061
transform 1 0 9200 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_84
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_88
timestamp 1586364061
transform 1 0 9200 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_96
timestamp 1586364061
transform 1 0 9936 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9384 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_100
timestamp 1586364061
transform 1 0 10304 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_105
timestamp 1586364061
transform 1 0 10764 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_101
timestamp 1586364061
transform 1 0 10396 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 10948 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_33_112
timestamp 1586364061
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_34_119
timestamp 1586364061
transform 1 0 12052 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_33_116
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 11040 0 -1 21216
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_34_125
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_132
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_142
timestamp 1586364061
transform 1 0 14168 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_138
timestamp 1586364061
transform 1 0 13800 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_136
timestamp 1586364061
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 13984 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12788 0 -1 21216
box -38 -48 1050 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 13984 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_149
timestamp 1586364061
transform 1 0 14812 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_146
timestamp 1586364061
transform 1 0 14536 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_149
timestamp 1586364061
transform 1 0 14812 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_156
timestamp 1586364061
transform 1 0 15456 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_33_153
timestamp 1586364061
transform 1 0 15180 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_34_169
timestamp 1586364061
transform 1 0 16652 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_165
timestamp 1586364061
transform 1 0 16284 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_168
timestamp 1586364061
transform 1 0 16560 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_173
timestamp 1586364061
transform 1 0 17020 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_176
timestamp 1586364061
transform 1 0 17296 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_172
timestamp 1586364061
transform 1 0 16928 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 16744 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 17112 0 1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 17112 0 -1 21216
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18676 0 -1 21216
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_180
timestamp 1586364061
transform 1 0 17664 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_195
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_183
timestamp 1586364061
transform 1 0 17940 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_34_188
timestamp 1586364061
transform 1 0 18400 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19872 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19872 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_199
timestamp 1586364061
transform 1 0 19412 0 1 20128
box -38 -48 314 592
use scs8hd_decap_6  FILLER_33_213
timestamp 1586364061
transform 1 0 20700 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_206
timestamp 1586364061
transform 1 0 20056 0 -1 21216
box -38 -48 774 592
use scs8hd_conb_1  _178_
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21436 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21252 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_230
timestamp 1586364061
transform 1 0 22264 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_34_218
timestamp 1586364061
transform 1 0 21160 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_222
timestamp 1586364061
transform 1 0 21528 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_242
timestamp 1586364061
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_234
timestamp 1586364061
transform 1 0 22632 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_246
timestamp 1586364061
transform 1 0 23736 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_258
timestamp 1586364061
transform 1 0 24840 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_4  FILLER_34_270
timestamp 1586364061
transform 1 0 25944 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_274
timestamp 1586364061
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 1 21216
box -38 -48 866 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3496 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3312 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_18
timestamp 1586364061
transform 1 0 2760 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_22
timestamp 1586364061
transform 1 0 3128 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_35
timestamp 1586364061
transform 1 0 4324 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 4508 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_71
timestamp 1586364061
transform 1 0 7636 0 1 21216
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_77
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_88
timestamp 1586364061
transform 1 0 9200 0 1 21216
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_92
timestamp 1586364061
transform 1 0 9568 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_95
timestamp 1586364061
transform 1 0 9844 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_105
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11500 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_111
timestamp 1586364061
transform 1 0 11316 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_115
timestamp 1586364061
transform 1 0 11684 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_119
timestamp 1586364061
transform 1 0 12052 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_132
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_136
timestamp 1586364061
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_140
timestamp 1586364061
transform 1 0 13984 0 1 21216
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14444 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_144
timestamp 1586364061
transform 1 0 14352 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_158
timestamp 1586364061
transform 1 0 15640 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 16376 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_162
timestamp 1586364061
transform 1 0 16008 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_175
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_179
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_195
timestamp 1586364061
transform 1 0 19044 0 1 21216
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_212
timestamp 1586364061
transform 1 0 20608 0 1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21804 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_217
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_223
timestamp 1586364061
transform 1 0 21620 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_227
timestamp 1586364061
transform 1 0 21988 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_239
timestamp 1586364061
transform 1 0 23092 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_243
timestamp 1586364061
transform 1 0 23460 0 1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_253
timestamp 1586364061
transform 1 0 24380 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_258
timestamp 1586364061
transform 1 0 24840 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_262
timestamp 1586364061
transform 1 0 25208 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_274
timestamp 1586364061
transform 1 0 26312 0 1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2668 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3496 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_19
timestamp 1586364061
transform 1 0 2852 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_23
timestamp 1586364061
transform 1 0 3220 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_36_28
timestamp 1586364061
transform 1 0 3680 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 406 592
use scs8hd_inv_8  _146_
timestamp 1586364061
transform 1 0 4416 0 -1 22304
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5980 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_45
timestamp 1586364061
transform 1 0 5244 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_49
timestamp 1586364061
transform 1 0 5612 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_8  FILLER_36_62
timestamp 1586364061
transform 1 0 6808 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  FILLER_36_70
timestamp 1586364061
transform 1 0 7544 0 -1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_84
timestamp 1586364061
transform 1 0 8832 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_96
timestamp 1586364061
transform 1 0 9936 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_100
timestamp 1586364061
transform 1 0 10304 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_3  FILLER_36_106
timestamp 1586364061
transform 1 0 10856 0 -1 22304
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 11132 0 -1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_120
timestamp 1586364061
transform 1 0 12144 0 -1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_137
timestamp 1586364061
transform 1 0 13708 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_149
timestamp 1586364061
transform 1 0 14812 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 130 592
use scs8hd_conb_1  _173_
timestamp 1586364061
transform 1 0 16928 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_164
timestamp 1586364061
transform 1 0 16192 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_168
timestamp 1586364061
transform 1 0 16560 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_8  FILLER_36_175
timestamp 1586364061
transform 1 0 17204 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_183
timestamp 1586364061
transform 1 0 17940 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_195
timestamp 1586364061
transform 1 0 19044 0 -1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_205
timestamp 1586364061
transform 1 0 19964 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_36_210
timestamp 1586364061
transform 1 0 20424 0 -1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_12  FILLER_36_224
timestamp 1586364061
transform 1 0 21712 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_236
timestamp 1586364061
transform 1 0 22816 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_248
timestamp 1586364061
transform 1 0 23920 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_260
timestamp 1586364061
transform 1 0 25024 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_272
timestamp 1586364061
transform 1 0 26128 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_inv_8  _144_
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_16
timestamp 1586364061
transform 1 0 2576 0 1 22304
box -38 -48 222 592
use scs8hd_buf_1  _158_
timestamp 1586364061
transform 1 0 3312 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2760 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 3772 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_20
timestamp 1586364061
transform 1 0 2944 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_31
timestamp 1586364061
transform 1 0 3956 0 1 22304
box -38 -48 774 592
use scs8hd_inv_8  _145_
timestamp 1586364061
transform 1 0 5152 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_41
timestamp 1586364061
transform 1 0 4876 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7176 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6992 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_69
timestamp 1586364061
transform 1 0 7452 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8188 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_73
timestamp 1586364061
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 10672 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 10488 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12052 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_113
timestamp 1586364061
transform 1 0 11500 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_117
timestamp 1586364061
transform 1 0 11868 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_121
timestamp 1586364061
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 13616 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 13984 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_132
timestamp 1586364061
transform 1 0 13248 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_138
timestamp 1586364061
transform 1 0 13800 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_142
timestamp 1586364061
transform 1 0 14168 0 1 22304
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_152
timestamp 1586364061
transform 1 0 15088 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_156
timestamp 1586364061
transform 1 0 15456 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_169
timestamp 1586364061
transform 1 0 16652 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_173
timestamp 1586364061
transform 1 0 17020 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_177
timestamp 1586364061
transform 1 0 17388 0 1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18216 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20056 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_197
timestamp 1586364061
transform 1 0 19228 0 1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_37_205
timestamp 1586364061
transform 1 0 19964 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21252 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21620 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_217
timestamp 1586364061
transform 1 0 21068 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_221
timestamp 1586364061
transform 1 0 21436 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_225
timestamp 1586364061
transform 1 0 21804 0 1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_37_231
timestamp 1586364061
transform 1 0 22356 0 1 22304
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_234
timestamp 1586364061
transform 1 0 22632 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_242
timestamp 1586364061
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_buf_2  _210_
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__210__A
timestamp 1586364061
transform 1 0 1932 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_7
timestamp 1586364061
transform 1 0 1748 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_11
timestamp 1586364061
transform 1 0 2116 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_18
timestamp 1586364061
transform 1 0 2760 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_30
timestamp 1586364061
transform 1 0 3864 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 590 592
use scs8hd_conb_1  _183_
timestamp 1586364061
transform 1 0 5704 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_38
timestamp 1586364061
transform 1 0 4600 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_42
timestamp 1586364061
transform 1 0 4968 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_46
timestamp 1586364061
transform 1 0 5336 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_38_53
timestamp 1586364061
transform 1 0 5980 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_61
timestamp 1586364061
transform 1 0 6716 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_65
timestamp 1586364061
transform 1 0 7084 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7820 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_76
timestamp 1586364061
transform 1 0 8096 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 774 592
use scs8hd_conb_1  _177_
timestamp 1586364061
transform 1 0 10396 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_8  FILLER_38_104
timestamp 1586364061
transform 1 0 10672 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_121
timestamp 1586364061
transform 1 0 12236 0 -1 23392
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 13616 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_125
timestamp 1586364061
transform 1 0 12604 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_135
timestamp 1586364061
transform 1 0 13524 0 -1 23392
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_163
timestamp 1586364061
transform 1 0 16100 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_167
timestamp 1586364061
transform 1 0 16468 0 -1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_180
timestamp 1586364061
transform 1 0 17664 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_38_191
timestamp 1586364061
transform 1 0 18676 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_195
timestamp 1586364061
transform 1 0 19044 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_38_207
timestamp 1586364061
transform 1 0 20148 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_213
timestamp 1586364061
transform 1 0 20700 0 -1 23392
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_38_224
timestamp 1586364061
transform 1 0 21712 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_235
timestamp 1586364061
transform 1 0 22724 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_247
timestamp 1586364061
transform 1 0 23828 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_259
timestamp 1586364061
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_271
timestamp 1586364061
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_6
timestamp 1586364061
transform 1 0 1656 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_7
timestamp 1586364061
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_11
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2300 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 314 592
use scs8hd_conb_1  _182_
timestamp 1586364061
transform 1 0 2392 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_17
timestamp 1586364061
transform 1 0 2668 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_39_22
timestamp 1586364061
transform 1 0 3128 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_18
timestamp 1586364061
transform 1 0 2760 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3496 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_29
timestamp 1586364061
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_29
timestamp 1586364061
transform 1 0 3772 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_33
timestamp 1586364061
transform 1 0 4140 0 1 23392
box -38 -48 1142 592
use scs8hd_buf_1  _110_
timestamp 1586364061
transform 1 0 5888 0 -1 24480
box -38 -48 314 592
use scs8hd_buf_2  _189_
timestamp 1586364061
transform 1 0 5612 0 1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_39_45
timestamp 1586364061
transform 1 0 5244 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_8  FILLER_40_55
timestamp 1586364061
transform 1 0 6164 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_57
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_71
timestamp 1586364061
transform 1 0 7636 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_66
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 6992 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7360 0 1 23392
box -38 -48 314 592
use scs8hd_buf_1  _136_
timestamp 1586364061
transform 1 0 6900 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_66
timestamp 1586364061
transform 1 0 7176 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_75
timestamp 1586364061
transform 1 0 8004 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_82
timestamp 1586364061
transform 1 0 8648 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_78
timestamp 1586364061
transform 1 0 8280 0 -1 24480
box -38 -48 1142 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 10488 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 10304 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 10488 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_90
timestamp 1586364061
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_101
timestamp 1586364061
transform 1 0 10396 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_104
timestamp 1586364061
transform 1 0 10672 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 11408 0 -1 24480
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_111
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_115
timestamp 1586364061
transform 1 0 11684 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_119
timestamp 1586364061
transform 1 0 12052 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_116
timestamp 1586364061
transform 1 0 11776 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_128
timestamp 1586364061
transform 1 0 12880 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_132
timestamp 1586364061
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _193_
timestamp 1586364061
transform 1 0 13248 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_140
timestamp 1586364061
transform 1 0 13984 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_136
timestamp 1586364061
transform 1 0 13616 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_3  FILLER_39_136
timestamp 1586364061
transform 1 0 13616 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 13892 0 1 23392
box -38 -48 222 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 14076 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_151
timestamp 1586364061
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_143
timestamp 1586364061
transform 1 0 14260 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_39_150
timestamp 1586364061
transform 1 0 14904 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_40_157
timestamp 1586364061
transform 1 0 15548 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_156
timestamp 1586364061
transform 1 0 15456 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 23392
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17296 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_169
timestamp 1586364061
transform 1 0 16652 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_173
timestamp 1586364061
transform 1 0 17020 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_178
timestamp 1586364061
transform 1 0 17480 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_40_162
timestamp 1586364061
transform 1 0 16008 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_168
timestamp 1586364061
transform 1 0 16560 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_188
timestamp 1586364061
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_192
timestamp 1586364061
transform 1 0 18768 0 1 23392
box -38 -48 774 592
use scs8hd_decap_8  FILLER_40_179
timestamp 1586364061
transform 1 0 17572 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 19688 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_200
timestamp 1586364061
transform 1 0 19504 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_206
timestamp 1586364061
transform 1 0 20056 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_210
timestamp 1586364061
transform 1 0 20424 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_214
timestamp 1586364061
transform 1 0 20792 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21712 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_218
timestamp 1586364061
transform 1 0 21160 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_222
timestamp 1586364061
transform 1 0 21528 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_226
timestamp 1586364061
transform 1 0 21896 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_218
timestamp 1586364061
transform 1 0 21160 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_230
timestamp 1586364061
transform 1 0 22264 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_39_238
timestamp 1586364061
transform 1 0 23000 0 1 23392
box -38 -48 590 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_242
timestamp 1586364061
transform 1 0 23368 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_258
timestamp 1586364061
transform 1 0 24840 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_262
timestamp 1586364061
transform 1 0 25208 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_254
timestamp 1586364061
transform 1 0 24472 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_266
timestamp 1586364061
transform 1 0 25576 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_274
timestamp 1586364061
transform 1 0 26312 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_274
timestamp 1586364061
transform 1 0 26312 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_6
timestamp 1586364061
transform 1 0 1656 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_10
timestamp 1586364061
transform 1 0 2024 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_22
timestamp 1586364061
transform 1 0 3128 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_34
timestamp 1586364061
transform 1 0 4232 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_46
timestamp 1586364061
transform 1 0 5336 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_41_58
timestamp 1586364061
transform 1 0 6440 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_114
timestamp 1586364061
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_118
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _200_
timestamp 1586364061
transform 1 0 12880 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 13432 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_127
timestamp 1586364061
transform 1 0 12788 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_132
timestamp 1586364061
transform 1 0 13248 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_136
timestamp 1586364061
transform 1 0 13616 0 1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14720 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15180 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_151
timestamp 1586364061
transform 1 0 14996 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_155
timestamp 1586364061
transform 1 0 15364 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_167
timestamp 1586364061
transform 1 0 16468 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_41_179
timestamp 1586364061
transform 1 0 17572 0 1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_42_112
timestamp 1586364061
transform 1 0 11408 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_116
timestamp 1586364061
transform 1 0 11776 0 -1 25568
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_128
timestamp 1586364061
transform 1 0 12880 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_140
timestamp 1586364061
transform 1 0 13984 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  FILLER_42_152
timestamp 1586364061
transform 1 0 15088 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 416 480 536 6 address[0]
port 0 nsew default input
rlabel metal2 s 570 27520 626 28000 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 1368 480 1488 6 address[2]
port 2 nsew default input
rlabel metal2 s 1766 27520 1822 28000 6 address[3]
port 3 nsew default input
rlabel metal3 s 0 2456 480 2576 6 address[4]
port 4 nsew default input
rlabel metal2 s 3054 27520 3110 28000 6 address[5]
port 5 nsew default input
rlabel metal2 s 4342 27520 4398 28000 6 address[6]
port 6 nsew default input
rlabel metal3 s 27520 552 28000 672 6 chanx_left_in[0]
port 7 nsew default input
rlabel metal3 s 0 3408 480 3528 6 chanx_left_in[1]
port 8 nsew default input
rlabel metal2 s 5630 27520 5686 28000 6 chanx_left_in[2]
port 9 nsew default input
rlabel metal2 s 5262 0 5318 480 6 chanx_left_in[3]
port 10 nsew default input
rlabel metal3 s 0 4496 480 4616 6 chanx_left_in[4]
port 11 nsew default input
rlabel metal3 s 27520 1776 28000 1896 6 chanx_left_in[5]
port 12 nsew default input
rlabel metal3 s 0 5584 480 5704 6 chanx_left_in[6]
port 13 nsew default input
rlabel metal2 s 7470 0 7526 480 6 chanx_left_in[7]
port 14 nsew default input
rlabel metal2 s 9586 0 9642 480 6 chanx_left_in[8]
port 15 nsew default input
rlabel metal2 s 11702 0 11758 480 6 chanx_left_out[0]
port 16 nsew default tristate
rlabel metal3 s 0 6536 480 6656 6 chanx_left_out[1]
port 17 nsew default tristate
rlabel metal3 s 27520 3136 28000 3256 6 chanx_left_out[2]
port 18 nsew default tristate
rlabel metal2 s 6918 27520 6974 28000 6 chanx_left_out[3]
port 19 nsew default tristate
rlabel metal3 s 27520 4496 28000 4616 6 chanx_left_out[4]
port 20 nsew default tristate
rlabel metal3 s 0 7624 480 7744 6 chanx_left_out[5]
port 21 nsew default tristate
rlabel metal3 s 27520 5856 28000 5976 6 chanx_left_out[6]
port 22 nsew default tristate
rlabel metal3 s 27520 7216 28000 7336 6 chanx_left_out[7]
port 23 nsew default tristate
rlabel metal3 s 0 8712 480 8832 6 chanx_left_out[8]
port 24 nsew default tristate
rlabel metal3 s 0 9664 480 9784 6 chanx_right_in[0]
port 25 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chanx_right_in[1]
port 26 nsew default input
rlabel metal2 s 8114 27520 8170 28000 6 chanx_right_in[2]
port 27 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_right_in[3]
port 28 nsew default input
rlabel metal2 s 9402 27520 9458 28000 6 chanx_right_in[4]
port 29 nsew default input
rlabel metal2 s 10690 27520 10746 28000 6 chanx_right_in[5]
port 30 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_right_in[6]
port 31 nsew default input
rlabel metal3 s 27520 8440 28000 8560 6 chanx_right_in[7]
port 32 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_right_in[8]
port 33 nsew default input
rlabel metal2 s 11978 27520 12034 28000 6 chanx_right_out[0]
port 34 nsew default tristate
rlabel metal2 s 13266 27520 13322 28000 6 chanx_right_out[1]
port 35 nsew default tristate
rlabel metal3 s 27520 9800 28000 9920 6 chanx_right_out[2]
port 36 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_right_out[3]
port 37 nsew default tristate
rlabel metal3 s 0 14832 480 14952 6 chanx_right_out[4]
port 38 nsew default tristate
rlabel metal3 s 27520 11160 28000 11280 6 chanx_right_out[5]
port 39 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_right_out[6]
port 40 nsew default tristate
rlabel metal2 s 16026 0 16082 480 6 chanx_right_out[7]
port 41 nsew default tristate
rlabel metal2 s 14554 27520 14610 28000 6 chanx_right_out[8]
port 42 nsew default tristate
rlabel metal3 s 0 17008 480 17128 6 chany_top_in[0]
port 43 nsew default input
rlabel metal3 s 0 17960 480 18080 6 chany_top_in[1]
port 44 nsew default input
rlabel metal3 s 27520 12520 28000 12640 6 chany_top_in[2]
port 45 nsew default input
rlabel metal2 s 15750 27520 15806 28000 6 chany_top_in[3]
port 46 nsew default input
rlabel metal3 s 0 19048 480 19168 6 chany_top_in[4]
port 47 nsew default input
rlabel metal2 s 17038 27520 17094 28000 6 chany_top_in[5]
port 48 nsew default input
rlabel metal2 s 18326 27520 18382 28000 6 chany_top_in[6]
port 49 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 chany_top_in[7]
port 50 nsew default input
rlabel metal2 s 18234 0 18290 480 6 chany_top_in[8]
port 51 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chany_top_out[0]
port 52 nsew default tristate
rlabel metal2 s 20350 0 20406 480 6 chany_top_out[1]
port 53 nsew default tristate
rlabel metal3 s 27520 15104 28000 15224 6 chany_top_out[2]
port 54 nsew default tristate
rlabel metal3 s 27520 16464 28000 16584 6 chany_top_out[3]
port 55 nsew default tristate
rlabel metal2 s 19614 27520 19670 28000 6 chany_top_out[4]
port 56 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chany_top_out[5]
port 57 nsew default tristate
rlabel metal2 s 20902 27520 20958 28000 6 chany_top_out[6]
port 58 nsew default tristate
rlabel metal3 s 27520 17824 28000 17944 6 chany_top_out[7]
port 59 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 chany_top_out[8]
port 60 nsew default tristate
rlabel metal2 s 3146 0 3202 480 6 data_in
port 61 nsew default input
rlabel metal2 s 1030 0 1086 480 6 enable
port 62 nsew default input
rlabel metal2 s 23386 27520 23442 28000 6 left_bottom_grid_pin_11_
port 63 nsew default input
rlabel metal3 s 27520 23128 28000 23248 6 left_bottom_grid_pin_13_
port 64 nsew default input
rlabel metal3 s 0 23128 480 23248 6 left_bottom_grid_pin_15_
port 65 nsew default input
rlabel metal3 s 27520 19184 28000 19304 6 left_bottom_grid_pin_1_
port 66 nsew default input
rlabel metal3 s 27520 20544 28000 20664 6 left_bottom_grid_pin_3_
port 67 nsew default input
rlabel metal2 s 22098 27520 22154 28000 6 left_bottom_grid_pin_5_
port 68 nsew default input
rlabel metal2 s 22466 0 22522 480 6 left_bottom_grid_pin_7_
port 69 nsew default input
rlabel metal3 s 27520 21768 28000 21888 6 left_bottom_grid_pin_9_
port 70 nsew default input
rlabel metal3 s 0 24216 480 24336 6 left_top_grid_pin_10_
port 71 nsew default input
rlabel metal3 s 0 26256 480 26376 6 right_bottom_grid_pin_11_
port 72 nsew default input
rlabel metal3 s 27520 25848 28000 25968 6 right_bottom_grid_pin_13_
port 73 nsew default input
rlabel metal3 s 27520 27208 28000 27328 6 right_bottom_grid_pin_15_
port 74 nsew default input
rlabel metal2 s 24674 27520 24730 28000 6 right_bottom_grid_pin_1_
port 75 nsew default input
rlabel metal2 s 24674 0 24730 480 6 right_bottom_grid_pin_3_
port 76 nsew default input
rlabel metal2 s 26790 0 26846 480 6 right_bottom_grid_pin_5_
port 77 nsew default input
rlabel metal3 s 27520 24488 28000 24608 6 right_bottom_grid_pin_7_
port 78 nsew default input
rlabel metal3 s 0 25304 480 25424 6 right_bottom_grid_pin_9_
port 79 nsew default input
rlabel metal2 s 25962 27520 26018 28000 6 right_top_grid_pin_10_
port 80 nsew default input
rlabel metal2 s 27250 27520 27306 28000 6 top_left_grid_pin_13_
port 81 nsew default input
rlabel metal3 s 0 27344 480 27464 6 top_right_grid_pin_11_
port 82 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 83 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 84 nsew default input
<< end >>
