* NGSPICE file created from sb_1__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

.subckt sb_1__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_left_grid_pin_13_ bottom_right_grid_pin_11_ chanx_left_in[0] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chanx_right_in[0] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chany_bottom_in[0]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_out[0] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] chany_top_in[0] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_out[0] chany_top_out[1] chany_top_out[2]
+ chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7]
+ chany_top_out[8] data_in enable left_bottom_grid_pin_12_ left_top_grid_pin_10_ right_bottom_grid_pin_12_
+ right_top_grid_pin_10_ top_left_grid_pin_13_ top_right_grid_pin_11_ vpwr vgnd
XFILLER_22_188 vpwr vgnd scs8hd_fill_2
XFILLER_22_144 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__203__B _199_/X vgnd vpwr scs8hd_diode_2
XFILLER_13_100 vgnd vpwr scs8hd_decap_3
XFILLER_9_159 vpwr vgnd scs8hd_fill_2
XFILLER_13_155 vgnd vpwr scs8hd_fill_1
XFILLER_13_199 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_203 vgnd vpwr scs8hd_decap_8
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_left_track_1.LATCH_6_.latch data_in mem_left_track_1.LATCH_6_.latch/Q _190_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_258 vgnd vpwr scs8hd_decap_4
XFILLER_27_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_114 vgnd vpwr scs8hd_decap_8
XFILLER_12_10 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _215_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__214__A _238_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_98 vpwr vgnd scs8hd_fill_2
XFILLER_37_73 vpwr vgnd scs8hd_fill_2
XFILLER_37_62 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_228 vpwr vgnd scs8hd_fill_2
XFILLER_33_217 vpwr vgnd scs8hd_fill_2
XFILLER_33_206 vpwr vgnd scs8hd_fill_2
XANTENNA__108__B _236_/A vgnd vpwr scs8hd_diode_2
X_277_ chany_top_in[0] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA__124__A _124_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_151 vgnd vpwr scs8hd_decap_3
XFILLER_5_173 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vpwr vgnd scs8hd_fill_2
XFILLER_5_195 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _241_/HI mem_bottom_track_17.LATCH_2_.latch/Q
+ mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_4_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_200_ _189_/A _199_/X _200_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__209__A _208_/X vgnd vpwr scs8hd_diode_2
XFILLER_15_228 vpwr vgnd scs8hd_fill_2
XFILLER_15_239 vgnd vpwr scs8hd_decap_3
X_131_ _131_/A _127_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_75 vgnd vpwr scs8hd_decap_3
XFILLER_2_154 vpwr vgnd scs8hd_fill_2
XFILLER_2_121 vgnd vpwr scs8hd_decap_4
XFILLER_0_79 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_11 vgnd vpwr scs8hd_decap_3
XFILLER_9_77 vgnd vpwr scs8hd_fill_1
XANTENNA__119__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_261 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _274_/A vgnd vpwr scs8hd_inv_1
Xmem_bottom_track_17.LATCH_2_.latch data_in mem_bottom_track_17.LATCH_2_.latch/Q _229_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_242 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__211__B _211_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_86 vgnd vpwr scs8hd_decap_4
XFILLER_7_213 vpwr vgnd scs8hd_fill_2
XFILLER_11_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
X_114_ _105_/A _238_/A _114_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_track_9.INVTX1_6_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_4_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_5_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__206__B _198_/X vgnd vpwr scs8hd_diode_2
XFILLER_29_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__222__A _238_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_87 vgnd vpwr scs8hd_decap_3
XFILLER_28_161 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[7] mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__132__A _109_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_150 vpwr vgnd scs8hd_fill_2
XFILLER_13_3 vpwr vgnd scs8hd_fill_2
XFILLER_34_197 vgnd vpwr scs8hd_decap_12
XFILLER_34_186 vgnd vpwr scs8hd_decap_8
XFILLER_34_175 vgnd vpwr scs8hd_decap_8
XFILLER_34_164 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_1_.latch data_in mem_right_track_8.LATCH_1_.latch/Q _161_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_153 vgnd vpwr scs8hd_decap_3
XFILLER_15_21 vpwr vgnd scs8hd_fill_2
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XFILLER_31_53 vpwr vgnd scs8hd_fill_2
XANTENNA__217__A _217_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_76 vgnd vpwr scs8hd_decap_3
XFILLER_0_263 vgnd vpwr scs8hd_decap_12
XFILLER_31_156 vgnd vpwr scs8hd_decap_4
XFILLER_31_134 vpwr vgnd scs8hd_fill_2
XANTENNA__127__A _127_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB _203_/Y vgnd vpwr scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_142 vgnd vpwr scs8hd_decap_4
XFILLER_16_175 vpwr vgnd scs8hd_fill_2
XFILLER_16_186 vgnd vpwr scs8hd_decap_3
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_track_8.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _241_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_123 vgnd vpwr scs8hd_decap_8
XFILLER_26_42 vpwr vgnd scs8hd_fill_2
XFILLER_13_123 vpwr vgnd scs8hd_fill_2
XFILLER_13_134 vpwr vgnd scs8hd_fill_2
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_127 vgnd vpwr scs8hd_decap_4
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_6_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_108 vgnd vpwr scs8hd_decap_6
XFILLER_10_137 vpwr vgnd scs8hd_fill_2
XFILLER_12_88 vgnd vpwr scs8hd_decap_4
XANTENNA__214__B _211_/B vgnd vpwr scs8hd_diode_2
XANTENNA__230__A _238_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_96 vpwr vgnd scs8hd_fill_2
XFILLER_37_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_41_262 vgnd vpwr scs8hd_decap_12
X_276_ chany_top_in[1] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_3_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _139_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_8.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[0] mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_6_.latch data_in mem_top_track_8.LATCH_6_.latch/Q _125_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_6_.latch data_in mem_right_track_0.LATCH_6_.latch/Q _143_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _251_/HI mem_top_track_8.LATCH_7_.latch/Q
+ mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_130_ _130_/A _131_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mem_right_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_98 vgnd vpwr scs8hd_decap_4
XANTENNA__225__A _225_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_36 vgnd vpwr scs8hd_decap_4
XFILLER_0_47 vgnd vpwr scs8hd_decap_4
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XANTENNA__135__A _135_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_259_ chanx_right_in[0] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_14_273 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_6_.latch_SLEEPB _167_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XFILLER_20_254 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_21 vpwr vgnd scs8hd_fill_2
XFILLER_34_64 vgnd vpwr scs8hd_decap_8
XFILLER_7_236 vpwr vgnd scs8hd_fill_2
X_113_ _134_/A _238_/A vgnd vpwr scs8hd_buf_1
XFILLER_11_254 vpwr vgnd scs8hd_fill_2
XFILLER_11_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _196_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_258 vpwr vgnd scs8hd_fill_2
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XFILLER_15_7 vgnd vpwr scs8hd_decap_3
Xmux_left_track_1.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[6] mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_8_.scs8hd_inv_1 chanx_left_in[8] mux_top_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__222__B _221_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_22 vpwr vgnd scs8hd_fill_2
XFILLER_4_206 vgnd vpwr scs8hd_decap_8
XFILLER_4_228 vpwr vgnd scs8hd_fill_2
XFILLER_29_53 vpwr vgnd scs8hd_fill_2
XFILLER_6_13 vgnd vpwr scs8hd_fill_1
XFILLER_34_110 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _223_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_184 vpwr vgnd scs8hd_fill_2
XFILLER_19_173 vpwr vgnd scs8hd_fill_2
XFILLER_34_154 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_187 vpwr vgnd scs8hd_fill_2
XFILLER_25_132 vpwr vgnd scs8hd_fill_2
XFILLER_31_10 vpwr vgnd scs8hd_fill_2
XFILLER_15_99 vpwr vgnd scs8hd_fill_2
XANTENNA__233__A _232_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_275 vpwr vgnd scs8hd_fill_2
XFILLER_16_121 vgnd vpwr scs8hd_decap_4
Xmux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_3_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_179 vpwr vgnd scs8hd_fill_2
XANTENNA__127__B _127_/B vgnd vpwr scs8hd_diode_2
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_154 vgnd vpwr scs8hd_fill_1
XFILLER_16_165 vgnd vpwr scs8hd_fill_1
XANTENNA__143__A _143_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_113 vgnd vpwr scs8hd_fill_1
XFILLER_22_102 vgnd vpwr scs8hd_decap_3
XFILLER_26_32 vpwr vgnd scs8hd_fill_2
XFILLER_26_65 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__228__A _236_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XFILLER_3_25 vpwr vgnd scs8hd_fill_2
XFILLER_3_14 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _270_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__138__A address[4] vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_7_.latch data_in mem_left_track_9.LATCH_7_.latch/Q _200_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_194 vpwr vgnd scs8hd_fill_2
XFILLER_27_227 vgnd vpwr scs8hd_decap_4
XFILLER_12_23 vgnd vpwr scs8hd_decap_4
XFILLER_12_45 vpwr vgnd scs8hd_fill_2
XFILLER_12_67 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__230__B _225_/X vgnd vpwr scs8hd_diode_2
XFILLER_37_31 vgnd vpwr scs8hd_decap_12
XFILLER_26_260 vgnd vpwr scs8hd_decap_12
XFILLER_41_274 vgnd vpwr scs8hd_decap_3
X_275_ chany_top_in[2] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_38_6 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_230 vgnd vpwr scs8hd_decap_4
Xmux_right_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[0] mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_263 vpwr vgnd scs8hd_fill_2
XFILLER_23_22 vpwr vgnd scs8hd_fill_2
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_167 vpwr vgnd scs8hd_fill_2
XANTENNA__135__B _135_/B vgnd vpwr scs8hd_diode_2
X_189_ _189_/A _191_/B _189_/Y vgnd vpwr scs8hd_nor2_4
X_258_ chanx_right_in[1] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_9_46 vpwr vgnd scs8hd_fill_2
XFILLER_9_57 vgnd vpwr scs8hd_fill_1
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA__151__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_20_266 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_34_43 vgnd vpwr scs8hd_decap_6
XFILLER_34_32 vgnd vpwr scs8hd_decap_8
XFILLER_18_66 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__236__A _236_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_211 vgnd vpwr scs8hd_decap_3
XFILLER_11_266 vpwr vgnd scs8hd_fill_2
X_112_ address[1] address[2] _084_/Y _134_/A vgnd vpwr scs8hd_or3_4
XFILLER_38_108 vgnd vpwr scs8hd_fill_1
XANTENNA__146__A _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_270 vgnd vpwr scs8hd_decap_4
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
XFILLER_37_130 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_6_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_32 vgnd vpwr scs8hd_decap_4
XFILLER_28_152 vgnd vpwr scs8hd_fill_1
XFILLER_34_122 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_177 vgnd vpwr scs8hd_decap_4
XFILLER_25_111 vpwr vgnd scs8hd_fill_2
XFILLER_0_232 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _240_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _147_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_11 vpwr vgnd scs8hd_fill_2
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_21_180 vgnd vpwr scs8hd_decap_3
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XANTENNA__228__B _225_/X vgnd vpwr scs8hd_diode_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_158 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_3_48 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__154__A _153_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_140 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_206 vpwr vgnd scs8hd_fill_2
XFILLER_5_7 vpwr vgnd scs8hd_fill_2
XFILLER_12_13 vgnd vpwr scs8hd_fill_1
XFILLER_18_206 vgnd vpwr scs8hd_decap_8
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_43 vgnd vpwr scs8hd_decap_12
XANTENNA__239__A _223_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_272 vgnd vpwr scs8hd_decap_3
XFILLER_18_239 vgnd vpwr scs8hd_decap_12
XFILLER_18_228 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_41_253 vpwr vgnd scs8hd_fill_2
X_274_ _274_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
Xmem_top_track_0.LATCH_0_.latch data_in mem_top_track_0.LATCH_0_.latch/Q _117_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__149__A _149_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_3_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_91 vgnd vpwr scs8hd_fill_1
Xmem_right_track_8.LATCH_7_.latch data_in mem_right_track_8.LATCH_7_.latch/Q _155_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_209 vpwr vgnd scs8hd_fill_2
XFILLER_23_275 vpwr vgnd scs8hd_fill_2
XFILLER_23_56 vgnd vpwr scs8hd_decap_3
XFILLER_2_179 vpwr vgnd scs8hd_fill_2
XFILLER_2_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_0_16 vgnd vpwr scs8hd_decap_4
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
Xmem_left_track_17.LATCH_3_.latch data_in mem_left_track_17.LATCH_3_.latch/Q _236_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_9_25 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_188_ _187_/X _191_/B vgnd vpwr scs8hd_buf_1
X_257_ chanx_right_in[2] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__151__B _150_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_234 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_3_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_45 vgnd vpwr scs8hd_fill_1
XANTENNA__236__B _236_/B vgnd vpwr scs8hd_diode_2
XANTENNA__252__A _252_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
X_111_ _105_/A _221_/A _111_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_205 vpwr vgnd scs8hd_fill_2
XANTENNA__146__B _147_/B vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _149_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_120 vpwr vgnd scs8hd_fill_2
XFILLER_37_175 vgnd vpwr scs8hd_decap_8
XFILLER_29_22 vgnd vpwr scs8hd_fill_1
XFILLER_29_11 vgnd vpwr scs8hd_decap_4
XFILLER_20_79 vpwr vgnd scs8hd_fill_2
XFILLER_20_68 vpwr vgnd scs8hd_fill_2
XFILLER_20_46 vgnd vpwr scs8hd_decap_3
XFILLER_28_142 vpwr vgnd scs8hd_fill_2
XFILLER_28_131 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_263 vgnd vpwr scs8hd_decap_12
XFILLER_3_252 vpwr vgnd scs8hd_fill_2
XFILLER_6_48 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__157__A _127_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_2_.latch data_in mem_bottom_track_1.LATCH_2_.latch/Q _171_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_31_78 vpwr vgnd scs8hd_fill_2
XFILLER_0_200 vgnd vpwr scs8hd_decap_4
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_259 vpwr vgnd scs8hd_fill_2
XFILLER_39_204 vgnd vpwr scs8hd_decap_12
XFILLER_22_148 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_192 vgnd vpwr scs8hd_decap_3
XFILLER_30_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_1_.latch data_in mem_left_track_1.LATCH_1_.latch/Q _195_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_23 vgnd vpwr scs8hd_decap_4
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XANTENNA__260__A _260_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_218 vgnd vpwr scs8hd_decap_12
XFILLER_8_152 vgnd vpwr scs8hd_fill_1
XFILLER_8_163 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__170__A _131_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_16.LATCH_2_.latch data_in mem_right_track_16.LATCH_2_.latch/Q _221_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_37_55 vgnd vpwr scs8hd_decap_6
XFILLER_18_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_37_77 vgnd vpwr scs8hd_decap_4
XANTENNA__239__B _236_/B vgnd vpwr scs8hd_diode_2
X_273_ chany_top_in[4] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_5_100 vpwr vgnd scs8hd_fill_2
XFILLER_5_111 vgnd vpwr scs8hd_decap_4
XANTENNA__255__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__149__B _149_/B vgnd vpwr scs8hd_diode_2
XFILLER_17_262 vpwr vgnd scs8hd_fill_2
XANTENNA__165__A _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_35 vpwr vgnd scs8hd_fill_2
XFILLER_2_125 vgnd vpwr scs8hd_fill_1
XFILLER_14_232 vgnd vpwr scs8hd_decap_3
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _187_/A _187_/X vgnd vpwr scs8hd_buf_1
X_256_ _256_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_110_ _109_/X _221_/A vgnd vpwr scs8hd_buf_1
XFILLER_11_235 vgnd vpwr scs8hd_decap_3
XFILLER_7_217 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_239_ _223_/A _236_/B _239_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA__162__B _153_/X vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_165 vpwr vgnd scs8hd_fill_2
XFILLER_28_154 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_9.LATCH_7_.latch_SLEEPB _177_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__263__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_3_275 vpwr vgnd scs8hd_fill_2
XFILLER_6_27 vpwr vgnd scs8hd_fill_2
XFILLER_19_154 vpwr vgnd scs8hd_fill_2
XFILLER_19_132 vgnd vpwr scs8hd_decap_3
XFILLER_20_8 vgnd vpwr scs8hd_fill_1
XFILLER_13_7 vpwr vgnd scs8hd_fill_2
XFILLER_34_168 vpwr vgnd scs8hd_fill_2
XFILLER_34_102 vgnd vpwr scs8hd_decap_8
XANTENNA__157__B _158_/B vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _149_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _206_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XANTENNA__083__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_15_25 vpwr vgnd scs8hd_fill_2
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
XFILLER_0_212 vgnd vpwr scs8hd_decap_3
XFILLER_31_138 vpwr vgnd scs8hd_fill_2
XANTENNA__258__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_102 vgnd vpwr scs8hd_decap_3
XFILLER_16_179 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_216 vgnd vpwr scs8hd_decap_12
XFILLER_21_90 vpwr vgnd scs8hd_fill_2
XANTENNA__168__A _127_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_92 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_271 vgnd vpwr scs8hd_decap_4
XFILLER_26_68 vpwr vgnd scs8hd_fill_2
XFILLER_26_46 vpwr vgnd scs8hd_fill_2
XFILLER_13_138 vpwr vgnd scs8hd_fill_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_0.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_160 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_90 vpwr vgnd scs8hd_fill_2
XANTENNA__170__B _165_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_241 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_89 vgnd vpwr scs8hd_decap_4
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_272_ chany_top_in[5] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
Xmem_right_track_0.LATCH_1_.latch data_in mem_right_track_0.LATCH_1_.latch/Q _148_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__271__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_1_.latch data_in mem_top_track_8.LATCH_1_.latch/Q _135_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_134 vpwr vgnd scs8hd_fill_2
XFILLER_5_156 vpwr vgnd scs8hd_fill_2
XFILLER_32_211 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_274 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__181__A _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vpwr vgnd scs8hd_fill_2
XANTENNA__091__A _119_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__266__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
X_255_ chanx_right_in[4] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_14_244 vpwr vgnd scs8hd_fill_2
X_186_ _152_/A _139_/B _152_/C _232_/D _187_/A vgnd vpwr scs8hd_or4_4
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[0] mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_1.INVTX1_6_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_25 vgnd vpwr scs8hd_decap_4
XANTENNA__086__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_258 vgnd vpwr scs8hd_decap_4
XFILLER_1_3 vgnd vpwr scs8hd_decap_6
Xmux_top_track_8.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[5] mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_238_ _238_/A _236_/B _238_/Y vgnd vpwr scs8hd_nor2_4
X_169_ _145_/A _165_/X _169_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_3 vgnd vpwr scs8hd_fill_1
XFILLER_37_100 vpwr vgnd scs8hd_fill_2
XFILLER_1_83 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_26 vpwr vgnd scs8hd_fill_2
XFILLER_29_79 vpwr vgnd scs8hd_fill_2
XFILLER_29_57 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB _210_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_243 vgnd vpwr scs8hd_fill_1
XFILLER_19_188 vgnd vpwr scs8hd_decap_4
XFILLER_19_177 vgnd vpwr scs8hd_decap_4
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
Xmem_top_track_0.LATCH_6_.latch data_in mem_top_track_0.LATCH_6_.latch/Q _099_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__173__B _165_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.LATCH_3_.latch data_in mem_bottom_track_9.LATCH_3_.latch/Q _181_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_117 vgnd vpwr scs8hd_decap_8
XFILLER_25_158 vpwr vgnd scs8hd_fill_2
XFILLER_25_136 vpwr vgnd scs8hd_fill_2
XFILLER_40_139 vgnd vpwr scs8hd_decap_12
XFILLER_40_128 vgnd vpwr scs8hd_decap_8
XFILLER_31_36 vpwr vgnd scs8hd_fill_2
XFILLER_31_25 vpwr vgnd scs8hd_fill_2
XFILLER_31_14 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__274__A _274_/A vgnd vpwr scs8hd_diode_2
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_158 vgnd vpwr scs8hd_decap_4
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_4_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_228 vgnd vpwr scs8hd_decap_12
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__184__A _149_/A vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_2_.latch data_in mem_left_track_9.LATCH_2_.latch/Q _205_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_3_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_36 vgnd vpwr scs8hd_decap_3
XANTENNA__094__A _093_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_172 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_7_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_8_.scs8hd_inv_1 left_bottom_grid_pin_12_ mux_left_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_29 vpwr vgnd scs8hd_fill_2
XFILLER_3_18 vpwr vgnd scs8hd_fill_2
XANTENNA__269__A _269_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_110 vpwr vgnd scs8hd_fill_2
XFILLER_8_198 vpwr vgnd scs8hd_fill_2
XANTENNA__179__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_27 vgnd vpwr scs8hd_fill_1
XFILLER_12_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB _227_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_68 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[1] mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_top_track_16.LATCH_3_.latch data_in mem_top_track_16.LATCH_3_.latch/Q _212_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__089__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_8
X_271_ chany_top_in[6] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__181__B _176_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_267 vgnd vpwr scs8hd_decap_8
XFILLER_23_245 vpwr vgnd scs8hd_fill_2
XFILLER_23_223 vgnd vpwr scs8hd_fill_1
XFILLER_3_7 vpwr vgnd scs8hd_fill_2
XFILLER_2_138 vgnd vpwr scs8hd_decap_4
XFILLER_2_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_14_201 vpwr vgnd scs8hd_fill_2
XANTENNA__282__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
X_254_ chanx_right_in[5] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_13_92 vpwr vgnd scs8hd_fill_2
X_185_ address[5] _150_/Y _232_/D vgnd vpwr scs8hd_or2_4
XANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_20_226 vgnd vpwr scs8hd_decap_6
XANTENNA__192__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_48 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_7_.latch data_in mem_left_track_1.LATCH_7_.latch/Q _189_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__277__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_8_.scs8hd_inv_1 chanx_left_in[4] mux_top_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_237_ _221_/A _236_/B _237_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_80 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_168_ _127_/A _165_/X _168_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_241 vgnd vpwr scs8hd_decap_4
XFILLER_6_274 vgnd vpwr scs8hd_fill_1
X_099_ _105_/A _124_/A _099_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_167 vpwr vgnd scs8hd_fill_2
XFILLER_37_156 vpwr vgnd scs8hd_fill_2
XFILLER_37_145 vpwr vgnd scs8hd_fill_2
XFILLER_37_134 vpwr vgnd scs8hd_fill_2
XFILLER_37_123 vgnd vpwr scs8hd_decap_4
XFILLER_37_112 vgnd vpwr scs8hd_decap_8
XANTENNA__187__A _187_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_95 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_6_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_112 vgnd vpwr scs8hd_decap_3
XFILLER_28_178 vpwr vgnd scs8hd_fill_2
XANTENNA__097__A _097_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_200 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_71 vpwr vgnd scs8hd_fill_2
XFILLER_19_112 vgnd vpwr scs8hd_fill_1
XFILLER_19_91 vpwr vgnd scs8hd_fill_2
XFILLER_35_90 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB _160_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_115 vgnd vpwr scs8hd_decap_4
XFILLER_15_38 vpwr vgnd scs8hd_fill_2
XFILLER_0_236 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_17.LATCH_3_.latch data_in mem_bottom_track_17.LATCH_3_.latch/Q _228_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_148 vgnd vpwr scs8hd_decap_4
XFILLER_31_118 vpwr vgnd scs8hd_fill_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_107 vgnd vpwr scs8hd_decap_6
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_7_50 vgnd vpwr scs8hd_fill_1
XFILLER_15_192 vpwr vgnd scs8hd_fill_2
XANTENNA__184__B _176_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_251 vgnd vpwr scs8hd_decap_4
XFILLER_26_15 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_59 vgnd vpwr scs8hd_decap_6
XFILLER_21_151 vgnd vpwr scs8hd_decap_3
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB _191_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_184 vgnd vpwr scs8hd_decap_4
XFILLER_29_251 vpwr vgnd scs8hd_fill_2
XANTENNA__285__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_12_184 vpwr vgnd scs8hd_fill_2
XFILLER_35_221 vgnd vpwr scs8hd_decap_12
XANTENNA__179__B _176_/X vgnd vpwr scs8hd_diode_2
XANTENNA__195__A _135_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_5_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_243 vpwr vgnd scs8hd_fill_2
XFILLER_26_232 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_2_.latch data_in mem_right_track_8.LATCH_2_.latch/Q _160_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_270_ _270_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB _218_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_243 vgnd vpwr scs8hd_fill_1
XFILLER_4_62 vpwr vgnd scs8hd_fill_2
XFILLER_4_191 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_128 vgnd vpwr scs8hd_fill_1
XFILLER_2_106 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[8] mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[5] mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_29 vpwr vgnd scs8hd_fill_2
XFILLER_14_213 vgnd vpwr scs8hd_fill_1
XFILLER_14_224 vgnd vpwr scs8hd_decap_8
X_253_ chanx_right_in[6] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_5_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_71 vgnd vpwr scs8hd_decap_3
X_184_ _149_/A _176_/A _184_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_7 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_6_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA__192__B _191_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_3_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_209 vpwr vgnd scs8hd_fill_2
XFILLER_11_216 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
X_236_ _236_/A _236_/B _236_/Y vgnd vpwr scs8hd_nor2_4
X_167_ _143_/A _165_/X _167_/Y vgnd vpwr scs8hd_nor2_4
X_098_ _097_/X _124_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_15 vgnd vpwr scs8hd_fill_1
XFILLER_28_146 vgnd vpwr scs8hd_decap_6
XFILLER_28_135 vpwr vgnd scs8hd_fill_2
XANTENNA__097__B _097_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB _236_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_7_.latch data_in mem_right_track_0.LATCH_7_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_7_.latch data_in mem_top_track_8.LATCH_7_.latch/Q _123_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_219_ _219_/A _221_/B _219_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_193 vpwr vgnd scs8hd_fill_2
XFILLER_33_160 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_149 vpwr vgnd scs8hd_fill_2
XFILLER_0_259 vpwr vgnd scs8hd_fill_2
XFILLER_0_226 vpwr vgnd scs8hd_fill_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_127 vpwr vgnd scs8hd_fill_2
XFILLER_16_138 vpwr vgnd scs8hd_fill_2
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _250_/HI mem_top_track_16.LATCH_2_.latch/Q
+ mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _245_/HI mem_left_track_9.LATCH_7_.latch/Q
+ mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_30_174 vgnd vpwr scs8hd_decap_4
XFILLER_30_141 vpwr vgnd scs8hd_fill_2
XFILLER_7_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _244_/HI mem_left_track_17.LATCH_2_.latch/Q
+ mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_29_263 vgnd vpwr scs8hd_fill_1
XFILLER_29_230 vgnd vpwr scs8hd_decap_6
XFILLER_29_274 vgnd vpwr scs8hd_decap_3
XFILLER_16_71 vpwr vgnd scs8hd_fill_2
XFILLER_16_82 vpwr vgnd scs8hd_fill_2
XFILLER_32_81 vgnd vpwr scs8hd_decap_3
XFILLER_8_123 vpwr vgnd scs8hd_fill_2
XFILLER_12_141 vgnd vpwr scs8hd_fill_1
XFILLER_12_152 vgnd vpwr scs8hd_fill_1
XFILLER_35_233 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__195__B _187_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_258 vpwr vgnd scs8hd_fill_2
XFILLER_5_104 vpwr vgnd scs8hd_fill_2
XFILLER_5_115 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_222 vpwr vgnd scs8hd_fill_2
XFILLER_32_203 vgnd vpwr scs8hd_decap_8
XFILLER_27_92 vgnd vpwr scs8hd_decap_3
XFILLER_17_266 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _260_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_4_85 vgnd vpwr scs8hd_decap_6
XFILLER_23_236 vpwr vgnd scs8hd_fill_2
XFILLER_23_203 vgnd vpwr scs8hd_decap_4
XFILLER_23_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_252_ _252_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_183_ _135_/A _176_/A _183_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_184 vpwr vgnd scs8hd_fill_2
XFILLER_1_173 vpwr vgnd scs8hd_fill_2
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_206 vgnd vpwr scs8hd_decap_6
XFILLER_9_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_235_ _219_/A _236_/B _235_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_93 vgnd vpwr scs8hd_decap_3
XFILLER_10_250 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_166_ _142_/A _165_/X _166_/Y vgnd vpwr scs8hd_nor2_4
X_097_ _097_/A _097_/B address[0] _097_/X vgnd vpwr scs8hd_or3_4
XFILLER_1_31 vpwr vgnd scs8hd_fill_2
XFILLER_1_42 vgnd vpwr scs8hd_decap_6
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XFILLER_1_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB _180_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_29_49 vpwr vgnd scs8hd_fill_2
XFILLER_29_38 vpwr vgnd scs8hd_fill_2
XFILLER_36_180 vgnd vpwr scs8hd_decap_8
XANTENNA__097__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_36_191 vgnd vpwr scs8hd_decap_12
XFILLER_3_235 vpwr vgnd scs8hd_fill_2
XFILLER_3_224 vpwr vgnd scs8hd_fill_2
XFILLER_3_213 vpwr vgnd scs8hd_fill_2
XFILLER_10_84 vgnd vpwr scs8hd_decap_4
XFILLER_34_139 vgnd vpwr scs8hd_decap_12
XFILLER_27_191 vpwr vgnd scs8hd_fill_2
XFILLER_19_169 vpwr vgnd scs8hd_fill_2
X_149_ _149_/A _149_/B _149_/Y vgnd vpwr scs8hd_nor2_4
X_218_ _218_/A _221_/B _218_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_249 vgnd vpwr scs8hd_decap_6
XFILLER_24_172 vgnd vpwr scs8hd_decap_4
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_94 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_7_96 vgnd vpwr scs8hd_fill_1
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_0.LATCH_6_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_60 vgnd vpwr scs8hd_decap_4
XFILLER_35_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_60 vgnd vpwr scs8hd_fill_1
XFILLER_17_245 vpwr vgnd scs8hd_fill_2
XFILLER_32_259 vgnd vpwr scs8hd_decap_12
XFILLER_32_248 vgnd vpwr scs8hd_decap_8
XFILLER_32_237 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _173_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_75 vpwr vgnd scs8hd_fill_2
XFILLER_23_226 vgnd vpwr scs8hd_fill_1
XFILLER_23_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_251_ _251_/HI _251_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_left_track_1.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_248 vpwr vgnd scs8hd_fill_2
X_182_ _147_/A _176_/X _182_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_141 vgnd vpwr scs8hd_decap_4
XANTENNA__100__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_270 vgnd vpwr scs8hd_decap_6
Xmux_top_track_8.INVTX1_2_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _240_/HI mem_bottom_track_1.LATCH_7_.latch/Q
+ mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_165_ _165_/A _165_/X vgnd vpwr scs8hd_buf_1
X_234_ _218_/A _236_/B _234_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_61 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB _213_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_222 vpwr vgnd scs8hd_fill_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
XFILLER_34_7 vgnd vpwr scs8hd_decap_12
X_096_ _094_/X _105_/A vgnd vpwr scs8hd_buf_1
Xmem_top_track_0.LATCH_1_.latch data_in mem_top_track_0.LATCH_1_.latch/Q _114_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_52 vgnd vpwr scs8hd_decap_4
XFILLER_10_96 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_19_137 vpwr vgnd scs8hd_fill_2
XFILLER_19_115 vpwr vgnd scs8hd_fill_2
XFILLER_19_104 vpwr vgnd scs8hd_fill_2
XFILLER_19_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_148_ _135_/A _149_/B _148_/Y vgnd vpwr scs8hd_nor2_4
X_217_ _217_/A _221_/B vgnd vpwr scs8hd_buf_1
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_192 vpwr vgnd scs8hd_fill_2
XFILLER_31_29 vgnd vpwr scs8hd_decap_4
Xmem_left_track_17.LATCH_4_.latch data_in mem_left_track_17.LATCH_4_.latch/Q _235_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_184 vgnd vpwr scs8hd_decap_4
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_107 vgnd vpwr scs8hd_decap_3
XFILLER_21_73 vpwr vgnd scs8hd_fill_2
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[0] mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_30_187 vgnd vpwr scs8hd_decap_3
XFILLER_30_154 vgnd vpwr scs8hd_decap_3
XPHY_4 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_9.INVTX1_8_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_184 vgnd vpwr scs8hd_fill_1
XFILLER_7_31 vpwr vgnd scs8hd_fill_2
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_7_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_29 vpwr vgnd scs8hd_fill_2
XFILLER_21_176 vpwr vgnd scs8hd_fill_2
XFILLER_12_121 vpwr vgnd scs8hd_fill_2
XFILLER_12_154 vpwr vgnd scs8hd_fill_2
XFILLER_12_165 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _230_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__103__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
XFILLER_35_213 vpwr vgnd scs8hd_fill_2
XFILLER_35_202 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_4_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_224 vgnd vpwr scs8hd_decap_8
XFILLER_26_202 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_3_.latch data_in mem_bottom_track_1.LATCH_3_.latch/Q _170_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_235 vpwr vgnd scs8hd_fill_2
XFILLER_17_202 vgnd vpwr scs8hd_decap_4
XFILLER_40_271 vgnd vpwr scs8hd_decap_4
XFILLER_4_54 vgnd vpwr scs8hd_decap_8
XFILLER_4_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_172 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_9.LATCH_6_.latch_SLEEPB _201_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_249 vgnd vpwr scs8hd_decap_3
XFILLER_14_205 vgnd vpwr scs8hd_decap_8
X_250_ _250_/HI _250_/LO vgnd vpwr scs8hd_conb_1
XFILLER_22_271 vgnd vpwr scs8hd_decap_4
X_181_ _131_/A _176_/X _181_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_13_41 vpwr vgnd scs8hd_fill_2
XFILLER_13_96 vpwr vgnd scs8hd_fill_2
Xmem_left_track_1.LATCH_2_.latch data_in mem_left_track_1.LATCH_2_.latch/Q _194_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_153 vgnd vpwr scs8hd_decap_3
XANTENNA__100__B _097_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[4] mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__201__A _124_/A vgnd vpwr scs8hd_diode_2
Xmem_right_track_16.LATCH_3_.latch data_in mem_right_track_16.LATCH_3_.latch/Q _220_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_233_ _232_/X _236_/B vgnd vpwr scs8hd_buf_1
X_164_ _163_/X _165_/A vgnd vpwr scs8hd_buf_1
XFILLER_24_84 vgnd vpwr scs8hd_decap_6
X_095_ _142_/A _094_/X _095_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_7 vpwr vgnd scs8hd_fill_2
XFILLER_37_149 vgnd vpwr scs8hd_decap_4
XFILLER_37_138 vgnd vpwr scs8hd_decap_4
XFILLER_1_11 vpwr vgnd scs8hd_fill_2
XFILLER_1_22 vpwr vgnd scs8hd_fill_2
XANTENNA__111__A _105_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_99 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_29_18 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[4] mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_259 vpwr vgnd scs8hd_fill_2
XFILLER_3_248 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_40 vpwr vgnd scs8hd_fill_2
X_147_ _147_/A _147_/B _147_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__106__A _097_/A vgnd vpwr scs8hd_diode_2
X_216_ _152_/A _139_/B _232_/C _152_/D _217_/A vgnd vpwr scs8hd_or4_4
XFILLER_18_3 vgnd vpwr scs8hd_decap_3
XFILLER_25_119 vgnd vpwr scs8hd_fill_1
XFILLER_18_171 vpwr vgnd scs8hd_fill_2
XFILLER_33_174 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_218 vgnd vpwr scs8hd_decap_8
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_52 vpwr vgnd scs8hd_fill_2
XFILLER_21_41 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_top_track_16.LATCH_3_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB _194_/Y vgnd vpwr scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_15_152 vgnd vpwr scs8hd_decap_3
XFILLER_7_10 vgnd vpwr scs8hd_fill_1
XFILLER_15_174 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_1.INVTX1_8_.scs8hd_inv_1 left_top_grid_pin_10_ mux_left_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_19 vgnd vpwr scs8hd_fill_1
XFILLER_21_111 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_266 vgnd vpwr scs8hd_decap_8
XFILLER_16_41 vpwr vgnd scs8hd_fill_2
XFILLER_16_52 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_3_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_148 vpwr vgnd scs8hd_fill_2
XFILLER_12_144 vpwr vgnd scs8hd_fill_2
XFILLER_12_188 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__103__B _097_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XFILLER_7_170 vpwr vgnd scs8hd_fill_2
XFILLER_7_181 vpwr vgnd scs8hd_fill_2
XFILLER_7_192 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB _221_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_247 vpwr vgnd scs8hd_fill_2
XFILLER_5_118 vpwr vgnd scs8hd_fill_2
XANTENNA__204__A _236_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_2_.scs8hd_inv_1 chany_top_in[7] mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__114__A _105_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_261 vgnd vpwr scs8hd_decap_12
XFILLER_31_250 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_20 vpwr vgnd scs8hd_fill_2
XFILLER_13_53 vgnd vpwr scs8hd_decap_4
X_180_ _145_/A _176_/X _180_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_198 vpwr vgnd scs8hd_fill_2
XANTENNA__100__C _084_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__109__A _097_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_254 vpwr vgnd scs8hd_fill_2
XFILLER_9_265 vpwr vgnd scs8hd_fill_2
XFILLER_34_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _243_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__201__B _199_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_232_ _139_/A _139_/B _232_/C _232_/D _232_/X vgnd vpwr scs8hd_or4_4
XFILLER_6_213 vgnd vpwr scs8hd_fill_1
X_094_ _093_/X _094_/X vgnd vpwr scs8hd_buf_1
X_163_ _232_/C _152_/D _139_/A _152_/B _163_/X vgnd vpwr scs8hd_or4_4
XANTENNA__111__B _221_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_2_.latch data_in mem_top_track_8.LATCH_2_.latch/Q _133_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _239_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_2_.latch data_in mem_right_track_0.LATCH_2_.latch/Q _147_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_117 vgnd vpwr scs8hd_decap_3
XFILLER_36_150 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_8.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_10 vpwr vgnd scs8hd_fill_2
XANTENNA__212__A _236_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_43 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_95 vgnd vpwr scs8hd_decap_3
XFILLER_35_73 vpwr vgnd scs8hd_fill_2
XFILLER_35_62 vpwr vgnd scs8hd_fill_2
X_215_ _223_/A _211_/B _215_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__122__A _135_/B vgnd vpwr scs8hd_diode_2
XANTENNA__106__B address[2] vgnd vpwr scs8hd_diode_2
X_146_ _131_/A _147_/B _146_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_6 vgnd vpwr scs8hd_decap_12
XFILLER_33_197 vgnd vpwr scs8hd_decap_6
XFILLER_33_164 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_0_208 vpwr vgnd scs8hd_fill_2
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__207__A _223_/A vgnd vpwr scs8hd_diode_2
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_30_145 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _094_/X vgnd vpwr scs8hd_diode_2
X_129_ _145_/A _127_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_99 vpwr vgnd scs8hd_fill_2
XFILLER_38_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_21_156 vgnd vpwr scs8hd_decap_4
XFILLER_21_134 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_4_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_4
Xmux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_75 vpwr vgnd scs8hd_fill_2
XFILLER_16_86 vpwr vgnd scs8hd_fill_2
XFILLER_32_96 vgnd vpwr scs8hd_decap_4
XFILLER_32_41 vpwr vgnd scs8hd_fill_2
XFILLER_8_127 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__103__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_37_19 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_7_.latch data_in mem_top_track_0.LATCH_7_.latch/Q _095_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__204__B _199_/X vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.LATCH_4_.latch data_in mem_bottom_track_9.LATCH_4_.latch/Q _180_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__220__A _236_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_52 vpwr vgnd scs8hd_fill_2
XFILLER_40_251 vgnd vpwr scs8hd_decap_4
XFILLER_32_218 vgnd vpwr scs8hd_decap_12
XANTENNA__114__B _238_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_23 vpwr vgnd scs8hd_fill_2
XFILLER_4_12 vpwr vgnd scs8hd_fill_2
XFILLER_4_152 vgnd vpwr scs8hd_fill_1
XANTENNA__130__A _130_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_7_.latch_SLEEPB _155_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_207 vgnd vpwr scs8hd_fill_1
XFILLER_31_273 vgnd vpwr scs8hd_decap_4
XANTENNA__215__A _223_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_76 vgnd vpwr scs8hd_decap_3
XFILLER_1_188 vgnd vpwr scs8hd_decap_4
XFILLER_1_177 vgnd vpwr scs8hd_decap_4
XFILLER_8_3 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_3_.latch data_in mem_left_track_9.LATCH_3_.latch/Q _204_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__109__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__125__A _143_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_6_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _183_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_192 vgnd vpwr scs8hd_decap_12
XFILLER_24_42 vpwr vgnd scs8hd_fill_2
X_162_ _149_/A _153_/X _162_/Y vgnd vpwr scs8hd_nor2_4
X_231_ _223_/A _225_/X _231_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_3_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_247 vpwr vgnd scs8hd_fill_2
XFILLER_6_258 vgnd vpwr scs8hd_decap_12
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
X_093_ _152_/A _152_/B _232_/C _139_/D _093_/X vgnd vpwr scs8hd_or4_4
Xmem_top_track_16.LATCH_4_.latch data_in mem_top_track_16.LATCH_4_.latch/Q _211_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XFILLER_1_79 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_239 vpwr vgnd scs8hd_fill_2
XFILLER_3_228 vpwr vgnd scs8hd_fill_2
XFILLER_3_217 vpwr vgnd scs8hd_fill_2
XFILLER_19_53 vgnd vpwr scs8hd_decap_4
XANTENNA__212__B _211_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_162 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_145_ _145_/A _147_/B _145_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_5_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_214_ _238_/A _211_/B _214_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__106__C _084_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_140 vgnd vpwr scs8hd_fill_1
XFILLER_33_143 vpwr vgnd scs8hd_fill_2
XFILLER_33_110 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_143 vpwr vgnd scs8hd_fill_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_4
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__207__B _198_/X vgnd vpwr scs8hd_diode_2
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__223__A _223_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_124 vpwr vgnd scs8hd_fill_2
XFILLER_30_102 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB _146_/Y vgnd vpwr scs8hd_diode_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XANTENNA__133__A _147_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_23 vpwr vgnd scs8hd_fill_2
XANTENNA__117__B _223_/A vgnd vpwr scs8hd_diode_2
X_128_ _103_/X _145_/A vgnd vpwr scs8hd_buf_1
Xmux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_213 vpwr vgnd scs8hd_fill_2
XANTENNA__218__A _218_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_102 vpwr vgnd scs8hd_fill_2
XFILLER_16_10 vpwr vgnd scs8hd_fill_2
XFILLER_32_86 vgnd vpwr scs8hd_decap_4
XFILLER_32_64 vgnd vpwr scs8hd_fill_1
XFILLER_8_106 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _103_/X vgnd vpwr scs8hd_diode_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__220__B _221_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_75 vpwr vgnd scs8hd_fill_2
XFILLER_17_249 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_27_97 vpwr vgnd scs8hd_fill_2
XFILLER_25_260 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_4_131 vpwr vgnd scs8hd_fill_2
XFILLER_4_142 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_79 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_17.LATCH_4_.latch data_in mem_bottom_track_17.LATCH_4_.latch/Q _227_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_219 vgnd vpwr scs8hd_decap_4
XFILLER_16_260 vgnd vpwr scs8hd_decap_4
XANTENNA__215__B _211_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_88 vpwr vgnd scs8hd_fill_2
XFILLER_38_30 vgnd vpwr scs8hd_fill_1
XFILLER_1_123 vgnd vpwr scs8hd_decap_3
XANTENNA__231__A _223_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_96 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__125__B _127_/B vgnd vpwr scs8hd_diode_2
XANTENNA__109__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_9_201 vpwr vgnd scs8hd_fill_2
XFILLER_9_223 vpwr vgnd scs8hd_fill_2
XFILLER_13_241 vgnd vpwr scs8hd_fill_1
XANTENNA__141__A _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _248_/HI mem_right_track_8.LATCH_7_.latch/Q
+ mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_24_76 vpwr vgnd scs8hd_fill_2
XFILLER_24_32 vgnd vpwr scs8hd_decap_3
XFILLER_6_215 vgnd vpwr scs8hd_decap_4
XFILLER_6_226 vgnd vpwr scs8hd_decap_4
XANTENNA__226__A _218_/A vgnd vpwr scs8hd_diode_2
X_161_ _135_/A _153_/X _161_/Y vgnd vpwr scs8hd_nor2_4
X_230_ _238_/A _225_/X _230_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_092_ address[5] address[6] _139_/D vgnd vpwr scs8hd_or2_4
XFILLER_37_108 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_3_.latch data_in mem_right_track_8.LATCH_3_.latch/Q _159_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__136__A _136_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_23 vpwr vgnd scs8hd_fill_2
XFILLER_10_67 vpwr vgnd scs8hd_fill_2
XFILLER_19_119 vgnd vpwr scs8hd_decap_3
XFILLER_19_108 vgnd vpwr scs8hd_decap_4
XFILLER_19_87 vpwr vgnd scs8hd_fill_2
XFILLER_19_65 vgnd vpwr scs8hd_decap_4
XFILLER_19_32 vpwr vgnd scs8hd_fill_2
XFILLER_35_53 vgnd vpwr scs8hd_decap_8
XFILLER_27_130 vgnd vpwr scs8hd_decap_3
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_144_ _127_/A _147_/B _144_/Y vgnd vpwr scs8hd_nor2_4
X_213_ _221_/A _211_/B _213_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_262 vgnd vpwr scs8hd_decap_12
XFILLER_2_251 vgnd vpwr scs8hd_decap_8
XFILLER_2_240 vgnd vpwr scs8hd_decap_8
XFILLER_18_196 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_5_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_9.INVTX1_2_.scs8hd_inv_1 chany_top_in[8] mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_188 vgnd vpwr scs8hd_fill_1
XFILLER_21_22 vpwr vgnd scs8hd_fill_2
XANTENNA__223__B _221_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_77 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_188 vpwr vgnd scs8hd_fill_2
X_127_ _127_/A _127_/B _127_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__133__B _127_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_13 vgnd vpwr scs8hd_fill_1
XFILLER_7_46 vgnd vpwr scs8hd_decap_4
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
XFILLER_7_79 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _278_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[5] mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_6_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA__218__B _221_/B vgnd vpwr scs8hd_diode_2
XFILLER_12_125 vgnd vpwr scs8hd_fill_1
XFILLER_12_169 vpwr vgnd scs8hd_fill_2
XFILLER_32_32 vgnd vpwr scs8hd_decap_6
XANTENNA__234__A _218_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_217 vpwr vgnd scs8hd_fill_2
XANTENNA__144__A _127_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_184 vgnd vpwr scs8hd_fill_1
XFILLER_26_206 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_3_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB _204_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_239 vpwr vgnd scs8hd_fill_2
XANTENNA__229__A _221_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_206 vgnd vpwr scs8hd_fill_1
XFILLER_25_272 vgnd vpwr scs8hd_decap_4
XFILLER_4_36 vgnd vpwr scs8hd_decap_3
XFILLER_4_154 vgnd vpwr scs8hd_decap_3
XFILLER_4_187 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _249_/HI mem_top_track_0.LATCH_7_.latch/Q
+ mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__139__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_242 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 chanx_right_in[5] mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__231__B _225_/X vgnd vpwr scs8hd_diode_2
XFILLER_13_231 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _249_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_3_.scs8hd_inv_1 right_bottom_grid_pin_12_ mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_205 vpwr vgnd scs8hd_fill_2
XANTENNA__226__B _225_/X vgnd vpwr scs8hd_diode_2
X_091_ _119_/A _232_/C vgnd vpwr scs8hd_buf_1
X_160_ _147_/A _158_/B _160_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__152__A _152_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_142 vgnd vpwr scs8hd_decap_8
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XANTENNA__237__A _221_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_175 vpwr vgnd scs8hd_fill_2
X_212_ _236_/A _211_/B _212_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
X_143_ _143_/A _147_/B _143_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_123 vgnd vpwr scs8hd_decap_4
XFILLER_18_175 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_178 vgnd vpwr scs8hd_decap_3
XFILLER_33_156 vpwr vgnd scs8hd_fill_2
XANTENNA__147__A _147_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_3_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_2_91 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[2] mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_1.INVTX1_8_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_56 vgnd vpwr scs8hd_decap_3
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_178 vgnd vpwr scs8hd_decap_3
Xmux_top_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_126_ _101_/A _127_/A vgnd vpwr scs8hd_buf_1
XFILLER_38_259 vgnd vpwr scs8hd_decap_12
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_38_204 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_29_259 vgnd vpwr scs8hd_decap_4
XFILLER_29_226 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _246_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XFILLER_12_137 vgnd vpwr scs8hd_decap_4
XFILLER_12_148 vgnd vpwr scs8hd_decap_4
XFILLER_16_45 vpwr vgnd scs8hd_fill_2
XFILLER_16_56 vpwr vgnd scs8hd_fill_2
XFILLER_32_77 vpwr vgnd scs8hd_fill_2
XANTENNA__234__B _236_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__144__B _147_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_174 vgnd vpwr scs8hd_decap_4
XFILLER_11_181 vpwr vgnd scs8hd_fill_2
X_109_ _097_/A address[2] address[0] _109_/X vgnd vpwr scs8hd_or3_4
XANTENNA__160__A _147_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_11 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_240 vpwr vgnd scs8hd_fill_2
XFILLER_17_218 vpwr vgnd scs8hd_fill_2
XANTENNA__229__B _225_/X vgnd vpwr scs8hd_diode_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_4_48 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_254 vgnd vpwr scs8hd_decap_4
XFILLER_31_232 vpwr vgnd scs8hd_fill_2
XFILLER_31_221 vpwr vgnd scs8hd_fill_2
XFILLER_31_210 vgnd vpwr scs8hd_decap_4
XANTENNA__139__B _139_/B vgnd vpwr scs8hd_diode_2
XANTENNA__155__A _142_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_13_24 vpwr vgnd scs8hd_fill_2
XFILLER_1_158 vpwr vgnd scs8hd_fill_2
XFILLER_1_114 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_1_169 vpwr vgnd scs8hd_fill_2
XFILLER_13_254 vpwr vgnd scs8hd_fill_2
XFILLER_13_276 vgnd vpwr scs8hd_fill_1
XFILLER_9_236 vpwr vgnd scs8hd_fill_2
XFILLER_9_258 vgnd vpwr scs8hd_decap_4
XFILLER_9_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_23 vgnd vpwr scs8hd_decap_4
XFILLER_24_12 vpwr vgnd scs8hd_fill_2
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_10_224 vgnd vpwr scs8hd_decap_3
XFILLER_10_246 vpwr vgnd scs8hd_fill_2
XFILLER_10_257 vgnd vpwr scs8hd_decap_12
X_090_ enable _119_/A vgnd vpwr scs8hd_inv_8
Xmux_right_track_0.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[7] mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_16 vgnd vpwr scs8hd_decap_4
XFILLER_1_27 vpwr vgnd scs8hd_fill_2
XFILLER_1_38 vpwr vgnd scs8hd_fill_2
XANTENNA__152__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_110 vgnd vpwr scs8hd_decap_8
XFILLER_36_154 vgnd vpwr scs8hd_fill_1
XFILLER_36_121 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_47 vgnd vpwr scs8hd_decap_3
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_154 vgnd vpwr scs8hd_fill_1
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XFILLER_35_77 vpwr vgnd scs8hd_fill_2
XFILLER_35_66 vgnd vpwr scs8hd_decap_4
XANTENNA__237__B _236_/B vgnd vpwr scs8hd_diode_2
X_142_ _142_/A _147_/B _142_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_187 vpwr vgnd scs8hd_fill_2
X_211_ _219_/A _211_/B _211_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__253__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_18_8 vpwr vgnd scs8hd_fill_2
XANTENNA__147__B _147_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_154 vgnd vpwr scs8hd_decap_4
XFILLER_18_143 vpwr vgnd scs8hd_fill_2
XANTENNA__163__A _232_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_179 vgnd vpwr scs8hd_decap_3
XFILLER_24_168 vpwr vgnd scs8hd_fill_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_135 vpwr vgnd scs8hd_fill_2
XFILLER_15_157 vgnd vpwr scs8hd_decap_4
XFILLER_30_149 vgnd vpwr scs8hd_decap_4
X_125_ _143_/A _127_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_7 vgnd vpwr scs8hd_decap_12
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XFILLER_21_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__158__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_238 vgnd vpwr scs8hd_decap_6
XFILLER_32_67 vgnd vpwr scs8hd_fill_1
XFILLER_32_45 vpwr vgnd scs8hd_fill_2
XFILLER_32_23 vgnd vpwr scs8hd_decap_8
Xmem_top_track_0.LATCH_2_.latch data_in mem_top_track_0.LATCH_2_.latch/Q _111_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_271 vgnd vpwr scs8hd_decap_4
X_108_ _105_/A _236_/A _108_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_3 vpwr vgnd scs8hd_fill_2
XANTENNA__160__B _158_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_230 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_274 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _283_/A vgnd vpwr scs8hd_inv_1
XFILLER_8_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.LATCH_5_.latch data_in mem_left_track_17.LATCH_5_.latch/Q _234_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_56 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_123 vpwr vgnd scs8hd_fill_2
XANTENNA__261__A _261_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_27 vpwr vgnd scs8hd_fill_2
XFILLER_4_16 vgnd vpwr scs8hd_decap_4
XANTENNA__139__C _152_/C vgnd vpwr scs8hd_diode_2
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__155__B _158_/B vgnd vpwr scs8hd_diode_2
XANTENNA__171__A _147_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_137 vpwr vgnd scs8hd_fill_2
XFILLER_8_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_7_.latch_SLEEPB _189_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__256__A _256_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_266 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_181 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__166__A _142_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_70 vpwr vgnd scs8hd_fill_2
XFILLER_39_163 vpwr vgnd scs8hd_fill_2
XFILLER_24_57 vpwr vgnd scs8hd_fill_2
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_10_269 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
X_287_ _287_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA__152__C _152_/C vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_4_.latch data_in mem_bottom_track_1.LATCH_4_.latch/Q _169_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A right_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_144 vpwr vgnd scs8hd_fill_2
X_141_ _149_/B _147_/B vgnd vpwr scs8hd_buf_1
X_210_ _218_/A _211_/B _210_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_210 vgnd vpwr scs8hd_decap_4
Xmux_right_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_4_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_114 vpwr vgnd scs8hd_fill_2
XFILLER_18_188 vpwr vgnd scs8hd_fill_2
XANTENNA__163__B _152_/D vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_3_.latch data_in mem_left_track_1.LATCH_3_.latch/Q _193_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_158 vgnd vpwr scs8hd_fill_1
XFILLER_24_147 vgnd vpwr scs8hd_decap_6
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_128 vgnd vpwr scs8hd_decap_4
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_124_ _124_/A _143_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_27 vpwr vgnd scs8hd_fill_2
XANTENNA__264__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_23_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_5_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__158__B _158_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_6 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.LATCH_4_.latch data_in mem_right_track_16.LATCH_4_.latch/Q _219_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__174__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_117 vpwr vgnd scs8hd_fill_2
XFILLER_20_161 vpwr vgnd scs8hd_fill_2
XANTENNA__084__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__259__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB _234_/Y vgnd vpwr scs8hd_diode_2
X_107_ _130_/A _236_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_110 vpwr vgnd scs8hd_fill_2
XFILLER_11_194 vpwr vgnd scs8hd_fill_2
XFILLER_34_242 vgnd vpwr scs8hd_decap_12
XFILLER_19_261 vpwr vgnd scs8hd_fill_2
XANTENNA__169__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_35 vpwr vgnd scs8hd_fill_2
XFILLER_27_24 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_27_79 vpwr vgnd scs8hd_fill_2
XFILLER_25_231 vgnd vpwr scs8hd_decap_3
XFILLER_4_146 vgnd vpwr scs8hd_decap_6
XFILLER_4_168 vpwr vgnd scs8hd_fill_2
XANTENNA__139__D _139_/D vgnd vpwr scs8hd_diode_2
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__171__B _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_37 vpwr vgnd scs8hd_fill_2
XFILLER_13_59 vpwr vgnd scs8hd_fill_2
XFILLER_1_149 vpwr vgnd scs8hd_fill_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_205 vgnd vpwr scs8hd_decap_3
XANTENNA__272__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__166__B _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr
+ scs8hd_diode_2
XANTENNA__182__A _147_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_153 vgnd vpwr scs8hd_decap_6
XFILLER_39_142 vpwr vgnd scs8hd_fill_2
XFILLER_39_131 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XANTENNA__092__A address[5] vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__267__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
X_286_ chany_bottom_in[0] chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_14_91 vgnd vpwr scs8hd_fill_1
XANTENNA__152__D _152_/D vgnd vpwr scs8hd_diode_2
XANTENNA__177__A _142_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vpwr vgnd scs8hd_fill_2
XFILLER_27_101 vpwr vgnd scs8hd_fill_2
XFILLER_19_69 vgnd vpwr scs8hd_fill_1
XFILLER_19_36 vpwr vgnd scs8hd_fill_2
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XANTENNA__087__A _189_/A vgnd vpwr scs8hd_diode_2
X_140_ _139_/X _149_/B vgnd vpwr scs8hd_buf_1
Xmux_bottom_track_9.INVTX1_2_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_233 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_4_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_269_ _269_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA__163__C _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_126 vgnd vpwr scs8hd_decap_6
XFILLER_2_83 vgnd vpwr scs8hd_decap_8
XFILLER_2_72 vpwr vgnd scs8hd_fill_2
XFILLER_21_37 vpwr vgnd scs8hd_fill_2
XFILLER_21_48 vpwr vgnd scs8hd_fill_2
XFILLER_30_107 vgnd vpwr scs8hd_decap_8
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_track_17.LATCH_4_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[2] mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_123_ _142_/A _127_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__280__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_11_81 vgnd vpwr scs8hd_decap_4
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XFILLER_21_107 vgnd vpwr scs8hd_decap_4
XANTENNA__174__B _139_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__190__A _143_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_6_.latch_SLEEPB _178_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_3_.latch data_in mem_top_track_8.LATCH_3_.latch/Q _131_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_right_track_0.LATCH_3_.latch data_in mem_right_track_0.LATCH_3_.latch/Q _146_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_195 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__275__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_11_151 vgnd vpwr scs8hd_decap_4
XFILLER_11_173 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _207_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_166 vpwr vgnd scs8hd_fill_2
XFILLER_7_188 vpwr vgnd scs8hd_fill_2
X_106_ _097_/A address[2] _084_/Y _130_/A vgnd vpwr scs8hd_or3_4
XFILLER_11_184 vgnd vpwr scs8hd_fill_1
XANTENNA__169__B _165_/X vgnd vpwr scs8hd_diode_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XFILLER_34_254 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_3_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__185__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_8_93 vgnd vpwr scs8hd_decap_4
XFILLER_25_210 vgnd vpwr scs8hd_decap_4
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XFILLER_25_276 vgnd vpwr scs8hd_fill_1
XANTENNA__095__A _142_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XFILLER_17_80 vpwr vgnd scs8hd_fill_2
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_224 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_49 vpwr vgnd scs8hd_fill_2
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__182__B _176_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_83 vpwr vgnd scs8hd_fill_2
XFILLER_6_209 vgnd vpwr scs8hd_decap_4
XFILLER_10_205 vpwr vgnd scs8hd_fill_2
XANTENNA__092__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_6_6 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__283__A _283_/A vgnd vpwr scs8hd_diode_2
X_285_ chany_bottom_in[1] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_14_70 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_5_.latch data_in mem_bottom_track_9.LATCH_5_.latch/Q _179_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__177__B _176_/X vgnd vpwr scs8hd_diode_2
XANTENNA__193__A _131_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XFILLER_19_15 vpwr vgnd scs8hd_fill_2
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_35_47 vgnd vpwr scs8hd_decap_3
XFILLER_27_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_201 vgnd vpwr scs8hd_decap_3
Xmux_left_track_1.INVTX1_2_.scs8hd_inv_1 chany_top_in[4] mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_127 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.INVTX1_5_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__278__A _278_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_102 vpwr vgnd scs8hd_fill_2
XFILLER_41_182 vgnd vpwr scs8hd_fill_1
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_25_91 vgnd vpwr scs8hd_decap_4
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_199_ _198_/X _199_/X vgnd vpwr scs8hd_buf_1
Xmem_left_track_9.LATCH_4_.latch data_in mem_left_track_9.LATCH_4_.latch/Q _203_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_268_ chanx_left_in[0] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA__163__D _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_3 vpwr vgnd scs8hd_fill_2
XANTENNA__188__A _187_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_5_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_8.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[1] mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__098__A _097_/X vgnd vpwr scs8hd_diode_2
XFILLER_23_171 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_122_ _135_/B _127_/B vgnd vpwr scs8hd_buf_1
Xmux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_60 vgnd vpwr scs8hd_fill_1
XFILLER_11_71 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB _211_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _242_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__174__C _152_/C vgnd vpwr scs8hd_diode_2
XANTENNA__190__B _191_/B vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_5_.latch data_in mem_top_track_16.LATCH_5_.latch/Q _210_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
XFILLER_28_252 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_134 vpwr vgnd scs8hd_fill_2
XFILLER_7_145 vpwr vgnd scs8hd_fill_2
X_105_ _105_/A _219_/A _105_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_178 vgnd vpwr scs8hd_fill_1
XFILLER_19_241 vgnd vpwr scs8hd_fill_1
XFILLER_34_266 vgnd vpwr scs8hd_decap_8
XANTENNA__185__B _150_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_72 vpwr vgnd scs8hd_fill_2
XFILLER_8_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__095__B _094_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_104 vpwr vgnd scs8hd_fill_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_236 vgnd vpwr scs8hd_decap_8
XFILLER_31_225 vgnd vpwr scs8hd_decap_4
XFILLER_31_214 vgnd vpwr scs8hd_fill_1
XANTENNA__286__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_16_211 vgnd vpwr scs8hd_decap_3
XFILLER_16_222 vgnd vpwr scs8hd_decap_4
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_track_0.LATCH_6_.latch_SLEEPB _099_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[4] mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__196__A _149_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_22_247 vgnd vpwr scs8hd_decap_3
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_214 vpwr vgnd scs8hd_fill_2
XFILLER_13_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_162 vpwr vgnd scs8hd_fill_2
XFILLER_0_173 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB _228_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_3_.scs8hd_inv_1 right_top_grid_pin_10_ mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_62 vgnd vpwr scs8hd_fill_1
XFILLER_8_262 vgnd vpwr scs8hd_decap_12
XFILLER_39_188 vpwr vgnd scs8hd_fill_2
XFILLER_24_38 vpwr vgnd scs8hd_fill_2
XFILLER_24_16 vpwr vgnd scs8hd_fill_2
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
X_284_ chany_bottom_in[2] chany_top_out[3] vgnd vpwr scs8hd_buf_2
Xmux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_6_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_70 vgnd vpwr scs8hd_decap_3
XFILLER_5_221 vpwr vgnd scs8hd_fill_2
XFILLER_5_254 vpwr vgnd scs8hd_fill_2
XFILLER_5_265 vgnd vpwr scs8hd_decap_12
XFILLER_14_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_169 vgnd vpwr scs8hd_decap_8
XFILLER_36_158 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__193__B _191_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_5_.latch data_in mem_bottom_track_17.LATCH_5_.latch/Q _226_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_158 vpwr vgnd scs8hd_fill_2
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_35_191 vpwr vgnd scs8hd_fill_2
XFILLER_33_139 vpwr vgnd scs8hd_fill_2
XFILLER_26_191 vgnd vpwr scs8hd_decap_4
XFILLER_18_147 vgnd vpwr scs8hd_decap_6
XFILLER_18_136 vgnd vpwr scs8hd_decap_4
XFILLER_18_125 vpwr vgnd scs8hd_fill_2
XFILLER_41_150 vgnd vpwr scs8hd_decap_12
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_267_ chanx_left_in[1] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
X_198_ _198_/A _198_/X vgnd vpwr scs8hd_buf_1
Xmux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_41 vpwr vgnd scs8hd_fill_2
XFILLER_32_183 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[3] mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_139 vpwr vgnd scs8hd_fill_2
XFILLER_23_150 vpwr vgnd scs8hd_fill_2
X_121_ _120_/X _135_/B vgnd vpwr scs8hd_buf_1
XANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_36_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__174__D _152_/D vgnd vpwr scs8hd_diode_2
XFILLER_29_209 vpwr vgnd scs8hd_fill_2
XANTENNA__199__A _198_/X vgnd vpwr scs8hd_diode_2
XFILLER_37_253 vpwr vgnd scs8hd_fill_2
XFILLER_37_220 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_4_.latch data_in mem_right_track_8.LATCH_4_.latch/Q _158_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.INVTX1_8_.scs8hd_inv_1 chanx_left_in[5] mux_right_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_8_.scs8hd_inv_1_A left_bottom_grid_pin_12_ vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_17.LATCH_0_.latch data_in mem_left_track_17.LATCH_0_.latch/Q _239_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_82 vpwr vgnd scs8hd_fill_2
X_104_ _103_/X _219_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mem_left_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_6 vgnd vpwr scs8hd_decap_4
XFILLER_8_40 vpwr vgnd scs8hd_fill_2
XFILLER_8_51 vpwr vgnd scs8hd_fill_2
XFILLER_6_190 vgnd vpwr scs8hd_decap_6
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_25_256 vpwr vgnd scs8hd_fill_2
XFILLER_40_259 vgnd vpwr scs8hd_decap_12
XFILLER_4_127 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_256 vpwr vgnd scs8hd_fill_2
XFILLER_16_267 vgnd vpwr scs8hd_decap_8
XFILLER_33_81 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB _192_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__196__B _187_/X vgnd vpwr scs8hd_diode_2
XFILLER_22_259 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_3_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_219 vpwr vgnd scs8hd_fill_2
XFILLER_13_237 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_196 vpwr vgnd scs8hd_fill_2
XFILLER_0_130 vpwr vgnd scs8hd_fill_2
XFILLER_28_81 vpwr vgnd scs8hd_fill_2
XFILLER_12_270 vgnd vpwr scs8hd_decap_4
XFILLER_8_274 vgnd vpwr scs8hd_fill_1
XFILLER_39_167 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB _219_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XFILLER_10_229 vgnd vpwr scs8hd_decap_4
X_283_ _283_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_14_83 vpwr vgnd scs8hd_fill_2
XFILLER_5_211 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[1] mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XFILLER_27_148 vgnd vpwr scs8hd_decap_6
XFILLER_27_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XFILLER_33_118 vpwr vgnd scs8hd_fill_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XFILLER_41_162 vgnd vpwr scs8hd_decap_12
X_266_ chanx_left_in[2] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_197_ _139_/A _152_/B _152_/C _232_/D _198_/A vgnd vpwr scs8hd_or4_4
XFILLER_24_107 vgnd vpwr scs8hd_decap_6
XFILLER_2_64 vpwr vgnd scs8hd_fill_2
XFILLER_2_53 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _279_/A vgnd vpwr scs8hd_inv_1
Xmux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _243_/HI mem_left_track_1.LATCH_7_.latch/Q
+ mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_17_181 vpwr vgnd scs8hd_fill_2
XFILLER_21_18 vpwr vgnd scs8hd_fill_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
XFILLER_23_184 vgnd vpwr scs8hd_decap_4
X_120_ _152_/A _139_/B _152_/C _139_/D _120_/X vgnd vpwr scs8hd_or4_4
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_184 vpwr vgnd scs8hd_fill_2
X_249_ _249_/HI _249_/LO vgnd vpwr scs8hd_conb_1
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB _237_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_165 vgnd vpwr scs8hd_decap_4
XFILLER_20_132 vpwr vgnd scs8hd_fill_2
XFILLER_28_232 vgnd vpwr scs8hd_fill_1
XFILLER_28_210 vgnd vpwr scs8hd_decap_4
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
XFILLER_11_198 vpwr vgnd scs8hd_fill_2
X_103_ address[1] _097_/B address[0] _103_/X vgnd vpwr scs8hd_or3_4
XFILLER_34_213 vgnd vpwr scs8hd_fill_1
XFILLER_19_265 vgnd vpwr scs8hd_decap_12
XFILLER_8_30 vgnd vpwr scs8hd_fill_1
XFILLER_27_39 vpwr vgnd scs8hd_fill_2
XFILLER_27_28 vpwr vgnd scs8hd_fill_2
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_25_268 vpwr vgnd scs8hd_fill_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_93 vpwr vgnd scs8hd_fill_2
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_271 vgnd vpwr scs8hd_decap_6
XFILLER_21_260 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XFILLER_28_93 vpwr vgnd scs8hd_fill_2
XFILLER_5_31 vpwr vgnd scs8hd_fill_2
XFILLER_39_179 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_282_ chany_bottom_in[4] chany_top_out[5] vgnd vpwr scs8hd_buf_2
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _265_/A vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_70 vgnd vpwr scs8hd_decap_12
XFILLER_36_138 vpwr vgnd scs8hd_fill_2
XANTENNA__101__A _101_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_35_39 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_83 vgnd vpwr scs8hd_decap_3
XFILLER_41_174 vgnd vpwr scs8hd_decap_8
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_25_72 vpwr vgnd scs8hd_fill_2
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
X_196_ _149_/A _187_/X _196_/Y vgnd vpwr scs8hd_nor2_4
X_265_ _265_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_32_163 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_130 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB _181_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_6
XFILLER_11_85 vgnd vpwr scs8hd_fill_1
XFILLER_36_60 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_141 vpwr vgnd scs8hd_fill_2
X_248_ _248_/HI _248_/LO vgnd vpwr scs8hd_conb_1
X_179_ _127_/A _176_/X _179_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_32_18 vpwr vgnd scs8hd_fill_2
XFILLER_20_199 vgnd vpwr scs8hd_decap_4
XFILLER_28_244 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_155 vgnd vpwr scs8hd_fill_1
X_102_ _105_/A _218_/A _102_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_177 vpwr vgnd scs8hd_fill_2
XFILLER_19_222 vpwr vgnd scs8hd_fill_2
XFILLER_19_233 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_214 vgnd vpwr scs8hd_fill_1
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_25_236 vpwr vgnd scs8hd_fill_2
XFILLER_31_217 vgnd vpwr scs8hd_fill_1
XFILLER_17_62 vgnd vpwr scs8hd_decap_3
XFILLER_17_84 vpwr vgnd scs8hd_fill_2
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_50 vpwr vgnd scs8hd_fill_2
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_184 vgnd vpwr scs8hd_decap_3
XANTENNA__104__A _103_/X vgnd vpwr scs8hd_diode_2
XFILLER_22_206 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_143 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_3_.latch data_in mem_top_track_0.LATCH_3_.latch/Q _108_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_210 vpwr vgnd scs8hd_fill_2
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_9.LATCH_0_.latch data_in mem_bottom_track_9.LATCH_0_.latch/Q _184_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_54 vpwr vgnd scs8hd_fill_2
XFILLER_5_87 vpwr vgnd scs8hd_fill_2
XFILLER_10_209 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_180 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_7_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
X_281_ chany_bottom_in[5] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_14_41 vgnd vpwr scs8hd_decap_4
XFILLER_14_52 vpwr vgnd scs8hd_fill_2
XFILLER_39_60 vgnd vpwr scs8hd_fill_1
XFILLER_30_84 vpwr vgnd scs8hd_fill_2
XFILLER_39_82 vgnd vpwr scs8hd_decap_12
XFILLER_36_106 vgnd vpwr scs8hd_fill_1
XFILLER_29_191 vgnd vpwr scs8hd_decap_4
XFILLER_29_180 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_2_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_19 vpwr vgnd scs8hd_fill_2
XANTENNA__202__A _218_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_7 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_106 vgnd vpwr scs8hd_decap_4
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_95 vgnd vpwr scs8hd_fill_1
XFILLER_25_62 vgnd vpwr scs8hd_fill_1
XFILLER_25_40 vpwr vgnd scs8hd_fill_2
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_264_ chanx_left_in[4] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
X_195_ _135_/A _187_/X _195_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_7 vgnd vpwr scs8hd_decap_12
XANTENNA__112__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_17_172 vgnd vpwr scs8hd_decap_3
XFILLER_32_186 vpwr vgnd scs8hd_fill_2
XFILLER_32_175 vgnd vpwr scs8hd_decap_8
XFILLER_32_142 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _214_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_175 vgnd vpwr scs8hd_fill_1
Xmem_top_track_16.LATCH_0_.latch data_in mem_top_track_16.LATCH_0_.latch/Q _215_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_42 vpwr vgnd scs8hd_fill_2
XFILLER_11_53 vgnd vpwr scs8hd_decap_4
XFILLER_11_97 vpwr vgnd scs8hd_fill_2
XFILLER_36_83 vpwr vgnd scs8hd_fill_2
XFILLER_36_72 vpwr vgnd scs8hd_fill_2
X_247_ _247_/HI _247_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__107__A _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_178_ _143_/A _176_/X _178_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_245 vgnd vpwr scs8hd_decap_8
XFILLER_28_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_178 vgnd vpwr scs8hd_decap_8
XFILLER_20_145 vgnd vpwr scs8hd_decap_6
Xmem_bottom_track_1.LATCH_5_.latch data_in mem_bottom_track_1.LATCH_5_.latch/Q _168_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_41 vpwr vgnd scs8hd_fill_2
XFILLER_7_138 vpwr vgnd scs8hd_fill_2
XFILLER_11_101 vpwr vgnd scs8hd_fill_2
XFILLER_11_134 vpwr vgnd scs8hd_fill_2
X_101_ _101_/A _218_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_149 vgnd vpwr scs8hd_decap_4
XFILLER_19_245 vpwr vgnd scs8hd_fill_2
XFILLER_8_32 vpwr vgnd scs8hd_fill_2
XFILLER_8_87 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_4_.scs8hd_inv_1 chanx_right_in[5] mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_left_track_1.LATCH_4_.latch data_in mem_left_track_1.LATCH_4_.latch/Q _192_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_108 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_9.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__210__A _218_/A vgnd vpwr scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_237 vgnd vpwr scs8hd_decap_8
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_73 vpwr vgnd scs8hd_fill_2
XFILLER_3_196 vpwr vgnd scs8hd_fill_2
XFILLER_3_174 vpwr vgnd scs8hd_fill_2
XFILLER_3_152 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_6 vgnd vpwr scs8hd_decap_4
XANTENNA__120__A _152_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_251 vpwr vgnd scs8hd_fill_2
XFILLER_22_229 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_4_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_38_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _231_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_right_track_16.LATCH_5_.latch data_in mem_right_track_16.LATCH_5_.latch/Q _218_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__205__A _221_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_62 vgnd vpwr scs8hd_decap_6
XFILLER_0_177 vpwr vgnd scs8hd_fill_2
XFILLER_12_251 vgnd vpwr scs8hd_decap_4
XFILLER_5_11 vgnd vpwr scs8hd_decap_3
XANTENNA__115__A address[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_0_.latch data_in mem_bottom_track_17.LATCH_0_.latch/Q _231_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_192 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB _202_/Y vgnd vpwr scs8hd_diode_2
X_280_ chany_bottom_in[6] chany_top_out[7] vgnd vpwr scs8hd_buf_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_5_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_5_236 vpwr vgnd scs8hd_fill_2
XFILLER_5_258 vgnd vpwr scs8hd_decap_4
XFILLER_14_97 vgnd vpwr scs8hd_fill_1
XFILLER_39_94 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__202__B _199_/X vgnd vpwr scs8hd_diode_2
XFILLER_2_206 vpwr vgnd scs8hd_fill_2
XFILLER_26_162 vgnd vpwr scs8hd_fill_1
XFILLER_26_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[0] mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_track_8.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_263_ chanx_left_in[5] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ _147_/A _191_/B _194_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_45 vgnd vpwr scs8hd_decap_8
XFILLER_2_23 vgnd vpwr scs8hd_decap_8
XFILLER_2_12 vgnd vpwr scs8hd_decap_8
XANTENNA__112__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_17_162 vgnd vpwr scs8hd_fill_1
XFILLER_17_184 vgnd vpwr scs8hd_decap_3
XFILLER_23_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__213__A _221_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[3] mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_154 vpwr vgnd scs8hd_fill_2
X_246_ _246_/HI _246_/LO vgnd vpwr scs8hd_conb_1
XFILLER_14_165 vpwr vgnd scs8hd_fill_2
XFILLER_14_176 vgnd vpwr scs8hd_decap_8
X_177_ _142_/A _176_/X _177_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__123__A _142_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XFILLER_20_157 vpwr vgnd scs8hd_fill_2
XFILLER_20_102 vpwr vgnd scs8hd_fill_2
XFILLER_9_180 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_224 vpwr vgnd scs8hd_fill_2
XFILLER_22_64 vpwr vgnd scs8hd_fill_2
XANTENNA__208__A _139_/A vgnd vpwr scs8hd_diode_2
X_100_ address[1] _097_/B _084_/Y _101_/A vgnd vpwr scs8hd_or3_4
XFILLER_22_86 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_1.LATCH_7_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_22 vpwr vgnd scs8hd_fill_2
XANTENNA__118__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_8_55 vpwr vgnd scs8hd_fill_2
X_229_ _221_/A _225_/X _229_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_227 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _195_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[8] mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__210__B _211_/B vgnd vpwr scs8hd_diode_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_260 vgnd vpwr scs8hd_decap_4
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_42 vpwr vgnd scs8hd_fill_2
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XFILLER_17_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _139_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_260 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__205__B _199_/X vgnd vpwr scs8hd_diode_2
XANTENNA__221__A _221_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _222_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_4
XFILLER_0_101 vgnd vpwr scs8hd_decap_4
XFILLER_28_85 vpwr vgnd scs8hd_fill_2
Xmem_right_track_0.LATCH_4_.latch data_in mem_right_track_0.LATCH_4_.latch/Q _145_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_top_track_8.LATCH_4_.latch data_in mem_top_track_8.LATCH_4_.latch/Q _129_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_245 vpwr vgnd scs8hd_fill_2
XFILLER_12_230 vgnd vpwr scs8hd_decap_4
XFILLER_12_274 vgnd vpwr scs8hd_fill_1
XANTENNA__115__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_39_149 vpwr vgnd scs8hd_fill_2
XFILLER_39_138 vpwr vgnd scs8hd_fill_2
XFILLER_39_127 vpwr vgnd scs8hd_fill_2
XANTENNA__131__A _131_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_2_.scs8hd_inv_1 chany_top_in[7] mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_10 vgnd vpwr scs8hd_fill_1
XFILLER_14_87 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_top_track_16.LATCH_5_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_5_215 vgnd vpwr scs8hd_decap_4
XANTENNA__216__A _152_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_40 vgnd vpwr scs8hd_fill_1
XANTENNA__126__A _101_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_229 vpwr vgnd scs8hd_fill_2
XFILLER_2_218 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
Xmux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_5_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_174 vpwr vgnd scs8hd_fill_2
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_18_119 vgnd vpwr scs8hd_decap_4
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
X_193_ _131_/A _191_/B _193_/Y vgnd vpwr scs8hd_nor2_4
X_262_ chanx_left_in[6] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__112__C _084_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_68 vpwr vgnd scs8hd_fill_2
XFILLER_32_199 vpwr vgnd scs8hd_fill_2
XFILLER_32_111 vgnd vpwr scs8hd_fill_1
XFILLER_32_100 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_199 vpwr vgnd scs8hd_fill_2
XANTENNA__213__B _211_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_77 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_track_1.LATCH_4_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_96 vgnd vpwr scs8hd_decap_8
Xmux_right_track_0.INVTX1_8_.scs8hd_inv_1 chanx_left_in[4] mux_right_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_111 vpwr vgnd scs8hd_fill_2
X_245_ _245_/HI _245_/LO vgnd vpwr scs8hd_conb_1
X_176_ _176_/A _176_/X vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__123__B _127_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_9.LATCH_6_.latch data_in mem_bottom_track_9.LATCH_6_.latch/Q _178_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__208__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XFILLER_11_158 vgnd vpwr scs8hd_decap_4
XANTENNA__224__A _152_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_159_ _131_/A _158_/B _159_/Y vgnd vpwr scs8hd_nor2_4
X_228_ _236_/A _225_/X _228_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__134__A _134_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_217 vgnd vpwr scs8hd_fill_1
Xmem_left_track_9.LATCH_5_.latch data_in mem_left_track_9.LATCH_5_.latch/Q _202_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _244_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_206 vgnd vpwr scs8hd_decap_3
XFILLER_17_21 vpwr vgnd scs8hd_fill_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__219__A _219_/A vgnd vpwr scs8hd_diode_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_97 vpwr vgnd scs8hd_fill_2
XANTENNA__120__C _152_/C vgnd vpwr scs8hd_diode_2
XANTENNA__129__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_272 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__221__B _221_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_97 vgnd vpwr scs8hd_decap_6
XANTENNA__131__B _127_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_35 vpwr vgnd scs8hd_fill_2
XANTENNA__115__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_39_106 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_3_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_6_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_66 vpwr vgnd scs8hd_fill_2
XANTENNA__216__B _139_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_43 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_4
XANTENNA__232__A _139_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _142_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_164 vpwr vgnd scs8hd_fill_2
XFILLER_35_153 vpwr vgnd scs8hd_fill_2
XFILLER_35_142 vpwr vgnd scs8hd_fill_2
XFILLER_35_120 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_6_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_175 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.INVTX1_5_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_197 vpwr vgnd scs8hd_fill_2
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_76 vpwr vgnd scs8hd_fill_2
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XANTENNA__227__A _219_/A vgnd vpwr scs8hd_diode_2
XPHY_32 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_261_ _261_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_25_98 vpwr vgnd scs8hd_fill_2
X_192_ _145_/A _191_/B _192_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_263 vpwr vgnd scs8hd_fill_2
XFILLER_1_252 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _184_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_142 vpwr vgnd scs8hd_fill_2
XFILLER_32_123 vpwr vgnd scs8hd_fill_2
XANTENNA__137__A _149_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_145 vgnd vpwr scs8hd_decap_3
XFILLER_23_178 vgnd vpwr scs8hd_decap_3
XFILLER_23_167 vpwr vgnd scs8hd_fill_2
XFILLER_11_12 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_64 vgnd vpwr scs8hd_decap_8
X_244_ _244_/HI _244_/LO vgnd vpwr scs8hd_conb_1
XFILLER_14_123 vpwr vgnd scs8hd_fill_2
XFILLER_14_145 vgnd vpwr scs8hd_decap_8
X_175_ _175_/A _176_/A vgnd vpwr scs8hd_buf_1
XFILLER_9_193 vpwr vgnd scs8hd_fill_2
XFILLER_28_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__208__C _232_/C vgnd vpwr scs8hd_diode_2
XFILLER_22_22 vgnd vpwr scs8hd_decap_4
XANTENNA__224__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_218 vgnd vpwr scs8hd_decap_12
XFILLER_27_270 vgnd vpwr scs8hd_decap_6
XFILLER_19_237 vgnd vpwr scs8hd_decap_4
XFILLER_19_226 vpwr vgnd scs8hd_fill_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XFILLER_8_68 vpwr vgnd scs8hd_fill_2
XFILLER_8_79 vpwr vgnd scs8hd_fill_2
X_227_ _219_/A _225_/X _227_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_152 vgnd vpwr scs8hd_fill_1
X_158_ _145_/A _158_/B _158_/Y vgnd vpwr scs8hd_nor2_4
X_089_ address[3] _152_/B vgnd vpwr scs8hd_buf_1
XANTENNA__150__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__219__B _221_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_218 vpwr vgnd scs8hd_fill_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_54 vgnd vpwr scs8hd_decap_4
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__235__A _219_/A vgnd vpwr scs8hd_diode_2
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__120__D _139_/D vgnd vpwr scs8hd_diode_2
XANTENNA__129__B _127_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_43 vpwr vgnd scs8hd_fill_2
XFILLER_28_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_147 vgnd vpwr scs8hd_decap_8
XFILLER_0_125 vgnd vpwr scs8hd_decap_3
Xmem_right_track_8.LATCH_5_.latch data_in mem_right_track_8.LATCH_5_.latch/Q _157_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _246_/HI mem_right_track_0.LATCH_7_.latch/Q
+ mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_8_203 vgnd vpwr scs8hd_decap_4
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_58 vgnd vpwr scs8hd_decap_3
XFILLER_39_118 vgnd vpwr scs8hd_decap_4
XFILLER_10_6 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_3_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_left_track_17.LATCH_1_.latch data_in mem_left_track_17.LATCH_1_.latch/Q _238_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__216__C _232_/C vgnd vpwr scs8hd_diode_2
XFILLER_14_23 vpwr vgnd scs8hd_fill_2
XFILLER_14_45 vgnd vpwr scs8hd_fill_1
XFILLER_14_56 vgnd vpwr scs8hd_fill_1
XFILLER_30_88 vgnd vpwr scs8hd_decap_4
XFILLER_30_66 vpwr vgnd scs8hd_fill_2
XANTENNA__232__B _139_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_173 vgnd vpwr scs8hd_decap_4
XFILLER_29_151 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _247_/HI mem_right_track_16.LATCH_2_.latch/Q
+ mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__142__B _147_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_198 vpwr vgnd scs8hd_fill_2
XFILLER_35_187 vpwr vgnd scs8hd_fill_2
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_154 vgnd vpwr scs8hd_decap_8
XFILLER_26_143 vgnd vpwr scs8hd_decap_8
XFILLER_25_11 vpwr vgnd scs8hd_fill_2
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_260_ _260_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XANTENNA__227__B _225_/X vgnd vpwr scs8hd_diode_2
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
X_191_ _127_/A _191_/B _191_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_1_275 vpwr vgnd scs8hd_fill_2
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XFILLER_32_157 vgnd vpwr scs8hd_decap_6
XFILLER_32_146 vgnd vpwr scs8hd_fill_1
XANTENNA__137__B _135_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_198 vpwr vgnd scs8hd_fill_2
XANTENNA__153__A _152_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_102 vgnd vpwr scs8hd_fill_1
XFILLER_11_24 vpwr vgnd scs8hd_fill_2
XFILLER_11_46 vpwr vgnd scs8hd_fill_2
XFILLER_11_57 vgnd vpwr scs8hd_fill_1
XFILLER_36_87 vgnd vpwr scs8hd_decap_4
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XANTENNA__238__A _238_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_0_.latch data_in mem_bottom_track_1.LATCH_0_.latch/Q _173_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_243_ _243_/HI _243_/LO vgnd vpwr scs8hd_conb_1
X_174_ _139_/A _139_/B _152_/C _152_/D _175_/A vgnd vpwr scs8hd_or4_4
XFILLER_28_7 vpwr vgnd scs8hd_fill_2
XANTENNA__148__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_116 vgnd vpwr scs8hd_fill_1
XFILLER_9_172 vpwr vgnd scs8hd_fill_2
XANTENNA__208__D _139_/D vgnd vpwr scs8hd_diode_2
XFILLER_11_138 vpwr vgnd scs8hd_fill_2
XFILLER_22_78 vpwr vgnd scs8hd_fill_2
XFILLER_22_45 vpwr vgnd scs8hd_fill_2
XANTENNA__224__C _232_/C vgnd vpwr scs8hd_diode_2
XFILLER_19_205 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_249 vgnd vpwr scs8hd_decap_3
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_157_ _127_/A _158_/B _157_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_8_36 vpwr vgnd scs8hd_fill_2
X_226_ _218_/A _225_/X _226_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_186 vpwr vgnd scs8hd_fill_2
X_088_ address[4] _152_/A vgnd vpwr scs8hd_buf_1
XFILLER_19_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_67 vpwr vgnd scs8hd_fill_2
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_77 vgnd vpwr scs8hd_decap_4
XFILLER_33_33 vpwr vgnd scs8hd_fill_2
XFILLER_33_11 vpwr vgnd scs8hd_fill_2
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_right_track_16.LATCH_0_.latch data_in mem_right_track_16.LATCH_0_.latch/Q _223_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__235__B _236_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_178 vgnd vpwr scs8hd_decap_3
XFILLER_3_156 vpwr vgnd scs8hd_fill_2
XFILLER_3_123 vgnd vpwr scs8hd_decap_3
XFILLER_3_101 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_5_.scs8hd_inv_1 chanx_left_in[1] mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__145__B _147_/B vgnd vpwr scs8hd_diode_2
X_209_ _208_/X _211_/B vgnd vpwr scs8hd_buf_1
XANTENNA__161__A _135_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_211 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_12_211 vgnd vpwr scs8hd_fill_1
XFILLER_8_226 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB _205_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_48 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__156__A _143_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_13 vgnd vpwr scs8hd_fill_1
XFILLER_30_23 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _245_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__216__D _152_/D vgnd vpwr scs8hd_diode_2
XFILLER_39_10 vgnd vpwr scs8hd_decap_12
XANTENNA__232__C _232_/C vgnd vpwr scs8hd_diode_2
XFILLER_4_251 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
X_190_ _143_/A _191_/B _190_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_23 vpwr vgnd scs8hd_fill_2
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XFILLER_1_210 vpwr vgnd scs8hd_fill_2
XFILLER_1_243 vgnd vpwr scs8hd_fill_1
XFILLER_1_232 vgnd vpwr scs8hd_decap_4
XFILLER_1_221 vgnd vpwr scs8hd_decap_4
XFILLER_32_103 vgnd vpwr scs8hd_decap_8
XFILLER_17_155 vgnd vpwr scs8hd_decap_4
XFILLER_17_177 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_2_.scs8hd_inv_1 chany_top_in[4] mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
XFILLER_36_77 vgnd vpwr scs8hd_decap_4
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XANTENNA__238__B _236_/B vgnd vpwr scs8hd_diode_2
X_242_ _242_/HI _242_/LO vgnd vpwr scs8hd_conb_1
XFILLER_22_180 vgnd vpwr scs8hd_decap_8
X_173_ _149_/A _165_/A _173_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__254__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__148__B _149_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_128 vpwr vgnd scs8hd_fill_2
XFILLER_20_106 vgnd vpwr scs8hd_decap_8
XANTENNA__164__A _163_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_92 vgnd vpwr scs8hd_decap_3
XFILLER_28_228 vgnd vpwr scs8hd_decap_4
XFILLER_28_206 vpwr vgnd scs8hd_fill_2
XFILLER_22_68 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__224__D _232_/D vgnd vpwr scs8hd_diode_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
XFILLER_34_209 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_225_ _225_/A _225_/X vgnd vpwr scs8hd_buf_1
X_087_ _189_/A _142_/A vgnd vpwr scs8hd_buf_1
Xmux_bottom_track_1.INVTX1_7_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_154 vpwr vgnd scs8hd_fill_2
X_156_ _143_/A _158_/B _156_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_8_26 vpwr vgnd scs8hd_fill_2
XFILLER_10_150 vgnd vpwr scs8hd_fill_1
XFILLER_10_194 vpwr vgnd scs8hd_fill_2
XANTENNA__159__A _131_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_6_.scs8hd_inv_1 chanx_left_in[2] mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_220 vpwr vgnd scs8hd_fill_2
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_135 vpwr vgnd scs8hd_fill_2
XFILLER_30_267 vgnd vpwr scs8hd_decap_8
XFILLER_30_256 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_139_ _139_/A _139_/B _152_/C _139_/D _139_/X vgnd vpwr scs8hd_or4_4
XANTENNA__161__B _153_/X vgnd vpwr scs8hd_diode_2
X_208_ _139_/A _152_/B _232_/C _139_/D _208_/X vgnd vpwr scs8hd_or4_4
XFILLER_2_190 vgnd vpwr scs8hd_decap_8
XFILLER_21_201 vpwr vgnd scs8hd_fill_2
XFILLER_0_71 vpwr vgnd scs8hd_fill_2
XFILLER_21_267 vpwr vgnd scs8hd_fill_2
XFILLER_21_256 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_91 vpwr vgnd scs8hd_fill_2
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_28_89 vgnd vpwr scs8hd_decap_3
XFILLER_28_23 vpwr vgnd scs8hd_fill_2
XFILLER_28_12 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_234 vgnd vpwr scs8hd_fill_1
XANTENNA__262__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_5_16 vgnd vpwr scs8hd_decap_4
XFILLER_8_249 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__156__B _158_/B vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _135_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__082__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_39_66 vpwr vgnd scs8hd_fill_2
XFILLER_39_44 vpwr vgnd scs8hd_fill_2
XFILLER_39_22 vgnd vpwr scs8hd_decap_12
XANTENNA__232__D _232_/D vgnd vpwr scs8hd_diode_2
XFILLER_29_197 vgnd vpwr scs8hd_decap_3
XANTENNA__257__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_112 vpwr vgnd scs8hd_fill_2
XFILLER_35_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_35_123 vgnd vpwr scs8hd_decap_4
XANTENNA__167__A _143_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_178 vgnd vpwr scs8hd_decap_4
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XFILLER_41_126 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_17_101 vpwr vgnd scs8hd_fill_2
XFILLER_17_123 vpwr vgnd scs8hd_fill_2
XFILLER_17_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB _226_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[5] mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_126 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_4_.latch data_in mem_top_track_0.LATCH_4_.latch/Q _105_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_bottom_track_9.LATCH_1_.latch data_in mem_bottom_track_9.LATCH_1_.latch/Q _183_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_4_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_56 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_137 vpwr vgnd scs8hd_fill_2
XFILLER_14_159 vgnd vpwr scs8hd_decap_4
X_241_ _241_/HI _241_/LO vgnd vpwr scs8hd_conb_1
XFILLER_22_192 vpwr vgnd scs8hd_fill_2
X_172_ _135_/A _165_/A _172_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__270__A _270_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_163 vpwr vgnd scs8hd_fill_2
XANTENNA__180__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_58 vgnd vpwr scs8hd_decap_4
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_0_.latch data_in mem_left_track_9.LATCH_0_.latch/Q _207_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__090__A enable vgnd vpwr scs8hd_diode_2
XFILLER_27_240 vpwr vgnd scs8hd_fill_2
XANTENNA__265__A _265_/A vgnd vpwr scs8hd_diode_2
X_224_ _152_/A _152_/B _232_/C _232_/D _225_/A vgnd vpwr scs8hd_or4_4
X_086_ _086_/A _189_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_144 vpwr vgnd scs8hd_fill_2
X_155_ _142_/A _158_/B _155_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_7 vpwr vgnd scs8hd_fill_2
XFILLER_33_232 vgnd vpwr scs8hd_decap_12
XFILLER_33_221 vpwr vgnd scs8hd_fill_2
XFILLER_33_210 vgnd vpwr scs8hd_decap_4
XFILLER_18_251 vgnd vpwr scs8hd_fill_1
XANTENNA__159__B _158_/B vgnd vpwr scs8hd_diode_2
XANTENNA__175__A _175_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_25 vpwr vgnd scs8hd_fill_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XFILLER_24_243 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__085__A _097_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_3_169 vgnd vpwr scs8hd_decap_3
Xmem_top_track_16.LATCH_1_.latch data_in mem_top_track_16.LATCH_1_.latch/Q _214_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_207_ _223_/A _198_/X _207_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_15_276 vgnd vpwr scs8hd_fill_1
X_138_ address[4] _139_/A vgnd vpwr scs8hd_inv_8
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_235 vpwr vgnd scs8hd_fill_2
XFILLER_21_224 vpwr vgnd scs8hd_fill_2
XFILLER_0_83 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_70 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_1.LATCH_6_.latch data_in mem_bottom_track_1.LATCH_6_.latch/Q _167_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__172__B _165_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_48 vpwr vgnd scs8hd_fill_2
XFILLER_30_58 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_34 vgnd vpwr scs8hd_decap_6
XFILLER_29_187 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__273__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_5_.latch data_in mem_left_track_1.LATCH_5_.latch/Q _191_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_17.INVTX1_2_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_146 vgnd vpwr scs8hd_decap_4
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_3_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_179 vpwr vgnd scs8hd_fill_2
XFILLER_35_168 vpwr vgnd scs8hd_fill_2
XFILLER_35_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_6_.latch_SLEEPB _190_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__167__B _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA__183__A _135_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_71 vpwr vgnd scs8hd_fill_2
XFILLER_6_93 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_4_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _287_/A vgnd vpwr scs8hd_inv_1
XFILLER_41_138 vgnd vpwr scs8hd_decap_12
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_124 vpwr vgnd scs8hd_fill_2
XFILLER_26_102 vgnd vpwr scs8hd_decap_3
XFILLER_25_36 vpwr vgnd scs8hd_fill_2
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__093__A _152_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_267 vgnd vpwr scs8hd_decap_8
XANTENNA__268__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_32_149 vgnd vpwr scs8hd_decap_4
XFILLER_32_127 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__178__A _143_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_193 vpwr vgnd scs8hd_fill_2
XFILLER_11_16 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A address[4] vgnd vpwr scs8hd_diode_2
X_240_ _240_/HI _240_/LO vgnd vpwr scs8hd_conb_1
XFILLER_14_127 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_171_ _147_/A _165_/X _171_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_17.LATCH_1_.latch data_in mem_bottom_track_17.LATCH_1_.latch/Q _230_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_142 vpwr vgnd scs8hd_fill_2
XFILLER_9_197 vpwr vgnd scs8hd_fill_2
XANTENNA__180__B _176_/X vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[2] mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[7] mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_274 vgnd vpwr scs8hd_fill_1
XFILLER_36_230 vgnd vpwr scs8hd_decap_12
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_223_ _223_/A _221_/B _223_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__281__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
X_154_ _153_/X _158_/B vgnd vpwr scs8hd_buf_1
XFILLER_10_163 vpwr vgnd scs8hd_fill_2
X_085_ _097_/A _097_/B _084_/Y _086_/A vgnd vpwr scs8hd_or3_4
XFILLER_26_7 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_track_9.LATCH_5_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
XANTENNA__191__A _127_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_200 vpwr vgnd scs8hd_fill_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_58 vgnd vpwr scs8hd_fill_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A right_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__085__B _097_/B vgnd vpwr scs8hd_diode_2
XANTENNA__276__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmem_right_track_8.LATCH_0_.latch data_in mem_right_track_8.LATCH_0_.latch/Q _162_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_91 vgnd vpwr scs8hd_decap_4
X_137_ _149_/A _135_/B _137_/Y vgnd vpwr scs8hd_nor2_4
X_206_ _238_/A _198_/X _206_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_60 vgnd vpwr scs8hd_fill_1
XANTENNA__186__A _152_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _252_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB _235_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_47 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__096__A _094_/X vgnd vpwr scs8hd_diode_2
XFILLER_12_203 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_6_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_8_207 vgnd vpwr scs8hd_fill_1
XFILLER_12_247 vpwr vgnd scs8hd_fill_2
XFILLER_12_258 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_27 vpwr vgnd scs8hd_fill_2
XFILLER_29_177 vgnd vpwr scs8hd_fill_1
XFILLER_29_155 vgnd vpwr scs8hd_fill_1
XFILLER_29_100 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _251_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_232 vgnd vpwr scs8hd_decap_4
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _256_/A vgnd vpwr scs8hd_inv_1
XANTENNA__183__B _176_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_61 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_25_15 vgnd vpwr scs8hd_fill_1
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__093__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_202 vgnd vpwr scs8hd_decap_4
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XANTENNA__284__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_25_191 vpwr vgnd scs8hd_fill_2
XFILLER_15_81 vgnd vpwr scs8hd_decap_3
XFILLER_31_91 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_5_.latch data_in mem_top_track_8.LATCH_5_.latch/Q _127_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__194__A _147_/A vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_5_.latch data_in mem_right_track_0.LATCH_5_.latch/Q _144_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__178__B _176_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_28 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_170_ _131_/A _165_/X _170_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__279__A _279_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_176 vpwr vgnd scs8hd_fill_2
XFILLER_36_242 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__189__A _189_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_209 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_3_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__099__A _105_/A vgnd vpwr scs8hd_diode_2
X_153_ _152_/X _153_/X vgnd vpwr scs8hd_buf_1
X_222_ _238_/A _221_/B _222_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _248_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_71 vpwr vgnd scs8hd_fill_2
XFILLER_12_93 vpwr vgnd scs8hd_fill_2
X_084_ address[0] _084_/Y vgnd vpwr scs8hd_inv_8
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 chanx_right_in[4] mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr
+ scs8hd_diode_2
XANTENNA__191__B _191_/B vgnd vpwr scs8hd_diode_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_212 vpwr vgnd scs8hd_fill_2
XFILLER_17_38 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _247_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_37 vpwr vgnd scs8hd_fill_2
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_267 vgnd vpwr scs8hd_decap_8
XFILLER_24_256 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__085__C _084_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_3_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB _179_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_215 vpwr vgnd scs8hd_fill_2
XFILLER_30_204 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_256 vpwr vgnd scs8hd_fill_2
X_205_ _221_/A _199_/X _205_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_136_ _136_/A _149_/A vgnd vpwr scs8hd_buf_1
XFILLER_31_6 vpwr vgnd scs8hd_fill_2
XFILLER_2_171 vgnd vpwr scs8hd_decap_8
XANTENNA__186__B _139_/B vgnd vpwr scs8hd_diode_2
XFILLER_12_215 vpwr vgnd scs8hd_fill_2
XFILLER_12_237 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_9.LATCH_7_.latch data_in mem_bottom_track_9.LATCH_7_.latch/Q _177_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__287__A _287_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_270 vgnd vpwr scs8hd_decap_6
X_119_ _119_/A _152_/C vgnd vpwr scs8hd_buf_1
XFILLER_38_145 vgnd vpwr scs8hd_decap_8
XFILLER_38_134 vgnd vpwr scs8hd_decap_8
XFILLER_38_123 vgnd vpwr scs8hd_decap_8
XFILLER_38_112 vgnd vpwr scs8hd_decap_8
XANTENNA__197__A _139_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_29_134 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_6_.latch data_in mem_left_track_9.LATCH_6_.latch/Q _201_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_7_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_84 vpwr vgnd scs8hd_fill_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XANTENNA__093__C _232_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_5_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_236 vgnd vpwr scs8hd_fill_1
XFILLER_1_225 vgnd vpwr scs8hd_fill_1
XFILLER_1_214 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_159 vgnd vpwr scs8hd_fill_1
XFILLER_40_151 vpwr vgnd scs8hd_fill_2
XFILLER_15_93 vgnd vpwr scs8hd_decap_4
XFILLER_31_151 vgnd vpwr scs8hd_decap_3
XANTENNA__194__B _191_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XFILLER_31_162 vpwr vgnd scs8hd_fill_2
XFILLER_39_240 vgnd vpwr scs8hd_decap_4
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_107 vpwr vgnd scs8hd_fill_2
XFILLER_14_118 vgnd vpwr scs8hd_decap_3
XFILLER_22_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _172_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_151 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_162 vpwr vgnd scs8hd_fill_2
XFILLER_13_184 vpwr vgnd scs8hd_fill_2
XFILLER_13_195 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XFILLER_36_254 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__189__B _191_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_28 vgnd vpwr scs8hd_decap_3
XFILLER_22_17 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_210 vpwr vgnd scs8hd_fill_2
XANTENNA__099__B _124_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_276 vgnd vpwr scs8hd_fill_1
XFILLER_27_254 vpwr vgnd scs8hd_fill_2
X_221_ _221_/A _221_/B _221_/Y vgnd vpwr scs8hd_nor2_4
X_152_ _152_/A _152_/B _152_/C _152_/D _152_/X vgnd vpwr scs8hd_or4_4
X_083_ address[2] _097_/B vgnd vpwr scs8hd_inv_8
Xmux_top_track_8.INVTX1_3_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_169 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_191 vpwr vgnd scs8hd_fill_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_235 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB _212_/Y vgnd vpwr scs8hd_diode_2
XFILLER_33_27 vgnd vpwr scs8hd_fill_1
XFILLER_3_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_204_ _236_/A _199_/X _204_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_15_224 vpwr vgnd scs8hd_fill_2
XFILLER_15_235 vpwr vgnd scs8hd_fill_2
XFILLER_15_268 vpwr vgnd scs8hd_fill_2
X_135_ _135_/A _135_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_0_97 vpwr vgnd scs8hd_fill_2
XANTENNA__186__C _152_/C vgnd vpwr scs8hd_diode_2
XFILLER_21_205 vgnd vpwr scs8hd_decap_4
XFILLER_9_62 vgnd vpwr scs8hd_decap_3
XFILLER_9_95 vgnd vpwr scs8hd_decap_4
XFILLER_28_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_7_231 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_118_ address[3] _139_/B vgnd vpwr scs8hd_inv_8
XFILLER_38_168 vgnd vpwr scs8hd_decap_12
XFILLER_38_157 vgnd vpwr scs8hd_decap_8
XFILLER_22_3 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _242_/HI mem_bottom_track_9.LATCH_7_.latch/Q
+ mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__197__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_39 vpwr vgnd scs8hd_fill_2
XFILLER_39_48 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB _102_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[3] mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_20_83 vpwr vgnd scs8hd_fill_2
XFILLER_20_72 vpwr vgnd scs8hd_fill_2
XFILLER_4_245 vgnd vpwr scs8hd_decap_4
XFILLER_35_116 vpwr vgnd scs8hd_fill_2
XFILLER_35_105 vpwr vgnd scs8hd_fill_2
XFILLER_28_190 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_39 vgnd vpwr scs8hd_decap_3
XANTENNA__093__D _139_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB _229_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_2_.scs8hd_inv_1 chany_top_in[8] mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_7 vpwr vgnd scs8hd_fill_2
XFILLER_1_259 vpwr vgnd scs8hd_fill_2
XFILLER_1_248 vpwr vgnd scs8hd_fill_2
XFILLER_17_138 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_6_.latch data_in mem_right_track_8.LATCH_6_.latch/Q _156_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_263 vgnd vpwr scs8hd_decap_12
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
Xmem_left_track_17.LATCH_2_.latch data_in mem_left_track_17.LATCH_2_.latch/Q _237_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_196 vgnd vpwr scs8hd_fill_1
XFILLER_22_163 vgnd vpwr scs8hd_decap_8
XFILLER_22_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_7_.latch_SLEEPB _200_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_101 vpwr vgnd scs8hd_fill_2
XFILLER_9_123 vpwr vgnd scs8hd_fill_2
XFILLER_9_167 vpwr vgnd scs8hd_fill_2
XFILLER_3_97 vpwr vgnd scs8hd_fill_2
XFILLER_3_75 vgnd vpwr scs8hd_decap_6
XFILLER_36_266 vgnd vpwr scs8hd_decap_8
XFILLER_36_211 vgnd vpwr scs8hd_decap_3
X_220_ _236_/A _221_/B _220_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_266 vpwr vgnd scs8hd_fill_2
X_151_ address[5] _150_/Y _152_/D vgnd vpwr scs8hd_nand2_4
XFILLER_6_148 vgnd vpwr scs8hd_decap_4
XFILLER_10_133 vpwr vgnd scs8hd_fill_2
XFILLER_10_144 vgnd vpwr scs8hd_decap_6
XFILLER_10_188 vgnd vpwr scs8hd_decap_4
XFILLER_12_84 vpwr vgnd scs8hd_fill_2
X_082_ address[1] _097_/A vgnd vpwr scs8hd_inv_8
Xmux_top_track_0.INVTX1_6_.scs8hd_inv_1 chanx_left_in[0] mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _250_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_81 vgnd vpwr scs8hd_fill_1
XFILLER_18_222 vgnd vpwr scs8hd_decap_4
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
XFILLER_30_228 vgnd vpwr scs8hd_decap_8
X_203_ _219_/A _199_/X _203_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[1] mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_134_ _134_/A _135_/A vgnd vpwr scs8hd_buf_1
Xmem_bottom_track_1.LATCH_1_.latch data_in mem_bottom_track_1.LATCH_1_.latch/Q _172_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_228 vpwr vgnd scs8hd_fill_2
XANTENNA__186__D _232_/D vgnd vpwr scs8hd_diode_2
XFILLER_0_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_43 vpwr vgnd scs8hd_fill_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_21_239 vgnd vpwr scs8hd_decap_3
XFILLER_9_74 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_60 vpwr vgnd scs8hd_fill_2
XFILLER_7_254 vpwr vgnd scs8hd_fill_2
XFILLER_7_265 vpwr vgnd scs8hd_fill_2
X_117_ _094_/X _223_/A _117_/Y vgnd vpwr scs8hd_nor2_4
Xmem_left_track_1.LATCH_0_.latch data_in mem_left_track_1.LATCH_0_.latch/Q _196_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__197__C _152_/C vgnd vpwr scs8hd_diode_2
XFILLER_15_3 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XFILLER_29_158 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB _193_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_8_.scs8hd_inv_1_A left_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_51 vgnd vpwr scs8hd_decap_4
XFILLER_4_224 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.LATCH_1_.latch data_in mem_right_track_16.LATCH_1_.latch/Q _222_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_128 vgnd vpwr scs8hd_decap_4
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_62 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB _220_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__102__A _105_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_197 vpwr vgnd scs8hd_fill_2
XFILLER_31_175 vpwr vgnd scs8hd_fill_2
XFILLER_39_275 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[6] mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[2] mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_72 vgnd vpwr scs8hd_decap_3
XFILLER_9_146 vpwr vgnd scs8hd_fill_2
XFILLER_13_175 vgnd vpwr scs8hd_decap_6
XFILLER_3_54 vgnd vpwr scs8hd_fill_1
XFILLER_8_190 vpwr vgnd scs8hd_fill_2
XFILLER_27_223 vpwr vgnd scs8hd_fill_2
X_150_ address[6] _150_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_127 vgnd vpwr scs8hd_decap_6
XFILLER_10_167 vgnd vpwr scs8hd_decap_8
XFILLER_12_30 vgnd vpwr scs8hd_fill_1
XFILLER_12_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_279_ _279_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_5_160 vpwr vgnd scs8hd_fill_2
XFILLER_24_215 vgnd vpwr scs8hd_decap_3
XFILLER_24_204 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _238_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__200__A _189_/A vgnd vpwr scs8hd_diode_2
X_133_ _147_/A _127_/B _133_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_95 vgnd vpwr scs8hd_fill_1
X_202_ _218_/A _199_/X _202_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__110__A _109_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_88 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_42 vpwr vgnd scs8hd_fill_2
XFILLER_9_53 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_207 vgnd vpwr scs8hd_decap_4
XFILLER_18_62 vpwr vgnd scs8hd_fill_2
XFILLER_34_72 vgnd vpwr scs8hd_decap_3
XANTENNA__105__A _105_/A vgnd vpwr scs8hd_diode_2
X_116_ _136_/A _223_/A vgnd vpwr scs8hd_buf_1
XFILLER_11_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__197__D _232_/D vgnd vpwr scs8hd_diode_2
XFILLER_30_19 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_1.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_41 vgnd vpwr scs8hd_decap_3
XFILLER_20_30 vgnd vpwr scs8hd_fill_1
XFILLER_35_129 vpwr vgnd scs8hd_fill_2
XFILLER_29_83 vpwr vgnd scs8hd_fill_2
XFILLER_6_10 vgnd vpwr scs8hd_fill_1
XFILLER_6_32 vgnd vpwr scs8hd_fill_1
XFILLER_34_151 vpwr vgnd scs8hd_fill_2
XFILLER_26_107 vgnd vpwr scs8hd_decap_6
XFILLER_25_19 vpwr vgnd scs8hd_fill_2
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_top_track_8.LATCH_0_.latch data_in mem_top_track_8.LATCH_0_.latch/Q _137_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_right_track_0.LATCH_0_.latch data_in mem_right_track_0.LATCH_0_.latch/Q _149_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_239 vgnd vpwr scs8hd_decap_4
XFILLER_1_228 vgnd vpwr scs8hd_fill_1
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_195 vpwr vgnd scs8hd_fill_2
XFILLER_25_173 vpwr vgnd scs8hd_fill_2
XFILLER_31_95 vgnd vpwr scs8hd_decap_4
XFILLER_31_62 vgnd vpwr scs8hd_decap_3
XFILLER_31_40 vpwr vgnd scs8hd_fill_2
XANTENNA__102__B _218_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_31_110 vpwr vgnd scs8hd_fill_2
XFILLER_16_162 vgnd vpwr scs8hd_fill_1
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__203__A _219_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_6 vgnd vpwr scs8hd_decap_4
XFILLER_26_84 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A _134_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_44 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_10_102 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _269_/A vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_17.INVTX1_7_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_53 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_278_ _278_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA__108__A _105_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB _182_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_271 vgnd vpwr scs8hd_decap_4
XANTENNA__200__B _199_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_208 vgnd vpwr scs8hd_decap_6
XFILLER_15_205 vpwr vgnd scs8hd_fill_2
XFILLER_23_52 vpwr vgnd scs8hd_fill_2
X_201_ _124_/A _199_/X _201_/Y vgnd vpwr scs8hd_nor2_4
X_132_ _109_/X _147_/A vgnd vpwr scs8hd_buf_1
Xmem_top_track_0.LATCH_5_.latch data_in mem_top_track_0.LATCH_5_.latch/Q _102_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_142 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_9.LATCH_2_.latch data_in mem_bottom_track_9.LATCH_2_.latch/Q _182_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _261_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_12 vpwr vgnd scs8hd_fill_2
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_67 vpwr vgnd scs8hd_fill_2
XFILLER_17_8 vpwr vgnd scs8hd_fill_2
XFILLER_9_87 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_20_274 vgnd vpwr scs8hd_fill_1
XFILLER_12_219 vpwr vgnd scs8hd_fill_2
XFILLER_18_52 vgnd vpwr scs8hd_fill_1
XFILLER_18_41 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__211__A _219_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_84 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__105__B _219_/A vgnd vpwr scs8hd_diode_2
X_115_ address[1] address[2] address[0] _136_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__121__A _120_/X vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_1_.latch data_in mem_left_track_9.LATCH_1_.latch/Q _206_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_160 vpwr vgnd scs8hd_fill_2
XFILLER_29_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB _145_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_171 vpwr vgnd scs8hd_fill_2
XANTENNA__206__A _238_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_62 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_4_259 vgnd vpwr scs8hd_decap_12
XFILLER_28_182 vgnd vpwr scs8hd_decap_8
XANTENNA__116__A _136_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_44 vpwr vgnd scs8hd_fill_2
XFILLER_6_66 vgnd vpwr scs8hd_decap_3
XFILLER_6_88 vgnd vpwr scs8hd_decap_4
XFILLER_20_3 vgnd vpwr scs8hd_decap_3
Xmem_top_track_16.LATCH_2_.latch data_in mem_top_track_16.LATCH_2_.latch/Q _213_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_5_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_15_42 vpwr vgnd scs8hd_fill_2
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_31_74 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_8.LATCH_6_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_152 vgnd vpwr scs8hd_fill_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_track_1.LATCH_7_.latch data_in mem_bottom_track_1.LATCH_7_.latch/Q _166_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
.ends

