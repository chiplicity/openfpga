* NGSPICE file created from sb_0__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

.subckt sb_0__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_left_grid_pin_11_ bottom_left_grid_pin_13_ bottom_left_grid_pin_15_
+ bottom_left_grid_pin_1_ bottom_left_grid_pin_3_ bottom_left_grid_pin_5_ bottom_left_grid_pin_7_
+ bottom_left_grid_pin_9_ bottom_right_grid_pin_11_ chanx_right_in[0] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_out[0] chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3]
+ chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7]
+ chany_bottom_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ right_bottom_grid_pin_12_ right_top_grid_pin_10_ top_left_grid_pin_11_ top_left_grid_pin_13_
+ top_left_grid_pin_15_ top_left_grid_pin_1_ top_left_grid_pin_3_ top_left_grid_pin_5_
+ top_left_grid_pin_7_ top_left_grid_pin_9_ top_right_grid_pin_11_ vpwr vgnd
XFILLER_39_233 vpwr vgnd scs8hd_fill_2
Xmem_right_track_12.LATCH_1_.latch data_in _181_/A _167_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_122 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_100 vgnd vpwr scs8hd_decap_3
XFILLER_13_199 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__113__B _110_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_3_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_269 vgnd vpwr scs8hd_decap_8
XFILLER_6_107 vgnd vpwr scs8hd_decap_3
XFILLER_10_103 vpwr vgnd scs8hd_fill_2
XFILLER_10_125 vpwr vgnd scs8hd_fill_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__214__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _181_/A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_37_62 vgnd vpwr scs8hd_decap_3
XFILLER_18_203 vgnd vpwr scs8hd_decap_8
XFILLER_18_247 vgnd vpwr scs8hd_decap_8
XANTENNA__108__B _110_/B vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _124_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _194_/HI _176_/Y mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_195 vgnd vpwr scs8hd_fill_1
XFILLER_24_239 vgnd vpwr scs8hd_decap_12
XFILLER_24_206 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _188_/HI mem_bottom_track_17.LATCH_2_.latch/Q
+ mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__209__A _209_/A vgnd vpwr scs8hd_diode_2
X_200_ _200_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
X_131_ _121_/A _134_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
XANTENNA__119__A _085_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_2_.latch data_in mem_bottom_track_17.LATCH_2_.latch/Q _151_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _213_/A vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_96 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
X_114_ address[4] _114_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__121__B _121_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_6_.scs8hd_inv_1 bottom_left_grid_pin_7_ mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_4_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_29_106 vgnd vpwr scs8hd_decap_3
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_20_32 vgnd vpwr scs8hd_decap_8
XANTENNA__222__A _222_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[6] mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__132__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_109 vgnd vpwr scs8hd_decap_6
XFILLER_13_3 vgnd vpwr scs8hd_decap_6
XFILLER_19_161 vgnd vpwr scs8hd_decap_4
Xmem_right_track_8.LATCH_1_.latch data_in _183_/A _169_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_53 vpwr vgnd scs8hd_fill_2
XFILLER_25_197 vpwr vgnd scs8hd_fill_2
XANTENNA__217__A _217_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_54 vgnd vpwr scs8hd_decap_4
Xmux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _178_/A mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_0_263 vgnd vpwr scs8hd_decap_12
XFILLER_31_123 vpwr vgnd scs8hd_fill_2
XANTENNA__127__A _083_/A vgnd vpwr scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _180_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _188_/HI vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _191_/HI _182_/Y mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_97 vgnd vpwr scs8hd_decap_3
XFILLER_26_64 vgnd vpwr scs8hd_decap_6
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_138 vpwr vgnd scs8hd_fill_2
XFILLER_13_178 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_182 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _195_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_18_259 vgnd vpwr scs8hd_decap_12
XANTENNA__124__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _109_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
X_130_ _109_/A _134_/B _130_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_15_218 vpwr vgnd scs8hd_fill_2
XANTENNA__225__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_23_87 vgnd vpwr scs8hd_decap_3
XFILLER_2_122 vgnd vpwr scs8hd_fill_1
XFILLER_2_111 vgnd vpwr scs8hd_decap_4
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
XANTENNA__119__B _121_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_23 vpwr vgnd scs8hd_fill_2
XANTENNA__135__A _103_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A top_left_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_210 vgnd vpwr scs8hd_decap_4
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_6
XFILLER_34_75 vgnd vpwr scs8hd_decap_6
XFILLER_34_42 vpwr vgnd scs8hd_fill_2
X_113_ _124_/A _110_/B _113_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_214 vgnd vpwr scs8hd_fill_1
XFILLER_38_129 vgnd vpwr scs8hd_decap_6
XFILLER_38_118 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _182_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _186_/A mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XFILLER_37_173 vgnd vpwr scs8hd_decap_3
XFILLER_37_162 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_20_77 vpwr vgnd scs8hd_fill_2
XFILLER_6_46 vgnd vpwr scs8hd_decap_12
XANTENNA__132__B _134_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_140 vpwr vgnd scs8hd_fill_2
XFILLER_19_184 vpwr vgnd scs8hd_fill_2
XFILLER_19_195 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_113 vgnd vpwr scs8hd_decap_12
XFILLER_25_154 vpwr vgnd scs8hd_fill_2
XFILLER_25_143 vpwr vgnd scs8hd_fill_2
XFILLER_25_132 vpwr vgnd scs8hd_fill_2
XFILLER_15_11 vpwr vgnd scs8hd_fill_2
XFILLER_15_22 vpwr vgnd scs8hd_fill_2
XFILLER_15_33 vpwr vgnd scs8hd_fill_2
XFILLER_40_157 vgnd vpwr scs8hd_decap_8
XFILLER_15_77 vpwr vgnd scs8hd_fill_2
XFILLER_15_88 vgnd vpwr scs8hd_decap_3
XFILLER_0_275 vpwr vgnd scs8hd_fill_2
XFILLER_31_146 vpwr vgnd scs8hd_fill_2
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B _168_/B vgnd vpwr scs8hd_diode_2
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _173_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_32 vgnd vpwr scs8hd_fill_1
XFILLER_9_117 vgnd vpwr scs8hd_decap_3
XFILLER_13_157 vpwr vgnd scs8hd_fill_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _180_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A bottom_left_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _209_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_2.INVTX1_2_.scs8hd_inv_1_A right_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A _137_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_150 vgnd vpwr scs8hd_fill_1
XFILLER_27_205 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_149 vpwr vgnd scs8hd_fill_2
XFILLER_12_67 vgnd vpwr scs8hd_decap_3
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XFILLER_5_175 vpwr vgnd scs8hd_fill_2
XFILLER_5_164 vgnd vpwr scs8hd_decap_6
XFILLER_5_153 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__140__B _138_/X vgnd vpwr scs8hd_diode_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_252 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr
+ scs8hd_diode_2
X_189_ _189_/HI _189_/LO vgnd vpwr scs8hd_conb_1
XFILLER_9_57 vgnd vpwr scs8hd_fill_1
XFILLER_9_79 vpwr vgnd scs8hd_fill_2
XANTENNA__135__B _114_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA__151__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_11 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_8
X_112_ _123_/A _110_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_259 vpwr vgnd scs8hd_fill_2
XANTENNA__146__A _170_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
XFILLER_37_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _175_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_207 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_5_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _173_/A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_98 vpwr vgnd scs8hd_fill_2
XFILLER_29_54 vgnd vpwr scs8hd_decap_4
XFILLER_28_163 vgnd vpwr scs8hd_fill_1
XFILLER_6_58 vgnd vpwr scs8hd_decap_3
XFILLER_3_240 vgnd vpwr scs8hd_decap_4
XFILLER_40_136 vgnd vpwr scs8hd_decap_4
XFILLER_40_125 vpwr vgnd scs8hd_fill_2
XFILLER_25_111 vpwr vgnd scs8hd_fill_2
XFILLER_40_169 vgnd vpwr scs8hd_decap_12
XFILLER_31_77 vpwr vgnd scs8hd_fill_2
XFILLER_0_232 vgnd vpwr scs8hd_decap_4
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__C _170_/C vgnd vpwr scs8hd_diode_2
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__143__B _138_/X vgnd vpwr scs8hd_diode_2
XFILLER_39_269 vgnd vpwr scs8hd_decap_8
XFILLER_39_225 vgnd vpwr scs8hd_decap_4
XFILLER_39_203 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_158 vpwr vgnd scs8hd_fill_2
XFILLER_22_103 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmem_right_track_4.LATCH_1_.latch data_in _175_/A _161_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _177_/Y mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__154__A _083_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_217 vgnd vpwr scs8hd_decap_12
Xmux_right_track_14.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_46 vpwr vgnd scs8hd_fill_2
XFILLER_12_57 vgnd vpwr scs8hd_decap_8
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_54 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_228 vgnd vpwr scs8hd_decap_4
Xmem_top_track_0.LATCH_0_.latch data_in mem_top_track_0.LATCH_0_.latch/Q _101_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_198 vpwr vgnd scs8hd_fill_2
XFILLER_5_187 vgnd vpwr scs8hd_decap_8
XFILLER_5_132 vpwr vgnd scs8hd_fill_2
XANTENNA__149__A _109_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_3_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_91 vgnd vpwr scs8hd_fill_1
XFILLER_23_264 vgnd vpwr scs8hd_decap_12
XFILLER_2_102 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_9_36 vpwr vgnd scs8hd_fill_2
XFILLER_14_242 vgnd vpwr scs8hd_decap_12
XANTENNA__135__C _115_/C vgnd vpwr scs8hd_diode_2
X_188_ _188_/HI _188_/LO vgnd vpwr scs8hd_conb_1
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XANTENNA__151__B _150_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _179_/A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_201 vgnd vpwr scs8hd_decap_3
Xmux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _193_/HI _174_/Y mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_23 vgnd vpwr scs8hd_decap_8
XFILLER_11_212 vgnd vpwr scs8hd_decap_3
X_111_ _122_/A _110_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_11_245 vpwr vgnd scs8hd_fill_2
XANTENNA__146__B _146_/B vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_77 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _196_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XFILLER_34_167 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__157__A _154_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_2_.latch data_in mem_bottom_track_1.LATCH_2_.latch/Q _132_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _192_/HI _185_/Y mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB _110_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_25_178 vgnd vpwr scs8hd_decap_3
XFILLER_15_46 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_244 vgnd vpwr scs8hd_decap_4
XFILLER_31_115 vpwr vgnd scs8hd_fill_2
XFILLER_16_112 vgnd vpwr scs8hd_decap_6
XFILLER_31_159 vpwr vgnd scs8hd_fill_2
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_237 vgnd vpwr scs8hd_decap_6
XFILLER_39_215 vpwr vgnd scs8hd_fill_2
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_181 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_89 vgnd vpwr scs8hd_decap_3
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_21_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _176_/A mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_163 vgnd vpwr scs8hd_decap_8
XANTENNA__170__A _170_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_229 vgnd vpwr scs8hd_decap_12
XFILLER_10_107 vpwr vgnd scs8hd_fill_2
XFILLER_10_129 vgnd vpwr scs8hd_decap_6
XFILLER_12_36 vgnd vpwr scs8hd_fill_1
XANTENNA__080__A enable vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_251 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _190_/HI _180_/Y mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__149__B _150_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_276 vgnd vpwr scs8hd_fill_1
XFILLER_23_79 vpwr vgnd scs8hd_fill_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XANTENNA__075__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_2_125 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.INVTX1_0_.scs8hd_inv_1 chany_top_in[6] mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_39 vpwr vgnd scs8hd_fill_2
XFILLER_9_15 vgnd vpwr scs8hd_decap_8
XFILLER_14_254 vgnd vpwr scs8hd_decap_12
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _187_/HI _187_/LO vgnd vpwr scs8hd_conb_1
Xmux_bottom_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _184_/Y mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_20_224 vgnd vpwr scs8hd_decap_12
XFILLER_18_68 vpwr vgnd scs8hd_fill_2
XFILLER_18_79 vgnd vpwr scs8hd_decap_4
X_110_ _121_/A _110_/B _110_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_257 vpwr vgnd scs8hd_fill_2
XFILLER_7_217 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _179_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__146__C _083_/C vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA__162__B _163_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_4_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_187 vgnd vpwr scs8hd_decap_12
XFILLER_28_176 vgnd vpwr scs8hd_decap_8
XFILLER_28_132 vgnd vpwr scs8hd_decap_4
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_3_253 vpwr vgnd scs8hd_fill_2
XFILLER_19_132 vpwr vgnd scs8hd_fill_2
XFILLER_34_179 vgnd vpwr scs8hd_decap_12
XFILLER_34_146 vgnd vpwr scs8hd_decap_4
XFILLER_34_102 vgnd vpwr scs8hd_decap_3
XANTENNA__157__B _163_/B vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _173_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_35 vgnd vpwr scs8hd_decap_3
XANTENNA__083__A _083_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _182_/A mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_15_58 vgnd vpwr scs8hd_fill_1
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
XFILLER_31_127 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_146 vpwr vgnd scs8hd_fill_2
XFILLER_16_157 vpwr vgnd scs8hd_fill_2
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__168__A _154_/X vgnd vpwr scs8hd_diode_2
XFILLER_22_149 vpwr vgnd scs8hd_fill_2
XFILLER_30_193 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_1_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__078__A _078_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_149 vpwr vgnd scs8hd_fill_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_3_39 vgnd vpwr scs8hd_decap_12
XFILLER_8_186 vgnd vpwr scs8hd_decap_4
XFILLER_12_182 vpwr vgnd scs8hd_fill_2
XANTENNA__170__B _170_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_89 vpwr vgnd scs8hd_fill_2
XFILLER_37_67 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[4] mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_263 vgnd vpwr scs8hd_decap_12
Xmem_top_track_8.LATCH_1_.latch data_in mem_top_track_8.LATCH_1_.latch/Q _112_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _181_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__165__B _170_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_60 vgnd vpwr scs8hd_decap_8
XANTENNA__181__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_47 vgnd vpwr scs8hd_fill_1
XANTENNA__091__A _090_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_211 vgnd vpwr scs8hd_decap_3
XFILLER_14_266 vgnd vpwr scs8hd_decap_8
X_186_ _186_/A _186_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _176_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_192 vgnd vpwr scs8hd_decap_12
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_236 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.INVTX1_6_.scs8hd_inv_1 bottom_left_grid_pin_5_ mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_46 vgnd vpwr scs8hd_decap_3
XFILLER_7_229 vgnd vpwr scs8hd_decap_12
XANTENNA__086__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_1_3 vgnd vpwr scs8hd_decap_8
Xmux_top_track_8.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_10.INVTX1_0_.scs8hd_inv_1 chany_top_in[5] mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_251 vgnd vpwr scs8hd_decap_12
X_169_ _170_/A _170_/B _170_/C _163_/D _169_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__162__C _083_/C vgnd vpwr scs8hd_diode_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_199 vgnd vpwr scs8hd_decap_12
XFILLER_28_166 vgnd vpwr scs8hd_fill_1
XFILLER_19_188 vpwr vgnd scs8hd_fill_2
XFILLER_19_199 vgnd vpwr scs8hd_decap_3
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XANTENNA__157__C _165_/C vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.LATCH_3_.latch data_in mem_bottom_track_9.LATCH_3_.latch/Q _141_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_25_158 vpwr vgnd scs8hd_fill_2
XFILLER_25_147 vgnd vpwr scs8hd_decap_4
XFILLER_25_136 vgnd vpwr scs8hd_decap_4
XANTENNA__083__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _174_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_80 vpwr vgnd scs8hd_fill_2
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _168_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_128 vpwr vgnd scs8hd_fill_2
XANTENNA__184__A _184_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_47 vgnd vpwr scs8hd_decap_6
XFILLER_26_36 vgnd vpwr scs8hd_decap_8
XANTENNA__094__A _093_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_121 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _178_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__170__C _170_/C vgnd vpwr scs8hd_diode_2
XANTENNA__179__A _179_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
Xmux_right_track_12.tap_buf4_0_.scs8hd_inv_1 mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _202_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_79 vgnd vpwr scs8hd_decap_8
Xmem_top_track_16.LATCH_3_.latch data_in mem_top_track_16.LATCH_3_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__089__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
XFILLER_5_102 vgnd vpwr scs8hd_fill_1
XFILLER_17_242 vpwr vgnd scs8hd_fill_2
XANTENNA__165__C _165_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _175_/Y mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_223 vgnd vpwr scs8hd_decap_12
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_13_81 vpwr vgnd scs8hd_fill_2
XFILLER_13_92 vpwr vgnd scs8hd_fill_2
X_185_ _185_/A _185_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_6.INVTX1_1_.scs8hd_inv_1 chany_top_in[8] mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_182 vgnd vpwr scs8hd_fill_1
XFILLER_20_248 vgnd vpwr scs8hd_decap_12
XANTENNA__086__B _086_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_58 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _176_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_91 vgnd vpwr scs8hd_fill_1
XFILLER_24_80 vgnd vpwr scs8hd_decap_4
XFILLER_6_263 vgnd vpwr scs8hd_decap_12
X_168_ _154_/X _168_/B _083_/C _164_/D _168_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__162__D _164_/D vgnd vpwr scs8hd_diode_2
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
X_099_ address[1] address[2] address[0] _100_/A vgnd vpwr scs8hd_or3_4
XFILLER_37_178 vgnd vpwr scs8hd_decap_4
XFILLER_37_134 vpwr vgnd scs8hd_fill_2
XFILLER_37_112 vpwr vgnd scs8hd_fill_2
XFILLER_1_73 vpwr vgnd scs8hd_fill_2
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_49 vgnd vpwr scs8hd_decap_12
XFILLER_29_58 vgnd vpwr scs8hd_fill_1
XFILLER_29_47 vgnd vpwr scs8hd_fill_1
XFILLER_28_145 vgnd vpwr scs8hd_decap_8
XFILLER_28_112 vgnd vpwr scs8hd_decap_4
XANTENNA__097__A _096_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_71 vpwr vgnd scs8hd_fill_2
XFILLER_10_93 vgnd vpwr scs8hd_fill_1
XFILLER_13_9 vgnd vpwr scs8hd_fill_1
XFILLER_19_167 vpwr vgnd scs8hd_fill_2
XFILLER_35_90 vgnd vpwr scs8hd_decap_6
XANTENNA__157__D _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_25_115 vpwr vgnd scs8hd_fill_2
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XANTENNA__083__C _083_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_203 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_17.LATCH_3_.latch data_in mem_bottom_track_17.LATCH_3_.latch/Q _150_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_137 vpwr vgnd scs8hd_fill_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_107 vpwr vgnd scs8hd_fill_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA__168__C _083_/C vgnd vpwr scs8hd_diode_2
XFILLER_30_140 vpwr vgnd scs8hd_fill_2
XFILLER_7_83 vpwr vgnd scs8hd_fill_2
XFILLER_7_94 vpwr vgnd scs8hd_fill_2
XFILLER_38_251 vgnd vpwr scs8hd_decap_12
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_6.tap_buf4_0_.scs8hd_inv_1 mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _205_/A vgnd vpwr scs8hd_inv_1
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _181_/Y mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_21_195 vpwr vgnd scs8hd_fill_2
XFILLER_16_70 vgnd vpwr scs8hd_decap_3
XFILLER_8_144 vgnd vpwr scs8hd_decap_6
XFILLER_8_199 vpwr vgnd scs8hd_fill_2
XANTENNA__170__D _164_/D vgnd vpwr scs8hd_diode_2
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XFILLER_37_58 vgnd vpwr scs8hd_fill_1
XFILLER_37_47 vgnd vpwr scs8hd_fill_1
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_136 vpwr vgnd scs8hd_fill_2
XFILLER_5_114 vpwr vgnd scs8hd_fill_2
XFILLER_32_213 vgnd vpwr scs8hd_fill_1
XANTENNA__165__D _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_23_235 vgnd vpwr scs8hd_decap_8
XFILLER_23_27 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _174_/A mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_14_202 vgnd vpwr scs8hd_decap_6
XFILLER_14_224 vpwr vgnd scs8hd_fill_2
X_184_ _184_/A _184_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_5_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_49 vgnd vpwr scs8hd_decap_8
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XANTENNA__086__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_11_249 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_098_ _085_/B _123_/A _098_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_271 vgnd vpwr scs8hd_decap_4
X_167_ _154_/X _168_/B _083_/C _163_/D _167_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_1_96 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.INVTX1_1_.scs8hd_inv_1 chany_top_in[7] mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_15 vgnd vpwr scs8hd_decap_12
XFILLER_28_157 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _178_/Y mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_8
XFILLER_3_212 vpwr vgnd scs8hd_fill_2
XFILLER_10_50 vpwr vgnd scs8hd_fill_2
XFILLER_19_113 vgnd vpwr scs8hd_decap_3
XFILLER_34_138 vgnd vpwr scs8hd_decap_6
XFILLER_19_81 vpwr vgnd scs8hd_fill_2
XFILLER_19_92 vpwr vgnd scs8hd_fill_2
XFILLER_19_179 vgnd vpwr scs8hd_decap_4
X_219_ chany_bottom_in[6] chany_top_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_33_182 vgnd vpwr scs8hd_fill_1
XFILLER_18_190 vpwr vgnd scs8hd_fill_2
XFILLER_31_27 vgnd vpwr scs8hd_decap_8
XFILLER_0_259 vpwr vgnd scs8hd_fill_2
XFILLER_0_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _198_/HI mem_top_track_16.LATCH_2_.latch/Q
+ mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_119 vgnd vpwr scs8hd_decap_3
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XANTENNA__168__D _164_/D vgnd vpwr scs8hd_diode_2
XFILLER_30_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_40 vpwr vgnd scs8hd_fill_2
XFILLER_7_62 vpwr vgnd scs8hd_fill_2
XFILLER_38_263 vgnd vpwr scs8hd_decap_12
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _182_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_174 vpwr vgnd scs8hd_fill_2
XFILLER_16_93 vpwr vgnd scs8hd_fill_2
Xmux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _180_/A mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_130 vpwr vgnd scs8hd_fill_2
XFILLER_12_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A top_left_grid_pin_7_ vgnd vpwr scs8hd_diode_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_4_96 vpwr vgnd scs8hd_fill_2
XFILLER_23_39 vgnd vpwr scs8hd_decap_8
XFILLER_2_129 vgnd vpwr scs8hd_decap_12
XFILLER_2_118 vgnd vpwr scs8hd_decap_4
XFILLER_2_107 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_236 vgnd vpwr scs8hd_decap_3
X_183_ _183_/A _183_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_262 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _186_/Y mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A bottom_left_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _180_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XFILLER_11_217 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 top_left_grid_pin_11_ mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_93 vpwr vgnd scs8hd_fill_2
XFILLER_10_250 vgnd vpwr scs8hd_decap_4
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_097_ _096_/X _123_/A vgnd vpwr scs8hd_buf_1
X_166_ _161_/A _170_/B _165_/C _164_/D _166_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_37_147 vgnd vpwr scs8hd_decap_6
XFILLER_37_169 vpwr vgnd scs8hd_fill_2
XFILLER_37_158 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _186_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_10_40 vgnd vpwr scs8hd_fill_1
XFILLER_10_84 vgnd vpwr scs8hd_decap_3
XFILLER_19_136 vpwr vgnd scs8hd_fill_2
XFILLER_34_117 vgnd vpwr scs8hd_decap_8
X_218_ _218_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
X_149_ _109_/A _150_/B _149_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_18 vpwr vgnd scs8hd_fill_2
XFILLER_15_29 vpwr vgnd scs8hd_fill_2
XFILLER_0_249 vgnd vpwr scs8hd_decap_6
Xmux_right_track_2.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_172 vgnd vpwr scs8hd_decap_4
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A bottom_left_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_150 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _189_/HI mem_bottom_track_9.LATCH_2_.latch/Q
+ mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_142 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_102 vpwr vgnd scs8hd_fill_2
XFILLER_32_93 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _175_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_186 vgnd vpwr scs8hd_decap_4
XFILLER_35_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _182_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XFILLER_5_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_234 vgnd vpwr scs8hd_decap_8
XFILLER_17_245 vgnd vpwr scs8hd_decap_12
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_248 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_182_ _182_/A _182_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_62 vpwr vgnd scs8hd_fill_2
XANTENNA__100__A _100_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_274 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_2_.scs8hd_inv_1 top_left_grid_pin_15_ mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_229 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _173_/Y mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_61 vgnd vpwr scs8hd_decap_3
X_165_ _161_/A _170_/B _165_/C _163_/D _165_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_40_71 vgnd vpwr scs8hd_decap_4
X_096_ address[1] address[2] _171_/D _096_/X vgnd vpwr scs8hd_or3_4
XFILLER_37_126 vpwr vgnd scs8hd_fill_2
XFILLER_37_104 vpwr vgnd scs8hd_fill_2
XFILLER_1_65 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_1_.latch data_in mem_top_track_0.LATCH_1_.latch/Q _098_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_39 vgnd vpwr scs8hd_decap_8
XFILLER_28_104 vpwr vgnd scs8hd_fill_2
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _177_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_140 vgnd vpwr scs8hd_decap_12
XFILLER_34_107 vgnd vpwr scs8hd_fill_1
X_217_ _217_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
X_148_ _085_/A _150_/B _148_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
X_079_ address[5] _083_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XFILLER_33_140 vpwr vgnd scs8hd_fill_2
XFILLER_0_228 vpwr vgnd scs8hd_fill_2
XFILLER_24_140 vgnd vpwr scs8hd_decap_8
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_62 vpwr vgnd scs8hd_fill_2
XFILLER_21_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_184 vpwr vgnd scs8hd_fill_2
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_29_232 vgnd vpwr scs8hd_decap_12
XFILLER_8_125 vgnd vpwr scs8hd_decap_4
XFILLER_12_165 vpwr vgnd scs8hd_fill_2
XFILLER_16_40 vpwr vgnd scs8hd_fill_2
XFILLER_16_51 vgnd vpwr scs8hd_decap_8
XFILLER_16_62 vpwr vgnd scs8hd_fill_2
XFILLER_16_84 vpwr vgnd scs8hd_fill_2
XFILLER_32_83 vgnd vpwr scs8hd_decap_4
XFILLER_32_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__103__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_4_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_39 vgnd vpwr scs8hd_decap_8
XFILLER_26_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_3_.latch data_in mem_bottom_track_1.LATCH_3_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_32_205 vgnd vpwr scs8hd_decap_8
XFILLER_27_83 vpwr vgnd scs8hd_fill_2
XFILLER_17_213 vpwr vgnd scs8hd_fill_2
XFILLER_17_257 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ _179_/Y mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_183 vgnd vpwr scs8hd_decap_12
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_87 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_22_260 vgnd vpwr scs8hd_decap_12
X_181_ _181_/A _181_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_52 vpwr vgnd scs8hd_fill_2
XFILLER_1_142 vgnd vpwr scs8hd_decap_12
XFILLER_13_85 vpwr vgnd scs8hd_fill_2
XFILLER_13_96 vpwr vgnd scs8hd_fill_2
Xmem_right_track_14.LATCH_0_.latch data_in _186_/A _172_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_93 vgnd vpwr scs8hd_decap_4
XFILLER_9_220 vgnd vpwr scs8hd_decap_12
XFILLER_9_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
X_095_ _085_/B _122_/A _095_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_84 vgnd vpwr scs8hd_fill_1
X_164_ _161_/A _163_/B _163_/C _164_/D _164_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_37_116 vgnd vpwr scs8hd_decap_6
XANTENNA__111__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_11 vgnd vpwr scs8hd_fill_1
XFILLER_1_77 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_28_116 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_160 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_62 vpwr vgnd scs8hd_fill_2
XFILLER_42_152 vgnd vpwr scs8hd_decap_3
XFILLER_27_193 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_147_ _146_/X _150_/B vgnd vpwr scs8hd_buf_1
X_216_ chany_top_in[0] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
X_078_ _078_/A _085_/A vgnd vpwr scs8hd_buf_1
XANTENNA__106__A _083_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_8
XFILLER_25_119 vgnd vpwr scs8hd_decap_3
XFILLER_18_182 vgnd vpwr scs8hd_decap_8
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_218 vgnd vpwr scs8hd_decap_6
XFILLER_0_207 vgnd vpwr scs8hd_decap_8
XFILLER_24_185 vpwr vgnd scs8hd_fill_2
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_3_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_30_144 vgnd vpwr scs8hd_decap_6
Xmux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _176_/Y mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_87 vpwr vgnd scs8hd_fill_2
XFILLER_7_98 vgnd vpwr scs8hd_decap_3
XFILLER_38_211 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_199 vpwr vgnd scs8hd_fill_2
XFILLER_32_51 vpwr vgnd scs8hd_fill_2
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_118 vpwr vgnd scs8hd_fill_2
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_62 vpwr vgnd scs8hd_fill_2
XFILLER_17_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB _164_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_195 vgnd vpwr scs8hd_decap_12
XFILLER_4_77 vgnd vpwr scs8hd_decap_8
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XANTENNA__114__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_228 vgnd vpwr scs8hd_decap_8
XFILLER_22_272 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_180_ _180_/A _180_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_20 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_121 vgnd vpwr scs8hd_fill_1
XFILLER_1_154 vgnd vpwr scs8hd_decap_12
XFILLER_38_61 vgnd vpwr scs8hd_decap_4
XANTENNA__109__A _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_232 vgnd vpwr scs8hd_decap_12
XFILLER_39_191 vpwr vgnd scs8hd_fill_2
XFILLER_40_84 vpwr vgnd scs8hd_fill_2
X_163_ _161_/A _163_/B _163_/C _163_/D _163_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_6_213 vgnd vpwr scs8hd_fill_1
X_094_ _093_/X _122_/A vgnd vpwr scs8hd_buf_1
XANTENNA__111__B _110_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _199_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_56 vgnd vpwr scs8hd_fill_1
XFILLER_1_89 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_2_.latch data_in mem_top_track_8.LATCH_2_.latch/Q _111_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_128 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _181_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _182_/Y mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_216 vgnd vpwr scs8hd_decap_12
XANTENNA__212__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_10_32 vgnd vpwr scs8hd_decap_8
XFILLER_10_54 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_85 vgnd vpwr scs8hd_decap_4
XFILLER_19_96 vpwr vgnd scs8hd_fill_2
XFILLER_35_73 vgnd vpwr scs8hd_decap_3
X_215_ chany_top_in[1] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA__122__A _122_/A vgnd vpwr scs8hd_diode_2
X_077_ address[1] _086_/B _171_/D _078_/A vgnd vpwr scs8hd_or3_4
XANTENNA__106__B _170_/B vgnd vpwr scs8hd_diode_2
X_146_ _170_/A _146_/B _083_/C _146_/X vgnd vpwr scs8hd_or3_4
XFILLER_33_164 vgnd vpwr scs8hd_decap_12
XFILLER_33_153 vpwr vgnd scs8hd_fill_2
XFILLER_18_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__207__A _207_/A vgnd vpwr scs8hd_diode_2
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _083_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_66 vgnd vpwr scs8hd_decap_4
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
X_129_ _085_/A _134_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_3_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_101 vpwr vgnd scs8hd_fill_2
XFILLER_21_123 vpwr vgnd scs8hd_fill_2
XFILLER_21_134 vpwr vgnd scs8hd_fill_2
XFILLER_21_145 vpwr vgnd scs8hd_fill_2
XFILLER_21_178 vgnd vpwr scs8hd_decap_3
XFILLER_29_245 vgnd vpwr scs8hd_decap_12
XFILLER_8_138 vgnd vpwr scs8hd_decap_4
XFILLER_12_112 vpwr vgnd scs8hd_fill_2
XFILLER_12_134 vgnd vpwr scs8hd_decap_4
XFILLER_12_145 vgnd vpwr scs8hd_decap_6
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_160 vgnd vpwr scs8hd_decap_4
XFILLER_7_193 vpwr vgnd scs8hd_fill_2
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_9.LATCH_4_.latch data_in mem_bottom_track_9.LATCH_4_.latch/Q _140_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__220__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _190_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_204 vpwr vgnd scs8hd_fill_2
XFILLER_40_251 vgnd vpwr scs8hd_decap_12
XFILLER_27_96 vpwr vgnd scs8hd_fill_2
XFILLER_4_141 vgnd vpwr scs8hd_decap_12
XFILLER_4_130 vpwr vgnd scs8hd_fill_2
XFILLER_4_163 vgnd vpwr scs8hd_decap_12
XFILLER_4_56 vgnd vpwr scs8hd_fill_1
XANTENNA__130__A _109_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _185_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__215__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_1_188 vpwr vgnd scs8hd_fill_2
XFILLER_1_100 vpwr vgnd scs8hd_fill_2
XFILLER_1_166 vgnd vpwr scs8hd_decap_12
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XANTENNA__109__B _110_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_266 vgnd vpwr scs8hd_decap_8
XANTENNA__125__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_6_.scs8hd_inv_1 bottom_left_grid_pin_9_ mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _178_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_97 vgnd vpwr scs8hd_decap_3
X_162_ _161_/A _163_/B _083_/C _164_/D _162_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_40_96 vpwr vgnd scs8hd_fill_2
XFILLER_40_30 vgnd vpwr scs8hd_fill_1
XFILLER_10_254 vgnd vpwr scs8hd_fill_1
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
X_093_ _093_/A address[2] address[0] _093_/X vgnd vpwr scs8hd_or3_4
Xmem_top_track_16.LATCH_4_.latch data_in mem_top_track_16.LATCH_4_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_right_track_10.LATCH_0_.latch data_in _180_/A _166_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_140 vpwr vgnd scs8hd_fill_2
XFILLER_3_228 vgnd vpwr scs8hd_decap_12
XFILLER_19_53 vpwr vgnd scs8hd_fill_2
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_27_173 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_214_ chany_top_in[2] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__106__C _163_/C vgnd vpwr scs8hd_diode_2
X_145_ address[5] _170_/A vgnd vpwr scs8hd_inv_8
XANTENNA__122__B _121_/B vgnd vpwr scs8hd_diode_2
X_076_ address[0] _171_/D vgnd vpwr scs8hd_inv_8
XFILLER_33_176 vgnd vpwr scs8hd_decap_6
XFILLER_33_110 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_3
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__223__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_30_102 vpwr vgnd scs8hd_fill_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_30_157 vgnd vpwr scs8hd_decap_12
XANTENNA__133__A _123_/A vgnd vpwr scs8hd_diode_2
X_128_ _127_/X _134_/B vgnd vpwr scs8hd_buf_1
XANTENNA__117__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _176_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
XANTENNA__218__A _218_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_6
XFILLER_8_106 vpwr vgnd scs8hd_fill_2
XANTENNA__128__A _127_/X vgnd vpwr scs8hd_diode_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_227 vgnd vpwr scs8hd_decap_12
XFILLER_26_205 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _184_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XFILLER_40_263 vgnd vpwr scs8hd_decap_12
XFILLER_4_175 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_17.LATCH_4_.latch data_in mem_bottom_track_17.LATCH_4_.latch/Q _149_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__130__B _134_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_219 vpwr vgnd scs8hd_fill_2
XFILLER_23_208 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_208 vgnd vpwr scs8hd_fill_1
XFILLER_13_66 vpwr vgnd scs8hd_fill_2
XFILLER_1_112 vgnd vpwr scs8hd_decap_3
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
XFILLER_1_178 vgnd vpwr scs8hd_decap_4
XFILLER_38_74 vgnd vpwr scs8hd_decap_12
XFILLER_9_201 vpwr vgnd scs8hd_fill_2
XFILLER_9_212 vpwr vgnd scs8hd_fill_2
XFILLER_9_245 vgnd vpwr scs8hd_decap_8
XFILLER_13_241 vgnd vpwr scs8hd_decap_3
XFILLER_13_263 vgnd vpwr scs8hd_decap_12
Xmem_right_track_6.LATCH_0_.latch data_in _178_/A _164_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__141__A _121_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__226__A _226_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_87 vgnd vpwr scs8hd_decap_4
XFILLER_24_32 vgnd vpwr scs8hd_decap_12
X_161_ _161_/A _163_/B _083_/C _163_/D _161_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
XFILLER_10_222 vpwr vgnd scs8hd_fill_2
X_092_ _085_/B _121_/A _092_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_108 vpwr vgnd scs8hd_fill_2
XFILLER_1_14 vgnd vpwr scs8hd_decap_12
XFILLER_1_69 vpwr vgnd scs8hd_fill_2
XANTENNA__136__A _135_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _178_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_163 vpwr vgnd scs8hd_fill_2
XFILLER_36_152 vgnd vpwr scs8hd_fill_1
XFILLER_28_108 vpwr vgnd scs8hd_fill_2
XFILLER_10_67 vpwr vgnd scs8hd_fill_2
XFILLER_10_89 vgnd vpwr scs8hd_decap_3
XFILLER_19_21 vgnd vpwr scs8hd_decap_4
XFILLER_19_32 vpwr vgnd scs8hd_fill_2
XFILLER_35_53 vpwr vgnd scs8hd_fill_2
XFILLER_35_42 vpwr vgnd scs8hd_fill_2
XFILLER_27_130 vgnd vpwr scs8hd_decap_3
Xmux_right_track_12.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[7] mux_right_track_12.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _199_/HI mem_top_track_8.LATCH_2_.latch/Q
+ mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_213_ _213_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
X_144_ _124_/A _138_/X _144_/Y vgnd vpwr scs8hd_nor2_4
X_075_ address[2] _086_/B vgnd vpwr scs8hd_inv_8
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.tap_buf4_0_.scs8hd_inv_1 mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _207_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _098_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_133 vgnd vpwr scs8hd_decap_4
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_9.INVTX1_5_.scs8hd_inv_1 bottom_left_grid_pin_1_ mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_44 vpwr vgnd scs8hd_fill_2
XFILLER_21_66 vgnd vpwr scs8hd_decap_3
XFILLER_30_169 vgnd vpwr scs8hd_decap_12
XFILLER_30_136 vpwr vgnd scs8hd_fill_2
XFILLER_30_125 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_188 vpwr vgnd scs8hd_fill_2
XANTENNA__117__C _170_/C vgnd vpwr scs8hd_diode_2
XFILLER_7_35 vgnd vpwr scs8hd_decap_3
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__133__B _134_/B vgnd vpwr scs8hd_diode_2
X_127_ _083_/A _168_/B _170_/C _127_/X vgnd vpwr scs8hd_or3_4
XFILLER_38_203 vgnd vpwr scs8hd_decap_8
XFILLER_16_3 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _217_/A vgnd vpwr scs8hd_inv_1
Xmux_top_track_16.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[2] mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
XFILLER_12_169 vgnd vpwr scs8hd_decap_4
XFILLER_16_66 vpwr vgnd scs8hd_fill_2
XFILLER_16_88 vgnd vpwr scs8hd_decap_4
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XANTENNA__144__A _124_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_151 vgnd vpwr scs8hd_decap_3
XFILLER_26_239 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _174_/Y mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_27_43 vpwr vgnd scs8hd_fill_2
XFILLER_17_217 vgnd vpwr scs8hd_decap_3
XFILLER_4_154 vgnd vpwr scs8hd_decap_4
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XANTENNA__139__A _085_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_12 vpwr vgnd scs8hd_fill_2
XFILLER_13_56 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_97 vgnd vpwr scs8hd_fill_1
XFILLER_38_86 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_253 vpwr vgnd scs8hd_fill_2
XFILLER_13_275 vpwr vgnd scs8hd_fill_2
XANTENNA__141__B _138_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_3
XFILLER_24_66 vgnd vpwr scs8hd_decap_3
XFILLER_24_44 vgnd vpwr scs8hd_decap_8
XFILLER_6_205 vgnd vpwr scs8hd_decap_8
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
XFILLER_10_201 vpwr vgnd scs8hd_fill_2
X_091_ _090_/X _121_/A vgnd vpwr scs8hd_buf_1
X_160_ _170_/A _161_/A vgnd vpwr scs8hd_buf_1
XFILLER_1_26 vgnd vpwr scs8hd_decap_12
XFILLER_1_48 vgnd vpwr scs8hd_decap_8
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XANTENNA__152__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_175 vgnd vpwr scs8hd_decap_12
XFILLER_27_153 vgnd vpwr scs8hd_fill_1
XFILLER_27_142 vpwr vgnd scs8hd_fill_2
XFILLER_19_11 vgnd vpwr scs8hd_decap_3
XFILLER_19_66 vgnd vpwr scs8hd_decap_4
XFILLER_19_109 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_42_123 vgnd vpwr scs8hd_fill_1
XFILLER_35_98 vpwr vgnd scs8hd_fill_2
X_212_ chany_top_in[4] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
X_143_ _123_/A _138_/X _143_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_123 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_120 vpwr vgnd scs8hd_fill_2
XANTENNA__147__A _146_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_189 vpwr vgnd scs8hd_fill_2
XFILLER_24_112 vpwr vgnd scs8hd_fill_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_9 vgnd vpwr scs8hd_decap_3
Xmux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _180_/Y mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_15_112 vgnd vpwr scs8hd_decap_4
XFILLER_15_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_156 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[5] mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_126_ _146_/B _168_/B vgnd vpwr scs8hd_buf_1
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[8] mux_right_track_10.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_16_12 vpwr vgnd scs8hd_fill_2
XFILLER_16_23 vgnd vpwr scs8hd_decap_8
XFILLER_32_66 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _186_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__144__B _138_/X vgnd vpwr scs8hd_diode_2
X_109_ _109_/A _110_/B _109_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__160__A _170_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_66 vpwr vgnd scs8hd_fill_2
XFILLER_17_229 vgnd vpwr scs8hd_decap_3
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_100 vgnd vpwr scs8hd_decap_4
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_232 vgnd vpwr scs8hd_decap_12
XANTENNA__139__B _138_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__155__A _170_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A bottom_left_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_13_35 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_258 vpwr vgnd scs8hd_fill_2
XFILLER_0_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_66 vgnd vpwr scs8hd_decap_3
XFILLER_6_239 vgnd vpwr scs8hd_decap_12
XFILLER_10_213 vgnd vpwr scs8hd_fill_1
X_090_ _093_/A address[2] _171_/D _090_/X vgnd vpwr scs8hd_or3_4
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_40_88 vgnd vpwr scs8hd_decap_4
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _182_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_38 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB _172_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__152__B _150_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_187 vgnd vpwr scs8hd_decap_12
Xmem_right_track_2.LATCH_0_.latch data_in _174_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_45 vpwr vgnd scs8hd_fill_2
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
X_211_ chany_top_in[5] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
X_142_ _122_/A _138_/X _142_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A bottom_left_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_157 vpwr vgnd scs8hd_fill_2
XFILLER_33_102 vpwr vgnd scs8hd_fill_2
XANTENNA__163__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_102 vgnd vpwr scs8hd_fill_1
XFILLER_24_168 vpwr vgnd scs8hd_fill_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
X_125_ address[6] _146_/B vgnd vpwr scs8hd_inv_8
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XANTENNA__158__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_21_138 vgnd vpwr scs8hd_decap_4
XFILLER_21_149 vpwr vgnd scs8hd_fill_2
XFILLER_32_89 vgnd vpwr scs8hd_decap_3
Xmem_top_track_0.LATCH_2_.latch data_in mem_top_track_0.LATCH_2_.latch/Q _095_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_116 vgnd vpwr scs8hd_decap_3
XFILLER_20_182 vpwr vgnd scs8hd_fill_2
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
X_108_ _085_/A _110_/B _108_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
XFILLER_7_197 vpwr vgnd scs8hd_fill_2
XFILLER_11_171 vpwr vgnd scs8hd_fill_2
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB _167_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _177_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _222_/A vgnd vpwr scs8hd_inv_1
XFILLER_17_208 vgnd vpwr scs8hd_decap_3
XFILLER_40_200 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _191_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_134 vgnd vpwr scs8hd_decap_4
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__171__A _154_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_104 vgnd vpwr scs8hd_decap_8
XANTENNA__081__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_233 vgnd vpwr scs8hd_decap_6
XANTENNA__166__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_163 vpwr vgnd scs8hd_fill_2
XANTENNA__076__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_5_262 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_1.LATCH_4_.latch data_in mem_bottom_track_1.LATCH_4_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_144 vpwr vgnd scs8hd_fill_2
XFILLER_36_111 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_199 vgnd vpwr scs8hd_decap_12
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_103 vpwr vgnd scs8hd_fill_2
XFILLER_27_177 vgnd vpwr scs8hd_decap_4
XFILLER_27_100 vgnd vpwr scs8hd_decap_3
XFILLER_19_57 vgnd vpwr scs8hd_decap_4
XFILLER_35_78 vgnd vpwr scs8hd_decap_3
X_210_ chany_top_in[6] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
X_141_ _121_/A _138_/X _141_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_3_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_136 vpwr vgnd scs8hd_fill_2
XFILLER_33_114 vpwr vgnd scs8hd_fill_2
XANTENNA__163__B _163_/B vgnd vpwr scs8hd_diode_2
Xmem_right_track_14.LATCH_1_.latch data_in _185_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _183_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_60 vgnd vpwr scs8hd_decap_6
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_58 vgnd vpwr scs8hd_decap_3
XFILLER_30_106 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_124_ _124_/A _121_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_191 vpwr vgnd scs8hd_fill_2
XFILLER_23_180 vgnd vpwr scs8hd_decap_3
XFILLER_7_27 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_5_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__174__A _174_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr
+ scs8hd_diode_2
XANTENNA__084__A _083_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
X_107_ _106_/X _110_/B vgnd vpwr scs8hd_buf_1
XFILLER_22_90 vpwr vgnd scs8hd_fill_2
XFILLER_14_3 vgnd vpwr scs8hd_decap_8
XANTENNA__169__A _170_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XANTENNA__079__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_40_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_27_79 vpwr vgnd scs8hd_fill_2
XFILLER_25_242 vpwr vgnd scs8hd_fill_2
XFILLER_4_113 vgnd vpwr scs8hd_decap_8
XFILLER_4_179 vgnd vpwr scs8hd_fill_1
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_12
XANTENNA__171__B _168_/B vgnd vpwr scs8hd_diode_2
XANTENNA__081__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_1_138 vpwr vgnd scs8hd_fill_2
XFILLER_9_205 vgnd vpwr scs8hd_decap_4
XFILLER_9_216 vpwr vgnd scs8hd_fill_2
XFILLER_13_212 vpwr vgnd scs8hd_fill_2
XFILLER_13_245 vgnd vpwr scs8hd_decap_8
XFILLER_0_171 vpwr vgnd scs8hd_fill_2
XANTENNA__166__B _170_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr
+ scs8hd_diode_2
XANTENNA__182__A _182_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_260 vgnd vpwr scs8hd_decap_12
XFILLER_39_175 vpwr vgnd scs8hd_fill_2
XFILLER_39_153 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_226 vgnd vpwr scs8hd_decap_12
XFILLER_10_259 vgnd vpwr scs8hd_decap_12
XANTENNA__092__A _085_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_274 vgnd vpwr scs8hd_decap_3
XFILLER_36_167 vgnd vpwr scs8hd_decap_4
XFILLER_36_123 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__177__A _177_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_35_57 vpwr vgnd scs8hd_fill_2
XFILLER_35_35 vgnd vpwr scs8hd_fill_1
XFILLER_27_156 vpwr vgnd scs8hd_fill_2
XANTENNA__087__A _086_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_140_ _109_/A _138_/X _140_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_16.LATCH_4_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_bottom_track_9.INVTX1_2_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_145 vpwr vgnd scs8hd_fill_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__163__C _163_/C vgnd vpwr scs8hd_diode_2
XFILLER_24_148 vgnd vpwr scs8hd_decap_3
XFILLER_2_83 vgnd vpwr scs8hd_fill_1
XFILLER_32_181 vgnd vpwr scs8hd_decap_12
XFILLER_21_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_48 vgnd vpwr scs8hd_decap_8
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_123_ _123_/A _121_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
Xmem_top_track_8.LATCH_3_.latch data_in mem_top_track_8.LATCH_3_.latch/Q _110_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_47 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_162 vgnd vpwr scs8hd_fill_1
XFILLER_28_251 vgnd vpwr scs8hd_decap_12
XFILLER_11_184 vgnd vpwr scs8hd_decap_6
XFILLER_11_195 vpwr vgnd scs8hd_fill_2
X_106_ _083_/A _170_/B _163_/C _106_/X vgnd vpwr scs8hd_or3_4
XANTENNA__169__B _170_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A _185_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_60 vgnd vpwr scs8hd_decap_3
XFILLER_8_82 vgnd vpwr scs8hd_decap_4
XFILLER_27_47 vgnd vpwr scs8hd_decap_3
XFILLER_25_210 vgnd vpwr scs8hd_decap_12
XANTENNA__095__A _085_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_158 vgnd vpwr scs8hd_fill_1
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XANTENNA__171__C _163_/C vgnd vpwr scs8hd_diode_2
XFILLER_22_224 vgnd vpwr scs8hd_decap_12
XFILLER_13_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__081__C _115_/C vgnd vpwr scs8hd_diode_2
XFILLER_38_57 vpwr vgnd scs8hd_fill_2
XFILLER_38_46 vpwr vgnd scs8hd_fill_2
XFILLER_1_117 vgnd vpwr scs8hd_decap_4
XFILLER_0_183 vgnd vpwr scs8hd_decap_3
XANTENNA__166__C _165_/C vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[4] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_272 vgnd vpwr scs8hd_decap_3
XFILLER_39_132 vpwr vgnd scs8hd_fill_2
XFILLER_5_94 vpwr vgnd scs8hd_fill_2
XFILLER_5_83 vpwr vgnd scs8hd_fill_2
XFILLER_39_187 vpwr vgnd scs8hd_fill_2
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XANTENNA__092__B _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_205 vgnd vpwr scs8hd_decap_8
XFILLER_10_238 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_253 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_5_.latch data_in mem_bottom_track_9.LATCH_5_.latch/Q _139_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_70 vgnd vpwr scs8hd_decap_3
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
XFILLER_30_91 vgnd vpwr scs8hd_fill_1
XFILLER_36_135 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _185_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_5_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_124 vpwr vgnd scs8hd_fill_2
XFILLER_18_157 vpwr vgnd scs8hd_fill_2
XFILLER_41_182 vgnd vpwr scs8hd_fill_1
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_199_ _199_/HI _199_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__163__D _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _192_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_116 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_4_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_32_193 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_4_.scs8hd_inv_1 chanx_right_in[5] mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_27 vgnd vpwr scs8hd_decap_6
XANTENNA__098__A _085_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_119 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_127 vgnd vpwr scs8hd_decap_4
X_122_ _122_/A _121_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_5_.latch data_in mem_top_track_16.LATCH_5_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_208 vgnd vpwr scs8hd_decap_12
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
Xmem_right_track_10.LATCH_1_.latch data_in _179_/A _165_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_141 vgnd vpwr scs8hd_fill_1
XFILLER_28_263 vgnd vpwr scs8hd_decap_12
XFILLER_22_70 vgnd vpwr scs8hd_decap_3
XFILLER_7_134 vpwr vgnd scs8hd_fill_2
XFILLER_7_156 vpwr vgnd scs8hd_fill_2
XFILLER_11_130 vpwr vgnd scs8hd_fill_2
X_105_ _105_/A _163_/C vgnd vpwr scs8hd_buf_1
XANTENNA__169__C _170_/C vgnd vpwr scs8hd_diode_2
XFILLER_34_211 vgnd vpwr scs8hd_decap_3
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
XFILLER_25_222 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__095__B _122_/A vgnd vpwr scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_222 vpwr vgnd scs8hd_fill_2
XFILLER_16_233 vgnd vpwr scs8hd_decap_8
XFILLER_16_244 vgnd vpwr scs8hd_decap_8
XFILLER_16_255 vgnd vpwr scs8hd_decap_12
XFILLER_17_92 vgnd vpwr scs8hd_decap_4
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
XANTENNA__171__D _171_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_236 vgnd vpwr scs8hd_decap_12
XFILLER_13_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_80 vgnd vpwr scs8hd_decap_6
XFILLER_0_195 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__166__D _164_/D vgnd vpwr scs8hd_diode_2
XFILLER_5_62 vpwr vgnd scs8hd_fill_2
XFILLER_5_51 vgnd vpwr scs8hd_decap_4
XFILLER_39_111 vpwr vgnd scs8hd_fill_2
XFILLER_39_199 vpwr vgnd scs8hd_fill_2
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _184_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_17.LATCH_5_.latch data_in mem_bottom_track_17.LATCH_5_.latch/Q _148_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_114 vgnd vpwr scs8hd_decap_3
XFILLER_19_49 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_128 vgnd vpwr scs8hd_decap_12
XFILLER_2_202 vgnd vpwr scs8hd_decap_12
XFILLER_33_106 vpwr vgnd scs8hd_fill_2
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XFILLER_25_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _187_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_198_ _198_/HI _198_/LO vgnd vpwr scs8hd_conb_1
Xmux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_180 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[4] mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_right_track_6.LATCH_1_.latch data_in _177_/A _163_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__098__B _123_/A vgnd vpwr scs8hd_diode_2
X_121_ _121_/A _121_/B _121_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_172 vpwr vgnd scs8hd_fill_2
XFILLER_23_150 vgnd vpwr scs8hd_decap_3
XFILLER_16_9 vgnd vpwr scs8hd_fill_1
XFILLER_36_91 vgnd vpwr scs8hd_fill_1
XFILLER_14_161 vgnd vpwr scs8hd_decap_3
XFILLER_14_183 vgnd vpwr scs8hd_decap_8
XFILLER_37_220 vgnd vpwr scs8hd_decap_12
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_120 vpwr vgnd scs8hd_fill_2
XFILLER_20_186 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _178_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_93 vgnd vpwr scs8hd_fill_1
XFILLER_22_82 vpwr vgnd scs8hd_fill_2
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
XFILLER_11_153 vgnd vpwr scs8hd_fill_1
XFILLER_11_175 vgnd vpwr scs8hd_decap_8
X_104_ _103_/Y address[4] _115_/C _105_/A vgnd vpwr scs8hd_or3_4
XANTENNA__169__D _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_8_40 vgnd vpwr scs8hd_fill_1
XFILLER_27_27 vgnd vpwr scs8hd_decap_12
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_25_245 vgnd vpwr scs8hd_decap_12
XFILLER_25_234 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_267 vgnd vpwr scs8hd_decap_8
XFILLER_3_182 vgnd vpwr scs8hd_fill_1
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_22_248 vgnd vpwr scs8hd_decap_12
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_13_259 vpwr vgnd scs8hd_fill_2
XFILLER_39_167 vpwr vgnd scs8hd_fill_2
XFILLER_39_156 vgnd vpwr scs8hd_decap_3
XFILLER_40_49 vgnd vpwr scs8hd_decap_8
XFILLER_40_38 vgnd vpwr scs8hd_decap_6
XFILLER_10_218 vpwr vgnd scs8hd_fill_2
XFILLER_36_148 vgnd vpwr scs8hd_decap_4
XFILLER_19_17 vpwr vgnd scs8hd_fill_2
XFILLER_19_28 vpwr vgnd scs8hd_fill_2
XFILLER_42_107 vgnd vpwr scs8hd_decap_12
XFILLER_35_38 vpwr vgnd scs8hd_fill_2
XFILLER_35_27 vgnd vpwr scs8hd_decap_8
XFILLER_27_126 vpwr vgnd scs8hd_fill_2
XFILLER_35_181 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.tap_buf4_0_.scs8hd_inv_1 mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _201_/A vgnd vpwr scs8hd_inv_1
XFILLER_41_140 vgnd vpwr scs8hd_decap_12
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XFILLER_33_118 vpwr vgnd scs8hd_fill_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XFILLER_41_162 vgnd vpwr scs8hd_decap_12
X_197_ _197_/HI _197_/LO vgnd vpwr scs8hd_conb_1
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _218_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_86 vgnd vpwr scs8hd_decap_6
XFILLER_24_129 vpwr vgnd scs8hd_fill_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
X_120_ _109_/A _121_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_195 vpwr vgnd scs8hd_fill_2
XFILLER_23_184 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_51 vpwr vgnd scs8hd_fill_2
XFILLER_11_62 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_154 vpwr vgnd scs8hd_fill_2
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
X_103_ address[3] _103_/Y vgnd vpwr scs8hd_inv_8
XFILLER_19_243 vgnd vpwr scs8hd_fill_1
XFILLER_8_74 vpwr vgnd scs8hd_fill_2
XFILLER_27_39 vpwr vgnd scs8hd_fill_2
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_25_257 vgnd vpwr scs8hd_decap_12
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_161 vgnd vpwr scs8hd_decap_12
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
XFILLER_13_216 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_175 vgnd vpwr scs8hd_decap_8
XFILLER_12_271 vgnd vpwr scs8hd_decap_4
XFILLER_39_179 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_51 vgnd vpwr scs8hd_decap_8
XFILLER_14_62 vpwr vgnd scs8hd_fill_2
XFILLER_14_84 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _204_/A vgnd vpwr scs8hd_inv_1
XFILLER_30_61 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_245 vgnd vpwr scs8hd_decap_8
XANTENNA__101__A _085_/B vgnd vpwr scs8hd_diode_2
XFILLER_42_119 vgnd vpwr scs8hd_decap_4
XFILLER_27_149 vgnd vpwr scs8hd_decap_4
XFILLER_27_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_215 vgnd vpwr scs8hd_decap_8
XFILLER_18_105 vpwr vgnd scs8hd_fill_2
XFILLER_18_116 vpwr vgnd scs8hd_fill_2
XFILLER_18_149 vgnd vpwr scs8hd_decap_4
XPHY_83 vgnd vpwr scs8hd_decap_3
XFILLER_41_174 vgnd vpwr scs8hd_decap_8
XFILLER_41_152 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_25_94 vpwr vgnd scs8hd_fill_2
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
XFILLER_41_82 vpwr vgnd scs8hd_fill_2
XFILLER_41_60 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
X_196_ _196_/HI _196_/LO vgnd vpwr scs8hd_conb_1
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_5_ mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_32_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _187_/HI mem_bottom_track_1.LATCH_2_.latch/Q
+ mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_8
XFILLER_11_74 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_93 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_141 vgnd vpwr scs8hd_decap_8
X_179_ _179_/A _179_/Y vgnd vpwr scs8hd_inv_8
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_20_133 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_211 vgnd vpwr scs8hd_decap_3
Xmem_right_track_2.LATCH_1_.latch data_in _173_/A _157_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_199 vpwr vgnd scs8hd_fill_2
X_102_ address[6] _170_/B vgnd vpwr scs8hd_buf_1
XFILLER_34_203 vgnd vpwr scs8hd_decap_8
XFILLER_8_86 vgnd vpwr scs8hd_fill_1
Xmux_right_track_2.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_192 vgnd vpwr scs8hd_decap_4
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_25_269 vgnd vpwr scs8hd_decap_8
XFILLER_17_51 vpwr vgnd scs8hd_fill_2
XFILLER_17_62 vpwr vgnd scs8hd_fill_2
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_83 vpwr vgnd scs8hd_fill_2
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XFILLER_3_173 vgnd vpwr scs8hd_decap_6
XFILLER_3_151 vgnd vpwr scs8hd_decap_8
XFILLER_3_140 vgnd vpwr scs8hd_decap_4
XANTENNA__104__A _103_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_206 vgnd vpwr scs8hd_decap_8
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_121 vgnd vpwr scs8hd_decap_3
XFILLER_28_50 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_3_.latch data_in mem_top_track_0.LATCH_3_.latch/Q _092_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_98 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_9.LATCH_0_.latch data_in mem_bottom_track_9.LATCH_0_.latch/Q _144_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_136 vpwr vgnd scs8hd_fill_2
XFILLER_40_18 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_191 vgnd vpwr scs8hd_decap_12
XFILLER_5_202 vgnd vpwr scs8hd_decap_12
XFILLER_14_96 vpwr vgnd scs8hd_fill_2
XFILLER_30_84 vgnd vpwr scs8hd_fill_1
XFILLER_39_93 vgnd vpwr scs8hd_decap_3
XFILLER_39_82 vpwr vgnd scs8hd_fill_2
XANTENNA__101__B _124_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_2_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 top_left_grid_pin_9_ mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_84 vgnd vpwr scs8hd_decap_3
XFILLER_41_131 vgnd vpwr scs8hd_fill_1
XFILLER_41_120 vpwr vgnd scs8hd_fill_2
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_194 vgnd vpwr scs8hd_decap_8
XFILLER_26_161 vpwr vgnd scs8hd_fill_2
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_73 vpwr vgnd scs8hd_fill_2
XFILLER_25_62 vpwr vgnd scs8hd_fill_2
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
X_195_ _195_/HI _195_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__112__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_77 vgnd vpwr scs8hd_decap_6
XFILLER_2_44 vpwr vgnd scs8hd_fill_2
XFILLER_2_11 vgnd vpwr scs8hd_fill_1
XFILLER_1_260 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_161 vgnd vpwr scs8hd_decap_4
XFILLER_17_172 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_0_.latch data_in mem_top_track_16.LATCH_0_.latch/Q _124_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_31 vgnd vpwr scs8hd_fill_1
XFILLER_11_97 vpwr vgnd scs8hd_fill_2
XFILLER_36_83 vgnd vpwr scs8hd_decap_8
XFILLER_36_72 vpwr vgnd scs8hd_fill_2
XANTENNA__107__A _106_/X vgnd vpwr scs8hd_diode_2
X_178_ _178_/A _178_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_245 vgnd vpwr scs8hd_decap_12
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_5_.latch data_in mem_bottom_track_1.LATCH_5_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_101_ _085_/B _124_/A _101_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_138 vpwr vgnd scs8hd_fill_2
XFILLER_11_112 vpwr vgnd scs8hd_fill_2
XFILLER_11_134 vpwr vgnd scs8hd_fill_2
XFILLER_11_156 vgnd vpwr scs8hd_decap_4
XFILLER_19_245 vgnd vpwr scs8hd_decap_12
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_32 vgnd vpwr scs8hd_decap_8
XFILLER_8_43 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB _092_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_7_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__210__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _183_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_215 vgnd vpwr scs8hd_decap_4
XFILLER_17_30 vpwr vgnd scs8hd_fill_2
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_4
XFILLER_3_196 vgnd vpwr scs8hd_decap_12
XANTENNA__104__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _153_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_229 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__205__A _205_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_73 vgnd vpwr scs8hd_decap_4
XFILLER_28_40 vgnd vpwr scs8hd_fill_1
XFILLER_8_211 vgnd vpwr scs8hd_decap_3
XFILLER_12_240 vgnd vpwr scs8hd_decap_4
XANTENNA__115__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_39_115 vgnd vpwr scs8hd_decap_4
XFILLER_5_77 vgnd vpwr scs8hd_decap_4
XFILLER_5_66 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_17.LATCH_0_.latch data_in mem_bottom_track_17.LATCH_0_.latch/Q _153_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_4_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_5_258 vpwr vgnd scs8hd_fill_2
XFILLER_5_214 vgnd vpwr scs8hd_decap_12
XFILLER_29_181 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_3_ vgnd vpwr scs8hd_diode_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XFILLER_35_173 vgnd vpwr scs8hd_decap_8
XFILLER_35_151 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr
+ scs8hd_diode_2
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_41_95 vpwr vgnd scs8hd_fill_2
XFILLER_41_73 vpwr vgnd scs8hd_fill_2
X_194_ _194_/HI _194_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__112__B _110_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_272 vgnd vpwr scs8hd_decap_4
XFILLER_17_140 vpwr vgnd scs8hd_fill_2
XFILLER_17_184 vgnd vpwr scs8hd_decap_3
XFILLER_23_176 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__213__A _213_/A vgnd vpwr scs8hd_diode_2
X_177_ _177_/A _177_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XFILLER_20_102 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A bottom_left_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__208__A right_top_grid_pin_10_ vgnd vpwr scs8hd_diode_2
X_100_ _100_/A _124_/A vgnd vpwr scs8hd_buf_1
XFILLER_22_86 vpwr vgnd scs8hd_fill_2
XFILLER_19_213 vpwr vgnd scs8hd_fill_2
XFILLER_19_224 vpwr vgnd scs8hd_fill_2
XFILLER_19_235 vpwr vgnd scs8hd_fill_2
XFILLER_19_257 vgnd vpwr scs8hd_decap_12
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _117_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_55 vgnd vpwr scs8hd_decap_3
XFILLER_10_190 vpwr vgnd scs8hd_fill_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_75 vpwr vgnd scs8hd_fill_2
XANTENNA__104__C _115_/C vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__221__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
Xmem_top_track_8.LATCH_4_.latch data_in mem_top_track_8.LATCH_4_.latch/Q _109_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__115__B _114_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_32 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_5_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_5_226 vgnd vpwr scs8hd_decap_12
XANTENNA__216__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_39_62 vgnd vpwr scs8hd_decap_4
XFILLER_39_40 vpwr vgnd scs8hd_fill_2
XANTENNA__126__A _146_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_119 vgnd vpwr scs8hd_decap_3
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_141 vgnd vpwr scs8hd_decap_12
XFILLER_26_130 vpwr vgnd scs8hd_fill_2
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_41_52 vgnd vpwr scs8hd_decap_8
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_193_ _193_/HI _193_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_251 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_55 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_track_1.LATCH_3_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_100 vpwr vgnd scs8hd_fill_2
XFILLER_14_122 vpwr vgnd scs8hd_fill_2
X_176_ _176_/A _176_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__B _121_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XFILLER_20_158 vgnd vpwr scs8hd_decap_4
XFILLER_9_181 vpwr vgnd scs8hd_fill_2
XANTENNA__224__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_65 vgnd vpwr scs8hd_decap_3
XFILLER_22_54 vpwr vgnd scs8hd_fill_2
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_19_269 vgnd vpwr scs8hd_decap_8
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_6_173 vgnd vpwr scs8hd_decap_6
XFILLER_8_78 vpwr vgnd scs8hd_fill_2
XFILLER_8_89 vgnd vpwr scs8hd_decap_3
X_159_ _154_/X _163_/B _165_/C _164_/D _159_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__134__A _124_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_206 vgnd vpwr scs8hd_decap_8
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__219__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_53 vpwr vgnd scs8hd_fill_2
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_98 vpwr vgnd scs8hd_fill_2
XFILLER_3_132 vgnd vpwr scs8hd_decap_6
XANTENNA__129__A _085_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_220 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_102 vgnd vpwr scs8hd_decap_4
XFILLER_0_113 vgnd vpwr scs8hd_decap_8
XFILLER_28_86 vgnd vpwr scs8hd_fill_1
XFILLER_8_224 vgnd vpwr scs8hd_decap_12
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XANTENNA__131__B _134_/B vgnd vpwr scs8hd_diode_2
XANTENNA__115__C _115_/C vgnd vpwr scs8hd_diode_2
XFILLER_14_11 vgnd vpwr scs8hd_decap_3
XFILLER_14_66 vpwr vgnd scs8hd_fill_2
XFILLER_14_88 vgnd vpwr scs8hd_decap_4
XFILLER_30_87 vgnd vpwr scs8hd_decap_4
XFILLER_30_65 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_238 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_271 vgnd vpwr scs8hd_decap_4
XANTENNA__142__A _122_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_bottom_track_9.LATCH_5_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_17.INVTX1_5_.scs8hd_inv_1 bottom_left_grid_pin_3_ mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_109 vpwr vgnd scs8hd_fill_2
XFILLER_41_123 vpwr vgnd scs8hd_fill_2
XFILLER_41_112 vgnd vpwr scs8hd_decap_8
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_43 vgnd vpwr scs8hd_fill_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_25_98 vpwr vgnd scs8hd_fill_2
X_192_ _192_/HI _192_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_230 vgnd vpwr scs8hd_decap_12
Xmux_right_track_14.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[3] mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_145 vgnd vpwr scs8hd_decap_8
XFILLER_32_134 vpwr vgnd scs8hd_fill_2
XANTENNA__137__A _083_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_123 vgnd vpwr scs8hd_decap_3
XFILLER_11_34 vpwr vgnd scs8hd_fill_2
XFILLER_11_78 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_53 vgnd vpwr scs8hd_decap_4
X_175_ _175_/A _175_/Y vgnd vpwr scs8hd_inv_8
XFILLER_20_137 vpwr vgnd scs8hd_fill_2
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_126 vpwr vgnd scs8hd_fill_2
XFILLER_22_44 vgnd vpwr scs8hd_fill_1
Xmux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_2_.scs8hd_inv_1/Y
+ _178_/A mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XFILLER_6_163 vgnd vpwr scs8hd_decap_8
X_089_ address[1] _093_/A vgnd vpwr scs8hd_inv_8
XANTENNA__134__B _134_/B vgnd vpwr scs8hd_diode_2
X_158_ address[0] _164_/D vgnd vpwr scs8hd_buf_1
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XANTENNA__150__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_55 vpwr vgnd scs8hd_fill_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vpwr vgnd scs8hd_fill_2
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_251 vgnd vpwr scs8hd_decap_12
XANTENNA__129__B _134_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_251 vgnd vpwr scs8hd_fill_1
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_0_91 vpwr vgnd scs8hd_fill_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_8
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
XFILLER_8_203 vgnd vpwr scs8hd_decap_8
XFILLER_8_236 vgnd vpwr scs8hd_decap_12
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_23 vgnd vpwr scs8hd_decap_8
XFILLER_39_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XFILLER_29_173 vgnd vpwr scs8hd_decap_8
XFILLER_29_151 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__B _138_/X vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _197_/HI mem_top_track_0.LATCH_2_.latch/Q
+ mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_165 vgnd vpwr scs8hd_decap_3
XFILLER_25_77 vpwr vgnd scs8hd_fill_2
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_41_65 vgnd vpwr scs8hd_decap_8
X_191_ _191_/HI _191_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_242 vpwr vgnd scs8hd_fill_2
XFILLER_17_176 vpwr vgnd scs8hd_fill_2
XFILLER_32_157 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__137__B _168_/B vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _124_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_146 vpwr vgnd scs8hd_fill_2
XFILLER_23_135 vpwr vgnd scs8hd_fill_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_1.LATCH_0_.latch data_in mem_bottom_track_1.LATCH_0_.latch/Q _134_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_157 vpwr vgnd scs8hd_fill_2
X_174_ _174_/A _174_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__148__A _085_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[1] mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_116 vpwr vgnd scs8hd_fill_2
XFILLER_20_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_227 vgnd vpwr scs8hd_decap_12
XFILLER_3_80 vpwr vgnd scs8hd_fill_2
XFILLER_11_116 vgnd vpwr scs8hd_decap_4
XFILLER_11_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_4_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_226_ _226_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
X_157_ _154_/X _163_/B _165_/C _163_/D _157_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_40_6 vgnd vpwr scs8hd_decap_12
X_088_ _085_/B _109_/A _088_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__150__B _150_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_8
XFILLER_18_271 vgnd vpwr scs8hd_decap_4
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_263 vgnd vpwr scs8hd_decap_12
XFILLER_16_219 vgnd vpwr scs8hd_fill_1
XFILLER_17_34 vpwr vgnd scs8hd_fill_2
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_101 vpwr vgnd scs8hd_fill_2
XFILLER_15_263 vgnd vpwr scs8hd_decap_12
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
X_209_ _209_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_137 vgnd vpwr scs8hd_decap_12
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_248 vgnd vpwr scs8hd_decap_12
XFILLER_39_119 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.tap_buf4_0_.scs8hd_inv_1 mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _203_/A vgnd vpwr scs8hd_inv_1
XANTENNA__156__A _171_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_21 vgnd vpwr scs8hd_decap_12
XFILLER_39_10 vpwr vgnd scs8hd_fill_2
XFILLER_30_78 vgnd vpwr scs8hd_decap_6
XFILLER_39_98 vpwr vgnd scs8hd_fill_2
XFILLER_29_196 vgnd vpwr scs8hd_decap_12
XFILLER_4_251 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 top_left_grid_pin_7_ mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_80 vgnd vpwr scs8hd_fill_1
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_158 vpwr vgnd scs8hd_fill_2
XFILLER_41_136 vpwr vgnd scs8hd_fill_2
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_177 vgnd vpwr scs8hd_decap_6
XPHY_45 vgnd vpwr scs8hd_decap_3
X_190_ _190_/HI _190_/LO vgnd vpwr scs8hd_conb_1
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XFILLER_41_99 vpwr vgnd scs8hd_fill_2
XFILLER_2_49 vgnd vpwr scs8hd_decap_8
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_276 vgnd vpwr scs8hd_fill_1
XFILLER_32_169 vgnd vpwr scs8hd_decap_12
XANTENNA__153__B _150_/B vgnd vpwr scs8hd_diode_2
XANTENNA__137__C _165_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _174_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
XFILLER_23_103 vpwr vgnd scs8hd_fill_2
XFILLER_36_99 vgnd vpwr scs8hd_fill_1
XFILLER_22_191 vpwr vgnd scs8hd_fill_2
X_173_ _173_/A _173_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__148__B _150_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_151 vpwr vgnd scs8hd_fill_2
XFILLER_9_184 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__164__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_239 vgnd vpwr scs8hd_decap_12
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XFILLER_19_217 vgnd vpwr scs8hd_decap_4
XFILLER_19_228 vgnd vpwr scs8hd_decap_4
XFILLER_19_239 vgnd vpwr scs8hd_decap_4
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
X_225_ chany_bottom_in[0] chany_top_out[1] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_1.INVTX1_7_.scs8hd_inv_1 bottom_left_grid_pin_11_ mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_194 vgnd vpwr scs8hd_decap_4
X_156_ _171_/D _163_/D vgnd vpwr scs8hd_buf_1
X_087_ _086_/X _109_/A vgnd vpwr scs8hd_buf_1
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
XANTENNA__159__A _154_/X vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[1] mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_13 vpwr vgnd scs8hd_fill_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_10.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[2] mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_79 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_179 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_275 vpwr vgnd scs8hd_fill_2
XANTENNA__161__B _163_/B vgnd vpwr scs8hd_diode_2
X_208_ right_top_grid_pin_10_ chanx_right_out[0] vgnd vpwr scs8hd_buf_2
X_139_ _085_/A _138_/X _139_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.tap_buf4_0_.scs8hd_inv_1 mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _206_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_190 vgnd vpwr scs8hd_decap_12
XFILLER_0_71 vgnd vpwr scs8hd_decap_12
XFILLER_21_245 vgnd vpwr scs8hd_decap_12
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_89 vgnd vpwr scs8hd_decap_3
XFILLER_12_201 vpwr vgnd scs8hd_fill_2
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _154_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_46 vgnd vpwr scs8hd_decap_6
XANTENNA__082__A _082_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_66 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_20_90 vpwr vgnd scs8hd_fill_2
XFILLER_35_156 vgnd vpwr scs8hd_decap_3
XFILLER_35_134 vpwr vgnd scs8hd_fill_2
XFILLER_35_123 vpwr vgnd scs8hd_fill_2
XANTENNA__167__A _154_/X vgnd vpwr scs8hd_diode_2
XFILLER_25_35 vgnd vpwr scs8hd_decap_8
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A address[1] vgnd vpwr scs8hd_diode_2
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XFILLER_25_46 vpwr vgnd scs8hd_fill_2
XFILLER_41_78 vpwr vgnd scs8hd_fill_2
XFILLER_1_222 vpwr vgnd scs8hd_fill_2
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_32_126 vpwr vgnd scs8hd_fill_2
XFILLER_17_123 vpwr vgnd scs8hd_fill_2
XFILLER_17_167 vpwr vgnd scs8hd_fill_2
XFILLER_17_189 vpwr vgnd scs8hd_fill_2
XFILLER_40_181 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_4_.latch data_in mem_top_track_0.LATCH_4_.latch/Q _088_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_59 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_1_.latch data_in mem_bottom_track_9.LATCH_1_.latch/Q _143_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _183_/A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_14_104 vpwr vgnd scs8hd_fill_2
XFILLER_14_137 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_172_ _154_/X _168_/B _163_/C address[0] _172_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _193_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_170 vpwr vgnd scs8hd_fill_2
XANTENNA__164__B _163_/B vgnd vpwr scs8hd_diode_2
XANTENNA__180__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_93 vpwr vgnd scs8hd_fill_2
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[5] mux_right_track_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__090__A _093_/A vgnd vpwr scs8hd_diode_2
X_224_ chany_bottom_in[1] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_6_133 vpwr vgnd scs8hd_fill_2
XFILLER_6_188 vpwr vgnd scs8hd_fill_2
X_086_ address[1] _086_/B address[0] _086_/X vgnd vpwr scs8hd_or3_4
X_155_ _170_/B _163_/B vgnd vpwr scs8hd_buf_1
XFILLER_33_232 vgnd vpwr scs8hd_decap_12
XANTENNA__159__B _163_/B vgnd vpwr scs8hd_diode_2
XANTENNA__175__A _175_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_47 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__085__A _085_/A vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_68 vpwr vgnd scs8hd_fill_2
XFILLER_33_57 vpwr vgnd scs8hd_fill_2
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_79 vpwr vgnd scs8hd_fill_2
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_3_147 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_1_.latch data_in mem_top_track_16.LATCH_1_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_243 vgnd vpwr scs8hd_fill_1
XFILLER_30_213 vgnd vpwr scs8hd_fill_1
X_207_ _207_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_15_254 vgnd vpwr scs8hd_fill_1
XANTENNA__161__C _083_/C vgnd vpwr scs8hd_diode_2
X_138_ _137_/X _138_/X vgnd vpwr scs8hd_buf_1
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_2_.scs8hd_inv_1/Y
+ _176_/A mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_61 vgnd vpwr scs8hd_fill_1
XFILLER_0_83 vgnd vpwr scs8hd_decap_8
XFILLER_0_94 vgnd vpwr scs8hd_fill_1
XFILLER_21_224 vgnd vpwr scs8hd_decap_12
XFILLER_21_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_213 vgnd vpwr scs8hd_fill_1
XFILLER_12_224 vpwr vgnd scs8hd_fill_2
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
Xmem_right_track_12.LATCH_0_.latch data_in _182_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__172__B _168_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_89 vpwr vgnd scs8hd_fill_2
XFILLER_39_78 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_2_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_102 vgnd vpwr scs8hd_decap_3
XFILLER_35_168 vgnd vpwr scs8hd_decap_3
XANTENNA__183__A _183_/A vgnd vpwr scs8hd_diode_2
XANTENNA__167__B _168_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _226_/A vgnd vpwr scs8hd_inv_1
XFILLER_41_127 vgnd vpwr scs8hd_decap_4
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_157 vpwr vgnd scs8hd_fill_2
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XANTENNA__077__B _086_/B vgnd vpwr scs8hd_diode_2
XPHY_36 vgnd vpwr scs8hd_decap_3
XANTENNA__093__A _093_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_256 vpwr vgnd scs8hd_fill_2
XFILLER_1_245 vgnd vpwr scs8hd_decap_6
XFILLER_17_102 vgnd vpwr scs8hd_decap_3
XANTENNA__178__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_27 vgnd vpwr scs8hd_decap_4
XFILLER_11_38 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A _085_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_79 vpwr vgnd scs8hd_fill_2
XFILLER_36_68 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_149 vpwr vgnd scs8hd_fill_2
X_171_ _154_/X _168_/B _163_/C _171_/D _171_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_17.LATCH_1_.latch data_in mem_bottom_track_17.LATCH_1_.latch/Q _152_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_142 vpwr vgnd scs8hd_fill_2
XFILLER_9_164 vpwr vgnd scs8hd_fill_2
XFILLER_9_175 vgnd vpwr scs8hd_decap_4
XANTENNA__164__C _163_/C vgnd vpwr scs8hd_diode_2
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XFILLER_22_48 vgnd vpwr scs8hd_decap_4
XANTENNA__090__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_27_241 vgnd vpwr scs8hd_decap_3
Xmux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_2_.scs8hd_inv_1/Y
+ _182_/A mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
X_223_ chany_bottom_in[2] chany_top_out[3] vgnd vpwr scs8hd_buf_2
X_085_ _085_/A _085_/B _085_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_123 vgnd vpwr scs8hd_fill_1
XFILLER_6_145 vgnd vpwr scs8hd_decap_8
XFILLER_10_163 vpwr vgnd scs8hd_fill_2
XFILLER_12_81 vgnd vpwr scs8hd_decap_3
X_154_ _083_/A _154_/X vgnd vpwr scs8hd_buf_1
Xmux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__159__C _165_/C vgnd vpwr scs8hd_diode_2
XFILLER_17_59 vpwr vgnd scs8hd_fill_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__B _085_/B vgnd vpwr scs8hd_diode_2
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_4.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[6] mux_right_track_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_222 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_0_.latch data_in _184_/A _170_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_206_ _206_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
X_137_ _083_/A _168_/B _165_/C _137_/X vgnd vpwr scs8hd_or3_4
XANTENNA__161__D _163_/D vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_60 vgnd vpwr scs8hd_fill_1
XANTENNA__186__A _186_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_203 vpwr vgnd scs8hd_fill_2
XFILLER_21_236 vgnd vpwr scs8hd_decap_8
XFILLER_21_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_69 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _180_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__096__A address[1] vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_5_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_12_247 vgnd vpwr scs8hd_decap_12
XFILLER_18_91 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__172__C _163_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A top_left_grid_pin_9_ vgnd vpwr scs8hd_diode_2
XFILLER_38_122 vgnd vpwr scs8hd_fill_1
XFILLER_14_38 vpwr vgnd scs8hd_fill_2
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XFILLER_39_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_114 vpwr vgnd scs8hd_fill_2
XANTENNA__167__C _083_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_72 vpwr vgnd scs8hd_fill_2
XFILLER_34_191 vgnd vpwr scs8hd_decap_12
XPHY_59 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XANTENNA__077__C _171_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__093__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_136 vpwr vgnd scs8hd_fill_2
XFILLER_40_150 vgnd vpwr scs8hd_decap_3
Xmem_top_track_8.LATCH_5_.latch data_in mem_top_track_8.LATCH_5_.latch/Q _108_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_139 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A bottom_left_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__088__B _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_183 vgnd vpwr scs8hd_decap_8
X_170_ _170_/A _170_/B _170_/C _164_/D _170_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__164__D _164_/D vgnd vpwr scs8hd_diode_2
XFILLER_3_62 vgnd vpwr scs8hd_decap_3
XFILLER_3_51 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__090__C _171_/D vgnd vpwr scs8hd_diode_2
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XANTENNA__099__A address[1] vgnd vpwr scs8hd_diode_2
X_222_ _222_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
X_153_ _124_/A _150_/B _153_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_102 vgnd vpwr scs8hd_decap_3
XFILLER_8_29 vpwr vgnd scs8hd_fill_2
XFILLER_10_120 vgnd vpwr scs8hd_decap_3
X_084_ _083_/X _085_/B vgnd vpwr scs8hd_buf_1
XFILLER_12_93 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__159__D _164_/D vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr
+ scs8hd_diode_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_6.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_201 vpwr vgnd scs8hd_fill_2
XFILLER_15_245 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_205_ _205_/A chanx_right_out[3] vgnd vpwr scs8hd_buf_2
X_136_ _135_/X _165_/C vgnd vpwr scs8hd_buf_1
XFILLER_0_30 vgnd vpwr scs8hd_fill_1
XFILLER_0_63 vgnd vpwr scs8hd_fill_1
XFILLER_9_83 vpwr vgnd scs8hd_fill_2
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XANTENNA__096__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _197_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_259 vgnd vpwr scs8hd_decap_12
XFILLER_34_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _173_/A vgnd vpwr
+ scs8hd_diode_2
X_119_ _085_/A _121_/B _119_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_241 vgnd vpwr scs8hd_decap_3
XFILLER_7_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__172__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_38_145 vgnd vpwr scs8hd_decap_8
XFILLER_38_101 vgnd vpwr scs8hd_decap_8
Xmux_right_track_2.INVTX1_2_.scs8hd_inv_1 right_bottom_grid_pin_12_ mux_right_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
XFILLER_39_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_156 vgnd vpwr scs8hd_decap_6
XFILLER_29_134 vpwr vgnd scs8hd_fill_2
XFILLER_20_93 vgnd vpwr scs8hd_fill_1
XANTENNA__167__D _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_6_84 vpwr vgnd scs8hd_fill_2
XFILLER_26_137 vpwr vgnd scs8hd_fill_2
XFILLER_26_126 vpwr vgnd scs8hd_fill_2
XFILLER_25_27 vgnd vpwr scs8hd_decap_6
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_41_48 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XANTENNA__093__C address[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_4_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_71 vgnd vpwr scs8hd_decap_4
XFILLER_15_93 vpwr vgnd scs8hd_fill_2
XFILLER_31_81 vpwr vgnd scs8hd_fill_2
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XFILLER_23_107 vpwr vgnd scs8hd_fill_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_118 vpwr vgnd scs8hd_fill_2
XFILLER_22_195 vpwr vgnd scs8hd_fill_2
XFILLER_22_162 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XFILLER_9_100 vpwr vgnd scs8hd_fill_2
XFILLER_9_188 vpwr vgnd scs8hd_fill_2
XFILLER_13_195 vpwr vgnd scs8hd_fill_2
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__099__B address[2] vgnd vpwr scs8hd_diode_2
X_221_ chany_bottom_in[4] chany_top_out[5] vgnd vpwr scs8hd_buf_2
Xmux_top_track_8.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_083_ _083_/A address[6] _083_/C _083_/X vgnd vpwr scs8hd_or3_4
XFILLER_12_50 vpwr vgnd scs8hd_fill_2
X_152_ _123_/A _150_/B _152_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
Xmux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _177_/A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_202 vpwr vgnd scs8hd_fill_2
XFILLER_17_17 vpwr vgnd scs8hd_fill_2
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
XFILLER_30_205 vgnd vpwr scs8hd_decap_8
X_204_ _204_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_15_235 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_135_ _103_/Y _114_/Y _115_/C _135_/X vgnd vpwr scs8hd_or3_4
XFILLER_9_40 vpwr vgnd scs8hd_fill_2
XFILLER_9_62 vgnd vpwr scs8hd_decap_4
XFILLER_21_216 vpwr vgnd scs8hd_fill_2
XFILLER_0_109 vpwr vgnd scs8hd_fill_2
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_205 vgnd vpwr scs8hd_decap_8
XANTENNA__096__C _171_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_260 vgnd vpwr scs8hd_decap_12
XFILLER_18_60 vgnd vpwr scs8hd_decap_6
XFILLER_18_93 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
X_118_ _117_/X _121_/B vgnd vpwr scs8hd_buf_1
XFILLER_7_253 vpwr vgnd scs8hd_fill_2
XFILLER_7_275 vpwr vgnd scs8hd_fill_2
XFILLER_38_179 vgnd vpwr scs8hd_decap_12
XFILLER_38_168 vgnd vpwr scs8hd_decap_8
XFILLER_38_157 vgnd vpwr scs8hd_decap_8
XFILLER_38_135 vgnd vpwr scs8hd_fill_1
Xmem_right_track_4.LATCH_0_.latch data_in _176_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
XFILLER_29_102 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ _174_/A mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_20_61 vgnd vpwr scs8hd_fill_1
XFILLER_35_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_1_204 vgnd vpwr scs8hd_decap_12
XFILLER_1_226 vpwr vgnd scs8hd_fill_2
XFILLER_25_193 vpwr vgnd scs8hd_fill_2
XFILLER_15_50 vpwr vgnd scs8hd_fill_2
XFILLER_31_163 vgnd vpwr scs8hd_decap_12
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
Xmux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _185_/A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_36_49 vpwr vgnd scs8hd_fill_2
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XFILLER_14_108 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_141 vgnd vpwr scs8hd_decap_6
Xmux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _195_/HI _178_/Y mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_93 vpwr vgnd scs8hd_fill_2
XFILLER_9_134 vpwr vgnd scs8hd_fill_2
XFILLER_13_174 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_97 vpwr vgnd scs8hd_fill_2
XFILLER_36_211 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _194_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__099__C address[0] vgnd vpwr scs8hd_diode_2
X_220_ chany_bottom_in[5] chany_top_out[6] vgnd vpwr scs8hd_buf_2
X_151_ _122_/A _150_/B _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_115 vgnd vpwr scs8hd_decap_8
XFILLER_6_137 vgnd vpwr scs8hd_decap_3
X_082_ _082_/A _083_/C vgnd vpwr scs8hd_buf_1
Xmux_top_track_0.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[0] mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _198_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_211 vgnd vpwr scs8hd_decap_3
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_39 vgnd vpwr scs8hd_decap_3
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_203_ _203_/A chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_23_83 vpwr vgnd scs8hd_fill_2
X_134_ _124_/A _134_/B _134_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_10 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_2_.scs8hd_inv_1/Y
+ _180_/A mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_1.LATCH_1_.latch data_in mem_bottom_track_1.LATCH_1_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_32 vgnd vpwr scs8hd_decap_4
XFILLER_0_43 vgnd vpwr scs8hd_decap_12
XFILLER_0_98 vpwr vgnd scs8hd_fill_2
XFILLER_9_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_228 vgnd vpwr scs8hd_decap_12
XFILLER_20_272 vgnd vpwr scs8hd_decap_3
XFILLER_7_210 vgnd vpwr scs8hd_decap_4
XFILLER_11_261 vgnd vpwr scs8hd_decap_12
X_117_ _083_/A address[6] _170_/C _117_/X vgnd vpwr scs8hd_or3_4
XFILLER_38_125 vpwr vgnd scs8hd_fill_2
XFILLER_15_3 vgnd vpwr scs8hd_decap_6
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _184_/A mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_213 vgnd vpwr scs8hd_fill_1
XFILLER_20_73 vpwr vgnd scs8hd_fill_2
XFILLER_20_84 vgnd vpwr scs8hd_decap_4
XFILLER_34_150 vgnd vpwr scs8hd_fill_1
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_6
XFILLER_1_216 vpwr vgnd scs8hd_fill_2
XFILLER_40_142 vgnd vpwr scs8hd_decap_8
XFILLER_32_109 vgnd vpwr scs8hd_decap_6
XFILLER_31_94 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__102__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_16_150 vgnd vpwr scs8hd_decap_3
XFILLER_31_175 vgnd vpwr scs8hd_decap_8
XFILLER_31_142 vpwr vgnd scs8hd_fill_2
XFILLER_16_161 vgnd vpwr scs8hd_decap_4
XFILLER_16_194 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB _163_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_72 vgnd vpwr scs8hd_decap_3
XFILLER_9_113 vpwr vgnd scs8hd_fill_2
XFILLER_13_153 vpwr vgnd scs8hd_fill_2
XFILLER_9_168 vpwr vgnd scs8hd_fill_2
XFILLER_3_76 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _179_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_245 vgnd vpwr scs8hd_decap_12
X_150_ _121_/A _150_/B _150_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_145 vpwr vgnd scs8hd_fill_2
XFILLER_10_167 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_081_ address[3] address[4] _115_/C _082_/A vgnd vpwr scs8hd_or3_4
XFILLER_5_160 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A top_left_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _174_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_259 vpwr vgnd scs8hd_fill_2
XFILLER_23_62 vgnd vpwr scs8hd_decap_4
X_133_ _123_/A _134_/B _133_/Y vgnd vpwr scs8hd_nor2_4
X_202_ _202_/A chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_2_141 vgnd vpwr scs8hd_decap_12
XANTENNA__110__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_22 vgnd vpwr scs8hd_decap_8
XFILLER_17_7 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_55 vgnd vpwr scs8hd_decap_6
XFILLER_9_53 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_83 vgnd vpwr scs8hd_decap_8
XFILLER_11_273 vgnd vpwr scs8hd_decap_4
X_116_ _115_/X _170_/C vgnd vpwr scs8hd_buf_1
XANTENNA__105__A _105_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_17 vpwr vgnd scs8hd_fill_2
XFILLER_35_118 vpwr vgnd scs8hd_fill_2
XFILLER_29_50 vpwr vgnd scs8hd_fill_2
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XFILLER_6_76 vpwr vgnd scs8hd_fill_2
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_top_track_8.LATCH_0_.latch data_in mem_top_track_8.LATCH_0_.latch/Q _113_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_25_162 vgnd vpwr scs8hd_fill_1
XFILLER_31_73 vpwr vgnd scs8hd_fill_2
XFILLER_31_40 vpwr vgnd scs8hd_fill_2
XFILLER_16_184 vgnd vpwr scs8hd_decap_8
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_243 vgnd vpwr scs8hd_fill_1
XFILLER_39_221 vpwr vgnd scs8hd_fill_2
XFILLER_22_154 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _176_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_84 vgnd vpwr scs8hd_decap_3
XFILLER_9_147 vpwr vgnd scs8hd_fill_2
XFILLER_13_132 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A _124_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_257 vgnd vpwr scs8hd_decap_12
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_10_135 vgnd vpwr scs8hd_fill_1
X_080_ enable _115_/C vgnd vpwr scs8hd_inv_8
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_7_.scs8hd_inv_1 bottom_left_grid_pin_15_ mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_86 vgnd vpwr scs8hd_decap_6
XFILLER_37_50 vpwr vgnd scs8hd_fill_2
XFILLER_18_224 vpwr vgnd scs8hd_fill_2
XFILLER_18_235 vgnd vpwr scs8hd_decap_12
XANTENNA__108__A _085_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_24_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_205 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_5_.latch data_in mem_top_track_0.LATCH_5_.latch/Q _085_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_132_ _122_/A _134_/B _132_/Y vgnd vpwr scs8hd_nor2_4
X_201_ _201_/A chanx_right_out[7] vgnd vpwr scs8hd_buf_2
Xmem_bottom_track_9.LATCH_2_.latch data_in mem_bottom_track_9.LATCH_2_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__110__B _110_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_67 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _175_/A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _174_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__211__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_85 vgnd vpwr scs8hd_decap_6
XFILLER_34_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_11_241 vgnd vpwr scs8hd_decap_3
XFILLER_7_245 vgnd vpwr scs8hd_decap_8
X_115_ address[3] _114_/Y _115_/C _115_/X vgnd vpwr scs8hd_or3_4
XANTENNA__121__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_138 vpwr vgnd scs8hd_fill_2
XFILLER_37_182 vgnd vpwr scs8hd_fill_1
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_4_259 vgnd vpwr scs8hd_decap_12
XFILLER_20_97 vgnd vpwr scs8hd_decap_3
XFILLER_29_73 vpwr vgnd scs8hd_fill_2
XANTENNA__116__A _115_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_88 vgnd vpwr scs8hd_decap_4
Xmem_top_track_16.LATCH_2_.latch data_in mem_top_track_16.LATCH_2_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_163 vpwr vgnd scs8hd_fill_2
XFILLER_19_171 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _196_/HI _183_/Y mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_40_188 vgnd vpwr scs8hd_decap_12
XFILLER_40_100 vpwr vgnd scs8hd_fill_2
XFILLER_25_174 vpwr vgnd scs8hd_fill_2
XFILLER_15_97 vpwr vgnd scs8hd_fill_2
XFILLER_0_240 vpwr vgnd scs8hd_fill_2
XFILLER_31_111 vpwr vgnd scs8hd_fill_2
XFILLER_31_100 vpwr vgnd scs8hd_fill_2
XFILLER_16_141 vgnd vpwr scs8hd_decap_3
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _189_/HI vgnd vpwr
+ scs8hd_diode_2
.ends

