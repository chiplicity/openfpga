* NGSPICE file created from grid_clb.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_dfbbp_1 abstract view
.subckt scs8hd_dfbbp_1 CLK D Q QN RESETB SETB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

.subckt grid_clb address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] address[7] address[8] address[9] bottom_width_0_height_0__pin_10_ bottom_width_0_height_0__pin_14_
+ bottom_width_0_height_0__pin_2_ bottom_width_0_height_0__pin_6_ clk data_in enable
+ left_width_0_height_0__pin_11_ left_width_0_height_0__pin_3_ left_width_0_height_0__pin_7_
+ reset right_width_0_height_0__pin_13_ right_width_0_height_0__pin_1_ right_width_0_height_0__pin_5_
+ right_width_0_height_0__pin_9_ set top_width_0_height_0__pin_0_ top_width_0_height_0__pin_12_
+ top_width_0_height_0__pin_4_ top_width_0_height_0__pin_8_ vpwr vgnd
XFILLER_79_391 vgnd vpwr scs8hd_decap_12
XFILLER_39_277 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_54_247 vpwr vgnd scs8hd_fill_2
XFILLER_35_461 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ _140_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_166 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_15 vgnd vpwr scs8hd_decap_12
XANTENNA__203__B _231_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_77_306 vgnd vpwr scs8hd_decap_12
XFILLER_77_59 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch_SLEEPB _354_/Y vgnd vpwr scs8hd_diode_2
XFILLER_73_501 vgnd vpwr scs8hd_decap_12
XFILLER_45_236 vpwr vgnd scs8hd_fill_2
XFILLER_33_409 vpwr vgnd scs8hd_fill_2
XFILLER_60_228 vgnd vpwr scs8hd_decap_4
XFILLER_60_206 vgnd vpwr scs8hd_decap_8
X_432_ _432_/HI _432_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _148_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_115 vgnd vpwr scs8hd_fill_1
X_363_ address[4] _362_/X _367_/B vgnd vpwr scs8hd_or2_4
X_294_ _276_/A _295_/B _294_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_486 vpwr vgnd scs8hd_fill_2
XFILLER_5_398 vpwr vgnd scs8hd_fill_2
XFILLER_5_387 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_328 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_361 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_247 vgnd vpwr scs8hd_decap_6
XFILLER_51_217 vpwr vgnd scs8hd_fill_2
XFILLER_17_461 vgnd vpwr scs8hd_decap_12
XFILLER_44_280 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__304__A _231_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch/Q ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_59_317 vgnd vpwr scs8hd_fill_1
XFILLER_55_501 vgnd vpwr scs8hd_decap_12
XFILLER_67_372 vpwr vgnd scs8hd_fill_2
XFILLER_27_225 vgnd vpwr scs8hd_decap_4
XFILLER_82_342 vgnd vpwr scs8hd_decap_12
XFILLER_27_258 vgnd vpwr scs8hd_decap_4
XFILLER_70_515 vgnd vpwr scs8hd_fill_1
XFILLER_63_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_82_397 vgnd vpwr scs8hd_decap_6
XFILLER_23_431 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ _147_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_50_261 vgnd vpwr scs8hd_decap_4
XFILLER_10_158 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XFILLER_10_169 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__214__A _178_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_346 vpwr vgnd scs8hd_fill_2
XFILLER_77_147 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ _379_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XFILLER_73_342 vgnd vpwr scs8hd_decap_12
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_14_431 vgnd vpwr scs8hd_decap_12
XFILLER_33_239 vgnd vpwr scs8hd_decap_3
X_415_ _371_/A _416_/B _415_/Y vgnd vpwr scs8hd_nor2_4
X_346_ _274_/A _352_/B _346_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_283 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _434_/HI ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_277_ _231_/A _280_/B _277_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__124__A address[0] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_195 vpwr vgnd scs8hd_fill_2
XFILLER_78_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_501 vgnd vpwr scs8hd_decap_12
XFILLER_64_331 vgnd vpwr scs8hd_decap_3
XFILLER_64_386 vpwr vgnd scs8hd_fill_2
XFILLER_52_515 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
+ _400_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_20_456 vpwr vgnd scs8hd_fill_2
XFILLER_74_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_74_27 vgnd vpwr scs8hd_decap_4
XFILLER_67_191 vpwr vgnd scs8hd_fill_2
XFILLER_55_342 vpwr vgnd scs8hd_fill_2
XFILLER_70_301 vpwr vgnd scs8hd_fill_2
XFILLER_55_386 vgnd vpwr scs8hd_decap_6
XFILLER_70_323 vgnd vpwr scs8hd_decap_12
XPHY_702 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_55_397 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch_SLEEPB _334_/Y vgnd vpwr scs8hd_diode_2
XPHY_735 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_724 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_713 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__209__A address[3] vgnd vpwr scs8hd_diode_2
XPHY_768 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_757 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_746 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_389 vgnd vpwr scs8hd_fill_1
XFILLER_11_412 vgnd vpwr scs8hd_decap_12
X_200_ _202_/A _200_/B _200_/Y vgnd vpwr scs8hd_nor2_4
XPHY_779 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_131_ _131_/A _131_/Y vgnd vpwr scs8hd_inv_8
XFILLER_11_489 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q
+ _350_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_143 vpwr vgnd scs8hd_fill_2
XFILLER_2_154 vgnd vpwr scs8hd_decap_8
XFILLER_78_434 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_501 vgnd vpwr scs8hd_decap_12
XFILLER_61_301 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q
+ _315_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_64_93 vgnd vpwr scs8hd_decap_12
XFILLER_61_367 vgnd vpwr scs8hd_decap_4
XFILLER_61_389 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_261 vpwr vgnd scs8hd_fill_2
XFILLER_9_88 vpwr vgnd scs8hd_fill_2
X_329_ _247_/A _326_/X _329_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_471 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q
+ _280_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_50_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__301__B _304_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_309 vpwr vgnd scs8hd_fill_2
XFILLER_69_489 vgnd vpwr scs8hd_decap_12
XFILLER_37_320 vgnd vpwr scs8hd_decap_8
XFILLER_49_191 vpwr vgnd scs8hd_fill_2
XFILLER_64_161 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_64_194 vpwr vgnd scs8hd_fill_2
XFILLER_52_323 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_345 vgnd vpwr scs8hd_fill_1
XFILLER_20_264 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch_SLEEPB _307_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__211__B _166_/X vgnd vpwr scs8hd_diode_2
XFILLER_75_415 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2/Z
+ _158_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_47_117 vgnd vpwr scs8hd_fill_1
XFILLER_28_331 vgnd vpwr scs8hd_decap_4
XFILLER_47_139 vgnd vpwr scs8hd_decap_3
XFILLER_16_515 vgnd vpwr scs8hd_fill_1
XFILLER_43_301 vpwr vgnd scs8hd_fill_2
XFILLER_18_97 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch/Q
+ _329_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_510 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/Y _151_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_521 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_378 vpwr vgnd scs8hd_fill_2
XPHY_532 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_543 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_587 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_576 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_231 vpwr vgnd scs8hd_fill_2
XPHY_554 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_565 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_598 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_297 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _144_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_452 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch/Q
+ _294_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__402__A _380_/A vgnd vpwr scs8hd_diode_2
XFILLER_66_459 vgnd vpwr scs8hd_decap_12
XFILLER_66_448 vgnd vpwr scs8hd_fill_1
XFILLER_19_353 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q
+ _259_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_507 vgnd vpwr scs8hd_decap_8
XFILLER_61_175 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q
+ _223_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__312__A _276_/A vgnd vpwr scs8hd_diode_2
XFILLER_69_242 vpwr vgnd scs8hd_fill_2
XFILLER_69_264 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_65_470 vgnd vpwr scs8hd_decap_12
XFILLER_25_301 vgnd vpwr scs8hd_decap_4
XFILLER_37_172 vpwr vgnd scs8hd_fill_2
XFILLER_25_367 vpwr vgnd scs8hd_fill_2
XFILLER_80_495 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch_SLEEPB _280_/Y vgnd vpwr scs8hd_diode_2
XFILLER_52_186 vpwr vgnd scs8hd_fill_2
XFILLER_52_175 vpwr vgnd scs8hd_fill_2
XFILLER_40_326 vgnd vpwr scs8hd_decap_6
XFILLER_71_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__206__B _377_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_238 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
XANTENNA__222__A _231_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_466 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ _405_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_75_245 vgnd vpwr scs8hd_decap_12
XFILLER_29_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
+ _197_/Y vgnd vpwr scs8hd_diode_2
XFILLER_56_481 vgnd vpwr scs8hd_decap_12
XFILLER_56_470 vgnd vpwr scs8hd_decap_8
XFILLER_71_440 vgnd vpwr scs8hd_decap_12
XFILLER_16_334 vpwr vgnd scs8hd_fill_2
XFILLER_16_356 vgnd vpwr scs8hd_decap_6
XFILLER_45_51 vgnd vpwr scs8hd_decap_8
XFILLER_45_62 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _154_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_389 vgnd vpwr scs8hd_decap_8
XPHY_340 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_351 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_337 vgnd vpwr scs8hd_fill_1
XPHY_362 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_373 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_384 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_395 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_94 vgnd vpwr scs8hd_decap_3
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XFILLER_3_260 vpwr vgnd scs8hd_fill_2
XANTENNA__132__A _132_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_66_201 vgnd vpwr scs8hd_decap_8
XFILLER_39_404 vpwr vgnd scs8hd_fill_2
XFILLER_66_223 vgnd vpwr scs8hd_fill_1
XFILLER_66_212 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_267 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _147_/Y vgnd vpwr scs8hd_diode_2
XFILLER_66_289 vgnd vpwr scs8hd_decap_8
XFILLER_34_131 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_304 vpwr vgnd scs8hd_fill_2
XFILLER_34_175 vpwr vgnd scs8hd_fill_2
XFILLER_62_495 vgnd vpwr scs8hd_decap_12
XFILLER_22_348 vgnd vpwr scs8hd_decap_8
XFILLER_34_186 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__307__A _280_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch_SLEEPB _252_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _140_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_57_245 vgnd vpwr scs8hd_decap_3
XFILLER_72_204 vgnd vpwr scs8hd_decap_8
XFILLER_57_267 vpwr vgnd scs8hd_fill_2
XFILLER_72_215 vgnd vpwr scs8hd_decap_6
XFILLER_82_27 vgnd vpwr scs8hd_decap_4
XFILLER_25_175 vpwr vgnd scs8hd_fill_2
XFILLER_25_197 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__217__A address[8] vgnd vpwr scs8hd_diode_2
XFILLER_15_98 vpwr vgnd scs8hd_fill_2
XFILLER_31_86 vgnd vpwr scs8hd_decap_8
XFILLER_31_97 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_267 vgnd vpwr scs8hd_decap_8
XFILLER_63_226 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch_SLEEPB _351_/Y vgnd vpwr scs8hd_diode_2
XFILLER_63_248 vpwr vgnd scs8hd_fill_2
XFILLER_31_101 vpwr vgnd scs8hd_fill_2
XFILLER_44_462 vgnd vpwr scs8hd_decap_3
XFILLER_44_473 vgnd vpwr scs8hd_decap_12
XFILLER_72_93 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_145 vgnd vpwr scs8hd_decap_8
XANTENNA__127__A enable vgnd vpwr scs8hd_diode_2
XFILLER_12_370 vgnd vpwr scs8hd_decap_4
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _134_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_201 vpwr vgnd scs8hd_fill_2
XFILLER_39_212 vpwr vgnd scs8hd_fill_2
XFILLER_54_215 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_54_237 vgnd vpwr scs8hd_decap_4
XFILLER_35_440 vgnd vpwr scs8hd_decap_4
XFILLER_62_281 vpwr vgnd scs8hd_fill_2
XFILLER_50_432 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_27 vgnd vpwr scs8hd_decap_12
XFILLER_77_318 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_513 vgnd vpwr scs8hd_decap_3
X_431_ _431_/HI _431_/LO vgnd vpwr scs8hd_conb_1
XFILLER_26_451 vgnd vpwr scs8hd_decap_4
XFILLER_13_112 vgnd vpwr scs8hd_decap_4
XFILLER_13_123 vgnd vpwr scs8hd_decap_4
X_362_ _263_/A address[7] _163_/X _272_/D _362_/X vgnd vpwr scs8hd_or4_4
XFILLER_13_167 vpwr vgnd scs8hd_fill_2
XFILLER_9_138 vpwr vgnd scs8hd_fill_2
X_293_ _247_/A _295_/B _293_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_300 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch_SLEEPB _324_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_377 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _158_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__410__A _176_/B vgnd vpwr scs8hd_diode_2
XFILLER_76_373 vgnd vpwr scs8hd_decap_12
XFILLER_36_204 vgnd vpwr scs8hd_decap_8
XFILLER_36_215 vpwr vgnd scs8hd_fill_2
XFILLER_36_226 vgnd vpwr scs8hd_decap_8
XFILLER_51_207 vgnd vpwr scs8hd_decap_4
XFILLER_17_473 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_80_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_160 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__304__B _304_/B vgnd vpwr scs8hd_diode_2
XFILLER_59_329 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__320__A _247_/A vgnd vpwr scs8hd_diode_2
XFILLER_55_513 vgnd vpwr scs8hd_decap_3
XFILLER_82_354 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_50_240 vgnd vpwr scs8hd_decap_8
XFILLER_50_284 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__214__B _214_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__230__A _276_/A vgnd vpwr scs8hd_diode_2
XFILLER_77_159 vgnd vpwr scs8hd_decap_12
XFILLER_18_215 vpwr vgnd scs8hd_fill_2
XFILLER_46_502 vgnd vpwr scs8hd_decap_12
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
XFILLER_73_354 vgnd vpwr scs8hd_decap_12
X_414_ _189_/B _416_/B _414_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_53_62 vgnd vpwr scs8hd_decap_12
XFILLER_53_51 vgnd vpwr scs8hd_decap_8
XFILLER_14_443 vgnd vpwr scs8hd_decap_12
XFILLER_41_240 vpwr vgnd scs8hd_fill_2
X_345_ _273_/A _352_/B _345_/Y vgnd vpwr scs8hd_nor2_4
X_276_ _276_/A _280_/B _276_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_295 vpwr vgnd scs8hd_fill_2
XANTENNA__405__A _178_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__140__A _140_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ _156_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_148 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ _214_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_513 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_395 vgnd vpwr scs8hd_decap_3
XFILLER_64_365 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_398 vgnd vpwr scs8hd_decap_6
XFILLER_17_281 vpwr vgnd scs8hd_fill_2
XFILLER_20_424 vgnd vpwr scs8hd_decap_12
XANTENNA__315__A _279_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
+ _383_/Y vgnd vpwr scs8hd_diode_2
XFILLER_59_159 vpwr vgnd scs8hd_fill_2
XFILLER_74_129 vgnd vpwr scs8hd_decap_12
XFILLER_55_310 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_321 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ _155_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_376 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_207 vgnd vpwr scs8hd_decap_4
XFILLER_70_335 vgnd vpwr scs8hd_fill_1
XPHY_736 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_725 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_714 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_703 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__209__B _280_/A vgnd vpwr scs8hd_diode_2
XPHY_769 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_758 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_747 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_424 vgnd vpwr scs8hd_decap_3
XFILLER_23_262 vpwr vgnd scs8hd_fill_2
XFILLER_7_406 vgnd vpwr scs8hd_decap_12
X_130_ address[7] _272_/B vgnd vpwr scs8hd_inv_8
XANTENNA__225__A _280_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_428 vgnd vpwr scs8hd_decap_12
XFILLER_78_446 vgnd vpwr scs8hd_decap_12
XFILLER_65_118 vpwr vgnd scs8hd_fill_2
XFILLER_19_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_310 vgnd vpwr scs8hd_decap_4
XFILLER_73_184 vgnd vpwr scs8hd_decap_12
XFILLER_61_313 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_78 vgnd vpwr scs8hd_fill_1
XFILLER_80_93 vgnd vpwr scs8hd_decap_12
XANTENNA__135__A _135_/A vgnd vpwr scs8hd_diode_2
X_328_ _274_/A _326_/X _328_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_259_ _231_/A _262_/B _259_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_483 vgnd vpwr scs8hd_decap_12
XFILLER_43_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_310 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_151 vpwr vgnd scs8hd_fill_2
XFILLER_37_365 vgnd vpwr scs8hd_fill_1
XFILLER_52_335 vgnd vpwr scs8hd_fill_1
XFILLER_52_313 vgnd vpwr scs8hd_fill_1
XFILLER_37_398 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_243 vgnd vpwr scs8hd_decap_4
XFILLER_20_287 vpwr vgnd scs8hd_fill_2
XFILLER_69_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/Y _142_/A vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
+ _170_/Y vgnd vpwr scs8hd_diode_2
XFILLER_55_140 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_28_398 vgnd vpwr scs8hd_fill_1
XFILLER_43_313 vpwr vgnd scs8hd_fill_2
XFILLER_70_154 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_500 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_187 vgnd vpwr scs8hd_decap_8
XFILLER_70_176 vgnd vpwr scs8hd_decap_8
XPHY_511 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_522 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_533 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_544 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_390 vpwr vgnd scs8hd_fill_2
XPHY_577 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ _151_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_555 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_566 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_599 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_588 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_276 vgnd vpwr scs8hd_decap_3
XFILLER_7_236 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _139_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _436_/HI ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__402__B _384_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_464 vgnd vpwr scs8hd_decap_12
XFILLER_78_276 vgnd vpwr scs8hd_decap_12
XFILLER_19_321 vpwr vgnd scs8hd_fill_2
XFILLER_74_471 vgnd vpwr scs8hd_decap_12
XFILLER_6_280 vpwr vgnd scs8hd_fill_2
XFILLER_69_210 vgnd vpwr scs8hd_decap_3
XANTENNA__312__B _314_/B vgnd vpwr scs8hd_diode_2
XFILLER_69_232 vpwr vgnd scs8hd_fill_2
XFILLER_69_276 vpwr vgnd scs8hd_fill_2
XFILLER_29_107 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_482 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_37_184 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_206 vpwr vgnd scs8hd_fill_2
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch_SLEEPB _255_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__222__B _225_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_478 vgnd vpwr scs8hd_decap_12
XFILLER_29_86 vpwr vgnd scs8hd_fill_2
XFILLER_75_257 vgnd vpwr scs8hd_decap_12
XFILLER_56_493 vgnd vpwr scs8hd_decap_12
XFILLER_28_151 vpwr vgnd scs8hd_fill_2
XFILLER_71_452 vgnd vpwr scs8hd_decap_12
XFILLER_43_110 vgnd vpwr scs8hd_decap_3
XFILLER_45_74 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/Y _160_/A vgnd vpwr scs8hd_inv_1
XPHY_330 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_341 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_352 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_327 vpwr vgnd scs8hd_fill_2
XFILLER_43_198 vpwr vgnd scs8hd_fill_2
XFILLER_61_51 vgnd vpwr scs8hd_decap_8
XPHY_363 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_374 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_385 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_62 vgnd vpwr scs8hd_decap_12
XPHY_396 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ _131_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
XANTENNA__413__A _391_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch/Q ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_438 vpwr vgnd scs8hd_fill_2
XFILLER_19_140 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_471 vpwr vgnd scs8hd_fill_2
XFILLER_19_184 vpwr vgnd scs8hd_fill_2
XFILLER_22_316 vgnd vpwr scs8hd_fill_1
XFILLER_34_154 vpwr vgnd scs8hd_fill_2
XFILLER_34_165 vgnd vpwr scs8hd_decap_8
XANTENNA__307__B _304_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_393 vgnd vpwr scs8hd_decap_4
XANTENNA__323__A _287_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_235 vpwr vgnd scs8hd_fill_2
XFILLER_57_224 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_471 vgnd vpwr scs8hd_decap_12
XFILLER_45_419 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch_SLEEPB _227_/Y vgnd vpwr scs8hd_diode_2
XFILLER_53_474 vgnd vpwr scs8hd_decap_3
XANTENNA__217__B _235_/B vgnd vpwr scs8hd_diode_2
XFILLER_40_146 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _433_/HI ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ _197_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
+ _392_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__233__A _279_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_231 vgnd vpwr scs8hd_decap_12
XFILLER_0_275 vpwr vgnd scs8hd_fill_2
XFILLER_48_202 vgnd vpwr scs8hd_fill_1
XFILLER_48_246 vgnd vpwr scs8hd_decap_8
XFILLER_36_419 vpwr vgnd scs8hd_fill_2
XFILLER_63_238 vgnd vpwr scs8hd_decap_4
XFILLER_56_290 vgnd vpwr scs8hd_decap_3
XFILLER_16_110 vgnd vpwr scs8hd_decap_12
XFILLER_16_154 vgnd vpwr scs8hd_decap_6
XFILLER_71_271 vgnd vpwr scs8hd_decap_6
XANTENNA__408__A _170_/B vgnd vpwr scs8hd_diode_2
XFILLER_44_485 vgnd vpwr scs8hd_decap_12
XPHY_160 vgnd vpwr scs8hd_decap_3
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_179 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__143__A _143_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_235 vpwr vgnd scs8hd_fill_2
XFILLER_27_419 vpwr vgnd scs8hd_fill_2
XFILLER_35_474 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__318__A _273_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_455 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
+ _405_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_146 vgnd vpwr scs8hd_fill_1
XFILLER_10_319 vpwr vgnd scs8hd_fill_2
XFILLER_22_179 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
+ set vgnd vpwr scs8hd_diode_2
XFILLER_2_507 vgnd vpwr scs8hd_decap_8
XFILLER_77_39 vgnd vpwr scs8hd_decap_12
XFILLER_58_511 vgnd vpwr scs8hd_decap_4
XFILLER_18_408 vpwr vgnd scs8hd_fill_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
XFILLER_26_430 vpwr vgnd scs8hd_fill_2
X_430_ _430_/HI _430_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__228__A _274_/A vgnd vpwr scs8hd_diode_2
XFILLER_53_271 vgnd vpwr scs8hd_decap_4
XFILLER_53_260 vpwr vgnd scs8hd_fill_2
X_361_ _280_/A _359_/B _361_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_146 vpwr vgnd scs8hd_fill_2
XFILLER_41_466 vpwr vgnd scs8hd_fill_2
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
X_292_ _274_/A _295_/B _292_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_5_356 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__410__B _416_/B vgnd vpwr scs8hd_diode_2
XFILLER_76_385 vgnd vpwr scs8hd_decap_12
XFILLER_17_485 vgnd vpwr scs8hd_decap_3
XFILLER_32_422 vpwr vgnd scs8hd_fill_2
XANTENNA__138__A _138_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ _142_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_44_293 vpwr vgnd scs8hd_fill_2
XFILLER_73_3 vgnd vpwr scs8hd_decap_12
XFILLER_8_183 vgnd vpwr scs8hd_fill_1
XANTENNA__320__B _325_/B vgnd vpwr scs8hd_diode_2
XFILLER_67_341 vpwr vgnd scs8hd_fill_2
XFILLER_82_311 vgnd vpwr scs8hd_decap_12
XFILLER_67_363 vgnd vpwr scs8hd_decap_3
XFILLER_82_366 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_208 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ _417_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_411 vpwr vgnd scs8hd_fill_2
XFILLER_23_422 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_260 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_455 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_127 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_56 vgnd vpwr scs8hd_decap_12
XANTENNA__230__B _231_/B vgnd vpwr scs8hd_diode_2
XFILLER_58_385 vpwr vgnd scs8hd_fill_2
XFILLER_46_514 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_249 vpwr vgnd scs8hd_fill_2
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
X_413_ _391_/A _416_/B _413_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_455 vgnd vpwr scs8hd_decap_3
XFILLER_53_74 vgnd vpwr scs8hd_decap_12
XFILLER_41_263 vpwr vgnd scs8hd_fill_2
X_344_ address[6] _272_/B _163_/X _272_/D _352_/B vgnd vpwr scs8hd_or4_4
X_275_ _247_/A _280_/B _275_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__405__B _402_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_153 vpwr vgnd scs8hd_fill_2
XFILLER_5_142 vpwr vgnd scs8hd_fill_2
XANTENNA__421__A _377_/A vgnd vpwr scs8hd_diode_2
XFILLER_78_93 vgnd vpwr scs8hd_decap_12
XFILLER_68_105 vgnd vpwr scs8hd_decap_12
XFILLER_49_363 vgnd vpwr scs8hd_fill_1
XFILLER_64_311 vgnd vpwr scs8hd_decap_3
XFILLER_17_260 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
+ _409_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_436 vgnd vpwr scs8hd_decap_12
XFILLER_32_285 vgnd vpwr scs8hd_decap_3
XFILLER_32_296 vpwr vgnd scs8hd_fill_2
XANTENNA__315__B _314_/B vgnd vpwr scs8hd_diode_2
XANTENNA__331__A _231_/A vgnd vpwr scs8hd_diode_2
XFILLER_59_127 vpwr vgnd scs8hd_fill_2
XFILLER_59_116 vgnd vpwr scs8hd_decap_4
XFILLER_59_138 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_503 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _131_/Y vgnd vpwr scs8hd_diode_2
XPHY_726 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_715 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_704 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_759 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_748 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_737 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_418 vgnd vpwr scs8hd_decap_8
XFILLER_23_88 vpwr vgnd scs8hd_fill_2
XANTENNA__225__B _225_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__241__A _287_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_73_196 vgnd vpwr scs8hd_decap_12
XANTENNA__416__A _194_/B vgnd vpwr scs8hd_diode_2
X_327_ _273_/A _326_/X _327_/Y vgnd vpwr scs8hd_nor2_4
X_258_ _276_/A _262_/B _258_/Y vgnd vpwr scs8hd_nor2_4
X_189_ _202_/A _189_/B _189_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_495 vgnd vpwr scs8hd_decap_12
XANTENNA__151__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_69_425 vpwr vgnd scs8hd_fill_2
XFILLER_69_403 vgnd vpwr scs8hd_fill_1
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ _395_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
+ _421_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_344 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_200 vgnd vpwr scs8hd_decap_8
XFILLER_20_211 vgnd vpwr scs8hd_decap_3
XANTENNA__326__A _263_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_75_428 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
XFILLER_28_377 vgnd vpwr scs8hd_decap_8
XFILLER_28_388 vpwr vgnd scs8hd_fill_2
XPHY_501 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_512 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_523 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_534 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__236__A _273_/A vgnd vpwr scs8hd_diode_2
XPHY_578 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_211 vgnd vpwr scs8hd_fill_1
XPHY_545 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_556 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_567 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_589 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_204 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_226 vgnd vpwr scs8hd_decap_3
XFILLER_3_410 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_59_62 vgnd vpwr scs8hd_decap_12
XFILLER_59_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_476 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_66_428 vgnd vpwr scs8hd_decap_3
XFILLER_78_288 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _149_/Y vgnd vpwr scs8hd_diode_2
XFILLER_74_483 vgnd vpwr scs8hd_decap_12
XFILLER_34_303 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_163 vgnd vpwr scs8hd_decap_8
XFILLER_34_369 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__146__A _146_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_439 vpwr vgnd scs8hd_fill_2
XFILLER_57_428 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
+ _427_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_25_347 vpwr vgnd scs8hd_fill_2
XFILLER_25_358 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _140_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_435 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_48_439 vpwr vgnd scs8hd_fill_2
XFILLER_75_269 vgnd vpwr scs8hd_decap_12
XFILLER_28_163 vgnd vpwr scs8hd_decap_3
XFILLER_71_464 vgnd vpwr scs8hd_decap_12
XFILLER_31_306 vgnd vpwr scs8hd_decap_4
XFILLER_43_144 vpwr vgnd scs8hd_fill_2
XFILLER_45_86 vgnd vpwr scs8hd_decap_4
XPHY_320 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_331 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_342 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_188 vgnd vpwr scs8hd_fill_1
XPHY_353 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_364 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ _132_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_375 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_386 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_61_74 vgnd vpwr scs8hd_decap_12
XPHY_397 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch_SLEEPB _224_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ _373_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__413__B _416_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_295 vgnd vpwr scs8hd_decap_4
XFILLER_39_417 vgnd vpwr scs8hd_decap_8
XFILLER_39_428 vgnd vpwr scs8hd_decap_3
XFILLER_54_409 vpwr vgnd scs8hd_fill_2
XFILLER_47_461 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_111 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_328 vgnd vpwr scs8hd_decap_8
XFILLER_30_361 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__323__B _325_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ _391_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_483 vgnd vpwr scs8hd_decap_12
XFILLER_65_291 vpwr vgnd scs8hd_fill_2
XFILLER_53_442 vgnd vpwr scs8hd_decap_4
XFILLER_53_431 vpwr vgnd scs8hd_fill_2
XFILLER_53_453 vpwr vgnd scs8hd_fill_2
XFILLER_13_306 vpwr vgnd scs8hd_fill_2
XFILLER_25_144 vgnd vpwr scs8hd_decap_4
XFILLER_40_103 vpwr vgnd scs8hd_fill_2
XFILLER_40_125 vgnd vpwr scs8hd_decap_3
XANTENNA__217__C _215_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_361 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__233__B _231_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_243 vgnd vpwr scs8hd_decap_4
XFILLER_63_206 vpwr vgnd scs8hd_fill_2
XFILLER_16_133 vgnd vpwr scs8hd_decap_4
XFILLER_16_144 vgnd vpwr scs8hd_decap_6
XANTENNA__408__B _416_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_114 vgnd vpwr scs8hd_decap_6
XFILLER_44_497 vgnd vpwr scs8hd_decap_12
XPHY_161 vgnd vpwr scs8hd_decap_3
XPHY_150 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ _139_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_31_158 vpwr vgnd scs8hd_fill_2
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_12_383 vpwr vgnd scs8hd_fill_2
XANTENNA__424__A _380_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_387 vpwr vgnd scs8hd_fill_2
XFILLER_8_376 vgnd vpwr scs8hd_decap_4
XFILLER_8_365 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch/Q
+ _309_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_67_501 vgnd vpwr scs8hd_decap_12
XFILLER_39_258 vgnd vpwr scs8hd_decap_12
XFILLER_82_515 vgnd vpwr scs8hd_fill_1
XFILLER_54_206 vpwr vgnd scs8hd_fill_2
XFILLER_35_431 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch/Q
+ _274_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch_SLEEPB _296_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_125 vgnd vpwr scs8hd_decap_6
XANTENNA__318__B _325_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_486 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__334__A _280_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_90 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch/Q
+ _238_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_44 vgnd vpwr scs8hd_decap_12
XANTENNA__228__B _231_/B vgnd vpwr scs8hd_diode_2
X_360_ _279_/A _359_/B _360_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_107 vpwr vgnd scs8hd_fill_2
XFILLER_41_456 vgnd vpwr scs8hd_decap_4
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
X_291_ _273_/A _295_/B _291_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_489 vgnd vpwr scs8hd_decap_12
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XANTENNA__244__A address[8] vgnd vpwr scs8hd_diode_2
XFILLER_5_335 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
+ _388_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XFILLER_67_51 vgnd vpwr scs8hd_decap_8
XFILLER_49_501 vgnd vpwr scs8hd_decap_12
XFILLER_3_59 vpwr vgnd scs8hd_fill_2
XFILLER_67_62 vgnd vpwr scs8hd_decap_12
XFILLER_64_515 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__419__A _202_/B vgnd vpwr scs8hd_diode_2
XFILLER_44_250 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_191 vpwr vgnd scs8hd_fill_2
XFILLER_8_151 vpwr vgnd scs8hd_fill_2
XANTENNA__154__A _154_/A vgnd vpwr scs8hd_diode_2
XFILLER_66_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _135_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_309 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch_SLEEPB _269_/Y vgnd vpwr scs8hd_diode_2
XFILLER_82_323 vgnd vpwr scs8hd_decap_12
XFILLER_70_507 vgnd vpwr scs8hd_decap_8
XANTENNA__329__A _247_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_489 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_305 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_206 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_367 vgnd vpwr scs8hd_decap_12
XANTENNA__239__A _276_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_412_ _183_/B _416_/B _412_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_250 vpwr vgnd scs8hd_fill_2
X_343_ _280_/A _343_/B _343_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_53_86 vgnd vpwr scs8hd_decap_12
X_274_ _274_/A _280_/B _274_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_176 vgnd vpwr scs8hd_decap_4
XANTENNA__421__B _416_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_68_117 vgnd vpwr scs8hd_decap_4
XFILLER_1_371 vgnd vpwr scs8hd_fill_1
XFILLER_49_353 vgnd vpwr scs8hd_decap_4
XANTENNA__149__A _149_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_294 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch_SLEEPB _241_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_253 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_448 vgnd vpwr scs8hd_decap_8
XFILLER_20_459 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
+ _214_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__331__B _326_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_55_301 vpwr vgnd scs8hd_fill_2
XFILLER_28_515 vgnd vpwr scs8hd_fill_1
XFILLER_70_337 vgnd vpwr scs8hd_decap_3
XPHY_727 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_716 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_705 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_231 vgnd vpwr scs8hd_decap_3
XPHY_749 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_738 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_404 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_297 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _141_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch_SLEEPB _340_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_113 vpwr vgnd scs8hd_fill_2
XANTENNA__241__B _243_/B vgnd vpwr scs8hd_diode_2
XFILLER_78_459 vgnd vpwr scs8hd_decap_12
XFILLER_48_97 vgnd vpwr scs8hd_decap_3
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XFILLER_46_367 vpwr vgnd scs8hd_fill_2
XFILLER_46_389 vgnd vpwr scs8hd_decap_6
XFILLER_61_337 vpwr vgnd scs8hd_fill_2
XFILLER_14_220 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__416__B _416_/B vgnd vpwr scs8hd_diode_2
X_326_ _263_/A _272_/B _163_/X _272_/D _326_/X vgnd vpwr scs8hd_or4_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_257_ _247_/A _262_/B _257_/Y vgnd vpwr scs8hd_nor2_4
X_188_ _122_/Y _279_/A _189_/B vgnd vpwr scs8hd_or2_4
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _132_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _157_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_367 vgnd vpwr scs8hd_decap_3
XFILLER_52_337 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__326__B _272_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _432_/HI ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_20_267 vgnd vpwr scs8hd_decap_6
XFILLER_9_290 vpwr vgnd scs8hd_fill_2
XANTENNA__342__A _279_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q
+ _360_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_301 vgnd vpwr scs8hd_decap_12
XFILLER_28_323 vpwr vgnd scs8hd_fill_2
XFILLER_16_507 vgnd vpwr scs8hd_decap_8
XFILLER_18_56 vgnd vpwr scs8hd_decap_12
XFILLER_55_175 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch_SLEEPB _313_/Y vgnd vpwr scs8hd_diode_2
XFILLER_70_145 vpwr vgnd scs8hd_fill_2
XFILLER_55_197 vpwr vgnd scs8hd_fill_2
XFILLER_43_337 vpwr vgnd scs8hd_fill_2
XFILLER_43_359 vgnd vpwr scs8hd_decap_4
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XPHY_502 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_513 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_524 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_535 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__236__B _243_/B vgnd vpwr scs8hd_diode_2
XPHY_546 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_557 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_568 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_579 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_245 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q
+ _325_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_50_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_249 vgnd vpwr scs8hd_decap_3
XANTENNA__252__A _280_/A vgnd vpwr scs8hd_diode_2
XFILLER_50_98 vpwr vgnd scs8hd_fill_2
XFILLER_3_422 vgnd vpwr scs8hd_decap_4
XFILLER_59_74 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/Y _148_/A vgnd vpwr scs8hd_inv_1
XFILLER_19_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_75_62 vgnd vpwr scs8hd_decap_12
XFILLER_75_51 vgnd vpwr scs8hd_decap_8
XFILLER_19_367 vpwr vgnd scs8hd_fill_2
XFILLER_19_378 vpwr vgnd scs8hd_fill_2
XFILLER_19_389 vpwr vgnd scs8hd_fill_2
XFILLER_74_495 vgnd vpwr scs8hd_decap_12
XFILLER_61_123 vgnd vpwr scs8hd_fill_1
XFILLER_34_348 vpwr vgnd scs8hd_fill_2
XFILLER_46_186 vpwr vgnd scs8hd_fill_2
XFILLER_61_156 vgnd vpwr scs8hd_decap_4
XANTENNA__427__A _178_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_510 vgnd vpwr scs8hd_decap_6
XFILLER_42_392 vpwr vgnd scs8hd_fill_2
X_309_ _273_/A _314_/B _309_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
+ _374_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_293 vgnd vpwr scs8hd_decap_6
XFILLER_69_245 vgnd vpwr scs8hd_decap_4
XFILLER_69_289 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_80_410 vgnd vpwr scs8hd_decap_12
XFILLER_37_164 vgnd vpwr scs8hd_decap_3
XFILLER_25_326 vgnd vpwr scs8hd_decap_6
XFILLER_52_145 vgnd vpwr scs8hd_decap_8
XANTENNA__337__A _274_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_370 vpwr vgnd scs8hd_fill_2
XFILLER_33_392 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch/Q
+ _339_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_219 vpwr vgnd scs8hd_fill_2
XFILLER_20_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch_SLEEPB _286_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _150_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_447 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q
+ _304_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_48_407 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_304 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_326 vgnd vpwr scs8hd_decap_8
XFILLER_28_186 vpwr vgnd scs8hd_fill_2
XFILLER_43_123 vpwr vgnd scs8hd_fill_2
XFILLER_71_476 vgnd vpwr scs8hd_decap_12
XANTENNA__247__A _247_/A vgnd vpwr scs8hd_diode_2
XPHY_310 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_321 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_332 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_343 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q
+ _269_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_354 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_365 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_376 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_86 vgnd vpwr scs8hd_decap_8
XPHY_387 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_398 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ _365_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_241 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q
+ _233_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_66_215 vgnd vpwr scs8hd_decap_8
XFILLER_19_164 vpwr vgnd scs8hd_fill_2
XFILLER_74_270 vgnd vpwr scs8hd_decap_4
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
XFILLER_34_101 vgnd vpwr scs8hd_fill_1
XFILLER_62_443 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__157__A _157_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_392 vgnd vpwr scs8hd_fill_1
XFILLER_30_340 vgnd vpwr scs8hd_decap_4
XFILLER_30_351 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_204 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
+ _367_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_451 vgnd vpwr scs8hd_decap_6
XFILLER_25_101 vpwr vgnd scs8hd_fill_2
XFILLER_25_123 vpwr vgnd scs8hd_fill_2
XFILLER_38_495 vgnd vpwr scs8hd_decap_12
XFILLER_80_251 vgnd vpwr scs8hd_decap_12
XFILLER_53_487 vgnd vpwr scs8hd_fill_1
XFILLER_13_329 vgnd vpwr scs8hd_decap_3
XFILLER_40_137 vgnd vpwr scs8hd_decap_6
XANTENNA__217__D _272_/D vgnd vpwr scs8hd_diode_2
XFILLER_21_351 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _155_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_200 vgnd vpwr scs8hd_decap_8
XFILLER_0_255 vpwr vgnd scs8hd_fill_2
XFILLER_48_215 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_97 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/Y _143_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_71_284 vpwr vgnd scs8hd_fill_2
XFILLER_16_178 vpwr vgnd scs8hd_fill_2
XPHY_151 vgnd vpwr scs8hd_decap_3
XPHY_140 vgnd vpwr scs8hd_decap_3
XFILLER_31_126 vgnd vpwr scs8hd_decap_4
XPHY_162 vgnd vpwr scs8hd_decap_3
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_395 vpwr vgnd scs8hd_fill_2
XFILLER_8_333 vgnd vpwr scs8hd_fill_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__424__B _406_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch_SLEEPB _357_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_513 vgnd vpwr scs8hd_decap_3
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__334__B _326_/X vgnd vpwr scs8hd_diode_2
XANTENNA__350__A _287_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ _148_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_56 vgnd vpwr scs8hd_decap_12
XFILLER_26_443 vgnd vpwr scs8hd_decap_6
XFILLER_53_284 vpwr vgnd scs8hd_fill_2
XFILLER_41_413 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
X_290_ _263_/A address[7] _272_/C _272_/D _295_/B vgnd vpwr scs8hd_or4_4
XFILLER_41_435 vpwr vgnd scs8hd_fill_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XANTENNA__244__B _235_/B vgnd vpwr scs8hd_diode_2
XFILLER_42_99 vpwr vgnd scs8hd_fill_2
XANTENNA__260__A _287_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
XFILLER_49_513 vgnd vpwr scs8hd_decap_3
XFILLER_67_74 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_76_398 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ _147_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__419__B _416_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_32_402 vgnd vpwr scs8hd_decap_3
XFILLER_32_435 vpwr vgnd scs8hd_fill_2
XFILLER_32_446 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_468 vgnd vpwr scs8hd_decap_8
XFILLER_32_479 vgnd vpwr scs8hd_decap_12
XFILLER_8_196 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_3 vgnd vpwr scs8hd_decap_12
XANTENNA__170__A _202_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_376 vpwr vgnd scs8hd_fill_2
XFILLER_67_354 vpwr vgnd scs8hd_fill_2
XFILLER_27_207 vgnd vpwr scs8hd_fill_1
XFILLER_82_335 vgnd vpwr scs8hd_decap_6
XANTENNA__329__B _326_/X vgnd vpwr scs8hd_diode_2
XFILLER_50_221 vpwr vgnd scs8hd_fill_2
XFILLER_23_435 vpwr vgnd scs8hd_fill_2
XFILLER_35_284 vpwr vgnd scs8hd_fill_2
XANTENNA__345__A _273_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_328 vgnd vpwr scs8hd_decap_8
XFILLER_58_365 vgnd vpwr scs8hd_decap_3
XFILLER_58_398 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__239__B _243_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_379 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _146_/Y vgnd vpwr scs8hd_diode_2
X_411_ _367_/A _416_/B _411_/Y vgnd vpwr scs8hd_nor2_4
X_342_ _279_/A _343_/B _342_/Y vgnd vpwr scs8hd_nor2_4
X_273_ _273_/A _280_/B _273_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_53_98 vgnd vpwr scs8hd_decap_3
XANTENNA__255__A _273_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_166 vgnd vpwr scs8hd_decap_4
XFILLER_5_199 vgnd vpwr scs8hd_decap_6
XFILLER_1_383 vgnd vpwr scs8hd_decap_6
XFILLER_49_321 vpwr vgnd scs8hd_fill_2
XFILLER_49_343 vgnd vpwr scs8hd_fill_1
XFILLER_49_376 vpwr vgnd scs8hd_fill_2
XFILLER_17_240 vpwr vgnd scs8hd_fill_2
XFILLER_32_210 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A _127_/Y vgnd vpwr scs8hd_diode_2
XFILLER_67_184 vgnd vpwr scs8hd_decap_4
XFILLER_55_357 vpwr vgnd scs8hd_fill_2
XFILLER_82_187 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_70_349 vgnd vpwr scs8hd_decap_8
XPHY_717 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_706 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_739 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_728 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_254 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_147 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_48_32 vgnd vpwr scs8hd_decap_12
XFILLER_73_110 vgnd vpwr scs8hd_decap_12
XFILLER_34_508 vgnd vpwr scs8hd_decap_8
XFILLER_46_346 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_379 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_210 vgnd vpwr scs8hd_decap_4
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_265 vgnd vpwr scs8hd_decap_8
XFILLER_9_59 vpwr vgnd scs8hd_fill_2
XFILLER_14_276 vpwr vgnd scs8hd_fill_2
X_325_ _280_/A _325_/B _325_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ _411_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_471 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
+ clk vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q
+ _334_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_256_ _274_/A _262_/B _256_/Y vgnd vpwr scs8hd_nor2_4
X_187_ address[2] _187_/B _279_/A vgnd vpwr scs8hd_or2_4
XFILLER_49_140 vgnd vpwr scs8hd_decap_6
XFILLER_37_302 vgnd vpwr scs8hd_fill_1
XFILLER_49_151 vpwr vgnd scs8hd_fill_2
XFILLER_49_195 vpwr vgnd scs8hd_fill_2
XFILLER_64_165 vgnd vpwr scs8hd_decap_3
XFILLER_37_379 vgnd vpwr scs8hd_decap_3
XFILLER_64_198 vpwr vgnd scs8hd_fill_2
XFILLER_52_327 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_224 vgnd vpwr scs8hd_decap_8
XFILLER_60_393 vpwr vgnd scs8hd_fill_2
XANTENNA__326__C _163_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__342__B _343_/B vgnd vpwr scs8hd_diode_2
XFILLER_68_471 vgnd vpwr scs8hd_decap_12
XFILLER_28_313 vgnd vpwr scs8hd_fill_1
XFILLER_55_132 vpwr vgnd scs8hd_fill_2
XFILLER_18_68 vgnd vpwr scs8hd_decap_12
XFILLER_28_335 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_503 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_514 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_525 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_382 vgnd vpwr scs8hd_decap_8
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
XPHY_536 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_547 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_558 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_569 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_235 vgnd vpwr scs8hd_decap_6
XFILLER_50_44 vgnd vpwr scs8hd_decap_12
XANTENNA__252__B _252_/B vgnd vpwr scs8hd_diode_2
XFILLER_78_202 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_86 vgnd vpwr scs8hd_decap_12
XFILLER_3_489 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_471 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_357 vgnd vpwr scs8hd_decap_6
XFILLER_46_121 vpwr vgnd scs8hd_fill_2
XFILLER_46_132 vpwr vgnd scs8hd_fill_2
XFILLER_75_74 vgnd vpwr scs8hd_decap_12
XFILLER_46_143 vgnd vpwr scs8hd_decap_8
XFILLER_61_135 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__427__B _424_/X vgnd vpwr scs8hd_diode_2
XFILLER_61_179 vgnd vpwr scs8hd_decap_4
XFILLER_42_360 vpwr vgnd scs8hd_fill_2
X_308_ address[6] address[7] _272_/C _272_/D _314_/B vgnd vpwr scs8hd_or4_4
X_239_ _276_/A _243_/B _239_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_290 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
+ _204_/Y vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_69_268 vpwr vgnd scs8hd_fill_2
XFILLER_57_408 vpwr vgnd scs8hd_fill_2
XFILLER_57_419 vpwr vgnd scs8hd_fill_2
XFILLER_65_441 vpwr vgnd scs8hd_fill_2
XFILLER_37_110 vpwr vgnd scs8hd_fill_2
XFILLER_80_422 vgnd vpwr scs8hd_decap_12
XFILLER_37_176 vpwr vgnd scs8hd_fill_2
XFILLER_52_168 vgnd vpwr scs8hd_decap_4
XFILLER_52_135 vgnd vpwr scs8hd_fill_1
XANTENNA__337__B _343_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__353__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_0_404 vgnd vpwr scs8hd_decap_12
XFILLER_0_459 vgnd vpwr scs8hd_decap_6
XFILLER_48_419 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__247__B _252_/B vgnd vpwr scs8hd_diode_2
XPHY_300 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_157 vgnd vpwr scs8hd_decap_3
XPHY_311 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_322 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_333 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _160_/Y vgnd vpwr scs8hd_diode_2
XPHY_344 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_355 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_366 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_393 vgnd vpwr scs8hd_decap_4
XPHY_377 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_515 vgnd vpwr scs8hd_fill_1
XPHY_388 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_399 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__263__A _263_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_10_80 vgnd vpwr scs8hd_fill_1
XFILLER_3_275 vpwr vgnd scs8hd_fill_2
XFILLER_3_264 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_81_208 vgnd vpwr scs8hd_decap_12
XFILLER_47_452 vgnd vpwr scs8hd_decap_3
XFILLER_62_422 vpwr vgnd scs8hd_fill_2
XFILLER_34_124 vgnd vpwr scs8hd_decap_4
XFILLER_34_135 vpwr vgnd scs8hd_fill_2
XFILLER_22_308 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_382 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__173__A _202_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__348__A _276_/A vgnd vpwr scs8hd_diode_2
XFILLER_80_263 vgnd vpwr scs8hd_decap_12
XFILLER_25_179 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2/Z
+ _134_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_341 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_56_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_289 vgnd vpwr scs8hd_decap_6
XFILLER_63_219 vgnd vpwr scs8hd_decap_4
XFILLER_29_441 vpwr vgnd scs8hd_fill_2
XFILLER_56_260 vpwr vgnd scs8hd_fill_2
XANTENNA__258__A _276_/A vgnd vpwr scs8hd_diode_2
XFILLER_71_241 vgnd vpwr scs8hd_fill_1
XPHY_152 vgnd vpwr scs8hd_decap_3
XPHY_141 vgnd vpwr scs8hd_decap_3
XPHY_130 vgnd vpwr scs8hd_decap_3
XPHY_163 vgnd vpwr scs8hd_decap_3
XFILLER_8_312 vgnd vpwr scs8hd_decap_4
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_90 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_79_330 vgnd vpwr scs8hd_decap_12
XFILLER_39_205 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_227 vpwr vgnd scs8hd_fill_2
XANTENNA__168__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_62_263 vgnd vpwr scs8hd_fill_1
XFILLER_62_285 vgnd vpwr scs8hd_decap_3
XFILLER_50_447 vgnd vpwr scs8hd_decap_8
XFILLER_22_149 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _156_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_160 vgnd vpwr scs8hd_decap_8
XFILLER_30_193 vpwr vgnd scs8hd_fill_2
XANTENNA__350__B _352_/B vgnd vpwr scs8hd_diode_2
XFILLER_45_219 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_455 vgnd vpwr scs8hd_fill_1
XFILLER_53_252 vpwr vgnd scs8hd_fill_2
XFILLER_26_68 vgnd vpwr scs8hd_decap_12
XFILLER_13_116 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_425 vpwr vgnd scs8hd_fill_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_12
XANTENNA__244__C _235_/C vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_315 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__260__B _262_/B vgnd vpwr scs8hd_diode_2
XFILLER_76_300 vgnd vpwr scs8hd_decap_12
XFILLER_3_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_67_86 vgnd vpwr scs8hd_decap_12
XFILLER_17_433 vpwr vgnd scs8hd_fill_2
XFILLER_32_414 vgnd vpwr scs8hd_decap_8
XFILLER_8_120 vgnd vpwr scs8hd_decap_3
XFILLER_40_480 vgnd vpwr scs8hd_decap_12
XFILLER_8_186 vgnd vpwr scs8hd_fill_1
XFILLER_8_164 vpwr vgnd scs8hd_fill_2
XFILLER_4_370 vgnd vpwr scs8hd_decap_8
XANTENNA__170__B _170_/B vgnd vpwr scs8hd_diode_2
XFILLER_79_171 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_399 vpwr vgnd scs8hd_fill_2
XFILLER_35_230 vgnd vpwr scs8hd_decap_4
XFILLER_50_200 vgnd vpwr scs8hd_decap_6
XFILLER_35_252 vpwr vgnd scs8hd_fill_2
XFILLER_35_274 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_50_288 vgnd vpwr scs8hd_decap_6
XANTENNA__345__B _352_/B vgnd vpwr scs8hd_diode_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ _156_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__361__A _280_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_318 vgnd vpwr scs8hd_fill_1
X_410_ _176_/B _416_/B _410_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_81_391 vgnd vpwr scs8hd_decap_12
X_341_ _287_/A _343_/B _341_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
X_272_ address[6] _272_/B _272_/C _272_/D _280_/B vgnd vpwr scs8hd_or4_4
XANTENNA__255__B _262_/B vgnd vpwr scs8hd_diode_2
XFILLER_41_299 vgnd vpwr scs8hd_decap_4
XANTENNA__271__A _280_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_123 vpwr vgnd scs8hd_fill_2
XFILLER_1_351 vpwr vgnd scs8hd_fill_2
XFILLER_1_362 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ _155_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_49_300 vgnd vpwr scs8hd_decap_3
XFILLER_76_141 vgnd vpwr scs8hd_decap_12
XFILLER_52_509 vgnd vpwr scs8hd_decap_6
XFILLER_72_380 vgnd vpwr scs8hd_decap_12
XANTENNA__165__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_9_440 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_71_3 vgnd vpwr scs8hd_decap_12
XANTENNA__181__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_6
XFILLER_55_325 vpwr vgnd scs8hd_fill_2
XFILLER_70_306 vgnd vpwr scs8hd_decap_8
XFILLER_82_199 vgnd vpwr scs8hd_decap_12
XPHY_718 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_707 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_63_380 vpwr vgnd scs8hd_fill_2
XANTENNA__356__A _247_/A vgnd vpwr scs8hd_diode_2
XPHY_729 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_428 vgnd vpwr scs8hd_decap_12
XFILLER_23_277 vpwr vgnd scs8hd_fill_2
XFILLER_23_288 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _152_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_48_44 vgnd vpwr scs8hd_decap_12
XFILLER_58_174 vgnd vpwr scs8hd_decap_8
XFILLER_58_163 vpwr vgnd scs8hd_fill_2
XFILLER_46_314 vgnd vpwr scs8hd_fill_1
XFILLER_58_185 vpwr vgnd scs8hd_fill_2
XFILLER_46_358 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_32 vgnd vpwr scs8hd_decap_12
XFILLER_61_317 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__266__A _247_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_27 vgnd vpwr scs8hd_decap_12
X_324_ _279_/A _325_/B _324_/Y vgnd vpwr scs8hd_nor2_4
X_255_ _273_/A _262_/B _255_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_483 vgnd vpwr scs8hd_decap_12
XFILLER_13_80 vpwr vgnd scs8hd_fill_2
X_186_ _202_/A _391_/A _186_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
+ _180_/Y vgnd vpwr scs8hd_diode_2
XFILLER_69_417 vgnd vpwr scs8hd_decap_8
XFILLER_69_406 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_69_428 vgnd vpwr scs8hd_decap_12
XFILLER_49_163 vgnd vpwr scs8hd_fill_1
XFILLER_64_111 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_358 vgnd vpwr scs8hd_decap_4
XFILLER_64_177 vpwr vgnd scs8hd_fill_2
XFILLER_52_306 vgnd vpwr scs8hd_decap_4
XANTENNA__176__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_60_372 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_247 vgnd vpwr scs8hd_fill_1
XANTENNA__326__D _272_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_483 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_144 vgnd vpwr scs8hd_fill_1
XFILLER_43_317 vgnd vpwr scs8hd_decap_3
XPHY_504 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_515 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_526 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_214 vpwr vgnd scs8hd_fill_2
XFILLER_11_203 vpwr vgnd scs8hd_fill_2
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XPHY_537 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_548 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_559 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_56 vgnd vpwr scs8hd_decap_12
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_66_409 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_59_98 vgnd vpwr scs8hd_decap_3
XFILLER_59_483 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_336 vpwr vgnd scs8hd_fill_2
XFILLER_75_86 vgnd vpwr scs8hd_decap_12
XFILLER_61_114 vpwr vgnd scs8hd_fill_2
XFILLER_61_103 vpwr vgnd scs8hd_fill_2
XFILLER_34_328 vgnd vpwr scs8hd_decap_8
XFILLER_46_199 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ _132_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch_SLEEPB _258_/Y vgnd vpwr scs8hd_diode_2
X_307_ _280_/A _304_/B _307_/Y vgnd vpwr scs8hd_nor2_4
X_238_ _247_/A _243_/B _238_/Y vgnd vpwr scs8hd_nor2_4
X_169_ _122_/Y _273_/A _170_/B vgnd vpwr scs8hd_or2_4
XFILLER_6_273 vpwr vgnd scs8hd_fill_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XFILLER_69_236 vgnd vpwr scs8hd_decap_4
XFILLER_65_420 vgnd vpwr scs8hd_decap_4
XFILLER_25_306 vgnd vpwr scs8hd_decap_3
XFILLER_37_144 vgnd vpwr scs8hd_decap_4
XFILLER_80_434 vgnd vpwr scs8hd_decap_12
XFILLER_52_125 vpwr vgnd scs8hd_fill_2
XFILLER_37_188 vgnd vpwr scs8hd_fill_1
XFILLER_18_391 vgnd vpwr scs8hd_decap_6
XFILLER_21_501 vgnd vpwr scs8hd_decap_12
XFILLER_40_309 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ _131_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__353__B _272_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XFILLER_0_416 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_56_431 vpwr vgnd scs8hd_fill_2
XFILLER_28_122 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_301 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _155_/Y vgnd vpwr scs8hd_diode_2
XFILLER_71_489 vgnd vpwr scs8hd_decap_12
XPHY_312 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_323 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_334 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_345 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_356 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_367 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_378 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_389 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_99 vpwr vgnd scs8hd_fill_2
XANTENNA__263__B _272_/B vgnd vpwr scs8hd_diode_2
XFILLER_79_501 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ _208_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch_SLEEPB _230_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_111 vgnd vpwr scs8hd_fill_1
XFILLER_19_90 vgnd vpwr scs8hd_decap_4
XFILLER_19_144 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_199 vpwr vgnd scs8hd_fill_2
XFILLER_47_475 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
+ _395_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__173__B _173_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_239 vgnd vpwr scs8hd_decap_4
XFILLER_57_228 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_423 vpwr vgnd scs8hd_fill_2
XFILLER_25_114 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch_SLEEPB _329_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__348__B _352_/B vgnd vpwr scs8hd_diode_2
XFILLER_25_158 vpwr vgnd scs8hd_fill_2
XFILLER_53_489 vgnd vpwr scs8hd_decap_12
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XFILLER_15_59 vpwr vgnd scs8hd_fill_2
XANTENNA__364__A _170_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_331 vgnd vpwr scs8hd_fill_1
XFILLER_21_386 vpwr vgnd scs8hd_fill_2
XFILLER_21_397 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_213 vpwr vgnd scs8hd_fill_2
XFILLER_76_515 vgnd vpwr scs8hd_fill_1
XFILLER_0_268 vgnd vpwr scs8hd_decap_4
XFILLER_48_206 vpwr vgnd scs8hd_fill_2
XFILLER_56_44 vgnd vpwr scs8hd_decap_12
XFILLER_29_464 vpwr vgnd scs8hd_fill_2
XANTENNA__258__B _262_/B vgnd vpwr scs8hd_diode_2
XFILLER_44_412 vpwr vgnd scs8hd_fill_2
XFILLER_71_231 vpwr vgnd scs8hd_fill_2
XFILLER_72_32 vgnd vpwr scs8hd_decap_12
XFILLER_71_253 vgnd vpwr scs8hd_decap_3
XFILLER_44_467 vgnd vpwr scs8hd_decap_3
XPHY_142 vgnd vpwr scs8hd_decap_3
XPHY_131 vgnd vpwr scs8hd_decap_3
XPHY_120 vgnd vpwr scs8hd_decap_3
XPHY_164 vgnd vpwr scs8hd_decap_3
XPHY_153 vgnd vpwr scs8hd_decap_3
XANTENNA__274__A _274_/A vgnd vpwr scs8hd_diode_2
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_79_342 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_239 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _181_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_423 vpwr vgnd scs8hd_fill_2
XFILLER_47_272 vgnd vpwr scs8hd_decap_4
XFILLER_47_283 vpwr vgnd scs8hd_fill_2
XFILLER_47_294 vpwr vgnd scs8hd_fill_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_478 vgnd vpwr scs8hd_decap_8
XFILLER_35_489 vgnd vpwr scs8hd_decap_12
XANTENNA__184__A address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _133_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch_SLEEPB _302_/Y vgnd vpwr scs8hd_diode_2
XFILLER_58_515 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__359__A _287_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_401 vpwr vgnd scs8hd_fill_2
XFILLER_38_250 vgnd vpwr scs8hd_decap_4
XFILLER_53_231 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ _173_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_283 vpwr vgnd scs8hd_fill_2
XFILLER_53_275 vgnd vpwr scs8hd_fill_1
XFILLER_53_297 vpwr vgnd scs8hd_fill_2
XFILLER_21_161 vpwr vgnd scs8hd_fill_2
XFILLER_42_68 vgnd vpwr scs8hd_decap_12
XANTENNA__244__D _263_/D vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ _422_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch/Q
+ _354_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_76_312 vgnd vpwr scs8hd_decap_12
XFILLER_67_98 vgnd vpwr scs8hd_decap_4
XFILLER_64_507 vgnd vpwr scs8hd_decap_8
XANTENNA__269__A _287_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch/Q
+ _319_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_423 vgnd vpwr scs8hd_decap_4
XFILLER_29_283 vgnd vpwr scs8hd_decap_3
XFILLER_17_489 vgnd vpwr scs8hd_decap_12
XFILLER_16_80 vgnd vpwr scs8hd_decap_12
XFILLER_44_297 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch/Q
+ _284_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_183 vgnd vpwr scs8hd_fill_1
XFILLER_8_154 vgnd vpwr scs8hd_decap_3
XFILLER_8_143 vgnd vpwr scs8hd_decap_8
XFILLER_8_132 vgnd vpwr scs8hd_decap_8
XFILLER_40_492 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_334 vgnd vpwr scs8hd_decap_4
XFILLER_67_301 vpwr vgnd scs8hd_fill_2
XFILLER_67_367 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch/Q
+ _248_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__179__A _122_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_82_304 vgnd vpwr scs8hd_decap_6
XFILLER_67_389 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch_SLEEPB _275_/Y vgnd vpwr scs8hd_diode_2
XFILLER_35_297 vpwr vgnd scs8hd_fill_2
XFILLER_50_267 vgnd vpwr scs8hd_decap_6
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
XANTENNA__361__B _359_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_308 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_323 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
+ _412_/Y vgnd vpwr scs8hd_diode_2
XFILLER_73_304 vgnd vpwr scs8hd_fill_1
XFILLER_58_389 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ _149_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_340_ _231_/A _343_/B _340_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_459 vgnd vpwr scs8hd_decap_12
XFILLER_41_245 vgnd vpwr scs8hd_decap_3
X_271_ _280_/A _269_/B _271_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_278 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_146 vgnd vpwr scs8hd_decap_4
XANTENNA__271__B _269_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_49_334 vgnd vpwr scs8hd_decap_3
XFILLER_64_348 vpwr vgnd scs8hd_fill_2
XFILLER_17_264 vpwr vgnd scs8hd_fill_2
XFILLER_27_90 vpwr vgnd scs8hd_fill_2
XFILLER_72_392 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_20_407 vpwr vgnd scs8hd_fill_2
XFILLER_32_267 vgnd vpwr scs8hd_decap_6
XFILLER_9_452 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch/Q
+ _227_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_64_3 vgnd vpwr scs8hd_decap_12
XANTENNA__181__B _181_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch_SLEEPB _247_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_67_142 vpwr vgnd scs8hd_fill_2
XFILLER_67_175 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_82_156 vgnd vpwr scs8hd_decap_12
XPHY_708 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ _400_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_212 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_719 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__356__B _359_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XFILLER_23_59 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__372__A _194_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_105 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_58_120 vgnd vpwr scs8hd_decap_3
XFILLER_48_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch_SLEEPB _346_/Y vgnd vpwr scs8hd_diode_2
XFILLER_64_44 vgnd vpwr scs8hd_decap_12
XFILLER_61_329 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__266__B _269_/B vgnd vpwr scs8hd_diode_2
XFILLER_80_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_39 vgnd vpwr scs8hd_decap_12
X_323_ _287_/A _325_/B _323_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_254_ _263_/A _272_/B _272_/C _272_/D _262_/B vgnd vpwr scs8hd_or4_4
XANTENNA__282__A _273_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_495 vgnd vpwr scs8hd_decap_12
X_185_ _122_/Y _287_/A _391_/A vgnd vpwr scs8hd_or2_4
XFILLER_77_440 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_49_175 vpwr vgnd scs8hd_fill_2
XFILLER_37_348 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_45_370 vgnd vpwr scs8hd_decap_6
XANTENNA__176__B _176_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_260 vgnd vpwr scs8hd_decap_4
XANTENNA__192__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_271 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _147_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
XFILLER_68_495 vgnd vpwr scs8hd_decap_12
XFILLER_28_348 vgnd vpwr scs8hd_fill_1
XFILLER_55_156 vpwr vgnd scs8hd_fill_2
XANTENNA__367__A _367_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_510 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XPHY_505 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_516 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_51_362 vgnd vpwr scs8hd_fill_1
XPHY_527 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_538 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_549 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_259 vpwr vgnd scs8hd_fill_2
XFILLER_7_208 vpwr vgnd scs8hd_fill_2
XFILLER_50_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch_SLEEPB _319_/Y vgnd vpwr scs8hd_diode_2
XFILLER_78_215 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_74_410 vgnd vpwr scs8hd_decap_12
XFILLER_75_98 vgnd vpwr scs8hd_decap_12
XANTENNA__277__A _231_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch/Q ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
X_306_ _279_/A _304_/B _306_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_80 vgnd vpwr scs8hd_decap_12
X_237_ _274_/A _243_/B _237_/Y vgnd vpwr scs8hd_nor2_4
X_168_ _178_/A _181_/B _181_/C _273_/A vgnd vpwr scs8hd_or3_4
XFILLER_6_241 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_215 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ _378_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
XFILLER_77_281 vgnd vpwr scs8hd_decap_12
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XFILLER_1_51 vgnd vpwr scs8hd_decap_8
XANTENNA__187__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_37_134 vgnd vpwr scs8hd_decap_8
XFILLER_1_84 vpwr vgnd scs8hd_fill_2
XFILLER_80_446 vgnd vpwr scs8hd_decap_12
XFILLER_21_513 vgnd vpwr scs8hd_decap_3
XFILLER_33_362 vpwr vgnd scs8hd_fill_2
XANTENNA__353__C _163_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_0_428 vgnd vpwr scs8hd_decap_6
XFILLER_16_318 vpwr vgnd scs8hd_fill_2
XFILLER_43_115 vpwr vgnd scs8hd_fill_2
XPHY_302 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_313 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_324 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_351 vgnd vpwr scs8hd_decap_6
XFILLER_51_181 vpwr vgnd scs8hd_fill_2
XPHY_335 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_346 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_357 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_368 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_379 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__263__C _272_/C vgnd vpwr scs8hd_diode_2
XFILLER_79_513 vgnd vpwr scs8hd_decap_3
XFILLER_10_93 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ _140_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_123 vpwr vgnd scs8hd_fill_2
XFILLER_47_421 vgnd vpwr scs8hd_decap_4
XFILLER_47_432 vgnd vpwr scs8hd_decap_3
XFILLER_59_292 vpwr vgnd scs8hd_fill_2
XFILLER_47_487 vgnd vpwr scs8hd_fill_1
XFILLER_62_457 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_362 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_398 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q
+ _349_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_443 vpwr vgnd scs8hd_fill_2
XFILLER_65_273 vgnd vpwr scs8hd_decap_3
XFILLER_53_402 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _156_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q
+ _314_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_295 vpwr vgnd scs8hd_fill_2
XFILLER_53_457 vpwr vgnd scs8hd_fill_2
XFILLER_53_446 vgnd vpwr scs8hd_fill_1
XFILLER_53_435 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ _139_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_148 vgnd vpwr scs8hd_fill_1
XFILLER_80_276 vgnd vpwr scs8hd_decap_12
XFILLER_53_479 vgnd vpwr scs8hd_decap_8
XFILLER_15_27 vgnd vpwr scs8hd_decap_12
XFILLER_40_107 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_321 vpwr vgnd scs8hd_fill_2
XFILLER_33_170 vpwr vgnd scs8hd_fill_2
XANTENNA__364__B _367_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_365 vgnd vpwr scs8hd_fill_1
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q
+ _279_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__380__A _380_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_247 vgnd vpwr scs8hd_fill_1
XFILLER_48_229 vpwr vgnd scs8hd_fill_2
XFILLER_56_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q
+ _243_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_56_273 vpwr vgnd scs8hd_fill_2
XFILLER_72_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_143 vgnd vpwr scs8hd_decap_3
XPHY_132 vgnd vpwr scs8hd_decap_3
XPHY_121 vgnd vpwr scs8hd_decap_3
XPHY_110 vgnd vpwr scs8hd_decap_3
XPHY_165 vgnd vpwr scs8hd_decap_3
XPHY_154 vgnd vpwr scs8hd_decap_3
XANTENNA__274__B _280_/B vgnd vpwr scs8hd_diode_2
XFILLER_12_354 vgnd vpwr scs8hd_fill_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_387 vgnd vpwr scs8hd_decap_8
XFILLER_8_325 vpwr vgnd scs8hd_fill_2
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__290__A _263_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_79_354 vgnd vpwr scs8hd_decap_12
XFILLER_35_402 vpwr vgnd scs8hd_fill_2
XANTENNA__168__C _181_/C vgnd vpwr scs8hd_diode_2
XFILLER_35_435 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch/Q
+ _328_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_35_457 vpwr vgnd scs8hd_fill_2
XFILLER_62_276 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
+ _391_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__184__B _181_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_391 vpwr vgnd scs8hd_fill_2
XFILLER_7_380 vgnd vpwr scs8hd_decap_4
XFILLER_7_94 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch/Q
+ _293_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__359__B _359_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
+ clk ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff/QN
+ reset set vgnd vpwr scs8hd_dfbbp_1
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _143_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XFILLER_26_413 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch/Q
+ _258_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_468 vgnd vpwr scs8hd_decap_12
XFILLER_13_129 vpwr vgnd scs8hd_fill_2
XANTENNA__375__A _202_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_140 vpwr vgnd scs8hd_fill_2
XFILLER_21_184 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q
+ _222_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_339 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_501 vgnd vpwr scs8hd_decap_12
XFILLER_76_324 vgnd vpwr scs8hd_decap_12
XANTENNA__269__B _269_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_240 vpwr vgnd scs8hd_fill_2
XFILLER_29_262 vpwr vgnd scs8hd_fill_2
XFILLER_44_210 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__285__A _276_/A vgnd vpwr scs8hd_diode_2
XFILLER_44_276 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_195 vgnd vpwr scs8hd_decap_4
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_79_184 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ _404_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__179__B _276_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_50_213 vgnd vpwr scs8hd_fill_1
XANTENNA__195__A _178_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_257 vpwr vgnd scs8hd_fill_2
XFILLER_50_279 vgnd vpwr scs8hd_decap_3
XFILLER_58_335 vgnd vpwr scs8hd_fill_1
XFILLER_66_390 vgnd vpwr scs8hd_decap_6
XFILLER_26_243 vpwr vgnd scs8hd_fill_2
XFILLER_26_254 vpwr vgnd scs8hd_fill_2
XFILLER_41_224 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_270_ _279_/A _269_/B _270_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_471 vgnd vpwr scs8hd_decap_12
XFILLER_5_114 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_154 vgnd vpwr scs8hd_decap_12
XFILLER_64_316 vpwr vgnd scs8hd_fill_2
XFILLER_64_327 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/Y _135_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _139_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_32_213 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch_SLEEPB _343_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_298 vpwr vgnd scs8hd_fill_2
XFILLER_32_224 vgnd vpwr scs8hd_decap_12
XFILLER_32_257 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
X_399_ _377_/A _391_/B _399_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_464 vgnd vpwr scs8hd_decap_12
XFILLER_57_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__181__C _181_/C vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_191 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_55_349 vgnd vpwr scs8hd_decap_8
XFILLER_55_338 vpwr vgnd scs8hd_fill_2
XFILLER_82_168 vgnd vpwr scs8hd_decap_12
XPHY_709 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_408 vpwr vgnd scs8hd_fill_2
XFILLER_23_27 vgnd vpwr scs8hd_decap_12
XANTENNA__372__B _367_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ _157_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_48_68 vgnd vpwr scs8hd_decap_12
XFILLER_73_135 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_64_56 vgnd vpwr scs8hd_decap_12
XFILLER_54_371 vpwr vgnd scs8hd_fill_2
XFILLER_54_360 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_224 vpwr vgnd scs8hd_fill_2
X_322_ _231_/A _325_/B _322_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_80_44 vgnd vpwr scs8hd_decap_12
X_253_ address[8] _235_/B _272_/C vgnd vpwr scs8hd_nand2_4
XANTENNA__282__B _286_/B vgnd vpwr scs8hd_diode_2
XFILLER_10_430 vgnd vpwr scs8hd_decap_12
XFILLER_6_401 vgnd vpwr scs8hd_decap_12
X_184_ address[2] _181_/B address[0] _287_/A vgnd vpwr scs8hd_or3_4
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch_SLEEPB _316_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_132 vpwr vgnd scs8hd_fill_2
XFILLER_77_452 vgnd vpwr scs8hd_decap_12
XFILLER_49_187 vpwr vgnd scs8hd_fill_2
XFILLER_64_157 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_341 vgnd vpwr scs8hd_decap_3
XFILLER_45_382 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__192__B _371_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_294 vpwr vgnd scs8hd_fill_2
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XFILLER_28_327 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _157_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__367__B _367_/B vgnd vpwr scs8hd_diode_2
XFILLER_70_105 vgnd vpwr scs8hd_decap_12
XFILLER_55_179 vpwr vgnd scs8hd_fill_2
XFILLER_70_149 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
+ _377_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XFILLER_36_393 vgnd vpwr scs8hd_decap_4
XPHY_506 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_517 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_528 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_539 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_227 vpwr vgnd scs8hd_fill_2
XANTENNA__383__A _178_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_426 vgnd vpwr scs8hd_fill_1
XFILLER_78_227 vgnd vpwr scs8hd_decap_12
XFILLER_74_422 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_102 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _153_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__277__B _280_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_382 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch_SLEEPB _289_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__293__A _247_/A vgnd vpwr scs8hd_diode_2
X_305_ _287_/A _304_/B _305_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_42_396 vgnd vpwr scs8hd_fill_1
X_236_ _273_/A _243_/B _236_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_260 vgnd vpwr scs8hd_decap_6
XFILLER_6_253 vgnd vpwr scs8hd_fill_1
XFILLER_6_231 vgnd vpwr scs8hd_fill_1
X_167_ address[4] _166_/X _202_/A vgnd vpwr scs8hd_or2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _148_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_65_400 vgnd vpwr scs8hd_decap_4
XFILLER_77_293 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_74 vgnd vpwr scs8hd_decap_8
XANTENNA__187__B _187_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_371 vpwr vgnd scs8hd_fill_2
XFILLER_52_138 vgnd vpwr scs8hd_decap_4
XFILLER_33_341 vpwr vgnd scs8hd_fill_2
XFILLER_33_374 vgnd vpwr scs8hd_decap_4
XFILLER_33_396 vpwr vgnd scs8hd_fill_2
XFILLER_60_193 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__353__D _263_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_15 vgnd vpwr scs8hd_decap_12
XFILLER_75_208 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ _213_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_59 vpwr vgnd scs8hd_fill_2
XANTENNA__378__A _208_/B vgnd vpwr scs8hd_diode_2
XFILLER_71_403 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_16_308 vgnd vpwr scs8hd_fill_1
XFILLER_28_168 vgnd vpwr scs8hd_decap_3
XFILLER_43_127 vpwr vgnd scs8hd_fill_2
XPHY_303 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_314 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_325 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_336 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_347 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_358 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_385 vpwr vgnd scs8hd_fill_2
XFILLER_8_507 vgnd vpwr scs8hd_decap_8
XPHY_369 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__263__D _263_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_256 vpwr vgnd scs8hd_fill_2
XANTENNA__288__A _279_/A vgnd vpwr scs8hd_diode_2
XFILLER_47_400 vpwr vgnd scs8hd_fill_2
XFILLER_74_274 vgnd vpwr scs8hd_fill_1
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ _133_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_311 vpwr vgnd scs8hd_fill_2
XFILLER_30_344 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_219_ _274_/A _225_/B _219_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_57_208 vgnd vpwr scs8hd_fill_1
XANTENNA__198__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_411 vpwr vgnd scs8hd_fill_2
XFILLER_65_252 vgnd vpwr scs8hd_decap_4
XFILLER_25_127 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch_SLEEPB _360_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_39 vgnd vpwr scs8hd_decap_12
XFILLER_80_288 vgnd vpwr scs8hd_decap_12
XFILLER_61_480 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_300 vgnd vpwr scs8hd_decap_3
XFILLER_33_193 vpwr vgnd scs8hd_fill_2
XFILLER_31_27 vgnd vpwr scs8hd_decap_12
XANTENNA__380__B _362_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_411 vpwr vgnd scs8hd_fill_2
XFILLER_56_68 vgnd vpwr scs8hd_decap_12
XFILLER_56_285 vgnd vpwr scs8hd_decap_3
XPHY_100 vgnd vpwr scs8hd_decap_3
XFILLER_72_56 vgnd vpwr scs8hd_decap_12
XFILLER_71_288 vgnd vpwr scs8hd_decap_12
XPHY_133 vgnd vpwr scs8hd_decap_3
XPHY_122 vgnd vpwr scs8hd_decap_3
XPHY_111 vgnd vpwr scs8hd_decap_3
XPHY_155 vgnd vpwr scs8hd_decap_3
XPHY_144 vgnd vpwr scs8hd_decap_3
XFILLER_12_333 vgnd vpwr scs8hd_decap_3
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_193 vpwr vgnd scs8hd_fill_2
XFILLER_12_366 vpwr vgnd scs8hd_fill_2
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_348 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__290__B address[7] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ _148_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
+ _416_/Y vgnd vpwr scs8hd_diode_2
XFILLER_82_509 vgnd vpwr scs8hd_decap_6
XFILLER_47_241 vgnd vpwr scs8hd_decap_3
XFILLER_62_255 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_428 vpwr vgnd scs8hd_fill_2
XFILLER_15_171 vpwr vgnd scs8hd_fill_2
XFILLER_22_108 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__184__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_30_152 vgnd vpwr scs8hd_fill_1
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XFILLER_7_51 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_263 vgnd vpwr scs8hd_decap_12
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XFILLER_26_425 vgnd vpwr scs8hd_decap_3
XFILLER_13_119 vgnd vpwr scs8hd_decap_3
XANTENNA__375__B _367_/B vgnd vpwr scs8hd_diode_2
XFILLER_41_417 vgnd vpwr scs8hd_decap_8
XFILLER_41_428 vpwr vgnd scs8hd_fill_2
XFILLER_41_439 vpwr vgnd scs8hd_fill_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA__391__A _391_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_174 vgnd vpwr scs8hd_decap_3
XFILLER_1_513 vgnd vpwr scs8hd_decap_3
XANTENNA__285__B _286_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_439 vpwr vgnd scs8hd_fill_2
XFILLER_16_93 vpwr vgnd scs8hd_fill_2
XFILLER_12_141 vgnd vpwr scs8hd_decap_12
XFILLER_40_450 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ _155_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_79_196 vgnd vpwr scs8hd_decap_12
XFILLER_67_358 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _144_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ _144_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_75_391 vgnd vpwr scs8hd_decap_12
XFILLER_35_200 vpwr vgnd scs8hd_fill_2
XFILLER_35_211 vpwr vgnd scs8hd_fill_2
XANTENNA__195__B _181_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_439 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_225 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_450 vpwr vgnd scs8hd_fill_2
XFILLER_31_461 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_73_306 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch/Q ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_222 vgnd vpwr scs8hd_decap_4
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__386__A _170_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_236 vpwr vgnd scs8hd_fill_2
XFILLER_22_483 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch_SLEEPB _219_/Y vgnd vpwr scs8hd_diode_2
XFILLER_78_44 vgnd vpwr scs8hd_decap_12
XFILLER_76_166 vgnd vpwr scs8hd_decap_12
XFILLER_64_306 vgnd vpwr scs8hd_decap_3
XFILLER_57_380 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_391 vpwr vgnd scs8hd_fill_2
XANTENNA__296__A _287_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_277 vpwr vgnd scs8hd_fill_2
XFILLER_32_236 vpwr vgnd scs8hd_fill_2
X_398_ _204_/B _391_/B _398_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_476 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ _194_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_155 vpwr vgnd scs8hd_fill_2
XFILLER_55_306 vpwr vgnd scs8hd_fill_2
XFILLER_82_125 vgnd vpwr scs8hd_decap_12
XFILLER_67_188 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_23_203 vgnd vpwr scs8hd_decap_3
XFILLER_63_394 vgnd vpwr scs8hd_decap_6
XFILLER_23_236 vgnd vpwr scs8hd_decap_6
XFILLER_23_258 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_58_133 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_317 vgnd vpwr scs8hd_decap_8
XFILLER_46_328 vgnd vpwr scs8hd_decap_8
XFILLER_73_147 vgnd vpwr scs8hd_decap_12
XFILLER_61_309 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_64_68 vgnd vpwr scs8hd_decap_12
XFILLER_14_247 vgnd vpwr scs8hd_decap_3
X_321_ _276_/A _325_/B _321_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_80_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
X_252_ _280_/A _252_/B _252_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_442 vgnd vpwr scs8hd_decap_12
X_183_ _202_/A _183_/B _183_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_413 vgnd vpwr scs8hd_decap_12
XFILLER_6_457 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_184 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_464 vgnd vpwr scs8hd_decap_12
XFILLER_37_306 vpwr vgnd scs8hd_fill_2
XFILLER_49_155 vpwr vgnd scs8hd_fill_2
XFILLER_37_328 vgnd vpwr scs8hd_fill_1
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XFILLER_49_199 vpwr vgnd scs8hd_fill_2
XFILLER_33_501 vgnd vpwr scs8hd_decap_12
XFILLER_72_191 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch_SLEEPB _291_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_240 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch/Q ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_114 vpwr vgnd scs8hd_fill_2
XFILLER_55_136 vpwr vgnd scs8hd_fill_2
XFILLER_70_117 vgnd vpwr scs8hd_decap_12
XFILLER_43_309 vpwr vgnd scs8hd_fill_2
XFILLER_63_180 vgnd vpwr scs8hd_fill_1
XFILLER_51_331 vgnd vpwr scs8hd_decap_8
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XPHY_507 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _210_/Y vgnd vpwr scs8hd_diode_2
XPHY_518 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_529 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__383__B _380_/X vgnd vpwr scs8hd_diode_2
XFILLER_50_15 vgnd vpwr scs8hd_decap_12
XFILLER_78_239 vgnd vpwr scs8hd_decap_12
XFILLER_19_317 vpwr vgnd scs8hd_fill_2
XFILLER_74_434 vgnd vpwr scs8hd_decap_12
XFILLER_46_125 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ _416_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_501 vgnd vpwr scs8hd_decap_12
XFILLER_61_139 vpwr vgnd scs8hd_fill_2
XFILLER_42_320 vgnd vpwr scs8hd_decap_4
XFILLER_42_364 vpwr vgnd scs8hd_fill_2
XANTENNA__293__B _295_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_304_ _231_/A _304_/B _304_/Y vgnd vpwr scs8hd_nor2_4
X_235_ address[8] _235_/B _235_/C _272_/D _243_/B vgnd vpwr scs8hd_or4_4
XFILLER_24_93 vgnd vpwr scs8hd_decap_3
X_166_ address[6] address[7] _163_/X _263_/D _166_/X vgnd vpwr scs8hd_or4_4
XFILLER_6_276 vpwr vgnd scs8hd_fill_2
XFILLER_6_265 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_206 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch_SLEEPB _264_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_471 vgnd vpwr scs8hd_decap_12
XFILLER_37_114 vpwr vgnd scs8hd_fill_2
XFILLER_65_445 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _158_/Y vgnd vpwr scs8hd_diode_2
XFILLER_65_489 vgnd vpwr scs8hd_decap_12
XFILLER_80_459 vgnd vpwr scs8hd_decap_12
XFILLER_60_172 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_27 vgnd vpwr scs8hd_decap_12
XFILLER_68_272 vgnd vpwr scs8hd_decap_3
XANTENNA__378__B _367_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_103 vpwr vgnd scs8hd_fill_2
XFILLER_56_456 vpwr vgnd scs8hd_fill_2
XFILLER_71_415 vgnd vpwr scs8hd_decap_12
XFILLER_43_106 vpwr vgnd scs8hd_fill_2
XFILLER_45_15 vgnd vpwr scs8hd_decap_12
XFILLER_45_59 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__394__A _194_/B vgnd vpwr scs8hd_diode_2
XPHY_304 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_315 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_515 vgnd vpwr scs8hd_fill_1
XPHY_326 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_337 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_348 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_359 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_84 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_209 vgnd vpwr scs8hd_fill_1
XANTENNA__288__B _286_/B vgnd vpwr scs8hd_diode_2
XFILLER_59_272 vgnd vpwr scs8hd_decap_4
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
XFILLER_47_489 vgnd vpwr scs8hd_decap_12
XFILLER_62_426 vgnd vpwr scs8hd_decap_4
XFILLER_34_128 vgnd vpwr scs8hd_fill_1
XFILLER_34_139 vgnd vpwr scs8hd_decap_12
XFILLER_62_459 vgnd vpwr scs8hd_decap_12
XFILLER_15_331 vgnd vpwr scs8hd_decap_3
XFILLER_15_353 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch_SLEEPB _236_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_386 vgnd vpwr scs8hd_decap_6
XFILLER_42_194 vgnd vpwr scs8hd_decap_3
XFILLER_30_378 vgnd vpwr scs8hd_decap_8
XFILLER_30_389 vpwr vgnd scs8hd_fill_2
X_218_ _273_/A _225_/B _218_/Y vgnd vpwr scs8hd_nor2_4
X_149_ _149_/A _149_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_290 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__198__B _181_/C vgnd vpwr scs8hd_diode_2
XFILLER_21_345 vgnd vpwr scs8hd_decap_6
XFILLER_21_367 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ _394_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_507 vgnd vpwr scs8hd_decap_8
XANTENNA__389__A _367_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_249 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
+ clk vgnd vpwr scs8hd_diode_2
XFILLER_29_423 vpwr vgnd scs8hd_fill_2
XFILLER_29_445 vgnd vpwr scs8hd_decap_8
XFILLER_29_489 vgnd vpwr scs8hd_decap_12
XFILLER_16_106 vpwr vgnd scs8hd_fill_2
XFILLER_44_437 vgnd vpwr scs8hd_decap_4
XFILLER_71_267 vpwr vgnd scs8hd_fill_2
XFILLER_72_68 vgnd vpwr scs8hd_decap_12
XPHY_134 vgnd vpwr scs8hd_decap_3
XPHY_123 vgnd vpwr scs8hd_decap_3
XPHY_112 vgnd vpwr scs8hd_decap_3
XPHY_101 vgnd vpwr scs8hd_decap_3
XFILLER_12_312 vgnd vpwr scs8hd_decap_4
XPHY_156 vgnd vpwr scs8hd_decap_3
XPHY_145 vgnd vpwr scs8hd_decap_3
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__290__C _272_/C vgnd vpwr scs8hd_diode_2
XFILLER_79_367 vgnd vpwr scs8hd_decap_12
XANTENNA__299__A _263_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_209 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_62_223 vpwr vgnd scs8hd_fill_2
XFILLER_62_212 vpwr vgnd scs8hd_fill_2
XFILLER_62_201 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2/Z
+ _141_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_62_234 vgnd vpwr scs8hd_decap_12
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_46_80 vgnd vpwr scs8hd_fill_1
XFILLER_62_267 vgnd vpwr scs8hd_decap_6
XFILLER_15_150 vpwr vgnd scs8hd_fill_2
XPHY_690 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_256 vpwr vgnd scs8hd_fill_2
XFILLER_53_278 vgnd vpwr scs8hd_decap_4
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__391__B _391_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_319 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_337 vgnd vpwr scs8hd_decap_12
XFILLER_17_415 vpwr vgnd scs8hd_fill_2
XFILLER_17_437 vgnd vpwr scs8hd_decap_12
XFILLER_29_275 vgnd vpwr scs8hd_decap_6
XFILLER_29_297 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_267 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ _156_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_179 vgnd vpwr scs8hd_decap_4
XFILLER_32_93 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_315 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _139_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_256 vpwr vgnd scs8hd_fill_2
XFILLER_50_215 vgnd vpwr scs8hd_decap_3
XANTENNA__195__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_23_407 vpwr vgnd scs8hd_fill_2
XFILLER_23_418 vpwr vgnd scs8hd_fill_2
XFILLER_35_278 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ _372_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _132_/Y vgnd vpwr scs8hd_diode_2
XFILLER_58_304 vgnd vpwr scs8hd_decap_4
XFILLER_58_348 vgnd vpwr scs8hd_decap_8
XFILLER_58_359 vgnd vpwr scs8hd_decap_4
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XFILLER_73_318 vgnd vpwr scs8hd_decap_12
XFILLER_26_201 vgnd vpwr scs8hd_decap_3
XFILLER_26_212 vpwr vgnd scs8hd_fill_2
XANTENNA__386__B _391_/B vgnd vpwr scs8hd_diode_2
XFILLER_53_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_407 vgnd vpwr scs8hd_decap_12
XFILLER_26_267 vgnd vpwr scs8hd_decap_8
XFILLER_26_289 vpwr vgnd scs8hd_fill_2
XFILLER_53_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_259 vpwr vgnd scs8hd_fill_2
XFILLER_22_495 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_127 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ _390_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_78_56 vgnd vpwr scs8hd_decap_12
XFILLER_1_311 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
+ _431_/HI ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_49_359 vgnd vpwr scs8hd_decap_4
XFILLER_76_178 vgnd vpwr scs8hd_decap_12
XFILLER_17_223 vpwr vgnd scs8hd_fill_2
XANTENNA__296__B _295_/B vgnd vpwr scs8hd_diode_2
XFILLER_17_256 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_440 vgnd vpwr scs8hd_decap_12
X_397_ _202_/B _391_/B _397_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_411 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_292 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_67_134 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_82_137 vgnd vpwr scs8hd_decap_12
XFILLER_63_362 vpwr vgnd scs8hd_fill_2
XFILLER_63_384 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_15 vgnd vpwr scs8hd_decap_12
XFILLER_58_101 vpwr vgnd scs8hd_fill_2
XFILLER_58_145 vpwr vgnd scs8hd_fill_2
XANTENNA__397__A _202_/B vgnd vpwr scs8hd_diode_2
XFILLER_58_189 vgnd vpwr scs8hd_decap_4
XFILLER_58_167 vpwr vgnd scs8hd_fill_2
XFILLER_73_159 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch/Q
+ _273_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_215 vpwr vgnd scs8hd_fill_2
X_320_ _247_/A _325_/B _320_/Y vgnd vpwr scs8hd_nor2_4
X_251_ _279_/A _252_/B _251_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_80_68 vgnd vpwr scs8hd_decap_12
XFILLER_13_51 vgnd vpwr scs8hd_decap_8
X_182_ _122_/Y _231_/A _183_/B vgnd vpwr scs8hd_or2_4
XFILLER_10_454 vgnd vpwr scs8hd_decap_4
XFILLER_6_425 vgnd vpwr scs8hd_decap_12
XFILLER_13_62 vgnd vpwr scs8hd_decap_12
XFILLER_13_84 vpwr vgnd scs8hd_fill_2
XFILLER_13_95 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch/Q
+ _237_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_130 vpwr vgnd scs8hd_fill_2
XFILLER_49_112 vpwr vgnd scs8hd_fill_2
XFILLER_77_476 vgnd vpwr scs8hd_decap_12
XFILLER_64_115 vgnd vpwr scs8hd_decap_4
XFILLER_33_513 vgnd vpwr scs8hd_decap_3
XFILLER_45_395 vgnd vpwr scs8hd_decap_3
XFILLER_54_80 vgnd vpwr scs8hd_decap_12
XFILLER_60_376 vgnd vpwr scs8hd_fill_1
XFILLER_13_281 vpwr vgnd scs8hd_fill_2
XFILLER_13_292 vgnd vpwr scs8hd_decap_4
XFILLER_62_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_432 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ _132_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch_SLEEPB _261_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_362 vgnd vpwr scs8hd_fill_1
XFILLER_70_129 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_63_170 vpwr vgnd scs8hd_fill_2
XFILLER_51_321 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_508 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_365 vgnd vpwr scs8hd_fill_1
XPHY_519 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_376 vgnd vpwr scs8hd_decap_4
XFILLER_11_207 vgnd vpwr scs8hd_decap_4
XFILLER_50_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_428 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_487 vgnd vpwr scs8hd_fill_1
XFILLER_74_446 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_362 vpwr vgnd scs8hd_fill_2
XFILLER_82_490 vgnd vpwr scs8hd_decap_6
XFILLER_61_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_513 vgnd vpwr scs8hd_decap_3
XFILLER_27_395 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ _131_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_354 vgnd vpwr scs8hd_decap_3
X_303_ _276_/A _304_/B _303_/Y vgnd vpwr scs8hd_nor2_4
X_234_ _280_/A _231_/B _234_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_200 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_165_ _127_/Y address[5] _263_/D vgnd vpwr scs8hd_or2_4
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_483 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_65_424 vgnd vpwr scs8hd_fill_1
XFILLER_37_148 vgnd vpwr scs8hd_fill_1
XFILLER_52_129 vgnd vpwr scs8hd_decap_6
XFILLER_33_310 vgnd vpwr scs8hd_fill_1
XFILLER_45_170 vpwr vgnd scs8hd_fill_2
XFILLER_33_332 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch_SLEEPB _233_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
+ _398_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_435 vpwr vgnd scs8hd_fill_2
XFILLER_28_126 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_27 vgnd vpwr scs8hd_decap_12
XANTENNA__394__B _391_/B vgnd vpwr scs8hd_diode_2
XPHY_305 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_316 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_15 vgnd vpwr scs8hd_decap_12
XFILLER_51_173 vpwr vgnd scs8hd_fill_2
XFILLER_51_162 vpwr vgnd scs8hd_fill_2
XPHY_327 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_338 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_349 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_59 vpwr vgnd scs8hd_fill_2
XFILLER_51_184 vpwr vgnd scs8hd_fill_2
XFILLER_24_398 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_236 vgnd vpwr scs8hd_decap_3
XFILLER_3_225 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_269 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch_SLEEPB _332_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_413 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_83 vpwr vgnd scs8hd_fill_2
XFILLER_19_159 vgnd vpwr scs8hd_decap_3
XFILLER_47_457 vpwr vgnd scs8hd_fill_2
XFILLER_74_276 vgnd vpwr scs8hd_decap_12
XFILLER_62_449 vgnd vpwr scs8hd_decap_8
XFILLER_27_170 vpwr vgnd scs8hd_fill_2
XFILLER_70_471 vgnd vpwr scs8hd_decap_12
XFILLER_15_376 vgnd vpwr scs8hd_decap_4
XFILLER_42_173 vgnd vpwr scs8hd_decap_8
XFILLER_15_398 vpwr vgnd scs8hd_fill_2
X_217_ address[8] _235_/B _215_/X _272_/D _225_/B vgnd vpwr scs8hd_or4_4
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_148_ _148_/A _148_/Y vgnd vpwr scs8hd_inv_8
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch/Q ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__198__C address[1] vgnd vpwr scs8hd_diode_2
XFILLER_38_424 vgnd vpwr scs8hd_decap_8
XFILLER_65_243 vgnd vpwr scs8hd_fill_1
XFILLER_38_457 vgnd vpwr scs8hd_fill_1
XFILLER_80_202 vgnd vpwr scs8hd_decap_12
XFILLER_65_287 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_53_449 vpwr vgnd scs8hd_fill_2
XFILLER_18_192 vpwr vgnd scs8hd_fill_2
XFILLER_46_490 vgnd vpwr scs8hd_decap_12
XFILLER_21_357 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__389__B _391_/B vgnd vpwr scs8hd_diode_2
XFILLER_56_221 vgnd vpwr scs8hd_decap_4
XFILLER_56_15 vgnd vpwr scs8hd_decap_12
XFILLER_56_265 vpwr vgnd scs8hd_fill_2
XFILLER_56_254 vgnd vpwr scs8hd_decap_4
XFILLER_29_468 vgnd vpwr scs8hd_decap_12
XFILLER_16_129 vpwr vgnd scs8hd_fill_2
XFILLER_44_416 vgnd vpwr scs8hd_decap_4
XFILLER_71_235 vgnd vpwr scs8hd_decap_6
XPHY_124 vgnd vpwr scs8hd_decap_3
XPHY_113 vgnd vpwr scs8hd_decap_3
XPHY_102 vgnd vpwr scs8hd_decap_3
XPHY_157 vgnd vpwr scs8hd_decap_3
XPHY_146 vgnd vpwr scs8hd_decap_3
XPHY_135 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch_SLEEPB _305_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_346 vgnd vpwr scs8hd_decap_8
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_51 vgnd vpwr scs8hd_decap_8
XFILLER_21_62 vgnd vpwr scs8hd_decap_12
XANTENNA__290__D _272_/D vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q
+ _359_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__299__B address[7] vgnd vpwr scs8hd_diode_2
XFILLER_79_379 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_287 vpwr vgnd scs8hd_fill_2
XFILLER_47_298 vgnd vpwr scs8hd_decap_4
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_184 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q
+ _324_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_482 vgnd vpwr scs8hd_decap_6
XPHY_680 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_62_80 vgnd vpwr scs8hd_decap_12
XFILLER_30_132 vgnd vpwr scs8hd_decap_3
XFILLER_30_154 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_691 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_86 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q
+ _289_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_213 vgnd vpwr scs8hd_fill_1
XFILLER_26_405 vpwr vgnd scs8hd_fill_2
XFILLER_38_287 vpwr vgnd scs8hd_fill_2
XFILLER_53_235 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _150_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch_SLEEPB _278_/Y vgnd vpwr scs8hd_diode_2
XFILLER_76_349 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_254 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_449 vgnd vpwr scs8hd_decap_12
XFILLER_25_471 vgnd vpwr scs8hd_decap_12
XFILLER_12_154 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch/Q
+ _338_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
+ _192_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_79_110 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch/Q ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch/Q
+ _303_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_67_338 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _149_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_471 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q
+ _268_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_43_290 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ _364_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q
+ _232_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_58_327 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
XFILLER_66_360 vgnd vpwr scs8hd_decap_8
XFILLER_81_330 vgnd vpwr scs8hd_decap_12
XFILLER_66_382 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_53_27 vgnd vpwr scs8hd_decap_12
XFILLER_14_419 vgnd vpwr scs8hd_decap_12
XFILLER_26_279 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch_SLEEPB _250_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_301 vpwr vgnd scs8hd_fill_2
XFILLER_1_334 vpwr vgnd scs8hd_fill_2
XFILLER_78_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_367 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _140_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_94 vpwr vgnd scs8hd_fill_2
XFILLER_72_396 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_452 vgnd vpwr scs8hd_decap_12
XFILLER_32_249 vpwr vgnd scs8hd_fill_2
X_396_ _200_/B _391_/B _396_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_489 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch_SLEEPB _349_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XFILLER_67_102 vgnd vpwr scs8hd_fill_1
XFILLER_67_179 vpwr vgnd scs8hd_fill_2
XFILLER_82_149 vgnd vpwr scs8hd_decap_6
XFILLER_48_393 vpwr vgnd scs8hd_fill_2
XFILLER_63_341 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_227 vpwr vgnd scs8hd_fill_2
XFILLER_31_260 vgnd vpwr scs8hd_decap_3
XFILLER_31_293 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_109 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_48_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__397__B _391_/B vgnd vpwr scs8hd_diode_2
XFILLER_64_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_81_171 vgnd vpwr scs8hd_decap_12
XFILLER_54_396 vgnd vpwr scs8hd_fill_1
X_250_ _287_/A _252_/B _250_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_181_ address[2] _181_/B _181_/C _231_/A vgnd vpwr scs8hd_or3_4
XFILLER_22_293 vpwr vgnd scs8hd_fill_2
XFILLER_13_74 vgnd vpwr scs8hd_decap_3
XFILLER_6_459 vgnd vpwr scs8hd_decap_12
XFILLER_6_437 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch/Q ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_175 vpwr vgnd scs8hd_fill_2
XFILLER_1_164 vpwr vgnd scs8hd_fill_2
XFILLER_49_179 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XFILLER_45_341 vpwr vgnd scs8hd_fill_2
XFILLER_72_171 vgnd vpwr scs8hd_decap_12
XFILLER_60_311 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch_SLEEPB _322_/Y vgnd vpwr scs8hd_diode_2
XFILLER_60_355 vgnd vpwr scs8hd_decap_8
XFILLER_20_208 vgnd vpwr scs8hd_fill_1
X_379_ _210_/B _367_/B _379_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_70_80 vgnd vpwr scs8hd_decap_12
XFILLER_9_275 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/Y _157_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_68_444 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_341 vgnd vpwr scs8hd_decap_4
XFILLER_51_344 vpwr vgnd scs8hd_fill_2
XPHY_509 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_59_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_59 vpwr vgnd scs8hd_fill_2
XFILLER_59_400 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_inv_1
XFILLER_59_455 vpwr vgnd scs8hd_fill_2
XFILLER_59_444 vpwr vgnd scs8hd_fill_2
XFILLER_59_433 vgnd vpwr scs8hd_decap_4
XANTENNA__201__A address[3] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_54_193 vpwr vgnd scs8hd_fill_2
XFILLER_54_182 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_333 vgnd vpwr scs8hd_fill_1
X_302_ _247_/A _304_/B _302_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_42_377 vgnd vpwr scs8hd_decap_8
XFILLER_42_388 vpwr vgnd scs8hd_fill_2
X_233_ _279_/A _231_/B _233_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
X_164_ address[6] address[7] _235_/C vgnd vpwr scs8hd_or2_4
XFILLER_10_285 vgnd vpwr scs8hd_decap_3
XFILLER_10_296 vgnd vpwr scs8hd_decap_8
XFILLER_69_219 vpwr vgnd scs8hd_fill_2
XFILLER_2_495 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_92 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_65_458 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_52_108 vgnd vpwr scs8hd_decap_8
XFILLER_45_193 vgnd vpwr scs8hd_decap_4
XFILLER_60_185 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _145_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ _140_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_56_414 vgnd vpwr scs8hd_decap_6
XFILLER_71_428 vgnd vpwr scs8hd_decap_12
XFILLER_36_171 vpwr vgnd scs8hd_fill_2
XFILLER_43_119 vgnd vpwr scs8hd_decap_3
XFILLER_45_39 vgnd vpwr scs8hd_decap_12
XPHY_306 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_36_182 vgnd vpwr scs8hd_decap_8
XFILLER_36_193 vpwr vgnd scs8hd_fill_2
XPHY_317 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_328 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_339 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
+ _381_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_204 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_74_222 vgnd vpwr scs8hd_decap_12
XFILLER_59_296 vpwr vgnd scs8hd_fill_2
XFILLER_19_51 vgnd vpwr scs8hd_decap_8
XFILLER_19_62 vgnd vpwr scs8hd_decap_12
XFILLER_19_127 vpwr vgnd scs8hd_fill_2
XFILLER_74_288 vgnd vpwr scs8hd_decap_12
XFILLER_62_439 vpwr vgnd scs8hd_fill_2
XFILLER_34_119 vpwr vgnd scs8hd_fill_2
XPHY_840 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_483 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_30_347 vpwr vgnd scs8hd_fill_2
X_216_ enable address[5] _272_/D vgnd vpwr scs8hd_nand2_4
X_147_ _147_/A _147_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_447 vpwr vgnd scs8hd_fill_2
XFILLER_53_406 vpwr vgnd scs8hd_fill_2
XFILLER_65_299 vgnd vpwr scs8hd_decap_6
XFILLER_21_325 vgnd vpwr scs8hd_decap_6
XFILLER_33_174 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ _410_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q
+ _333_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ _147_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_218 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_211 vgnd vpwr scs8hd_decap_3
XFILLER_56_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q
+ _298_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_71_214 vpwr vgnd scs8hd_fill_2
XFILLER_72_15 vgnd vpwr scs8hd_decap_12
XPHY_125 vgnd vpwr scs8hd_decap_3
XPHY_114 vgnd vpwr scs8hd_decap_3
XFILLER_52_450 vgnd vpwr scs8hd_decap_8
XPHY_103 vgnd vpwr scs8hd_decap_3
XPHY_158 vgnd vpwr scs8hd_decap_3
XPHY_147 vgnd vpwr scs8hd_decap_3
XPHY_136 vgnd vpwr scs8hd_decap_3
XFILLER_52_472 vgnd vpwr scs8hd_decap_4
XFILLER_12_325 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/Y _146_/A vgnd vpwr scs8hd_inv_1
XFILLER_24_163 vgnd vpwr scs8hd_decap_3
XFILLER_24_174 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_329 vgnd vpwr scs8hd_decap_4
XFILLER_21_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _141_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__299__C _272_/C vgnd vpwr scs8hd_diode_2
XFILLER_47_200 vgnd vpwr scs8hd_decap_3
XFILLER_47_233 vpwr vgnd scs8hd_fill_2
XFILLER_47_255 vpwr vgnd scs8hd_fill_2
XFILLER_35_406 vpwr vgnd scs8hd_fill_2
XFILLER_28_491 vgnd vpwr scs8hd_decap_12
XFILLER_46_93 vpwr vgnd scs8hd_fill_2
XFILLER_50_409 vgnd vpwr scs8hd_decap_8
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_15_130 vpwr vgnd scs8hd_fill_2
XFILLER_43_450 vgnd vpwr scs8hd_decap_4
XFILLER_43_461 vpwr vgnd scs8hd_fill_2
XPHY_670 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_144 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XPHY_692 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_681 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_177 vgnd vpwr scs8hd_decap_6
XFILLER_30_188 vgnd vpwr scs8hd_decap_3
XFILLER_11_380 vpwr vgnd scs8hd_fill_2
XFILLER_7_362 vpwr vgnd scs8hd_fill_2
XFILLER_81_501 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_409 vpwr vgnd scs8hd_fill_2
XFILLER_61_280 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _132_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_472 vgnd vpwr scs8hd_decap_12
XFILLER_21_144 vpwr vgnd scs8hd_fill_2
XFILLER_21_199 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_69_380 vpwr vgnd scs8hd_fill_2
XFILLER_67_59 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_222 vgnd vpwr scs8hd_decap_3
XFILLER_17_428 vgnd vpwr scs8hd_decap_3
XFILLER_25_461 vgnd vpwr scs8hd_decap_3
XFILLER_25_483 vgnd vpwr scs8hd_decap_4
XFILLER_52_291 vpwr vgnd scs8hd_fill_2
XFILLER_4_398 vgnd vpwr scs8hd_decap_3
XFILLER_63_501 vgnd vpwr scs8hd_decap_12
XFILLER_35_236 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_206 vgnd vpwr scs8hd_fill_1
XFILLER_16_483 vgnd vpwr scs8hd_decap_12
XFILLER_31_475 vgnd vpwr scs8hd_fill_1
XFILLER_31_486 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _159_/Y vgnd vpwr scs8hd_diode_2
XFILLER_81_342 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_53_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ _158_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_118 vgnd vpwr scs8hd_decap_4
XANTENNA__204__A _202_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_49_317 vpwr vgnd scs8hd_fill_2
XFILLER_49_339 vpwr vgnd scs8hd_fill_2
XFILLER_45_501 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_236 vpwr vgnd scs8hd_fill_2
XFILLER_27_51 vgnd vpwr scs8hd_decap_8
XFILLER_27_62 vgnd vpwr scs8hd_decap_12
XFILLER_60_515 vgnd vpwr scs8hd_fill_1
XFILLER_32_206 vgnd vpwr scs8hd_decap_4
XFILLER_13_464 vgnd vpwr scs8hd_decap_12
X_395_ _197_/B _391_/B _395_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_94 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_195 vgnd vpwr scs8hd_decap_4
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XFILLER_68_80 vgnd vpwr scs8hd_decap_12
XFILLER_67_114 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_99 vgnd vpwr scs8hd_fill_1
XFILLER_82_106 vgnd vpwr scs8hd_decap_12
XFILLER_63_320 vpwr vgnd scs8hd_fill_2
XFILLER_48_383 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_272 vgnd vpwr scs8hd_decap_4
XFILLER_58_125 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
+ _403_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_501 vgnd vpwr scs8hd_decap_12
XFILLER_66_180 vgnd vpwr scs8hd_decap_8
XFILLER_64_27 vgnd vpwr scs8hd_decap_4
XFILLER_54_320 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_383 vpwr vgnd scs8hd_fill_2
XFILLER_54_331 vgnd vpwr scs8hd_decap_4
XFILLER_54_375 vgnd vpwr scs8hd_decap_4
XFILLER_14_206 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_239 vgnd vpwr scs8hd_decap_6
XFILLER_80_15 vgnd vpwr scs8hd_decap_12
X_180_ _202_/A _367_/A _180_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_449 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _155_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch/Q ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_49_136 vpwr vgnd scs8hd_fill_2
XFILLER_77_489 vgnd vpwr scs8hd_decap_12
XFILLER_64_139 vgnd vpwr scs8hd_decap_12
XFILLER_64_128 vgnd vpwr scs8hd_decap_8
XFILLER_60_301 vgnd vpwr scs8hd_fill_1
XFILLER_72_183 vgnd vpwr scs8hd_decap_8
XFILLER_54_93 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_389 vpwr vgnd scs8hd_fill_2
X_447_ _447_/HI _447_/LO vgnd vpwr scs8hd_conb_1
XFILLER_9_221 vpwr vgnd scs8hd_fill_2
X_378_ _208_/B _367_/B _378_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_298 vgnd vpwr scs8hd_decap_4
XFILLER_48_3 vgnd vpwr scs8hd_decap_12
XFILLER_68_456 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_161 vpwr vgnd scs8hd_fill_2
XFILLER_51_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_27 vgnd vpwr scs8hd_decap_12
XFILLER_59_423 vpwr vgnd scs8hd_fill_2
XFILLER_75_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_489 vgnd vpwr scs8hd_decap_12
XANTENNA__201__B _276_/A vgnd vpwr scs8hd_diode_2
XFILLER_75_59 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_320 vgnd vpwr scs8hd_decap_4
XFILLER_46_117 vpwr vgnd scs8hd_fill_2
XFILLER_74_459 vgnd vpwr scs8hd_decap_12
XFILLER_54_172 vgnd vpwr scs8hd_fill_1
X_301_ _274_/A _304_/B _301_/Y vgnd vpwr scs8hd_nor2_4
X_232_ _287_/A _231_/B _232_/Y vgnd vpwr scs8hd_nor2_4
X_163_ address[8] address[9] _163_/X vgnd vpwr scs8hd_or2_4
XFILLER_6_224 vgnd vpwr scs8hd_decap_4
XFILLER_77_220 vgnd vpwr scs8hd_decap_12
XFILLER_65_404 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_301 vpwr vgnd scs8hd_fill_2
XFILLER_33_345 vpwr vgnd scs8hd_fill_2
XFILLER_60_142 vgnd vpwr scs8hd_fill_1
XFILLER_33_378 vgnd vpwr scs8hd_fill_1
XANTENNA__302__A _247_/A vgnd vpwr scs8hd_diode_2
XFILLER_68_264 vgnd vpwr scs8hd_decap_8
XFILLER_56_448 vgnd vpwr scs8hd_decap_8
XFILLER_28_139 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ _133_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_307 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_312 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_507 vgnd vpwr scs8hd_decap_8
XPHY_318 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_329 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_389 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch/Q ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__212__A _171_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_74 vpwr vgnd scs8hd_fill_2
XFILLER_74_234 vgnd vpwr scs8hd_decap_12
XFILLER_19_96 vpwr vgnd scs8hd_fill_2
XFILLER_47_448 vpwr vgnd scs8hd_fill_2
XFILLER_62_407 vgnd vpwr scs8hd_decap_12
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XFILLER_42_120 vgnd vpwr scs8hd_fill_1
XFILLER_70_451 vgnd vpwr scs8hd_decap_6
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
XPHY_841 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_830 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_495 vgnd vpwr scs8hd_decap_12
XFILLER_30_315 vpwr vgnd scs8hd_fill_2
X_215_ _263_/A address[7] _215_/X vgnd vpwr scs8hd_or2_4
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
X_146_ _146_/A _146_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__122__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_271 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_223 vpwr vgnd scs8hd_fill_2
XFILLER_76_80 vgnd vpwr scs8hd_decap_12
XFILLER_65_234 vpwr vgnd scs8hd_fill_2
XFILLER_38_459 vgnd vpwr scs8hd_decap_12
XFILLER_80_215 vgnd vpwr scs8hd_decap_12
XFILLER_33_142 vgnd vpwr scs8hd_decap_4
XFILLER_33_153 vpwr vgnd scs8hd_fill_2
XFILLER_21_315 vgnd vpwr scs8hd_decap_4
XFILLER_21_337 vpwr vgnd scs8hd_fill_2
XFILLER_33_197 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
+ _419_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ _148_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_208 vgnd vpwr scs8hd_decap_3
XFILLER_29_415 vgnd vpwr scs8hd_decap_6
XFILLER_29_437 vpwr vgnd scs8hd_fill_2
XFILLER_44_429 vgnd vpwr scs8hd_decap_6
XFILLER_71_248 vgnd vpwr scs8hd_decap_3
XFILLER_72_27 vgnd vpwr scs8hd_decap_4
XPHY_115 vgnd vpwr scs8hd_decap_3
XPHY_104 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XPHY_148 vgnd vpwr scs8hd_decap_3
XPHY_137 vgnd vpwr scs8hd_decap_3
XPHY_126 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_159 vgnd vpwr scs8hd_decap_3
XFILLER_8_308 vpwr vgnd scs8hd_fill_2
XFILLER_24_197 vgnd vpwr scs8hd_decap_4
XANTENNA__207__A _181_/C vgnd vpwr scs8hd_diode_2
XFILLER_21_86 vpwr vgnd scs8hd_fill_2
XANTENNA__299__D _263_/D vgnd vpwr scs8hd_diode_2
XFILLER_47_223 vpwr vgnd scs8hd_fill_2
XFILLER_47_245 vgnd vpwr scs8hd_decap_4
XFILLER_62_215 vgnd vpwr scs8hd_decap_8
XFILLER_47_278 vpwr vgnd scs8hd_fill_2
XFILLER_62_259 vgnd vpwr scs8hd_decap_4
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XFILLER_30_112 vgnd vpwr scs8hd_decap_6
XPHY_671 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_660 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_693 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_682 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_62_93 vgnd vpwr scs8hd_decap_8
X_129_ address[6] _263_/A vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
XFILLER_81_513 vgnd vpwr scs8hd_decap_3
XFILLER_34_484 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_123 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ _155_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
+ _425_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_189 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch/Q ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_67_27 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_44_215 vpwr vgnd scs8hd_fill_2
XFILLER_12_112 vgnd vpwr scs8hd_decap_4
XFILLER_40_443 vpwr vgnd scs8hd_fill_2
XFILLER_12_167 vgnd vpwr scs8hd_decap_12
XFILLER_8_105 vpwr vgnd scs8hd_fill_2
XFILLER_4_366 vpwr vgnd scs8hd_fill_2
XFILLER_79_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__400__A _208_/B vgnd vpwr scs8hd_diode_2
XFILLER_63_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch_SLEEPB _222_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_204 vgnd vpwr scs8hd_decap_4
XFILLER_35_226 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_248 vpwr vgnd scs8hd_fill_2
XFILLER_16_495 vgnd vpwr scs8hd_decap_12
XFILLER_31_454 vpwr vgnd scs8hd_fill_2
XFILLER_31_465 vpwr vgnd scs8hd_fill_2
XFILLER_78_3 vgnd vpwr scs8hd_decap_12
XPHY_490 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_193 vpwr vgnd scs8hd_fill_2
XFILLER_7_171 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ _206_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__310__A _274_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_215 vpwr vgnd scs8hd_fill_2
XFILLER_26_226 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_81_354 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_218 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_15 vgnd vpwr scs8hd_decap_12
XANTENNA__204__B _204_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _151_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_1_347 vpwr vgnd scs8hd_fill_2
XFILLER_1_358 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__220__A _247_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_57_395 vpwr vgnd scs8hd_fill_2
XFILLER_57_384 vpwr vgnd scs8hd_fill_2
XFILLER_57_373 vgnd vpwr scs8hd_fill_1
XFILLER_45_513 vgnd vpwr scs8hd_decap_3
XFILLER_27_74 vgnd vpwr scs8hd_decap_12
XFILLER_72_398 vgnd vpwr scs8hd_decap_12
XFILLER_25_281 vgnd vpwr scs8hd_decap_4
XFILLER_9_425 vpwr vgnd scs8hd_fill_2
X_394_ _194_/B _391_/B _394_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_476 vgnd vpwr scs8hd_decap_12
XFILLER_40_262 vgnd vpwr scs8hd_decap_4
XFILLER_43_51 vgnd vpwr scs8hd_decap_8
XFILLER_43_62 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _160_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_141 vpwr vgnd scs8hd_fill_2
XFILLER_4_174 vgnd vpwr scs8hd_decap_6
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
XANTENNA__130__A address[7] vgnd vpwr scs8hd_diode_2
XFILLER_67_159 vgnd vpwr scs8hd_decap_3
XFILLER_48_362 vgnd vpwr scs8hd_decap_4
XFILLER_82_118 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_63_354 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_63_376 vpwr vgnd scs8hd_fill_2
XFILLER_16_270 vgnd vpwr scs8hd_decap_4
XFILLER_31_240 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch/Q ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__305__A _287_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch_SLEEPB _294_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_170 vgnd vpwr scs8hd_fill_1
XFILLER_27_513 vgnd vpwr scs8hd_decap_3
XFILLER_81_184 vgnd vpwr scs8hd_decap_12
XFILLER_54_398 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_80_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
+ set vgnd vpwr scs8hd_diode_2
XANTENNA__215__A _263_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_188 vgnd vpwr scs8hd_decap_3
XFILLER_64_107 vgnd vpwr scs8hd_fill_1
XFILLER_49_159 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ _131_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_45_310 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ _170_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
+ _386_/Y vgnd vpwr scs8hd_diode_2
X_446_ _446_/HI _446_/LO vgnd vpwr scs8hd_conb_1
XFILLER_60_379 vgnd vpwr scs8hd_fill_1
XFILLER_9_211 vgnd vpwr scs8hd_fill_1
X_377_ _377_/A _367_/B _377_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ _421_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_70_93 vgnd vpwr scs8hd_decap_12
XANTENNA__125__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch/Q
+ _318_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_55_118 vpwr vgnd scs8hd_fill_2
XFILLER_36_310 vgnd vpwr scs8hd_fill_1
XFILLER_51_313 vpwr vgnd scs8hd_fill_2
XFILLER_36_365 vpwr vgnd scs8hd_fill_2
XFILLER_63_184 vgnd vpwr scs8hd_decap_4
XFILLER_36_398 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch/Q
+ _283_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch_SLEEPB _267_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _156_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch/Q
+ _247_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_75_27 vgnd vpwr scs8hd_decap_12
XFILLER_46_129 vgnd vpwr scs8hd_fill_1
X_300_ _273_/A _304_/B _300_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_42_324 vgnd vpwr scs8hd_fill_1
XFILLER_42_346 vgnd vpwr scs8hd_decap_8
X_231_ _231_/A _231_/B _231_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_243 vpwr vgnd scs8hd_fill_2
X_162_ _162_/A _162_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_77_232 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_416 vpwr vgnd scs8hd_fill_2
XFILLER_37_118 vpwr vgnd scs8hd_fill_2
XFILLER_18_365 vgnd vpwr scs8hd_decap_4
XFILLER_18_376 vgnd vpwr scs8hd_decap_8
XFILLER_45_140 vgnd vpwr scs8hd_decap_8
XFILLER_60_121 vpwr vgnd scs8hd_fill_2
XFILLER_18_387 vpwr vgnd scs8hd_fill_2
XFILLER_18_398 vpwr vgnd scs8hd_fill_2
XFILLER_33_324 vpwr vgnd scs8hd_fill_2
XFILLER_60_154 vgnd vpwr scs8hd_decap_3
X_429_ _429_/HI _429_/LO vgnd vpwr scs8hd_conb_1
XFILLER_60_3 vgnd vpwr scs8hd_decap_12
XANTENNA__302__B _304_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch_SLEEPB _239_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_276 vgnd vpwr scs8hd_decap_4
XFILLER_28_107 vgnd vpwr scs8hd_decap_6
XFILLER_64_471 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
+ _212_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_140 vgnd vpwr scs8hd_decap_6
XFILLER_51_132 vpwr vgnd scs8hd_fill_2
XPHY_308 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_319 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_368 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_10_44 vgnd vpwr scs8hd_decap_12
XFILLER_10_99 vpwr vgnd scs8hd_fill_2
XANTENNA__212__B _214_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/Y _134_/A vgnd vpwr scs8hd_inv_1
XFILLER_74_202 vgnd vpwr scs8hd_decap_12
XFILLER_59_276 vgnd vpwr scs8hd_fill_1
XFILLER_19_107 vgnd vpwr scs8hd_decap_4
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_74_246 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ _399_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_140 vpwr vgnd scs8hd_fill_2
XFILLER_15_313 vgnd vpwr scs8hd_decap_4
XFILLER_27_195 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch_SLEEPB _338_/Y vgnd vpwr scs8hd_diode_2
XPHY_820 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_42_132 vpwr vgnd scs8hd_fill_2
XPHY_842 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_831 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_42_165 vpwr vgnd scs8hd_fill_2
X_214_ _178_/B _214_/B _214_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_51_62 vgnd vpwr scs8hd_decap_12
XFILLER_51_51 vgnd vpwr scs8hd_decap_8
XFILLER_7_501 vgnd vpwr scs8hd_decap_12
XFILLER_51_95 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_145_ _145_/A _145_/Y vgnd vpwr scs8hd_inv_8
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ _142_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__403__A _171_/X vgnd vpwr scs8hd_diode_2
XFILLER_2_283 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_419 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_80_227 vgnd vpwr scs8hd_decap_12
XFILLER_18_173 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _134_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__313__A _231_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_56_235 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_116 vgnd vpwr scs8hd_decap_3
XPHY_105 vgnd vpwr scs8hd_decap_3
XPHY_149 vgnd vpwr scs8hd_decap_3
XPHY_138 vgnd vpwr scs8hd_decap_3
XPHY_127 vgnd vpwr scs8hd_decap_3
XFILLER_52_485 vgnd vpwr scs8hd_decap_12
XANTENNA__207__B address[1] vgnd vpwr scs8hd_diode_2
XFILLER_4_515 vgnd vpwr scs8hd_fill_1
XANTENNA__223__A _287_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch_SLEEPB _311_/Y vgnd vpwr scs8hd_diode_2
XFILLER_62_205 vgnd vpwr scs8hd_decap_4
XFILLER_35_419 vpwr vgnd scs8hd_fill_2
XFILLER_46_84 vgnd vpwr scs8hd_decap_8
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_154 vpwr vgnd scs8hd_fill_2
XFILLER_43_474 vpwr vgnd scs8hd_fill_2
XPHY_661 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_650 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_694 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_683 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_672 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/Y _152_/A vgnd vpwr scs8hd_inv_1
XFILLER_11_393 vgnd vpwr scs8hd_decap_4
X_128_ address[9] _235_/B vgnd vpwr scs8hd_inv_8
XANTENNA__133__A _133_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_202 vgnd vpwr scs8hd_decap_12
XFILLER_38_224 vgnd vpwr scs8hd_decap_12
XFILLER_38_246 vpwr vgnd scs8hd_fill_2
XFILLER_38_279 vpwr vgnd scs8hd_fill_2
XFILLER_53_227 vpwr vgnd scs8hd_fill_2
XFILLER_53_216 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
+ _372_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_496 vgnd vpwr scs8hd_decap_12
XANTENNA__308__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_21_157 vpwr vgnd scs8hd_fill_2
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_67_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ _377_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_69_371 vgnd vpwr scs8hd_decap_6
XFILLER_29_213 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_419 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_227 vgnd vpwr scs8hd_fill_1
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch_SLEEPB _284_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_411 vgnd vpwr scs8hd_decap_12
XANTENNA__218__A _273_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_124 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_117 vgnd vpwr scs8hd_fill_1
XFILLER_12_179 vgnd vpwr scs8hd_decap_4
XFILLER_4_389 vgnd vpwr scs8hd_decap_8
XFILLER_79_135 vgnd vpwr scs8hd_decap_12
XFILLER_75_330 vgnd vpwr scs8hd_decap_12
XANTENNA__400__B _391_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_290 vpwr vgnd scs8hd_fill_2
XANTENNA__128__A address[9] vgnd vpwr scs8hd_diode_2
XFILLER_31_433 vpwr vgnd scs8hd_fill_2
XPHY_480 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_491 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_58_319 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__310__B _314_/B vgnd vpwr scs8hd_diode_2
XFILLER_78_190 vgnd vpwr scs8hd_decap_12
XFILLER_66_396 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
+ _365_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch/Q
+ _348_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_78_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_315 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_105 vgnd vpwr scs8hd_decap_12
XANTENNA__220__B _225_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_341 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_205 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q
+ _313_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_72_344 vgnd vpwr scs8hd_decap_12
XFILLER_72_333 vgnd vpwr scs8hd_decap_3
XFILLER_27_86 vpwr vgnd scs8hd_fill_2
XFILLER_25_260 vpwr vgnd scs8hd_fill_2
X_393_ _371_/A _391_/B _393_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_43_74 vgnd vpwr scs8hd_decap_12
XFILLER_40_285 vgnd vpwr scs8hd_fill_1
XFILLER_40_296 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q
+ _278_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _155_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_131 vgnd vpwr scs8hd_fill_1
XFILLER_4_120 vpwr vgnd scs8hd_fill_2
XANTENNA__411__A _367_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_68 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_68_93 vgnd vpwr scs8hd_decap_12
XFILLER_67_138 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q
+ _242_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_48_330 vgnd vpwr scs8hd_decap_4
XFILLER_48_341 vgnd vpwr scs8hd_decap_3
XFILLER_75_171 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch_SLEEPB _355_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_208 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _148_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_230 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
+ clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__305__B _304_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch/Q ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_58_105 vpwr vgnd scs8hd_fill_2
XANTENNA__321__A _276_/A vgnd vpwr scs8hd_diode_2
XFILLER_58_149 vgnd vpwr scs8hd_decap_4
XFILLER_39_352 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_363 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch/Q
+ _327_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_54_388 vgnd vpwr scs8hd_decap_8
XFILLER_81_196 vgnd vpwr scs8hd_decap_12
XFILLER_22_241 vgnd vpwr scs8hd_decap_4
XFILLER_22_252 vgnd vpwr scs8hd_decap_6
XFILLER_22_285 vgnd vpwr scs8hd_decap_8
XANTENNA__215__B address[7] vgnd vpwr scs8hd_diode_2
XFILLER_13_99 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch/Q
+ _292_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_134 vpwr vgnd scs8hd_fill_2
XFILLER_1_123 vpwr vgnd scs8hd_fill_2
XFILLER_77_403 vgnd vpwr scs8hd_decap_12
XANTENNA__231__A _231_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ _132_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch/Q ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_49_116 vgnd vpwr scs8hd_decap_4
XFILLER_57_160 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch/Q
+ _257_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_45_300 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_72_141 vgnd vpwr scs8hd_decap_12
XFILLER_72_196 vpwr vgnd scs8hd_fill_2
X_445_ _445_/HI _445_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_263 vgnd vpwr scs8hd_decap_6
XFILLER_13_285 vpwr vgnd scs8hd_fill_2
X_376_ _204_/B _367_/B _376_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_267 vpwr vgnd scs8hd_fill_2
XFILLER_9_256 vpwr vgnd scs8hd_fill_2
XANTENNA__406__A address[6] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch/Q
+ _221_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_440 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__141__A _141_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_333 vgnd vpwr scs8hd_decap_3
XFILLER_63_174 vgnd vpwr scs8hd_decap_6
XFILLER_51_358 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__316__A _280_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ _403_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_39 vgnd vpwr scs8hd_decap_12
XFILLER_27_300 vpwr vgnd scs8hd_fill_2
XFILLER_39_160 vpwr vgnd scs8hd_fill_2
XFILLER_39_171 vpwr vgnd scs8hd_fill_2
XFILLER_54_163 vgnd vpwr scs8hd_decap_3
XFILLER_42_303 vgnd vpwr scs8hd_decap_3
XFILLER_24_32 vgnd vpwr scs8hd_decap_12
X_230_ _276_/A _231_/B _230_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__226__A address[8] vgnd vpwr scs8hd_diode_2
X_161_ _161_/A _161_/Y vgnd vpwr scs8hd_inv_8
XFILLER_10_266 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _401_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ _139_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_49_51 vgnd vpwr scs8hd_decap_8
XFILLER_49_62 vgnd vpwr scs8hd_decap_12
XFILLER_49_95 vpwr vgnd scs8hd_fill_2
XFILLER_65_428 vpwr vgnd scs8hd_fill_2
XFILLER_45_163 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_45_174 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_358 vpwr vgnd scs8hd_fill_2
X_428_ _428_/HI _428_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__136__A _136_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_380 vpwr vgnd scs8hd_fill_2
XFILLER_41_391 vgnd vpwr scs8hd_fill_1
X_359_ _287_/A _359_/B _359_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch/Q ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_270 vpwr vgnd scs8hd_fill_2
XFILLER_68_200 vpwr vgnd scs8hd_fill_2
XFILLER_68_233 vgnd vpwr scs8hd_decap_12
XFILLER_49_480 vgnd vpwr scs8hd_decap_8
XFILLER_64_450 vgnd vpwr scs8hd_decap_8
XFILLER_64_483 vgnd vpwr scs8hd_decap_12
XFILLER_36_163 vgnd vpwr scs8hd_decap_8
XPHY_309 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_188 vpwr vgnd scs8hd_fill_2
XFILLER_51_177 vpwr vgnd scs8hd_fill_2
XFILLER_51_166 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_229 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_56 vgnd vpwr scs8hd_decap_12
XFILLER_59_222 vpwr vgnd scs8hd_fill_2
XFILLER_59_255 vpwr vgnd scs8hd_fill_2
XFILLER_47_417 vpwr vgnd scs8hd_fill_2
XFILLER_47_428 vpwr vgnd scs8hd_fill_2
XFILLER_74_258 vgnd vpwr scs8hd_decap_12
XFILLER_82_280 vgnd vpwr scs8hd_decap_12
XFILLER_55_472 vpwr vgnd scs8hd_fill_2
XFILLER_15_336 vpwr vgnd scs8hd_fill_2
XFILLER_27_174 vpwr vgnd scs8hd_fill_2
XPHY_810 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_843 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_832 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_821 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_328 vgnd vpwr scs8hd_decap_8
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
X_213_ _187_/B _214_/B _213_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_380 vpwr vgnd scs8hd_fill_2
XFILLER_42_199 vpwr vgnd scs8hd_fill_2
XFILLER_7_513 vgnd vpwr scs8hd_decap_3
XFILLER_51_74 vgnd vpwr scs8hd_decap_12
X_144_ _144_/A _144_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__403__B _402_/X vgnd vpwr scs8hd_diode_2
XFILLER_76_93 vgnd vpwr scs8hd_decap_12
XFILLER_65_269 vpwr vgnd scs8hd_fill_2
XFILLER_18_152 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_450 vgnd vpwr scs8hd_decap_8
XFILLER_80_239 vgnd vpwr scs8hd_decap_12
XFILLER_33_100 vpwr vgnd scs8hd_fill_2
XFILLER_18_196 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_33_166 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/Y _149_/A vgnd vpwr scs8hd_buf_1
XANTENNA__313__B _314_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_56_203 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_56_225 vgnd vpwr scs8hd_fill_1
XFILLER_71_206 vgnd vpwr scs8hd_decap_6
XFILLER_56_269 vpwr vgnd scs8hd_fill_2
XFILLER_2_90 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_442 vgnd vpwr scs8hd_decap_4
XPHY_106 vgnd vpwr scs8hd_decap_3
XFILLER_24_133 vpwr vgnd scs8hd_fill_2
XPHY_139 vgnd vpwr scs8hd_decap_3
XPHY_128 vgnd vpwr scs8hd_decap_3
XPHY_117 vgnd vpwr scs8hd_decap_3
XFILLER_52_497 vgnd vpwr scs8hd_decap_12
XANTENNA__207__C address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__223__B _225_/B vgnd vpwr scs8hd_diode_2
XFILLER_79_306 vgnd vpwr scs8hd_decap_12
XFILLER_75_501 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_55_280 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XPHY_662 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_651 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_640 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch/Q ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_188 vpwr vgnd scs8hd_fill_2
XFILLER_15_199 vpwr vgnd scs8hd_fill_2
XPHY_695 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_684 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_673 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ _150_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__414__A _189_/B vgnd vpwr scs8hd_diode_2
X_127_ enable _127_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_398 vpwr vgnd scs8hd_fill_2
XFILLER_7_387 vpwr vgnd scs8hd_fill_2
XFILLER_7_376 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q
+ _343_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_361 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_236 vgnd vpwr scs8hd_fill_1
XFILLER_26_409 vpwr vgnd scs8hd_fill_2
XFILLER_53_239 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_280 vgnd vpwr scs8hd_decap_4
XFILLER_21_103 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
+ _200_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
XANTENNA__308__B address[7] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__324__A _279_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ _369_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_69_350 vgnd vpwr scs8hd_decap_6
XFILLER_57_501 vgnd vpwr scs8hd_decap_12
XFILLER_29_203 vgnd vpwr scs8hd_fill_1
XFILLER_29_236 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _147_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_258 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_72_515 vgnd vpwr scs8hd_fill_1
XFILLER_44_206 vpwr vgnd scs8hd_fill_2
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XFILLER_37_280 vgnd vpwr scs8hd_decap_3
XFILLER_44_239 vgnd vpwr scs8hd_decap_8
XANTENNA__218__B _225_/B vgnd vpwr scs8hd_diode_2
XFILLER_40_423 vgnd vpwr scs8hd_decap_4
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XANTENNA__234__A _280_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_98 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_79_147 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ _212_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_57_62 vgnd vpwr scs8hd_decap_12
XFILLER_57_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_342 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__409__A _173_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_280 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_209 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_423 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_31_478 vgnd vpwr scs8hd_decap_8
XPHY_470 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_489 vgnd vpwr scs8hd_decap_12
XPHY_481 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_492 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__144__A _144_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _146_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_501 vgnd vpwr scs8hd_decap_12
XFILLER_66_353 vgnd vpwr scs8hd_decap_4
XFILLER_54_504 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_386 vpwr vgnd scs8hd_fill_2
XFILLER_26_206 vgnd vpwr scs8hd_decap_4
XANTENNA__319__A _274_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_239 vpwr vgnd scs8hd_fill_2
XFILLER_81_367 vgnd vpwr scs8hd_decap_12
XFILLER_34_250 vgnd vpwr scs8hd_decap_4
XFILLER_22_434 vgnd vpwr scs8hd_fill_1
XFILLER_34_272 vgnd vpwr scs8hd_decap_3
XFILLER_34_283 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch_SLEEPB _352_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_117 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_72_356 vgnd vpwr scs8hd_decap_12
XFILLER_60_507 vgnd vpwr scs8hd_decap_8
XANTENNA__229__A _247_/A vgnd vpwr scs8hd_diode_2
X_392_ _189_/B _391_/B _392_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_40_242 vgnd vpwr scs8hd_decap_3
XFILLER_13_489 vgnd vpwr scs8hd_decap_12
XFILLER_43_86 vgnd vpwr scs8hd_decap_8
XFILLER_4_154 vgnd vpwr scs8hd_decap_3
XANTENNA__411__B _416_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_382 vpwr vgnd scs8hd_fill_2
XFILLER_0_393 vpwr vgnd scs8hd_fill_2
XFILLER_36_504 vgnd vpwr scs8hd_decap_12
XFILLER_48_375 vgnd vpwr scs8hd_decap_8
XANTENNA__139__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_297 vpwr vgnd scs8hd_fill_2
XFILLER_8_471 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__321__B _325_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch_SLEEPB _325_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_320 vpwr vgnd scs8hd_fill_2
XFILLER_39_331 vpwr vgnd scs8hd_fill_2
XFILLER_10_459 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _156_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__231__B _231_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_415 vgnd vpwr scs8hd_decap_12
XFILLER_1_179 vpwr vgnd scs8hd_fill_2
XFILLER_1_168 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_515 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_45_345 vpwr vgnd scs8hd_fill_2
XFILLER_45_378 vpwr vgnd scs8hd_fill_2
X_444_ _444_/HI _444_/LO vgnd vpwr scs8hd_conb_1
XFILLER_60_337 vpwr vgnd scs8hd_fill_2
XFILLER_13_231 vpwr vgnd scs8hd_fill_2
X_375_ _202_/B _367_/B _375_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__406__B address[7] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_452 vgnd vpwr scs8hd_decap_12
XANTENNA__422__A _208_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
+ _430_/HI ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_459 vgnd vpwr scs8hd_decap_12
XFILLER_36_345 vgnd vpwr scs8hd_fill_1
XFILLER_48_183 vpwr vgnd scs8hd_fill_2
XFILLER_48_194 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_131 vpwr vgnd scs8hd_fill_2
XFILLER_36_378 vgnd vpwr scs8hd_decap_8
XFILLER_36_389 vpwr vgnd scs8hd_fill_2
XFILLER_51_348 vgnd vpwr scs8hd_fill_1
XANTENNA__316__B _314_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_290 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__332__A _287_/A vgnd vpwr scs8hd_diode_2
XFILLER_59_404 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_59_459 vgnd vpwr scs8hd_decap_12
XFILLER_59_448 vgnd vpwr scs8hd_decap_4
XFILLER_67_470 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_27_345 vpwr vgnd scs8hd_fill_2
XFILLER_27_367 vpwr vgnd scs8hd_fill_2
XFILLER_27_378 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_50_370 vpwr vgnd scs8hd_fill_2
XFILLER_24_44 vgnd vpwr scs8hd_decap_12
XANTENNA__226__B _235_/B vgnd vpwr scs8hd_diode_2
XFILLER_50_392 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _143_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_99 vgnd vpwr scs8hd_decap_6
X_160_ _160_/A _160_/Y vgnd vpwr scs8hd_inv_8
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XANTENNA__242__A _279_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_77_245 vgnd vpwr scs8hd_decap_12
XFILLER_49_74 vgnd vpwr scs8hd_decap_12
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XFILLER_65_51 vgnd vpwr scs8hd_decap_8
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XFILLER_73_440 vgnd vpwr scs8hd_decap_12
XFILLER_65_62 vgnd vpwr scs8hd_decap_12
XFILLER_60_145 vpwr vgnd scs8hd_fill_2
XFILLER_45_197 vgnd vpwr scs8hd_fill_1
X_427_ _178_/B _424_/X _427_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__417__A _197_/B vgnd vpwr scs8hd_diode_2
X_358_ _231_/A _359_/B _358_/Y vgnd vpwr scs8hd_nor2_4
X_289_ _280_/A _286_/B _289_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__152__A _152_/A vgnd vpwr scs8hd_diode_2
XFILLER_46_3 vgnd vpwr scs8hd_decap_12
XFILLER_68_223 vgnd vpwr scs8hd_fill_1
XFILLER_68_289 vgnd vpwr scs8hd_decap_12
XFILLER_64_495 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_145 vpwr vgnd scs8hd_fill_2
XFILLER_51_123 vpwr vgnd scs8hd_fill_2
XFILLER_24_337 vgnd vpwr scs8hd_decap_3
XFILLER_36_197 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ _148_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__327__A _273_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ _192_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_208 vgnd vpwr scs8hd_decap_4
XFILLER_10_68 vgnd vpwr scs8hd_decap_12
XFILLER_59_212 vgnd vpwr scs8hd_decap_3
XFILLER_59_245 vgnd vpwr scs8hd_fill_1
XFILLER_74_215 vgnd vpwr scs8hd_decap_4
XFILLER_27_153 vpwr vgnd scs8hd_fill_2
XFILLER_42_112 vgnd vpwr scs8hd_decap_8
XFILLER_82_292 vgnd vpwr scs8hd_decap_12
XPHY_811 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_800 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_359 vgnd vpwr scs8hd_fill_1
XFILLER_42_145 vpwr vgnd scs8hd_fill_2
XPHY_844 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_833 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_822 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__237__A _274_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_98 vgnd vpwr scs8hd_decap_8
X_212_ _171_/X _214_/B _212_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_51_86 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ _147_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_143_ _143_/A _143_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_252 vgnd vpwr scs8hd_decap_4
XFILLER_65_204 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/Y _140_/A vgnd vpwr scs8hd_inv_1
XFILLER_38_407 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_248 vpwr vgnd scs8hd_fill_2
XFILLER_46_473 vgnd vpwr scs8hd_decap_8
XFILLER_61_443 vpwr vgnd scs8hd_fill_2
XFILLER_61_421 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
+ _173_/Y vgnd vpwr scs8hd_diode_2
XFILLER_33_123 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__147__A _147_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _161_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _139_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_215 vgnd vpwr scs8hd_decap_4
XFILLER_2_80 vgnd vpwr scs8hd_decap_8
XFILLER_37_451 vpwr vgnd scs8hd_fill_2
XFILLER_71_218 vpwr vgnd scs8hd_fill_2
XFILLER_37_462 vpwr vgnd scs8hd_fill_2
XPHY_107 vgnd vpwr scs8hd_decap_3
XPHY_129 vgnd vpwr scs8hd_decap_3
XPHY_118 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_178 vgnd vpwr scs8hd_decap_4
XANTENNA__207__D address[2] vgnd vpwr scs8hd_diode_2
XFILLER_20_340 vgnd vpwr scs8hd_decap_8
XFILLER_20_351 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_373 vpwr vgnd scs8hd_fill_2
XFILLER_79_318 vgnd vpwr scs8hd_decap_12
XFILLER_75_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_237 vpwr vgnd scs8hd_fill_2
XFILLER_47_259 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_134 vgnd vpwr scs8hd_decap_3
XPHY_652 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_641 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_630 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_30_104 vpwr vgnd scs8hd_fill_2
XPHY_696 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_685 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_674 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_663 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_362 vpwr vgnd scs8hd_fill_2
XANTENNA__414__B _416_/B vgnd vpwr scs8hd_diode_2
X_126_ address[4] _380_/A vgnd vpwr scs8hd_inv_8
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ _143_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch_SLEEPB _256_/Y vgnd vpwr scs8hd_diode_2
XFILLER_78_373 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ _415_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_440 vgnd vpwr scs8hd_decap_12
XFILLER_61_240 vpwr vgnd scs8hd_fill_2
XFILLER_61_284 vpwr vgnd scs8hd_fill_2
XANTENNA__308__C _272_/C vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/Y _158_/A vgnd vpwr scs8hd_inv_1
XANTENNA__324__B _325_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch/Q ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__340__A _231_/A vgnd vpwr scs8hd_diode_2
XFILLER_69_384 vgnd vpwr scs8hd_decap_4
XFILLER_57_513 vgnd vpwr scs8hd_decap_3
XFILLER_25_443 vpwr vgnd scs8hd_fill_2
XFILLER_52_251 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_56 vgnd vpwr scs8hd_decap_12
XFILLER_52_295 vpwr vgnd scs8hd_fill_2
XFILLER_25_487 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_468 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _157_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XANTENNA__234__B _231_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_192 vgnd vpwr scs8hd_fill_1
XANTENNA__250__A _287_/A vgnd vpwr scs8hd_diode_2
XFILLER_79_159 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_354 vgnd vpwr scs8hd_decap_12
XFILLER_57_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_62 vgnd vpwr scs8hd_decap_12
XFILLER_73_51 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__409__B _416_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_402 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _432_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_273 vpwr vgnd scs8hd_fill_2
XPHY_460 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_471 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch_SLEEPB _228_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__425__A _171_/X vgnd vpwr scs8hd_diode_2
XPHY_482 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_493 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_170 vpwr vgnd scs8hd_fill_2
XFILLER_7_141 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_380 vpwr vgnd scs8hd_fill_2
XANTENNA__160__A _160_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
+ _393_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _148_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_281 vgnd vpwr scs8hd_decap_4
XFILLER_26_229 vgnd vpwr scs8hd_fill_1
XFILLER_81_379 vgnd vpwr scs8hd_decap_12
XANTENNA__319__B _325_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_446 vgnd vpwr scs8hd_decap_12
XANTENNA__335__A _263_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_306 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch_SLEEPB _327_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_328 vgnd vpwr scs8hd_decap_4
XFILLER_76_129 vgnd vpwr scs8hd_decap_12
XFILLER_57_354 vpwr vgnd scs8hd_fill_2
XFILLER_72_313 vgnd vpwr scs8hd_decap_12
XFILLER_57_376 vgnd vpwr scs8hd_fill_1
XFILLER_72_368 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__229__B _231_/B vgnd vpwr scs8hd_diode_2
XFILLER_25_240 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_402 vpwr vgnd scs8hd_fill_2
XFILLER_13_413 vpwr vgnd scs8hd_fill_2
X_391_ _391_/A _391_/B _391_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_417 vgnd vpwr scs8hd_decap_8
XANTENNA__245__A _273_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_428 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch/Q ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ _393_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_67_118 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_184 vgnd vpwr scs8hd_decap_12
XFILLER_63_324 vpwr vgnd scs8hd_fill_2
XFILLER_48_398 vpwr vgnd scs8hd_fill_2
XFILLER_51_508 vgnd vpwr scs8hd_decap_8
XFILLER_16_262 vgnd vpwr scs8hd_decap_6
XFILLER_31_210 vpwr vgnd scs8hd_fill_2
XFILLER_31_221 vpwr vgnd scs8hd_fill_2
XFILLER_31_254 vgnd vpwr scs8hd_decap_4
XANTENNA__155__A _155_/A vgnd vpwr scs8hd_diode_2
XFILLER_76_3 vgnd vpwr scs8hd_decap_12
XPHY_290 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_483 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch/Q ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_310 vgnd vpwr scs8hd_fill_1
XFILLER_66_140 vgnd vpwr scs8hd_decap_6
XFILLER_54_302 vgnd vpwr scs8hd_decap_4
XFILLER_81_110 vgnd vpwr scs8hd_decap_12
XFILLER_54_335 vgnd vpwr scs8hd_fill_1
XFILLER_54_324 vgnd vpwr scs8hd_decap_4
XFILLER_39_387 vpwr vgnd scs8hd_fill_2
XFILLER_42_508 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch_SLEEPB _300_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_114 vgnd vpwr scs8hd_decap_3
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_57_184 vgnd vpwr scs8hd_decap_3
XFILLER_45_324 vpwr vgnd scs8hd_fill_2
XFILLER_72_154 vgnd vpwr scs8hd_decap_12
X_443_ _443_/HI _443_/LO vgnd vpwr scs8hd_conb_1
XFILLER_9_203 vpwr vgnd scs8hd_fill_2
X_374_ _200_/B _367_/B _374_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_236 vpwr vgnd scs8hd_fill_2
XFILLER_13_298 vpwr vgnd scs8hd_fill_2
XANTENNA__406__C _163_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_464 vgnd vpwr scs8hd_decap_12
XANTENNA__422__B _416_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_76_471 vgnd vpwr scs8hd_decap_12
XFILLER_63_121 vgnd vpwr scs8hd_fill_1
XFILLER_63_110 vgnd vpwr scs8hd_fill_1
XFILLER_36_313 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_165 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ _134_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__332__B _326_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch_SLEEPB _273_/Y vgnd vpwr scs8hd_diode_2
XFILLER_67_482 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_54_110 vpwr vgnd scs8hd_fill_2
XFILLER_27_313 vgnd vpwr scs8hd_fill_1
XFILLER_27_335 vgnd vpwr scs8hd_decap_8
XFILLER_39_184 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_187 vgnd vpwr scs8hd_decap_4
XFILLER_42_327 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch/Q ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_56 vgnd vpwr scs8hd_decap_12
XANTENNA__226__C _215_/X vgnd vpwr scs8hd_diode_2
XFILLER_10_224 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ _371_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_228 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
+ _410_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XANTENNA__242__B _243_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_401 vgnd vpwr scs8hd_decap_12
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XFILLER_49_86 vgnd vpwr scs8hd_decap_6
XFILLER_77_257 vgnd vpwr scs8hd_decap_12
XFILLER_1_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_45_110 vpwr vgnd scs8hd_fill_2
XFILLER_73_452 vgnd vpwr scs8hd_decap_12
XFILLER_65_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_132 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_81_62 vgnd vpwr scs8hd_decap_12
XFILLER_81_51 vgnd vpwr scs8hd_decap_8
XFILLER_60_168 vpwr vgnd scs8hd_fill_2
XANTENNA__417__B _416_/B vgnd vpwr scs8hd_diode_2
X_426_ _187_/B _424_/X _426_/Y vgnd vpwr scs8hd_nor2_4
X_357_ _276_/A _359_/B _357_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_288_ _279_/A _286_/B _288_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ _389_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_39_3 vgnd vpwr scs8hd_decap_12
XFILLER_36_121 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch_SLEEPB _245_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__327__B _326_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__343__A _280_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_235 vpwr vgnd scs8hd_fill_2
XFILLER_59_279 vpwr vgnd scs8hd_fill_2
XFILLER_27_132 vpwr vgnd scs8hd_fill_2
XFILLER_70_411 vpwr vgnd scs8hd_fill_2
XPHY_801 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
+ _422_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_349 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XPHY_845 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_834 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_823 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_812 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__237__B _243_/B vgnd vpwr scs8hd_diode_2
X_211_ _380_/A _166_/X _214_/B vgnd vpwr scs8hd_or2_4
X_142_ _142_/A _142_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__253__A address[8] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_65_238 vgnd vpwr scs8hd_decap_3
XFILLER_65_227 vpwr vgnd scs8hd_fill_2
XFILLER_18_110 vgnd vpwr scs8hd_decap_12
XFILLER_46_430 vgnd vpwr scs8hd_decap_4
XFILLER_73_260 vgnd vpwr scs8hd_decap_12
XFILLER_61_411 vpwr vgnd scs8hd_fill_2
XFILLER_61_400 vpwr vgnd scs8hd_fill_2
XFILLER_18_154 vpwr vgnd scs8hd_fill_2
XFILLER_33_113 vgnd vpwr scs8hd_decap_6
XFILLER_33_179 vpwr vgnd scs8hd_fill_2
X_409_ _173_/B _416_/B _409_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__163__A address[8] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch/Q
+ _236_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ _156_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__338__A _247_/A vgnd vpwr scs8hd_diode_2
XPHY_119 vgnd vpwr scs8hd_decap_3
XPHY_108 vgnd vpwr scs8hd_decap_3
XFILLER_12_308 vpwr vgnd scs8hd_fill_2
XFILLER_24_168 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_190 vgnd vpwr scs8hd_fill_1
XFILLER_20_363 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_4_507 vgnd vpwr scs8hd_decap_8
XFILLER_20_396 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_205 vgnd vpwr scs8hd_decap_3
XFILLER_47_227 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_32 vgnd vpwr scs8hd_decap_12
XFILLER_47_249 vgnd vpwr scs8hd_fill_1
XANTENNA__248__A _276_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_113 vgnd vpwr scs8hd_decap_3
XFILLER_43_433 vpwr vgnd scs8hd_fill_2
XFILLER_46_98 vpwr vgnd scs8hd_fill_2
XPHY_620 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ _155_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_653 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_642 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_631 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
XFILLER_30_127 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_686 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_675 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_664 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_341 vpwr vgnd scs8hd_fill_2
XFILLER_11_330 vpwr vgnd scs8hd_fill_2
XPHY_697 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_301 vpwr vgnd scs8hd_fill_2
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_345 vpwr vgnd scs8hd_fill_2
X_125_ address[1] _181_/B vgnd vpwr scs8hd_inv_8
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_78_385 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ right_width_0_height_0__pin_13_ vgnd vpwr scs8hd_inv_1
XFILLER_19_452 vgnd vpwr scs8hd_decap_12
XANTENNA__158__A _158_/A vgnd vpwr scs8hd_diode_2
XFILLER_46_293 vpwr vgnd scs8hd_fill_2
XFILLER_61_263 vpwr vgnd scs8hd_fill_2
XFILLER_21_127 vpwr vgnd scs8hd_fill_2
XANTENNA__308__D _272_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch_SLEEPB _225_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__340__B _343_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
+ clk ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff/QN
+ reset set vgnd vpwr scs8hd_dfbbp_1
XFILLER_25_400 vpwr vgnd scs8hd_fill_2
XFILLER_44_219 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_411 vgnd vpwr scs8hd_decap_4
XFILLER_25_422 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_68 vgnd vpwr scs8hd_decap_12
XFILLER_12_116 vgnd vpwr scs8hd_fill_1
XFILLER_8_109 vgnd vpwr scs8hd_decap_8
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_315 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_337 vgnd vpwr scs8hd_decap_3
XANTENNA__250__B _252_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_57_86 vgnd vpwr scs8hd_decap_12
XFILLER_35_208 vgnd vpwr scs8hd_fill_1
XFILLER_73_74 vgnd vpwr scs8hd_decap_12
XFILLER_31_469 vgnd vpwr scs8hd_decap_6
XPHY_450 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_461 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__425__B _424_/X vgnd vpwr scs8hd_diode_2
XPHY_472 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_483 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_494 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
XFILLER_7_197 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_300 vgnd vpwr scs8hd_decap_6
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_414 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _158_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__335__B _272_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_80 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__351__A _279_/A vgnd vpwr scs8hd_diode_2
XFILLER_69_193 vpwr vgnd scs8hd_fill_2
XFILLER_17_219 vpwr vgnd scs8hd_fill_2
XFILLER_72_325 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_425 vpwr vgnd scs8hd_fill_2
X_390_ _183_/B _391_/B _390_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_285 vgnd vpwr scs8hd_fill_1
XFILLER_9_407 vpwr vgnd scs8hd_fill_2
XANTENNA__245__B _252_/B vgnd vpwr scs8hd_diode_2
XFILLER_40_266 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch_SLEEPB _297_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_288 vpwr vgnd scs8hd_fill_2
XFILLER_4_145 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__261__A _279_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XFILLER_0_351 vgnd vpwr scs8hd_decap_3
XFILLER_0_362 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_48_322 vpwr vgnd scs8hd_fill_2
XFILLER_75_196 vgnd vpwr scs8hd_decap_12
XFILLER_63_358 vpwr vgnd scs8hd_fill_2
XFILLER_16_274 vgnd vpwr scs8hd_fill_1
XFILLER_71_391 vgnd vpwr scs8hd_decap_12
XFILLER_16_285 vpwr vgnd scs8hd_fill_2
XFILLER_16_296 vgnd vpwr scs8hd_decap_8
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_291 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ _186_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_69_3 vgnd vpwr scs8hd_decap_12
XFILLER_8_495 vgnd vpwr scs8hd_decap_12
XANTENNA__171__A address[0] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q
+ _358_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
+ _389_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ _131_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_66_163 vgnd vpwr scs8hd_decap_4
XFILLER_66_152 vgnd vpwr scs8hd_fill_1
XFILLER_39_355 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q
+ _323_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__346__A _274_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q
+ _288_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_77_428 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_108 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch_SLEEPB _270_/Y vgnd vpwr scs8hd_diode_2
XFILLER_45_303 vpwr vgnd scs8hd_fill_2
XFILLER_57_196 vpwr vgnd scs8hd_fill_2
XFILLER_54_32 vgnd vpwr scs8hd_decap_12
XFILLER_45_358 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q
+ _252_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_60_328 vgnd vpwr scs8hd_decap_8
X_442_ _442_/HI _442_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__256__A _274_/A vgnd vpwr scs8hd_diode_2
X_373_ _197_/B _367_/B _373_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__406__D _272_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_79_62 vgnd vpwr scs8hd_decap_12
XFILLER_79_51 vgnd vpwr scs8hd_decap_8
XFILLER_5_476 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _136_/Y vgnd vpwr scs8hd_diode_2
XFILLER_68_417 vgnd vpwr scs8hd_decap_12
XFILLER_68_406 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _436_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_483 vgnd vpwr scs8hd_decap_12
XFILLER_48_163 vgnd vpwr scs8hd_decap_3
XFILLER_63_144 vpwr vgnd scs8hd_fill_2
XFILLER_36_358 vgnd vpwr scs8hd_decap_4
XFILLER_63_188 vgnd vpwr scs8hd_fill_1
XFILLER_51_317 vpwr vgnd scs8hd_fill_2
XFILLER_51_306 vgnd vpwr scs8hd_decap_4
XFILLER_51_339 vgnd vpwr scs8hd_decap_3
XANTENNA__166__A address[6] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch/Q
+ _337_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch/Q
+ _302_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_59_428 vpwr vgnd scs8hd_fill_2
XFILLER_59_439 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_122 vpwr vgnd scs8hd_fill_2
XFILLER_27_358 vpwr vgnd scs8hd_fill_2
XFILLER_82_497 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch/Q
+ _267_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
+ reset vgnd vpwr scs8hd_diode_2
XFILLER_35_380 vpwr vgnd scs8hd_fill_2
XANTENNA__226__D _263_/D vgnd vpwr scs8hd_diode_2
XFILLER_24_68 vgnd vpwr scs8hd_decap_12
XFILLER_10_247 vpwr vgnd scs8hd_fill_2
XFILLER_10_269 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch_SLEEPB _242_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_2_413 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q
+ _231_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_457 vgnd vpwr scs8hd_fill_1
XFILLER_77_269 vgnd vpwr scs8hd_decap_12
XFILLER_58_450 vgnd vpwr scs8hd_decap_8
XFILLER_1_39 vgnd vpwr scs8hd_decap_12
XFILLER_18_314 vgnd vpwr scs8hd_decap_3
XFILLER_73_464 vgnd vpwr scs8hd_decap_12
XFILLER_65_86 vgnd vpwr scs8hd_decap_12
XFILLER_60_103 vgnd vpwr scs8hd_decap_3
XFILLER_33_306 vgnd vpwr scs8hd_decap_4
XFILLER_33_328 vpwr vgnd scs8hd_fill_2
XFILLER_60_136 vgnd vpwr scs8hd_decap_6
X_425_ _171_/X _424_/X _425_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_81_74 vgnd vpwr scs8hd_decap_12
X_356_ _247_/A _359_/B _356_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_394 vpwr vgnd scs8hd_fill_2
X_287_ _287_/A _286_/B _287_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_5_251 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch/Q ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch_SLEEPB _341_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_247 vgnd vpwr scs8hd_fill_1
XFILLER_56_409 vgnd vpwr scs8hd_decap_3
XFILLER_49_472 vpwr vgnd scs8hd_fill_2
XFILLER_49_461 vpwr vgnd scs8hd_fill_2
XFILLER_36_111 vgnd vpwr scs8hd_fill_1
XFILLER_24_306 vgnd vpwr scs8hd_decap_4
XFILLER_24_317 vpwr vgnd scs8hd_fill_2
XFILLER_51_114 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _139_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_380 vgnd vpwr scs8hd_fill_1
XFILLER_24_328 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__343__B _343_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_79 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _132_/Y vgnd vpwr scs8hd_diode_2
XFILLER_55_442 vpwr vgnd scs8hd_fill_2
XFILLER_82_261 vgnd vpwr scs8hd_decap_12
XFILLER_15_317 vgnd vpwr scs8hd_fill_1
XPHY_802 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_27_199 vgnd vpwr scs8hd_decap_8
XFILLER_42_136 vgnd vpwr scs8hd_decap_6
XPHY_835 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_824 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_813 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_350 vpwr vgnd scs8hd_fill_2
XFILLER_42_169 vpwr vgnd scs8hd_fill_2
XFILLER_11_501 vgnd vpwr scs8hd_decap_12
X_210_ _202_/A _210_/B _210_/Y vgnd vpwr scs8hd_nor2_4
X_141_ _141_/A _141_/Y vgnd vpwr scs8hd_inv_8
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__253__B _235_/B vgnd vpwr scs8hd_diode_2
XFILLER_51_99 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_232 vgnd vpwr scs8hd_fill_1
XFILLER_2_287 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_280 vgnd vpwr scs8hd_fill_1
XFILLER_18_122 vpwr vgnd scs8hd_fill_2
XFILLER_73_272 vgnd vpwr scs8hd_decap_12
XFILLER_61_456 vgnd vpwr scs8hd_decap_12
XFILLER_61_489 vgnd vpwr scs8hd_decap_12
X_408_ _170_/B _416_/B _408_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_372 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch_SLEEPB _314_/Y vgnd vpwr scs8hd_diode_2
X_339_ _276_/A _343_/B _339_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__163__B address[9] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_3 vgnd vpwr scs8hd_decap_12
XFILLER_69_501 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XFILLER_37_431 vpwr vgnd scs8hd_fill_2
XFILLER_49_291 vgnd vpwr scs8hd_decap_3
XFILLER_52_434 vpwr vgnd scs8hd_fill_2
XFILLER_37_486 vpwr vgnd scs8hd_fill_2
XANTENNA__338__B _343_/B vgnd vpwr scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_decap_3
XANTENNA__354__A _273_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _149_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
+ _375_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_431 vgnd vpwr scs8hd_decap_4
XFILLER_62_209 vgnd vpwr scs8hd_fill_1
XFILLER_46_44 vgnd vpwr scs8hd_decap_12
XANTENNA__248__B _252_/B vgnd vpwr scs8hd_diode_2
XFILLER_43_423 vpwr vgnd scs8hd_fill_2
XPHY_610 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_158 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_62_32 vgnd vpwr scs8hd_decap_12
XPHY_643 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_632 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_621 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_478 vpwr vgnd scs8hd_fill_2
XFILLER_43_489 vgnd vpwr scs8hd_decap_12
XPHY_687 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_676 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_665 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_654 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__264__A _273_/A vgnd vpwr scs8hd_diode_2
XPHY_698 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_397 vgnd vpwr scs8hd_fill_1
X_124_ address[0] _181_/C vgnd vpwr scs8hd_inv_8
XFILLER_7_335 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch/Q ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_80 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _150_/Y vgnd vpwr scs8hd_diode_2
XFILLER_66_515 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch_SLEEPB _287_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_53_209 vgnd vpwr scs8hd_decap_4
XFILLER_19_464 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_412 vgnd vpwr scs8hd_decap_3
XFILLER_34_445 vpwr vgnd scs8hd_fill_2
XFILLER_61_297 vpwr vgnd scs8hd_fill_2
XANTENNA__174__A _181_/C vgnd vpwr scs8hd_diode_2
XFILLER_14_191 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_72_507 vgnd vpwr scs8hd_decap_8
XANTENNA__349__A _231_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_294 vpwr vgnd scs8hd_fill_2
XFILLER_52_231 vgnd vpwr scs8hd_decap_4
XFILLER_25_456 vgnd vpwr scs8hd_decap_3
XFILLER_25_467 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_489 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_128 vpwr vgnd scs8hd_fill_2
XFILLER_20_150 vgnd vpwr scs8hd_decap_3
XFILLER_20_161 vgnd vpwr scs8hd_decap_6
XFILLER_20_183 vgnd vpwr scs8hd_decap_6
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_349 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_48_515 vgnd vpwr scs8hd_fill_1
XFILLER_75_367 vgnd vpwr scs8hd_decap_12
XFILLER_57_98 vgnd vpwr scs8hd_decap_3
XANTENNA__259__A _231_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
+ _368_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_456 vpwr vgnd scs8hd_fill_2
XFILLER_73_86 vgnd vpwr scs8hd_decap_12
XFILLER_31_426 vgnd vpwr scs8hd_fill_1
XFILLER_43_253 vgnd vpwr scs8hd_fill_1
XFILLER_43_286 vpwr vgnd scs8hd_fill_2
XFILLER_31_437 vpwr vgnd scs8hd_fill_2
XPHY_440 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_451 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_462 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_297 vpwr vgnd scs8hd_fill_2
XPHY_473 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_484 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_495 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_132 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _433_/HI
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_154 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_393 vgnd vpwr scs8hd_decap_6
XFILLER_66_323 vpwr vgnd scs8hd_fill_2
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__169__A _122_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_22_404 vgnd vpwr scs8hd_fill_1
XFILLER_22_426 vgnd vpwr scs8hd_decap_8
XFILLER_34_264 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch/Q ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_459 vgnd vpwr scs8hd_decap_12
XFILLER_34_286 vpwr vgnd scs8hd_fill_2
XANTENNA__335__C _163_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/Y _141_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__351__B _352_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch_SLEEPB _358_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_57_301 vpwr vgnd scs8hd_fill_2
XFILLER_57_323 vgnd vpwr scs8hd_fill_1
XFILLER_72_304 vgnd vpwr scs8hd_decap_6
XFILLER_57_367 vgnd vpwr scs8hd_decap_6
XFILLER_72_337 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ _160_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_264 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ _409_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_25_297 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch/Q ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q
+ _332_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_124 vgnd vpwr scs8hd_decap_4
XFILLER_4_113 vgnd vpwr scs8hd_decap_4
XANTENNA__261__B _262_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q
+ _297_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_63_337 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_389 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_234 vgnd vpwr scs8hd_decap_4
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q
+ _262_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_292 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_278 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
+ _414_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__171__B _181_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
+ reset vgnd vpwr scs8hd_diode_2
XFILLER_58_109 vgnd vpwr scs8hd_decap_8
XFILLER_39_367 vgnd vpwr scs8hd_decap_3
XFILLER_81_123 vgnd vpwr scs8hd_decap_12
XFILLER_66_197 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_348 vgnd vpwr scs8hd_decap_12
XFILLER_62_392 vgnd vpwr scs8hd_decap_4
XANTENNA__346__B _352_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_407 vgnd vpwr scs8hd_decap_8
XFILLER_22_267 vgnd vpwr scs8hd_decap_8
XFILLER_10_418 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_59 vpwr vgnd scs8hd_fill_2
XANTENNA__362__A _263_/A vgnd vpwr scs8hd_diode_2
XFILLER_57_142 vgnd vpwr scs8hd_decap_3
XFILLER_18_507 vgnd vpwr scs8hd_decap_8
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XFILLER_57_175 vpwr vgnd scs8hd_fill_2
XFILLER_57_164 vgnd vpwr scs8hd_decap_8
XFILLER_45_337 vpwr vgnd scs8hd_fill_2
X_441_ _441_/HI _441_/LO vgnd vpwr scs8hd_conb_1
XFILLER_54_44 vgnd vpwr scs8hd_decap_12
XFILLER_53_381 vgnd vpwr scs8hd_decap_4
XFILLER_13_201 vpwr vgnd scs8hd_fill_2
XFILLER_13_212 vpwr vgnd scs8hd_fill_2
X_372_ _194_/B _367_/B _372_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__256__B _262_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ _140_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_245 vgnd vpwr scs8hd_decap_3
XFILLER_70_32 vgnd vpwr scs8hd_decap_12
XANTENNA__272__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_79_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _131_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_160 vpwr vgnd scs8hd_fill_2
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
XFILLER_76_495 vgnd vpwr scs8hd_decap_12
XFILLER_36_304 vgnd vpwr scs8hd_decap_6
XFILLER_63_123 vgnd vpwr scs8hd_fill_1
XFILLER_36_337 vgnd vpwr scs8hd_fill_1
XFILLER_36_348 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__166__B address[7] vgnd vpwr scs8hd_diode_2
XFILLER_44_392 vgnd vpwr scs8hd_decap_3
XFILLER_81_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_271 vpwr vgnd scs8hd_fill_2
XANTENNA__182__A _122_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ _139_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_304 vgnd vpwr scs8hd_fill_1
XFILLER_39_164 vgnd vpwr scs8hd_decap_4
XFILLER_39_175 vpwr vgnd scs8hd_fill_2
XANTENNA__357__A _276_/A vgnd vpwr scs8hd_diode_2
XFILLER_50_351 vpwr vgnd scs8hd_fill_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XFILLER_2_425 vgnd vpwr scs8hd_decap_12
XFILLER_18_337 vpwr vgnd scs8hd_fill_2
XFILLER_18_348 vgnd vpwr scs8hd_decap_8
XFILLER_73_476 vgnd vpwr scs8hd_decap_12
XFILLER_65_98 vgnd vpwr scs8hd_decap_4
XANTENNA__267__A _276_/A vgnd vpwr scs8hd_diode_2
XFILLER_45_178 vgnd vpwr scs8hd_decap_3
X_424_ _380_/A _406_/X _424_/X vgnd vpwr scs8hd_or2_4
XFILLER_81_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_355_ _274_/A _359_/B _355_/Y vgnd vpwr scs8hd_nor2_4
X_286_ _231_/A _286_/B _286_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_296 vpwr vgnd scs8hd_fill_2
XFILLER_5_285 vpwr vgnd scs8hd_fill_2
XFILLER_68_204 vpwr vgnd scs8hd_fill_2
XFILLER_68_215 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_68_259 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__177__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_351 vpwr vgnd scs8hd_fill_2
XFILLER_32_362 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_259 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_55_476 vgnd vpwr scs8hd_decap_12
XFILLER_82_273 vgnd vpwr scs8hd_decap_6
XFILLER_27_178 vgnd vpwr scs8hd_decap_3
XPHY_836 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_825 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_814 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_803 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_457 vgnd vpwr scs8hd_fill_1
XFILLER_11_513 vgnd vpwr scs8hd_decap_3
XFILLER_23_362 vpwr vgnd scs8hd_fill_2
XFILLER_23_384 vgnd vpwr scs8hd_decap_3
X_140_ _140_/A _140_/Y vgnd vpwr scs8hd_inv_8
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_211 vgnd vpwr scs8hd_fill_1
XFILLER_2_244 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
+ clk vgnd vpwr scs8hd_diode_2
XFILLER_58_292 vgnd vpwr scs8hd_decap_12
XFILLER_73_284 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_468 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_407_ address[4] _406_/X _416_/B vgnd vpwr scs8hd_or2_4
XFILLER_25_90 vpwr vgnd scs8hd_fill_2
XPHY_90 vgnd vpwr scs8hd_decap_3
X_338_ _247_/A _343_/B _338_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_170 vgnd vpwr scs8hd_decap_3
X_269_ _287_/A _269_/B _269_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _440_/HI
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_3 vgnd vpwr scs8hd_decap_12
XFILLER_69_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_37_421 vgnd vpwr scs8hd_decap_6
XFILLER_37_443 vgnd vpwr scs8hd_decap_4
XFILLER_52_402 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_262 vpwr vgnd scs8hd_fill_2
XFILLER_52_413 vgnd vpwr scs8hd_decap_12
XFILLER_52_468 vpwr vgnd scs8hd_fill_2
XFILLER_52_446 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_137 vgnd vpwr scs8hd_decap_12
XFILLER_20_310 vgnd vpwr scs8hd_decap_4
XANTENNA__354__B _359_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_59 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__370__A _189_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
+ _206_/Y vgnd vpwr scs8hd_diode_2
XFILLER_55_240 vpwr vgnd scs8hd_fill_2
XFILLER_28_454 vpwr vgnd scs8hd_fill_2
XFILLER_46_56 vgnd vpwr scs8hd_decap_12
XFILLER_55_284 vpwr vgnd scs8hd_fill_2
XFILLER_55_273 vgnd vpwr scs8hd_decap_4
XFILLER_70_243 vgnd vpwr scs8hd_decap_12
XFILLER_70_232 vgnd vpwr scs8hd_decap_8
XPHY_611 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_600 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_446 vpwr vgnd scs8hd_fill_2
XFILLER_43_457 vpwr vgnd scs8hd_fill_2
XFILLER_70_276 vgnd vpwr scs8hd_decap_4
XFILLER_62_44 vgnd vpwr scs8hd_decap_12
XPHY_644 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_633 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_622 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_677 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_666 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_655 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_699 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_688 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__264__B _269_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_376 vpwr vgnd scs8hd_fill_2
X_123_ address[2] _178_/A vgnd vpwr scs8hd_inv_8
XFILLER_7_39 vgnd vpwr scs8hd_decap_12
XFILLER_7_358 vpwr vgnd scs8hd_fill_2
XANTENNA__280__A _280_/A vgnd vpwr scs8hd_diode_2
XFILLER_78_398 vgnd vpwr scs8hd_decap_12
XFILLER_19_476 vgnd vpwr scs8hd_decap_12
XFILLER_34_424 vgnd vpwr scs8hd_decap_12
XFILLER_61_221 vpwr vgnd scs8hd_fill_2
XFILLER_34_457 vgnd vpwr scs8hd_fill_1
XFILLER_34_468 vpwr vgnd scs8hd_fill_2
XFILLER_21_107 vpwr vgnd scs8hd_fill_2
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_181 vgnd vpwr scs8hd_decap_3
XANTENNA__174__B address[1] vgnd vpwr scs8hd_diode_2
XANTENNA__190__A address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_69_310 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_69_365 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA__349__B _352_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ _157_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_276 vgnd vpwr scs8hd_decap_6
XFILLER_52_265 vpwr vgnd scs8hd_fill_2
XANTENNA__365__A _173_/B vgnd vpwr scs8hd_diode_2
XFILLER_40_427 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_328 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
+ reset vgnd vpwr scs8hd_diode_2
XFILLER_75_379 vgnd vpwr scs8hd_decap_12
XANTENNA__259__B _262_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_424 vgnd vpwr scs8hd_decap_12
XFILLER_28_284 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_43_232 vpwr vgnd scs8hd_fill_2
XFILLER_73_98 vgnd vpwr scs8hd_decap_12
XANTENNA__275__A _247_/A vgnd vpwr scs8hd_diode_2
XPHY_430 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_441 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_452 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_463 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_474 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_485 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_496 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_184 vpwr vgnd scs8hd_fill_2
XFILLER_22_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_335 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_66_368 vgnd vpwr scs8hd_decap_3
XANTENNA__169__B _273_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_240 vpwr vgnd scs8hd_fill_2
XFILLER_19_262 vpwr vgnd scs8hd_fill_2
XANTENNA__185__A _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_254 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__335__D _263_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_93 vgnd vpwr scs8hd_decap_3
XFILLER_69_162 vpwr vgnd scs8hd_fill_2
XFILLER_69_184 vpwr vgnd scs8hd_fill_2
XFILLER_65_390 vgnd vpwr scs8hd_decap_4
XFILLER_25_221 vgnd vpwr scs8hd_decap_4
XFILLER_40_213 vgnd vpwr scs8hd_fill_1
XFILLER_40_224 vgnd vpwr scs8hd_decap_3
XFILLER_40_235 vgnd vpwr scs8hd_decap_4
XFILLER_40_279 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch/Q ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_320 vpwr vgnd scs8hd_fill_2
XFILLER_75_110 vgnd vpwr scs8hd_decap_12
XFILLER_0_386 vgnd vpwr scs8hd_decap_4
XFILLER_0_397 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_346 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_471 vgnd vpwr scs8hd_decap_12
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_431 vgnd vpwr scs8hd_decap_12
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_293 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_302 vgnd vpwr scs8hd_decap_3
XFILLER_39_324 vgnd vpwr scs8hd_decap_4
XFILLER_39_335 vpwr vgnd scs8hd_fill_2
XFILLER_39_379 vpwr vgnd scs8hd_fill_2
XFILLER_81_135 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_224 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_290 vgnd vpwr scs8hd_decap_12
XANTENNA__362__B address[7] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ _383_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_57_132 vgnd vpwr scs8hd_decap_4
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
X_440_ _440_/HI _440_/LO vgnd vpwr scs8hd_conb_1
XFILLER_54_56 vgnd vpwr scs8hd_decap_12
X_371_ _371_/A _367_/B _371_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_80_190 vgnd vpwr scs8hd_decap_12
XFILLER_13_235 vpwr vgnd scs8hd_fill_2
XFILLER_70_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_217 vpwr vgnd scs8hd_fill_2
XANTENNA__272__B _272_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_489 vgnd vpwr scs8hd_decap_12
XFILLER_79_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _141_/Y vgnd vpwr scs8hd_diode_2
XFILLER_48_187 vgnd vpwr scs8hd_decap_4
XANTENNA__166__C _163_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _437_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_360 vgnd vpwr scs8hd_decap_6
XFILLER_74_3 vgnd vpwr scs8hd_decap_12
XFILLER_12_290 vpwr vgnd scs8hd_fill_2
XANTENNA__182__B _231_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_59_419 vpwr vgnd scs8hd_fill_2
XFILLER_39_132 vpwr vgnd scs8hd_fill_2
XFILLER_39_143 vpwr vgnd scs8hd_fill_2
XFILLER_27_316 vpwr vgnd scs8hd_fill_2
XFILLER_82_466 vgnd vpwr scs8hd_decap_12
XFILLER_54_168 vpwr vgnd scs8hd_fill_2
XANTENNA__357__B _359_/B vgnd vpwr scs8hd_diode_2
XFILLER_42_308 vgnd vpwr scs8hd_decap_3
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_396 vgnd vpwr scs8hd_fill_1
XANTENNA__373__A _197_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch/Q ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _132_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_437 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ _204_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_459 vgnd vpwr scs8hd_decap_12
XFILLER_58_463 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ _148_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__267__B _269_/B vgnd vpwr scs8hd_diode_2
X_423_ _210_/B _416_/B _423_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_26_371 vpwr vgnd scs8hd_fill_2
XFILLER_60_149 vgnd vpwr scs8hd_decap_4
XFILLER_26_393 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_341 vpwr vgnd scs8hd_fill_2
X_354_ _273_/A _359_/B _354_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_352 vgnd vpwr scs8hd_decap_4
XFILLER_41_363 vgnd vpwr scs8hd_fill_1
XFILLER_81_98 vgnd vpwr scs8hd_decap_12
XANTENNA__283__A _274_/A vgnd vpwr scs8hd_diode_2
X_285_ _276_/A _286_/B _285_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_242 vpwr vgnd scs8hd_fill_2
XFILLER_30_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_441 vpwr vgnd scs8hd_fill_2
XFILLER_64_433 vpwr vgnd scs8hd_fill_2
XANTENNA__177__B address[1] vgnd vpwr scs8hd_diode_2
XFILLER_36_146 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_51_149 vpwr vgnd scs8hd_fill_2
XFILLER_32_341 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ _147_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_32_374 vpwr vgnd scs8hd_fill_2
XANTENNA__193__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
+ _183_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XFILLER_55_422 vpwr vgnd scs8hd_fill_2
XANTENNA__368__A _183_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _159_/Y vgnd vpwr scs8hd_diode_2
XFILLER_82_230 vgnd vpwr scs8hd_decap_12
XFILLER_55_455 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_157 vpwr vgnd scs8hd_fill_2
XPHY_826 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_815 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_804 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_42_149 vpwr vgnd scs8hd_fill_2
XPHY_837 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_50_171 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ top_width_0_height_0__pin_12_ vgnd vpwr scs8hd_inv_1
XFILLER_23_396 vgnd vpwr scs8hd_decap_6
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_267 vpwr vgnd scs8hd_fill_2
XFILLER_76_32 vgnd vpwr scs8hd_decap_12
XANTENNA__278__A _287_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_135 vpwr vgnd scs8hd_fill_2
XFILLER_73_296 vgnd vpwr scs8hd_decap_8
XFILLER_33_127 vpwr vgnd scs8hd_fill_2
XFILLER_33_138 vpwr vgnd scs8hd_fill_2
XFILLER_33_149 vpwr vgnd scs8hd_fill_2
X_406_ address[6] address[7] _163_/X _272_/D _406_/X vgnd vpwr scs8hd_or4_4
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _144_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_41_193 vpwr vgnd scs8hd_fill_2
X_337_ _274_/A _343_/B _337_/Y vgnd vpwr scs8hd_nor2_4
X_268_ _231_/A _269_/B _268_/Y vgnd vpwr scs8hd_nor2_4
X_199_ address[3] _247_/A _200_/B vgnd vpwr scs8hd_or2_4
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__188__A _122_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_37_466 vgnd vpwr scs8hd_decap_12
XFILLER_37_455 vgnd vpwr scs8hd_decap_4
XFILLER_64_274 vgnd vpwr scs8hd_fill_1
XFILLER_24_116 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_149 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ _420_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
+ reset vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch/Q ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_32_171 vgnd vpwr scs8hd_fill_1
XFILLER_32_193 vpwr vgnd scs8hd_fill_2
XFILLER_20_388 vgnd vpwr scs8hd_decap_8
XFILLER_21_27 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch_SLEEPB _259_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__370__B _367_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_219 vpwr vgnd scs8hd_fill_2
XFILLER_46_68 vgnd vpwr scs8hd_decap_12
XFILLER_43_403 vgnd vpwr scs8hd_decap_4
XPHY_601 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_634 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_623 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_612 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_108 vpwr vgnd scs8hd_fill_2
XPHY_678 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_62_56 vgnd vpwr scs8hd_decap_12
XPHY_667 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_656 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_645 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch/Q
+ _282_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_51_480 vpwr vgnd scs8hd_fill_2
XFILLER_11_311 vpwr vgnd scs8hd_fill_2
XFILLER_23_160 vpwr vgnd scs8hd_fill_2
XFILLER_23_171 vpwr vgnd scs8hd_fill_2
XPHY_689 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_315 vpwr vgnd scs8hd_fill_2
X_122_ address[3] _122_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__280__B _280_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_93 vpwr vgnd scs8hd_fill_2
XFILLER_78_300 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch/Q
+ _246_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ _427_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_46_263 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _155_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_160 vpwr vgnd scs8hd_fill_2
XANTENNA__190__B _178_/B vgnd vpwr scs8hd_diode_2
XFILLER_69_333 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_69_399 vgnd vpwr scs8hd_decap_4
XFILLER_29_219 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch_SLEEPB _231_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_252 vpwr vgnd scs8hd_fill_2
XFILLER_52_244 vgnd vpwr scs8hd_decap_4
XFILLER_52_211 vgnd vpwr scs8hd_decap_3
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
XFILLER_52_255 vgnd vpwr scs8hd_fill_1
XFILLER_12_108 vpwr vgnd scs8hd_fill_2
XANTENNA__365__B _367_/B vgnd vpwr scs8hd_diode_2
XFILLER_52_299 vgnd vpwr scs8hd_decap_4
XFILLER_40_439 vpwr vgnd scs8hd_fill_2
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
+ _396_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__381__A _171_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_230 vgnd vpwr scs8hd_decap_8
XFILLER_16_436 vgnd vpwr scs8hd_decap_12
XANTENNA__275__B _280_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_406 vpwr vgnd scs8hd_fill_2
XPHY_420 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_428 vpwr vgnd scs8hd_fill_2
XPHY_431 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_442 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_453 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_141 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch_SLEEPB _330_/Y vgnd vpwr scs8hd_diode_2
XPHY_464 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_475 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_486 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_174 vpwr vgnd scs8hd_fill_2
XPHY_497 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__291__A _273_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _434_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_141 vgnd vpwr scs8hd_decap_12
XFILLER_81_306 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ _398_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_285 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch/Q ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _444_/HI
+ vgnd vpwr scs8hd_diode_2
XANTENNA__185__B _287_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_299 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_69_141 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_358 vgnd vpwr scs8hd_decap_8
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_59 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__376__A _204_/B vgnd vpwr scs8hd_diode_2
XFILLER_80_361 vgnd vpwr scs8hd_decap_12
XFILLER_13_406 vgnd vpwr scs8hd_decap_4
XFILLER_13_417 vgnd vpwr scs8hd_decap_8
XFILLER_13_428 vgnd vpwr scs8hd_decap_12
XFILLER_25_277 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_258 vpwr vgnd scs8hd_fill_2
XFILLER_40_269 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_159 vpwr vgnd scs8hd_fill_2
XFILLER_68_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch_SLEEPB _303_/Y vgnd vpwr scs8hd_diode_2
XFILLER_48_303 vgnd vpwr scs8hd_decap_3
XFILLER_48_358 vpwr vgnd scs8hd_fill_2
XFILLER_63_306 vgnd vpwr scs8hd_decap_3
XANTENNA__286__A _231_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_222 vgnd vpwr scs8hd_decap_4
XFILLER_17_92 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_225 vpwr vgnd scs8hd_fill_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_294 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_483 vgnd vpwr scs8hd_decap_12
XFILLER_8_443 vgnd vpwr scs8hd_decap_12
XFILLER_66_111 vgnd vpwr scs8hd_fill_1
XFILLER_54_328 vgnd vpwr scs8hd_fill_1
XFILLER_81_147 vgnd vpwr scs8hd_decap_12
XANTENNA__196__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_47_380 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_247 vgnd vpwr scs8hd_decap_3
XFILLER_13_39 vgnd vpwr scs8hd_decap_12
XFILLER_30_280 vgnd vpwr scs8hd_fill_1
XANTENNA__362__C _163_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_45_306 vpwr vgnd scs8hd_fill_2
XFILLER_45_328 vgnd vpwr scs8hd_decap_4
XFILLER_54_68 vgnd vpwr scs8hd_decap_12
X_370_ _189_/B _367_/B _370_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_501 vgnd vpwr scs8hd_decap_12
XFILLER_9_207 vgnd vpwr scs8hd_decap_4
XFILLER_13_269 vgnd vpwr scs8hd_fill_1
XFILLER_70_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch_SLEEPB _276_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__272__C _272_/C vgnd vpwr scs8hd_diode_2
XFILLER_5_402 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ _376_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_79_98 vgnd vpwr scs8hd_decap_12
XFILLER_0_151 vgnd vpwr scs8hd_decap_4
XFILLER_0_140 vpwr vgnd scs8hd_fill_2
XFILLER_36_317 vgnd vpwr scs8hd_decap_8
XFILLER_63_114 vgnd vpwr scs8hd_decap_4
XFILLER_28_80 vgnd vpwr scs8hd_decap_12
XFILLER_36_328 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
+ _413_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__166__D _263_/D vgnd vpwr scs8hd_diode_2
XFILLER_67_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_5_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_95 vpwr vgnd scs8hd_fill_2
XFILLER_67_442 vpwr vgnd scs8hd_fill_2
XFILLER_67_431 vpwr vgnd scs8hd_fill_2
XFILLER_67_420 vgnd vpwr scs8hd_decap_6
XFILLER_39_111 vpwr vgnd scs8hd_fill_2
XFILLER_54_114 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_188 vpwr vgnd scs8hd_fill_2
XFILLER_82_478 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_501 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_206 vgnd vpwr scs8hd_decap_8
XFILLER_10_228 vgnd vpwr scs8hd_decap_6
XANTENNA__373__B _367_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_2_449 vgnd vpwr scs8hd_decap_8
XFILLER_58_475 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch_SLEEPB _248_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_328 vgnd vpwr scs8hd_decap_8
XFILLER_45_114 vgnd vpwr scs8hd_decap_6
XFILLER_45_136 vpwr vgnd scs8hd_fill_2
XFILLER_73_489 vgnd vpwr scs8hd_decap_12
XFILLER_60_117 vpwr vgnd scs8hd_fill_2
X_422_ _208_/B _416_/B _422_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_26_361 vgnd vpwr scs8hd_decap_8
X_353_ address[6] _272_/B _163_/X _263_/D _359_/B vgnd vpwr scs8hd_or4_4
XANTENNA__283__B _286_/B vgnd vpwr scs8hd_diode_2
X_284_ _247_/A _286_/B _284_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_93 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ _141_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch/Q
+ _347_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_221 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch/Q
+ _312_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_125 vgnd vpwr scs8hd_decap_4
XFILLER_51_128 vpwr vgnd scs8hd_fill_2
XFILLER_17_383 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch_SLEEPB _347_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_515 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__193__B _273_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q
+ _277_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
+ _429_/HI ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_59_217 vgnd vpwr scs8hd_decap_3
XFILLER_59_239 vgnd vpwr scs8hd_decap_3
XFILLER_19_27 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q
+ _241_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_55_401 vpwr vgnd scs8hd_fill_2
XFILLER_67_294 vgnd vpwr scs8hd_fill_1
XANTENNA__368__B _367_/B vgnd vpwr scs8hd_diode_2
XFILLER_82_242 vgnd vpwr scs8hd_decap_6
XFILLER_27_136 vpwr vgnd scs8hd_fill_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_70_415 vgnd vpwr scs8hd_decap_12
XFILLER_55_489 vgnd vpwr scs8hd_decap_12
XFILLER_15_309 vpwr vgnd scs8hd_fill_2
XPHY_827 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_816 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_805 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_459 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_331 vpwr vgnd scs8hd_fill_2
XANTENNA__384__A _263_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_838 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_50_183 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _147_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_224 vpwr vgnd scs8hd_fill_2
XFILLER_78_515 vgnd vpwr scs8hd_fill_1
XFILLER_2_279 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ _156_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_76_44 vgnd vpwr scs8hd_decap_12
XFILLER_58_250 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__278__B _280_/B vgnd vpwr scs8hd_diode_2
XFILLER_46_434 vgnd vpwr scs8hd_fill_1
XFILLER_73_231 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_147 vgnd vpwr scs8hd_decap_3
XFILLER_18_158 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_61_415 vgnd vpwr scs8hd_decap_4
XFILLER_26_180 vgnd vpwr scs8hd_decap_4
X_405_ _178_/B _402_/X _405_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__294__A _276_/A vgnd vpwr scs8hd_diode_2
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_decap_3
X_336_ _273_/A _343_/B _336_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch/Q
+ _291_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_267_ _276_/A _269_/B _267_/Y vgnd vpwr scs8hd_nor2_4
X_198_ _178_/A _181_/C address[1] _247_/A vgnd vpwr scs8hd_or3_4
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch_SLEEPB _320_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _441_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_250 vpwr vgnd scs8hd_fill_2
XANTENNA__188__B _279_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch/Q
+ _256_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_478 vgnd vpwr scs8hd_decap_8
XFILLER_37_489 vgnd vpwr scs8hd_decap_12
XFILLER_17_180 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/Y _161_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch/Q
+ _220_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_390 vpwr vgnd scs8hd_fill_2
XFILLER_21_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__379__A _210_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_412 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_297 vpwr vgnd scs8hd_fill_2
XPHY_602 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_139 vpwr vgnd scs8hd_fill_2
XFILLER_70_267 vgnd vpwr scs8hd_decap_8
XPHY_635 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_624 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_613 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_289 vgnd vpwr scs8hd_decap_12
XFILLER_62_68 vgnd vpwr scs8hd_decap_12
XPHY_668 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_657 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_646 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_492 vpwr vgnd scs8hd_fill_2
XFILLER_11_301 vpwr vgnd scs8hd_fill_2
XPHY_679 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_345 vpwr vgnd scs8hd_fill_2
XFILLER_11_334 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_11_83 vgnd vpwr scs8hd_decap_4
XFILLER_78_312 vgnd vpwr scs8hd_decap_12
XFILLER_66_507 vgnd vpwr scs8hd_decap_8
XANTENNA__289__A _280_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_423 vpwr vgnd scs8hd_fill_2
XFILLER_19_489 vgnd vpwr scs8hd_decap_12
XFILLER_61_234 vgnd vpwr scs8hd_decap_4
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XFILLER_46_297 vgnd vpwr scs8hd_decap_4
XFILLER_61_267 vpwr vgnd scs8hd_fill_2
XFILLER_61_245 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_319_ _274_/A _325_/B _319_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_69_301 vpwr vgnd scs8hd_fill_2
XFILLER_69_323 vpwr vgnd scs8hd_fill_2
XFILLER_69_367 vpwr vgnd scs8hd_fill_2
XFILLER_69_356 vgnd vpwr scs8hd_fill_1
XANTENNA__199__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_37_231 vgnd vpwr scs8hd_decap_6
XFILLER_25_415 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_142 vgnd vpwr scs8hd_decap_6
XANTENNA__381__B _380_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_319 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _156_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_448 vgnd vpwr scs8hd_decap_8
XFILLER_16_459 vgnd vpwr scs8hd_decap_12
XPHY_410 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_245 vpwr vgnd scs8hd_fill_2
XFILLER_43_256 vpwr vgnd scs8hd_fill_2
XPHY_421 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_432 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_443 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _138_/Y vgnd vpwr scs8hd_diode_2
XPHY_454 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_465 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_476 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_153 vpwr vgnd scs8hd_fill_2
XPHY_487 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_498 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__291__B _295_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
XFILLER_22_93 vpwr vgnd scs8hd_fill_2
XFILLER_3_363 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_337 vgnd vpwr scs8hd_decap_3
XFILLER_81_318 vgnd vpwr scs8hd_decap_12
XFILLER_19_253 vpwr vgnd scs8hd_fill_2
XFILLER_47_90 vgnd vpwr scs8hd_fill_1
XFILLER_19_297 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ _132_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_462 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch/Q ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_69_131 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_175 vpwr vgnd scs8hd_fill_2
XFILLER_57_315 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_57_337 vpwr vgnd scs8hd_fill_2
XFILLER_27_27 vgnd vpwr scs8hd_decap_12
XANTENNA__376__B _367_/B vgnd vpwr scs8hd_diode_2
XFILLER_25_201 vgnd vpwr scs8hd_fill_1
XFILLER_25_245 vgnd vpwr scs8hd_decap_4
XFILLER_80_373 vgnd vpwr scs8hd_decap_12
XFILLER_43_15 vgnd vpwr scs8hd_decap_12
XFILLER_43_59 vpwr vgnd scs8hd_fill_2
XANTENNA__392__A _189_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_149 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ _131_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch/Q ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_300 vgnd vpwr scs8hd_decap_4
XFILLER_68_56 vgnd vpwr scs8hd_decap_12
XFILLER_0_333 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_0_366 vgnd vpwr scs8hd_decap_4
XFILLER_48_326 vpwr vgnd scs8hd_fill_2
XFILLER_75_123 vgnd vpwr scs8hd_decap_12
XFILLER_48_337 vpwr vgnd scs8hd_fill_2
XANTENNA__286__B _286_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_212 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_245 vpwr vgnd scs8hd_fill_2
XFILLER_16_289 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_295 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_495 vgnd vpwr scs8hd_decap_12
XFILLER_8_455 vgnd vpwr scs8hd_decap_3
XFILLER_33_92 vgnd vpwr scs8hd_fill_1
XFILLER_79_440 vgnd vpwr scs8hd_decap_12
XFILLER_3_193 vpwr vgnd scs8hd_fill_2
XFILLER_66_123 vpwr vgnd scs8hd_fill_2
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_39_348 vgnd vpwr scs8hd_decap_4
XFILLER_39_359 vgnd vpwr scs8hd_decap_4
XFILLER_66_167 vgnd vpwr scs8hd_fill_1
XANTENNA__196__B _274_/A vgnd vpwr scs8hd_diode_2
XFILLER_81_159 vgnd vpwr scs8hd_decap_12
XFILLER_62_373 vgnd vpwr scs8hd_fill_1
XFILLER_50_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _134_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__362__D _272_/D vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q
+ _342_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_119 vgnd vpwr scs8hd_decap_3
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_57_112 vgnd vpwr scs8hd_decap_4
XFILLER_57_156 vpwr vgnd scs8hd_fill_2
XANTENNA__387__A _173_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q
+ _307_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_53_362 vpwr vgnd scs8hd_fill_2
XFILLER_41_513 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_259 vpwr vgnd scs8hd_fill_2
XFILLER_70_68 vgnd vpwr scs8hd_decap_12
XANTENNA__272__D _272_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ _368_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_76_410 vgnd vpwr scs8hd_decap_12
XANTENNA__297__A _279_/A vgnd vpwr scs8hd_diode_2
XFILLER_48_145 vgnd vpwr scs8hd_decap_6
XFILLER_29_370 vpwr vgnd scs8hd_fill_2
XFILLER_63_148 vpwr vgnd scs8hd_fill_2
XFILLER_44_351 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch/Q ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_44_80 vgnd vpwr scs8hd_decap_12
XFILLER_8_263 vgnd vpwr scs8hd_decap_8
XFILLER_8_252 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _438_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_285 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
XFILLER_79_281 vgnd vpwr scs8hd_decap_12
XFILLER_82_435 vgnd vpwr scs8hd_decap_12
XFILLER_54_126 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_513 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/Y _133_/A vgnd vpwr scs8hd_buf_1
XFILLER_35_384 vpwr vgnd scs8hd_fill_2
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_432 vgnd vpwr scs8hd_decap_4
XFILLER_58_421 vgnd vpwr scs8hd_decap_6
XFILLER_58_487 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_159 vpwr vgnd scs8hd_fill_2
X_421_ _377_/A _416_/B _421_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_26_351 vgnd vpwr scs8hd_fill_1
XFILLER_53_192 vpwr vgnd scs8hd_fill_2
X_352_ _280_/A _352_/B _352_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_376 vpwr vgnd scs8hd_fill_2
X_283_ _274_/A _286_/B _283_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_387 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _152_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_266 vpwr vgnd scs8hd_fill_2
XFILLER_30_93 vgnd vpwr scs8hd_decap_8
XFILLER_76_251 vgnd vpwr scs8hd_decap_12
XFILLER_49_476 vpwr vgnd scs8hd_fill_2
XFILLER_49_454 vgnd vpwr scs8hd_decap_4
XFILLER_51_118 vpwr vgnd scs8hd_fill_2
XFILLER_17_351 vgnd vpwr scs8hd_decap_4
XFILLER_17_362 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_192 vpwr vgnd scs8hd_fill_2
XFILLER_32_398 vpwr vgnd scs8hd_fill_2
XFILLER_67_240 vpwr vgnd scs8hd_fill_2
XFILLER_19_39 vgnd vpwr scs8hd_decap_12
XFILLER_67_284 vpwr vgnd scs8hd_fill_2
XFILLER_67_273 vpwr vgnd scs8hd_fill_2
XFILLER_27_115 vgnd vpwr scs8hd_decap_4
XFILLER_55_446 vgnd vpwr scs8hd_decap_4
XFILLER_70_427 vgnd vpwr scs8hd_decap_12
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XPHY_817 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_806 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_35_181 vpwr vgnd scs8hd_fill_2
XPHY_839 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_828 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_50_140 vgnd vpwr scs8hd_decap_8
XFILLER_23_354 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__384__B address[7] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_51_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_376 vpwr vgnd scs8hd_fill_2
XFILLER_51_59 vpwr vgnd scs8hd_fill_2
XFILLER_2_203 vgnd vpwr scs8hd_decap_8
XFILLER_76_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_46_413 vgnd vpwr scs8hd_decap_4
XFILLER_73_243 vgnd vpwr scs8hd_fill_1
XFILLER_46_446 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch/Q ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ _149_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_404_ _187_/B _402_/X _404_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__294__B _295_/B vgnd vpwr scs8hd_diode_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_82 vgnd vpwr scs8hd_decap_3
XFILLER_41_140 vpwr vgnd scs8hd_fill_2
X_335_ _263_/A _272_/B _163_/X _263_/D _343_/B vgnd vpwr scs8hd_or4_4
XFILLER_14_376 vgnd vpwr scs8hd_decap_4
XPHY_93 vgnd vpwr scs8hd_decap_3
X_266_ _247_/A _269_/B _266_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
+ _378_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
X_197_ _202_/A _197_/B _197_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _155_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_280 vpwr vgnd scs8hd_fill_2
XFILLER_37_402 vpwr vgnd scs8hd_fill_2
XFILLER_37_413 vpwr vgnd scs8hd_fill_2
XFILLER_64_243 vgnd vpwr scs8hd_decap_6
XFILLER_37_435 vpwr vgnd scs8hd_fill_2
XFILLER_64_276 vpwr vgnd scs8hd_fill_2
XFILLER_52_438 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_60_471 vgnd vpwr scs8hd_decap_12
XFILLER_32_151 vpwr vgnd scs8hd_fill_2
XFILLER_20_335 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _148_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__379__B _367_/B vgnd vpwr scs8hd_diode_2
XFILLER_46_15 vgnd vpwr scs8hd_decap_12
XFILLER_55_232 vpwr vgnd scs8hd_fill_2
XFILLER_55_210 vgnd vpwr scs8hd_decap_3
XFILLER_28_446 vgnd vpwr scs8hd_decap_8
XFILLER_55_254 vpwr vgnd scs8hd_fill_2
XANTENNA__395__A _197_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_468 vgnd vpwr scs8hd_decap_8
XFILLER_28_479 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
XFILLER_70_257 vgnd vpwr scs8hd_fill_1
XPHY_625 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_614 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_603 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_140 vgnd vpwr scs8hd_decap_4
XPHY_669 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_658 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_647 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_636 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_184 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_339 vgnd vpwr scs8hd_decap_4
XFILLER_11_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_501 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_62 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_324 vgnd vpwr scs8hd_decap_12
XANTENNA__289__B _286_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_402 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_46_243 vpwr vgnd scs8hd_fill_2
XFILLER_46_276 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_449 vgnd vpwr scs8hd_decap_8
XFILLER_14_173 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_80 vgnd vpwr scs8hd_decap_12
X_318_ _273_/A _325_/B _318_/Y vgnd vpwr scs8hd_nor2_4
X_249_ _231_/A _252_/B _249_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _145_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_350 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_372 vgnd vpwr scs8hd_decap_3
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XANTENNA__199__B _247_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_243 vgnd vpwr scs8hd_fill_1
XFILLER_37_265 vpwr vgnd scs8hd_fill_2
XFILLER_37_276 vpwr vgnd scs8hd_fill_2
XFILLER_37_298 vgnd vpwr scs8hd_decap_4
XFILLER_33_460 vpwr vgnd scs8hd_fill_2
XFILLER_33_471 vgnd vpwr scs8hd_decap_12
XFILLER_20_121 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_515 vgnd vpwr scs8hd_fill_1
XFILLER_28_210 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_265 vpwr vgnd scs8hd_fill_2
XFILLER_28_276 vgnd vpwr scs8hd_decap_4
XFILLER_43_202 vpwr vgnd scs8hd_fill_2
XPHY_400 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_411 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_422 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_419 vgnd vpwr scs8hd_decap_4
XPHY_433 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_444 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_290 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ _189_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_455 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_466 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_477 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch_SLEEPB _361_/Y vgnd vpwr scs8hd_diode_2
XPHY_488 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_499 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_158 vpwr vgnd scs8hd_fill_2
XFILLER_3_353 vgnd vpwr scs8hd_decap_4
XFILLER_78_154 vgnd vpwr scs8hd_decap_12
XFILLER_66_327 vgnd vpwr scs8hd_decap_8
XFILLER_66_349 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _435_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_224 vpwr vgnd scs8hd_fill_2
XFILLER_34_246 vpwr vgnd scs8hd_fill_2
XFILLER_34_279 vgnd vpwr scs8hd_decap_4
XFILLER_30_430 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_474 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _445_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
+ _417_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_213 vgnd vpwr scs8hd_decap_6
XFILLER_80_385 vgnd vpwr scs8hd_decap_12
XFILLER_40_205 vpwr vgnd scs8hd_fill_2
XFILLER_43_27 vgnd vpwr scs8hd_decap_12
XANTENNA__392__B _391_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_441 vgnd vpwr scs8hd_decap_12
XFILLER_21_485 vgnd vpwr scs8hd_decap_3
XFILLER_4_128 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_68 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_356 vgnd vpwr scs8hd_decap_3
XFILLER_75_135 vgnd vpwr scs8hd_decap_12
XFILLER_71_352 vpwr vgnd scs8hd_fill_2
XFILLER_71_341 vpwr vgnd scs8hd_fill_2
XFILLER_71_330 vpwr vgnd scs8hd_fill_2
XFILLER_16_235 vgnd vpwr scs8hd_fill_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_290 vpwr vgnd scs8hd_fill_2
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_296 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_79_452 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_308 vgnd vpwr scs8hd_decap_3
XFILLER_74_190 vgnd vpwr scs8hd_decap_12
XFILLER_62_341 vgnd vpwr scs8hd_decap_3
XFILLER_62_330 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ _140_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_62_396 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ _414_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__387__B _391_/B vgnd vpwr scs8hd_diode_2
XFILLER_72_105 vgnd vpwr scs8hd_decap_12
XFILLER_57_179 vpwr vgnd scs8hd_fill_2
XFILLER_38_360 vgnd vpwr scs8hd_decap_3
XFILLER_65_190 vgnd vpwr scs8hd_decap_3
XFILLER_54_15 vgnd vpwr scs8hd_decap_12
XFILLER_38_393 vgnd vpwr scs8hd_decap_4
XFILLER_13_216 vpwr vgnd scs8hd_fill_2
XFILLER_53_385 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_426 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XFILLER_76_422 vgnd vpwr scs8hd_decap_12
XFILLER_0_175 vgnd vpwr scs8hd_decap_4
XFILLER_48_113 vgnd vpwr scs8hd_decap_4
XANTENNA__297__B _295_/B vgnd vpwr scs8hd_diode_2
XFILLER_48_168 vgnd vpwr scs8hd_decap_6
XFILLER_63_127 vpwr vgnd scs8hd_fill_2
XFILLER_28_93 vgnd vpwr scs8hd_fill_1
XFILLER_29_382 vgnd vpwr scs8hd_fill_1
XFILLER_32_503 vgnd vpwr scs8hd_decap_12
XFILLER_71_193 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_271 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_60_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch_SLEEPB _220_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ left_width_0_height_0__pin_11_ vgnd vpwr scs8hd_inv_1
XFILLER_5_86 vgnd vpwr scs8hd_decap_6
XFILLER_79_293 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_179 vpwr vgnd scs8hd_fill_2
XFILLER_82_447 vgnd vpwr scs8hd_decap_12
XFILLER_54_149 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ _147_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_363 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_366 vpwr vgnd scs8hd_fill_2
XFILLER_50_355 vpwr vgnd scs8hd_fill_2
XFILLER_50_388 vpwr vgnd scs8hd_fill_2
XFILLER_50_377 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ _136_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_49_15 vgnd vpwr scs8hd_decap_12
XFILLER_77_208 vgnd vpwr scs8hd_decap_12
XFILLER_49_59 vpwr vgnd scs8hd_fill_2
XANTENNA__398__A _204_/B vgnd vpwr scs8hd_diode_2
XFILLER_73_403 vgnd vpwr scs8hd_decap_12
XFILLER_58_499 vgnd vpwr scs8hd_decap_12
X_420_ _204_/B _416_/B _420_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_53_160 vgnd vpwr scs8hd_decap_4
X_351_ _279_/A _352_/B _351_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
X_282_ _273_/A _286_/B _282_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _147_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_245 vgnd vpwr scs8hd_decap_4
XFILLER_5_234 vpwr vgnd scs8hd_fill_2
XFILLER_5_289 vpwr vgnd scs8hd_fill_2
XFILLER_68_208 vgnd vpwr scs8hd_decap_6
XFILLER_1_440 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_400 vgnd vpwr scs8hd_decap_3
XFILLER_76_263 vgnd vpwr scs8hd_decap_12
XFILLER_64_414 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_105 vgnd vpwr scs8hd_decap_6
XFILLER_36_149 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_300 vgnd vpwr scs8hd_decap_8
XFILLER_32_311 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_72_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ _392_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_82_211 vgnd vpwr scs8hd_decap_6
XFILLER_55_414 vpwr vgnd scs8hd_fill_2
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XPHY_818 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_807 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_439 vgnd vpwr scs8hd_decap_12
XPHY_829 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__384__C _163_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_27 vgnd vpwr scs8hd_decap_12
XFILLER_50_163 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch_SLEEPB _292_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_248 vpwr vgnd scs8hd_fill_2
XFILLER_76_68 vgnd vpwr scs8hd_decap_12
XFILLER_61_439 vpwr vgnd scs8hd_fill_2
XFILLER_61_428 vpwr vgnd scs8hd_fill_2
XFILLER_54_480 vgnd vpwr scs8hd_decap_12
X_403_ _171_/X _402_/X _403_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_119 vgnd vpwr scs8hd_fill_1
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_decap_3
X_334_ _280_/A _326_/X _334_/Y vgnd vpwr scs8hd_nor2_4
XPHY_94 vgnd vpwr scs8hd_decap_3
X_265_ _274_/A _269_/B _265_/Y vgnd vpwr scs8hd_nor2_4
X_196_ address[3] _274_/A _197_/B vgnd vpwr scs8hd_or2_4
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_49_274 vpwr vgnd scs8hd_fill_2
XFILLER_64_233 vgnd vpwr scs8hd_decap_8
XFILLER_37_447 vgnd vpwr scs8hd_fill_1
XFILLER_49_296 vpwr vgnd scs8hd_fill_2
XFILLER_64_266 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _442_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_480 vgnd vpwr scs8hd_fill_1
XFILLER_60_483 vgnd vpwr scs8hd_decap_12
XFILLER_32_163 vpwr vgnd scs8hd_fill_2
XFILLER_9_370 vpwr vgnd scs8hd_fill_2
XFILLER_20_369 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch/Q ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ _158_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch_SLEEPB _265_/Y vgnd vpwr scs8hd_diode_2
XFILLER_46_27 vgnd vpwr scs8hd_decap_4
XFILLER_55_277 vgnd vpwr scs8hd_fill_1
XANTENNA__395__B _391_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_480 vgnd vpwr scs8hd_decap_12
XFILLER_43_428 vgnd vpwr scs8hd_decap_3
XFILLER_62_15 vgnd vpwr scs8hd_decap_12
XPHY_626 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_615 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_604 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_659 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_648 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_637 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_472 vpwr vgnd scs8hd_fill_2
XFILLER_11_358 vpwr vgnd scs8hd_fill_2
XFILLER_11_74 vgnd vpwr scs8hd_decap_6
XFILLER_3_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_46_255 vgnd vpwr scs8hd_fill_1
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XFILLER_14_141 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ _370_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_317_ address[6] address[7] _272_/C _263_/D _325_/B vgnd vpwr scs8hd_or4_4
X_248_ _276_/A _252_/B _248_/Y vgnd vpwr scs8hd_nor2_4
X_179_ _122_/Y _276_/A _367_/A vgnd vpwr scs8hd_or2_4
XFILLER_6_384 vgnd vpwr scs8hd_decap_12
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_77_391 vgnd vpwr scs8hd_decap_12
XFILLER_37_200 vpwr vgnd scs8hd_fill_2
XFILLER_52_203 vpwr vgnd scs8hd_fill_2
XFILLER_25_439 vpwr vgnd scs8hd_fill_2
XFILLER_52_269 vgnd vpwr scs8hd_decap_6
XFILLER_60_291 vpwr vgnd scs8hd_fill_2
XFILLER_20_111 vgnd vpwr scs8hd_fill_1
XFILLER_33_483 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch_SLEEPB _237_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ _388_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_57_15 vgnd vpwr scs8hd_decap_12
XFILLER_48_509 vgnd vpwr scs8hd_decap_6
XFILLER_75_306 vgnd vpwr scs8hd_decap_12
XFILLER_57_59 vpwr vgnd scs8hd_fill_2
XFILLER_71_501 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XPHY_401 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_236 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch/Q ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_412 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_423 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_434 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_269 vpwr vgnd scs8hd_fill_2
XPHY_445 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_456 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_467 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_478 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_489 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_199 vpwr vgnd scs8hd_fill_2
XFILLER_11_188 vpwr vgnd scs8hd_fill_2
XFILLER_7_115 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/Y _138_/A vgnd vpwr scs8hd_inv_1
XFILLER_3_332 vpwr vgnd scs8hd_fill_2
XFILLER_3_376 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch_SLEEPB _336_/Y vgnd vpwr scs8hd_diode_2
XFILLER_78_166 vgnd vpwr scs8hd_decap_12
XFILLER_19_211 vpwr vgnd scs8hd_fill_2
XFILLER_74_361 vgnd vpwr scs8hd_decap_12
XFILLER_19_277 vpwr vgnd scs8hd_fill_2
XFILLER_34_236 vgnd vpwr scs8hd_fill_1
XFILLER_42_280 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_486 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch/Q ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_69_144 vpwr vgnd scs8hd_fill_2
XFILLER_69_155 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_501 vgnd vpwr scs8hd_decap_12
XFILLER_25_236 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_431 vgnd vpwr scs8hd_decap_4
XFILLER_33_280 vpwr vgnd scs8hd_fill_2
XFILLER_40_239 vgnd vpwr scs8hd_fill_1
XFILLER_43_39 vgnd vpwr scs8hd_decap_12
XFILLER_21_453 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_324 vpwr vgnd scs8hd_fill_2
XFILLER_75_147 vgnd vpwr scs8hd_decap_12
XFILLER_56_350 vgnd vpwr scs8hd_decap_8
XFILLER_17_51 vgnd vpwr scs8hd_decap_8
XFILLER_17_62 vgnd vpwr scs8hd_decap_12
XFILLER_71_364 vpwr vgnd scs8hd_fill_2
XFILLER_31_206 vpwr vgnd scs8hd_fill_2
XFILLER_31_217 vpwr vgnd scs8hd_fill_2
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch_SLEEPB _309_/Y vgnd vpwr scs8hd_diode_2
XPHY_286 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_431 vgnd vpwr scs8hd_decap_12
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_297 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_79_464 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_306 vpwr vgnd scs8hd_fill_2
XFILLER_58_80 vgnd vpwr scs8hd_decap_12
XFILLER_39_328 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_501 vgnd vpwr scs8hd_decap_12
XFILLER_62_320 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_364 vgnd vpwr scs8hd_decap_3
XFILLER_62_353 vgnd vpwr scs8hd_decap_8
XFILLER_30_261 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ _133_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
+ _370_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _139_/Y vgnd vpwr scs8hd_diode_2
XFILLER_72_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch/Q ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_54_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_53_397 vgnd vpwr scs8hd_decap_3
XFILLER_13_239 vgnd vpwr scs8hd_decap_3
XFILLER_70_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_261 vpwr vgnd scs8hd_fill_2
XFILLER_21_272 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch_SLEEPB _282_/Y vgnd vpwr scs8hd_diode_2
XFILLER_76_434 vgnd vpwr scs8hd_decap_12
XFILLER_0_187 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_106 vpwr vgnd scs8hd_fill_2
XFILLER_17_501 vgnd vpwr scs8hd_decap_12
XFILLER_29_394 vpwr vgnd scs8hd_fill_2
XFILLER_32_515 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_93 vgnd vpwr scs8hd_decap_4
XFILLER_12_294 vgnd vpwr scs8hd_decap_4
XFILLER_8_298 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_471 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _439_/HI
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ _148_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_136 vgnd vpwr scs8hd_decap_4
XFILLER_39_147 vpwr vgnd scs8hd_fill_2
XFILLER_82_404 vgnd vpwr scs8hd_decap_12
XFILLER_67_489 vgnd vpwr scs8hd_decap_12
XFILLER_27_309 vgnd vpwr scs8hd_decap_4
XFILLER_82_459 vgnd vpwr scs8hd_decap_6
XFILLER_54_139 vgnd vpwr scs8hd_decap_8
XFILLER_35_331 vpwr vgnd scs8hd_fill_2
XFILLER_35_342 vpwr vgnd scs8hd_fill_2
XFILLER_35_397 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__398__B _391_/B vgnd vpwr scs8hd_diode_2
XFILLER_65_15 vgnd vpwr scs8hd_decap_12
XFILLER_73_415 vgnd vpwr scs8hd_decap_12
XFILLER_18_309 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_106 vpwr vgnd scs8hd_fill_2
XFILLER_65_59 vpwr vgnd scs8hd_fill_2
XFILLER_14_515 vgnd vpwr scs8hd_fill_1
XFILLER_26_375 vgnd vpwr scs8hd_decap_3
X_350_ _287_/A _352_/B _350_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_345 vpwr vgnd scs8hd_fill_2
XFILLER_41_356 vgnd vpwr scs8hd_fill_1
X_281_ address[6] _272_/B _272_/C _263_/D _286_/B vgnd vpwr scs8hd_or4_4
Xltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_1_452 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _157_/Y vgnd vpwr scs8hd_diode_2
XFILLER_49_423 vpwr vgnd scs8hd_fill_2
XFILLER_49_412 vgnd vpwr scs8hd_decap_4
XFILLER_64_404 vgnd vpwr scs8hd_fill_1
XFILLER_49_489 vgnd vpwr scs8hd_decap_12
XFILLER_64_459 vgnd vpwr scs8hd_decap_12
XFILLER_64_437 vgnd vpwr scs8hd_decap_4
XFILLER_29_191 vpwr vgnd scs8hd_fill_2
XFILLER_32_345 vgnd vpwr scs8hd_decap_4
XFILLER_20_507 vgnd vpwr scs8hd_decap_8
XFILLER_32_378 vpwr vgnd scs8hd_fill_2
XFILLER_32_389 vgnd vpwr scs8hd_decap_8
XFILLER_65_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ _155_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_67_297 vpwr vgnd scs8hd_fill_2
XFILLER_55_459 vpwr vgnd scs8hd_fill_2
XFILLER_55_426 vgnd vpwr scs8hd_fill_1
XFILLER_70_407 vpwr vgnd scs8hd_fill_2
XPHY_808 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_301 vpwr vgnd scs8hd_fill_2
XPHY_819 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _148_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__384__D _263_/D vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ _183_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_51_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch/Q
+ _357_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_78_507 vgnd vpwr scs8hd_decap_8
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_223 vpwr vgnd scs8hd_fill_2
XFILLER_18_139 vgnd vpwr scs8hd_decap_8
XFILLER_46_426 vpwr vgnd scs8hd_fill_2
XFILLER_46_459 vgnd vpwr scs8hd_decap_3
XFILLER_73_256 vpwr vgnd scs8hd_fill_2
XFILLER_73_245 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_402_ _380_/A _384_/X _402_/X vgnd vpwr scs8hd_or2_4
XPHY_40 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q
+ _322_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch_SLEEPB _262_/Y vgnd vpwr scs8hd_diode_2
XFILLER_54_492 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
+ set vgnd vpwr scs8hd_diode_2
XFILLER_25_51 vgnd vpwr scs8hd_decap_8
XFILLER_25_62 vgnd vpwr scs8hd_decap_12
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XFILLER_14_389 vgnd vpwr scs8hd_decap_8
X_333_ _279_/A _326_/X _333_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_153 vpwr vgnd scs8hd_fill_2
XFILLER_41_175 vpwr vgnd scs8hd_fill_2
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
X_264_ _273_/A _269_/B _264_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_197 vgnd vpwr scs8hd_decap_8
X_195_ _178_/A _181_/B address[0] _274_/A vgnd vpwr scs8hd_or3_4
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_94 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q
+ _287_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XFILLER_49_220 vpwr vgnd scs8hd_fill_2
XFILLER_66_80 vgnd vpwr scs8hd_decap_12
XFILLER_64_223 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q
+ _251_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_64_289 vgnd vpwr scs8hd_decap_8
XFILLER_17_161 vpwr vgnd scs8hd_fill_2
XFILLER_17_172 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_60_495 vgnd vpwr scs8hd_decap_12
XFILLER_32_175 vpwr vgnd scs8hd_fill_2
XFILLER_32_186 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_407 vgnd vpwr scs8hd_fill_1
XFILLER_70_215 vgnd vpwr scs8hd_decap_8
XFILLER_15_109 vpwr vgnd scs8hd_fill_2
XFILLER_62_27 vgnd vpwr scs8hd_decap_4
XPHY_616 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_605 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_131 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _135_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_492 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch/Q
+ _336_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_649 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_638 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_627 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_484 vgnd vpwr scs8hd_decap_4
XFILLER_11_315 vpwr vgnd scs8hd_fill_2
XFILLER_23_175 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_319 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch_SLEEPB _234_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch/Q
+ _301_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_78_337 vgnd vpwr scs8hd_decap_12
XFILLER_46_212 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
+ _399_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_407 vgnd vpwr scs8hd_decap_3
XFILLER_46_267 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch/Q
+ _266_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_481 vgnd vpwr scs8hd_decap_6
XFILLER_42_473 vgnd vpwr scs8hd_decap_8
X_316_ _280_/A _314_/B _316_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_42_484 vgnd vpwr scs8hd_decap_12
XFILLER_52_93 vgnd vpwr scs8hd_decap_6
X_247_ _247_/A _252_/B _247_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
X_178_ _178_/A _178_/B _276_/A vgnd vpwr scs8hd_or2_4
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch/Q
+ _230_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_396 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_359 vgnd vpwr scs8hd_decap_6
XFILLER_69_337 vpwr vgnd scs8hd_fill_2
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch_SLEEPB _333_/Y vgnd vpwr scs8hd_diode_2
XFILLER_52_215 vgnd vpwr scs8hd_decap_3
XFILLER_25_418 vpwr vgnd scs8hd_fill_2
XFILLER_52_248 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_167 vgnd vpwr scs8hd_fill_1
XFILLER_20_189 vgnd vpwr scs8hd_fill_1
XFILLER_75_318 vgnd vpwr scs8hd_decap_12
XFILLER_57_27 vgnd vpwr scs8hd_decap_12
XFILLER_28_201 vgnd vpwr scs8hd_decap_3
XFILLER_73_15 vgnd vpwr scs8hd_decap_12
XFILLER_71_513 vgnd vpwr scs8hd_decap_3
XFILLER_16_407 vgnd vpwr scs8hd_decap_8
XFILLER_43_215 vgnd vpwr scs8hd_decap_6
XFILLER_73_59 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_462 vgnd vpwr scs8hd_decap_12
XPHY_402 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_413 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_424 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_435 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_11_123 vgnd vpwr scs8hd_decap_3
XFILLER_11_112 vgnd vpwr scs8hd_fill_1
XPHY_446 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_457 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_468 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_145 vgnd vpwr scs8hd_decap_6
XPHY_479 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_178 vgnd vpwr scs8hd_decap_3
XFILLER_7_138 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_178 vgnd vpwr scs8hd_decap_12
XFILLER_74_373 vgnd vpwr scs8hd_decap_12
XFILLER_15_440 vgnd vpwr scs8hd_decap_12
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_498 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch_SLEEPB _306_/Y vgnd vpwr scs8hd_diode_2
XFILLER_69_123 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _446_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_189 vpwr vgnd scs8hd_fill_2
XANTENNA__300__A _273_/A vgnd vpwr scs8hd_diode_2
XFILLER_65_373 vpwr vgnd scs8hd_fill_2
XFILLER_53_513 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/Y _153_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_80_398 vgnd vpwr scs8hd_decap_12
XFILLER_40_229 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_465 vgnd vpwr scs8hd_decap_12
XFILLER_68_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _162_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__210__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_75_159 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_362 vgnd vpwr scs8hd_decap_4
XFILLER_71_321 vgnd vpwr scs8hd_decap_6
XFILLER_16_226 vgnd vpwr scs8hd_fill_1
XFILLER_17_74 vgnd vpwr scs8hd_decap_12
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_96 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_270 vgnd vpwr scs8hd_decap_4
XFILLER_12_443 vgnd vpwr scs8hd_decap_12
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_51 vgnd vpwr scs8hd_decap_8
XPHY_287 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_298 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_130 vpwr vgnd scs8hd_fill_2
XFILLER_79_476 vgnd vpwr scs8hd_decap_12
XFILLER_66_148 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch_SLEEPB _279_/Y vgnd vpwr scs8hd_diode_2
XFILLER_35_513 vgnd vpwr scs8hd_decap_3
XFILLER_47_362 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_74_80 vgnd vpwr scs8hd_decap_12
XFILLER_62_376 vgnd vpwr scs8hd_fill_1
XFILLER_50_505 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_292 vgnd vpwr scs8hd_fill_1
XFILLER_30_240 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
+ _194_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_72_129 vgnd vpwr scs8hd_decap_12
XFILLER_53_321 vpwr vgnd scs8hd_fill_2
XFILLER_53_376 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _149_/Y vgnd vpwr scs8hd_diode_2
XFILLER_70_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_240 vpwr vgnd scs8hd_fill_2
XFILLER_5_428 vgnd vpwr scs8hd_decap_12
XFILLER_5_406 vgnd vpwr scs8hd_decap_12
XANTENNA__205__A address[0] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_76_446 vgnd vpwr scs8hd_decap_12
XFILLER_63_118 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _142_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_513 vgnd vpwr scs8hd_decap_3
XFILLER_29_351 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_56_181 vpwr vgnd scs8hd_fill_2
XFILLER_71_151 vgnd vpwr scs8hd_decap_12
XFILLER_71_184 vpwr vgnd scs8hd_fill_2
XFILLER_44_398 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch_SLEEPB _251_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch/Q ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_60_93 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_483 vgnd vpwr scs8hd_decap_12
XFILLER_5_99 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _140_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q
+ _352_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_115 vgnd vpwr scs8hd_decap_4
XFILLER_67_446 vgnd vpwr scs8hd_decap_12
XFILLER_67_435 vpwr vgnd scs8hd_fill_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XFILLER_82_416 vgnd vpwr scs8hd_decap_12
XFILLER_54_118 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_321 vgnd vpwr scs8hd_fill_1
XFILLER_35_376 vpwr vgnd scs8hd_fill_2
XFILLER_50_346 vgnd vpwr scs8hd_decap_3
XFILLER_50_335 vgnd vpwr scs8hd_fill_1
XFILLER_49_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch_SLEEPB _350_/Y vgnd vpwr scs8hd_diode_2
XFILLER_65_27 vgnd vpwr scs8hd_decap_12
XFILLER_38_181 vgnd vpwr scs8hd_decap_8
XFILLER_53_140 vgnd vpwr scs8hd_decap_4
XFILLER_81_15 vgnd vpwr scs8hd_decap_12
XFILLER_53_184 vgnd vpwr scs8hd_fill_1
XFILLER_81_59 vpwr vgnd scs8hd_fill_2
X_280_ _280_/A _280_/B _280_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_464 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_76_276 vgnd vpwr scs8hd_decap_12
XFILLER_17_321 vpwr vgnd scs8hd_fill_2
XFILLER_72_471 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ _408_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_376 vgnd vpwr scs8hd_decap_4
XFILLER_17_398 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q
+ _331_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_58_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q
+ _296_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_67_232 vpwr vgnd scs8hd_fill_2
XFILLER_67_221 vgnd vpwr scs8hd_decap_3
XFILLER_67_254 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_809 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_35_162 vpwr vgnd scs8hd_fill_2
XFILLER_35_173 vpwr vgnd scs8hd_fill_2
XFILLER_23_335 vpwr vgnd scs8hd_fill_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q
+ _261_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_50_187 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch_SLEEPB _323_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_228 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _158_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q
+ _225_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_76_15 vgnd vpwr scs8hd_decap_12
XANTENNA__202__B _202_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/Y _155_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_58_232 vpwr vgnd scs8hd_fill_2
XFILLER_58_276 vgnd vpwr scs8hd_decap_4
XFILLER_58_254 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_401_ _210_/B _391_/B _401_/Y vgnd vpwr scs8hd_nor2_4
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_74 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vpwr vgnd scs8hd_fill_2
XFILLER_14_368 vpwr vgnd scs8hd_fill_2
XFILLER_25_74 vgnd vpwr scs8hd_decap_12
X_332_ _287_/A _326_/X _332_/Y vgnd vpwr scs8hd_nor2_4
XPHY_85 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_decap_3
X_263_ _263_/A _272_/B _272_/C _263_/D _269_/B vgnd vpwr scs8hd_or4_4
Xltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch/Q ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_194_ _202_/A _194_/B _194_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_49_243 vgnd vpwr scs8hd_fill_1
XFILLER_64_202 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_17_140 vgnd vpwr scs8hd_decap_8
XFILLER_17_184 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_32_143 vgnd vpwr scs8hd_decap_8
XFILLER_20_327 vgnd vpwr scs8hd_decap_8
XFILLER_9_361 vpwr vgnd scs8hd_fill_2
XFILLER_13_390 vgnd vpwr scs8hd_fill_1
XFILLER_9_394 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _443_/HI
+ vgnd vpwr scs8hd_diode_2
XANTENNA__303__A _276_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_427 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_43_419 vpwr vgnd scs8hd_fill_2
XPHY_617 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_606 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_121 vgnd vpwr scs8hd_fill_1
XPHY_639 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_628 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_51_496 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__213__A _187_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_78_349 vgnd vpwr scs8hd_decap_12
XFILLER_27_460 vpwr vgnd scs8hd_fill_2
XFILLER_61_249 vgnd vpwr scs8hd_fill_1
XFILLER_14_154 vgnd vpwr scs8hd_decap_4
XFILLER_42_463 vgnd vpwr scs8hd_fill_1
XFILLER_42_496 vgnd vpwr scs8hd_decap_12
X_315_ _279_/A _314_/B _315_/Y vgnd vpwr scs8hd_nor2_4
X_246_ _274_/A _252_/B _246_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
+ _382_/Y vgnd vpwr scs8hd_diode_2
X_177_ address[0] address[1] _178_/B vgnd vpwr scs8hd_or2_4
XFILLER_6_364 vgnd vpwr scs8hd_decap_8
XANTENNA__123__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_69_327 vgnd vpwr scs8hd_decap_4
XFILLER_37_213 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch/Q ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_471 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _136_/Y vgnd vpwr scs8hd_diode_2
XFILLER_52_227 vpwr vgnd scs8hd_fill_2
XFILLER_20_157 vpwr vgnd scs8hd_fill_2
XFILLER_20_179 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_57_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ _159_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_73_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch/Q ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ _132_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_43_249 vgnd vpwr scs8hd_decap_4
XFILLER_24_441 vgnd vpwr scs8hd_fill_1
XPHY_403 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_414 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_425 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_36_290 vgnd vpwr scs8hd_decap_3
XFILLER_51_282 vpwr vgnd scs8hd_fill_2
XANTENNA__208__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_474 vgnd vpwr scs8hd_decap_12
XPHY_436 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_447 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_458 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_469 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_157 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_66_308 vgnd vpwr scs8hd_decap_6
XFILLER_59_382 vgnd vpwr scs8hd_decap_3
XFILLER_19_257 vgnd vpwr scs8hd_decap_3
XFILLER_47_94 vpwr vgnd scs8hd_fill_2
XFILLER_74_385 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_15_452 vgnd vpwr scs8hd_decap_12
XFILLER_30_411 vpwr vgnd scs8hd_fill_2
XFILLER_42_271 vgnd vpwr scs8hd_decap_4
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
X_229_ _247_/A _231_/B _229_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_8_88 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/Y _144_/A vgnd vpwr scs8hd_inv_1
XFILLER_6_150 vgnd vpwr scs8hd_decap_3
XFILLER_6_183 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XFILLER_69_135 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_179 vpwr vgnd scs8hd_fill_2
XFILLER_57_319 vgnd vpwr scs8hd_decap_4
XANTENNA__300__B _304_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_80_300 vgnd vpwr scs8hd_decap_12
XFILLER_65_352 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_396 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_477 vgnd vpwr scs8hd_decap_8
XFILLER_4_109 vpwr vgnd scs8hd_fill_2
XFILLER_68_27 vgnd vpwr scs8hd_decap_4
XFILLER_0_337 vpwr vgnd scs8hd_fill_2
XFILLER_48_308 vgnd vpwr scs8hd_decap_3
XANTENNA__210__B _210_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _154_/Y vgnd vpwr scs8hd_diode_2
XFILLER_71_300 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ _139_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_width_0_height_0__pin_10_ vgnd vpwr scs8hd_inv_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_249 vpwr vgnd scs8hd_fill_2
XFILLER_17_86 vgnd vpwr scs8hd_decap_4
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _132_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_455 vgnd vpwr scs8hd_decap_3
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_288 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_299 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XFILLER_8_459 vgnd vpwr scs8hd_decap_12
XFILLER_33_96 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_175 vpwr vgnd scs8hd_fill_2
XFILLER_3_164 vpwr vgnd scs8hd_fill_2
XANTENNA__401__A _210_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_197 vpwr vgnd scs8hd_fill_2
XFILLER_66_127 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_58_93 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_47_352 vpwr vgnd scs8hd_fill_2
XFILLER_47_396 vpwr vgnd scs8hd_fill_2
XFILLER_62_388 vpwr vgnd scs8hd_fill_2
XFILLER_22_208 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__311__A _247_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_116 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_138 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/Y _162_/A vgnd vpwr scs8hd_inv_1
XFILLER_53_333 vpwr vgnd scs8hd_fill_2
XFILLER_38_374 vpwr vgnd scs8hd_fill_2
XFILLER_38_385 vgnd vpwr scs8hd_decap_6
XFILLER_80_141 vgnd vpwr scs8hd_decap_12
XFILLER_21_230 vgnd vpwr scs8hd_fill_1
XFILLER_21_285 vpwr vgnd scs8hd_fill_2
XFILLER_21_296 vpwr vgnd scs8hd_fill_2
XFILLER_5_418 vgnd vpwr scs8hd_decap_8
XFILLER_79_15 vgnd vpwr scs8hd_decap_12
XANTENNA__205__B _181_/B vgnd vpwr scs8hd_diode_2
XFILLER_79_59 vpwr vgnd scs8hd_fill_2
XANTENNA__221__A _276_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_156 vpwr vgnd scs8hd_fill_2
XFILLER_48_127 vgnd vpwr scs8hd_decap_12
XFILLER_29_363 vgnd vpwr scs8hd_fill_1
XFILLER_29_374 vpwr vgnd scs8hd_fill_2
XFILLER_71_163 vgnd vpwr scs8hd_fill_1
XFILLER_44_377 vgnd vpwr scs8hd_decap_8
XFILLER_44_388 vpwr vgnd scs8hd_fill_2
XFILLER_8_201 vgnd vpwr scs8hd_decap_12
XFILLER_12_274 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_256 vgnd vpwr scs8hd_decap_4
XFILLER_4_451 vgnd vpwr scs8hd_decap_6
XFILLER_4_495 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__131__A _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_67_403 vpwr vgnd scs8hd_fill_2
XFILLER_67_458 vgnd vpwr scs8hd_decap_12
XFILLER_82_428 vgnd vpwr scs8hd_decap_6
XFILLER_47_160 vpwr vgnd scs8hd_fill_2
XFILLER_62_141 vgnd vpwr scs8hd_fill_1
XFILLER_35_355 vpwr vgnd scs8hd_fill_2
XFILLER_50_303 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _150_/Y vgnd vpwr scs8hd_diode_2
XFILLER_50_325 vpwr vgnd scs8hd_fill_2
XANTENNA__306__A _279_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_58_436 vgnd vpwr scs8hd_fill_1
XFILLER_65_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_428 vgnd vpwr scs8hd_decap_12
XFILLER_38_171 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_344 vgnd vpwr scs8hd_decap_4
XFILLER_81_27 vgnd vpwr scs8hd_decap_12
XFILLER_53_152 vpwr vgnd scs8hd_fill_2
XFILLER_53_196 vpwr vgnd scs8hd_fill_2
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__216__A enable vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_476 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2/Z
+ _150_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_51 vgnd vpwr scs8hd_decap_8
XFILLER_49_458 vgnd vpwr scs8hd_fill_1
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XFILLER_76_288 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
+ _404_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_355 vgnd vpwr scs8hd_fill_1
XFILLER_72_483 vgnd vpwr scs8hd_decap_12
XFILLER_55_94 vgnd vpwr scs8hd_decap_3
XFILLER_44_152 vgnd vpwr scs8hd_fill_1
XFILLER_44_196 vgnd vpwr scs8hd_fill_1
XANTENNA__126__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_67_288 vgnd vpwr scs8hd_decap_6
XFILLER_67_277 vpwr vgnd scs8hd_fill_2
XFILLER_55_428 vgnd vpwr scs8hd_decap_3
XFILLER_27_119 vgnd vpwr scs8hd_fill_1
XFILLER_63_461 vgnd vpwr scs8hd_decap_12
XFILLER_23_314 vpwr vgnd scs8hd_fill_2
XFILLER_23_358 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_27 vgnd vpwr scs8hd_decap_4
XFILLER_58_244 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_450 vgnd vpwr scs8hd_decap_8
XPHY_20 vgnd vpwr scs8hd_decap_3
X_400_ _208_/B _391_/B _400_/Y vgnd vpwr scs8hd_nor2_4
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_26_141 vgnd vpwr scs8hd_fill_1
XFILLER_26_163 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_decap_3
X_331_ _231_/A _326_/X _331_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_86 vpwr vgnd scs8hd_fill_2
XFILLER_25_97 vpwr vgnd scs8hd_fill_2
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_decap_3
X_262_ _280_/A _262_/B _262_/Y vgnd vpwr scs8hd_nor2_4
X_193_ address[3] _273_/A _194_/B vgnd vpwr scs8hd_or2_4
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ _382_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_273 vpwr vgnd scs8hd_fill_2
XFILLER_1_284 vpwr vgnd scs8hd_fill_2
XFILLER_49_233 vpwr vgnd scs8hd_fill_2
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_37_417 vpwr vgnd scs8hd_fill_2
XFILLER_37_439 vpwr vgnd scs8hd_fill_2
XFILLER_66_93 vgnd vpwr scs8hd_decap_12
XFILLER_64_258 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_72_280 vgnd vpwr scs8hd_decap_12
XFILLER_45_483 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_306 vpwr vgnd scs8hd_fill_2
XFILLER_20_317 vgnd vpwr scs8hd_decap_8
XFILLER_70_3 vgnd vpwr scs8hd_decap_12
XANTENNA__303__B _304_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_55_258 vpwr vgnd scs8hd_fill_2
XFILLER_55_236 vpwr vgnd scs8hd_fill_2
XFILLER_70_206 vgnd vpwr scs8hd_decap_8
XPHY_607 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_420 vgnd vpwr scs8hd_decap_4
XFILLER_23_111 vpwr vgnd scs8hd_fill_2
XPHY_629 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_618 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_144 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_306 vgnd vpwr scs8hd_decap_3
XFILLER_23_199 vpwr vgnd scs8hd_fill_2
XANTENNA__213__B _214_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
+ _428_/HI ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_406 vpwr vgnd scs8hd_fill_2
XFILLER_19_428 vgnd vpwr scs8hd_decap_12
XFILLER_46_203 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
+ _408_/Y vgnd vpwr scs8hd_diode_2
XFILLER_46_247 vgnd vpwr scs8hd_decap_8
XFILLER_61_217 vpwr vgnd scs8hd_fill_2
XFILLER_42_431 vgnd vpwr scs8hd_decap_6
X_314_ _287_/A _314_/B _314_/Y vgnd vpwr scs8hd_nor2_4
X_245_ _273_/A _252_/B _245_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_176_ _202_/A _176_/B _176_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_354 vgnd vpwr scs8hd_fill_1
XANTENNA__404__A _187_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ _202_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_69_306 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_501 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
+ clk ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff/QN
+ reset set vgnd vpwr scs8hd_dfbbp_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_80_515 vgnd vpwr scs8hd_fill_1
XFILLER_37_269 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_483 vgnd vpwr scs8hd_decap_12
XFILLER_20_103 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__314__A _287_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_269 vgnd vpwr scs8hd_decap_6
XFILLER_73_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XPHY_404 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_415 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_426 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__208__B _208_/B vgnd vpwr scs8hd_diode_2
XFILLER_24_486 vgnd vpwr scs8hd_decap_12
XPHY_437 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_448 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_459 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XFILLER_7_107 vgnd vpwr scs8hd_decap_8
XFILLER_22_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch/Q ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__224__A _279_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
+ _420_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_203 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_501 vgnd vpwr scs8hd_decap_12
XFILLER_59_394 vgnd vpwr scs8hd_decap_4
XFILLER_19_236 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_47_51 vgnd vpwr scs8hd_decap_8
XFILLER_47_62 vgnd vpwr scs8hd_decap_12
XFILLER_62_515 vgnd vpwr scs8hd_fill_1
XFILLER_34_206 vgnd vpwr scs8hd_decap_8
XFILLER_27_280 vgnd vpwr scs8hd_fill_1
XFILLER_34_228 vgnd vpwr scs8hd_decap_8
XFILLER_15_464 vgnd vpwr scs8hd_decap_12
XFILLER_30_423 vgnd vpwr scs8hd_fill_1
XFILLER_8_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_228_ _274_/A _231_/B _228_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__134__A _134_/A vgnd vpwr scs8hd_diode_2
X_159_ _159_/A _159_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
XFILLER_80_312 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _447_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_280 vgnd vpwr scs8hd_decap_3
XANTENNA__309__A _273_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_401 vpwr vgnd scs8hd_fill_2
XFILLER_40_209 vgnd vpwr scs8hd_decap_4
XFILLER_21_489 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_501 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ _140_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_206 vgnd vpwr scs8hd_decap_4
XFILLER_44_515 vgnd vpwr scs8hd_fill_1
XFILLER_71_334 vgnd vpwr scs8hd_decap_4
XFILLER_71_367 vgnd vpwr scs8hd_decap_12
XFILLER_71_356 vgnd vpwr scs8hd_decap_8
XFILLER_71_345 vpwr vgnd scs8hd_fill_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__219__A _274_/A vgnd vpwr scs8hd_diode_2
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_261 vpwr vgnd scs8hd_fill_2
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ _419_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_24_294 vgnd vpwr scs8hd_fill_1
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_289 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
+ _426_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__401__B _391_/B vgnd vpwr scs8hd_diode_2
XFILLER_79_489 vgnd vpwr scs8hd_decap_12
XFILLER_59_191 vgnd vpwr scs8hd_decap_4
XFILLER_62_301 vpwr vgnd scs8hd_fill_2
XFILLER_74_93 vgnd vpwr scs8hd_decap_12
XANTENNA__129__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_790 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch/Q
+ _245_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__311__B _314_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ _426_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_504 vgnd vpwr scs8hd_decap_12
XFILLER_53_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch_SLEEPB _223_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_90 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch/Q ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_79_27 vgnd vpwr scs8hd_decap_12
XANTENNA__205__C address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__221__B _225_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_179 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ _147_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_48_117 vgnd vpwr scs8hd_fill_1
XFILLER_76_459 vgnd vpwr scs8hd_decap_12
XFILLER_48_139 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_71_175 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_235 vpwr vgnd scs8hd_fill_2
XFILLER_8_213 vgnd vpwr scs8hd_fill_1
XANTENNA__412__A _183_/B vgnd vpwr scs8hd_diode_2
XFILLER_79_220 vgnd vpwr scs8hd_decap_12
XFILLER_39_106 vgnd vpwr scs8hd_decap_3
XFILLER_67_426 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_301 vpwr vgnd scs8hd_fill_2
XANTENNA__306__B _304_/B vgnd vpwr scs8hd_diode_2
XANTENNA__322__A _231_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_404 vpwr vgnd scs8hd_fill_2
XFILLER_58_459 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ _397_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_81_440 vgnd vpwr scs8hd_decap_12
XFILLER_53_175 vpwr vgnd scs8hd_fill_2
XFILLER_14_507 vgnd vpwr scs8hd_decap_8
XFILLER_26_389 vpwr vgnd scs8hd_fill_2
XFILLER_41_315 vpwr vgnd scs8hd_fill_2
XFILLER_81_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_14_44 vgnd vpwr scs8hd_decap_12
XFILLER_41_359 vgnd vpwr scs8hd_decap_4
XFILLER_14_99 vgnd vpwr scs8hd_decap_3
XANTENNA__216__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_5_205 vgnd vpwr scs8hd_fill_1
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_238 vpwr vgnd scs8hd_fill_2
XANTENNA__232__A _287_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_400 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_49_437 vpwr vgnd scs8hd_fill_2
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XFILLER_57_470 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch_SLEEPB _295_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_62 vgnd vpwr scs8hd_decap_12
XFILLER_55_51 vgnd vpwr scs8hd_decap_8
XFILLER_17_334 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _143_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_72_495 vgnd vpwr scs8hd_decap_12
XFILLER_32_315 vgnd vpwr scs8hd_decap_4
XFILLER_32_337 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_175 vgnd vpwr scs8hd_decap_3
XANTENNA__407__A address[4] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _142_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_418 vpwr vgnd scs8hd_fill_2
XFILLER_27_109 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_473 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch/Q ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__317__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
+ _387_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_370 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_58_267 vgnd vpwr scs8hd_decap_8
XFILLER_54_473 vgnd vpwr scs8hd_decap_4
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XFILLER_81_281 vgnd vpwr scs8hd_decap_12
XFILLER_14_337 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_26_186 vgnd vpwr scs8hd_decap_4
XPHY_65 vgnd vpwr scs8hd_decap_3
X_330_ _276_/A _326_/X _330_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_123 vpwr vgnd scs8hd_fill_2
XANTENNA__227__A _273_/A vgnd vpwr scs8hd_diode_2
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_decap_3
X_261_ _279_/A _262_/B _261_/Y vgnd vpwr scs8hd_nor2_4
X_192_ _202_/A _371_/A _192_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch_SLEEPB _268_/Y vgnd vpwr scs8hd_diode_2
XFILLER_41_86 vgnd vpwr scs8hd_decap_8
XFILLER_41_97 vpwr vgnd scs8hd_fill_2
XFILLER_1_252 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_49_245 vgnd vpwr scs8hd_decap_3
XFILLER_64_215 vgnd vpwr scs8hd_decap_8
XFILLER_49_278 vpwr vgnd scs8hd_fill_2
XFILLER_72_292 vgnd vpwr scs8hd_decap_12
XANTENNA__137__A _137_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_167 vgnd vpwr scs8hd_decap_4
XFILLER_9_330 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_374 vgnd vpwr scs8hd_decap_4
XFILLER_63_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ _375_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_55_215 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_451 vgnd vpwr scs8hd_decap_6
XPHY_608 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_63_292 vgnd vpwr scs8hd_decap_4
XPHY_619 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_432 vgnd vpwr scs8hd_fill_1
XFILLER_23_123 vpwr vgnd scs8hd_fill_2
XFILLER_23_156 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_476 vpwr vgnd scs8hd_fill_2
XFILLER_23_167 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_89 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_215 vpwr vgnd scs8hd_fill_2
XFILLER_46_226 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch_SLEEPB _240_/Y vgnd vpwr scs8hd_diode_2
XFILLER_46_259 vpwr vgnd scs8hd_fill_2
XFILLER_54_270 vgnd vpwr scs8hd_decap_3
XFILLER_14_145 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
+ _213_/Y vgnd vpwr scs8hd_diode_2
X_313_ _231_/A _314_/B _313_/Y vgnd vpwr scs8hd_nor2_4
X_244_ address[8] _235_/B _235_/C _263_/D _252_/B vgnd vpwr scs8hd_or4_4
XFILLER_10_351 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_333 vgnd vpwr scs8hd_fill_1
X_175_ _122_/Y _178_/A _181_/C address[1] _176_/B vgnd vpwr scs8hd_or4_4
XANTENNA__404__B _402_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__420__A _204_/B vgnd vpwr scs8hd_diode_2
XFILLER_65_513 vgnd vpwr scs8hd_decap_3
XFILLER_37_204 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch/Q ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_248 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_207 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/Y _132_/A vgnd vpwr scs8hd_inv_1
XFILLER_18_495 vgnd vpwr scs8hd_decap_12
XFILLER_33_421 vgnd vpwr scs8hd_decap_6
XFILLER_33_432 vpwr vgnd scs8hd_fill_2
XFILLER_60_273 vpwr vgnd scs8hd_fill_2
XFILLER_33_487 vgnd vpwr scs8hd_fill_1
XFILLER_60_295 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch_SLEEPB _339_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _141_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch/Q
+ _346_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_171 vgnd vpwr scs8hd_fill_1
XANTENNA__314__B _314_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_509 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__330__A _276_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch/Q
+ _311_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_56_513 vgnd vpwr scs8hd_decap_3
XFILLER_28_226 vpwr vgnd scs8hd_fill_2
XFILLER_28_248 vgnd vpwr scs8hd_decap_8
XFILLER_51_240 vpwr vgnd scs8hd_fill_2
XPHY_405 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_416 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_427 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_438 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_449 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch/Q
+ _276_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_115 vpwr vgnd scs8hd_fill_2
XFILLER_24_498 vgnd vpwr scs8hd_decap_12
XFILLER_22_44 vgnd vpwr scs8hd_decap_12
XANTENNA__224__B _225_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_336 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__240__A _231_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q
+ _240_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_59_362 vpwr vgnd scs8hd_fill_2
XFILLER_47_513 vgnd vpwr scs8hd_decap_3
XFILLER_19_226 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _132_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_248 vgnd vpwr scs8hd_decap_3
XFILLER_47_74 vgnd vpwr scs8hd_decap_12
XFILLER_74_398 vgnd vpwr scs8hd_decap_12
XFILLER_63_51 vgnd vpwr scs8hd_decap_8
XFILLER_15_421 vgnd vpwr scs8hd_decap_6
XFILLER_63_62 vgnd vpwr scs8hd_decap_12
XFILLER_15_476 vgnd vpwr scs8hd_decap_12
XFILLER_42_284 vpwr vgnd scs8hd_fill_2
XFILLER_30_457 vgnd vpwr scs8hd_fill_1
X_227_ _273_/A _231_/B _227_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__415__A _371_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_68 vgnd vpwr scs8hd_decap_12
X_158_ _158_/A _158_/Y vgnd vpwr scs8hd_inv_8
XFILLER_69_159 vgnd vpwr scs8hd_fill_1
XANTENNA__150__A _150_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch_SLEEPB _312_/Y vgnd vpwr scs8hd_diode_2
XFILLER_65_310 vpwr vgnd scs8hd_fill_2
XFILLER_65_365 vgnd vpwr scs8hd_fill_1
XFILLER_80_324 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ _134_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_292 vgnd vpwr scs8hd_decap_3
XANTENNA__309__B _314_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_424 vgnd vpwr scs8hd_fill_1
XFILLER_33_273 vgnd vpwr scs8hd_decap_4
XFILLER_33_284 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__325__A _280_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/Y _150_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_306 vpwr vgnd scs8hd_fill_2
XFILLER_0_328 vpwr vgnd scs8hd_fill_2
XFILLER_29_513 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch/Q
+ _255_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_71_313 vpwr vgnd scs8hd_fill_2
XFILLER_16_229 vgnd vpwr scs8hd_decap_4
XANTENNA__219__B _225_/B vgnd vpwr scs8hd_diode_2
XFILLER_71_379 vgnd vpwr scs8hd_decap_12
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
+ _373_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch/Q
+ _219_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__235__A address[8] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_66_107 vgnd vpwr scs8hd_decap_4
XFILLER_47_321 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_324 vgnd vpwr scs8hd_decap_4
XFILLER_47_376 vpwr vgnd scs8hd_fill_2
XFILLER_15_240 vpwr vgnd scs8hd_fill_2
XFILLER_15_273 vpwr vgnd scs8hd_fill_2
XFILLER_15_295 vgnd vpwr scs8hd_decap_8
XPHY_780 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_791 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch_SLEEPB _285_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__145__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_265 vpwr vgnd scs8hd_fill_2
XFILLER_30_276 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_140 vpwr vgnd scs8hd_fill_2
XFILLER_65_173 vpwr vgnd scs8hd_fill_2
XFILLER_65_162 vpwr vgnd scs8hd_fill_2
XFILLER_65_184 vgnd vpwr scs8hd_decap_4
XFILLER_80_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__205__D address[2] vgnd vpwr scs8hd_diode_2
XFILLER_79_39 vgnd vpwr scs8hd_decap_12
XFILLER_0_136 vpwr vgnd scs8hd_fill_2
XFILLER_0_125 vpwr vgnd scs8hd_fill_2
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
XFILLER_29_332 vgnd vpwr scs8hd_decap_4
XFILLER_71_110 vgnd vpwr scs8hd_decap_12
XFILLER_29_398 vpwr vgnd scs8hd_fill_2
XFILLER_44_324 vgnd vpwr scs8hd_fill_1
XFILLER_44_346 vgnd vpwr scs8hd_decap_3
XFILLER_71_143 vgnd vpwr scs8hd_fill_1
XFILLER_12_210 vgnd vpwr scs8hd_decap_4
XFILLER_52_390 vgnd vpwr scs8hd_decap_6
XFILLER_12_276 vgnd vpwr scs8hd_decap_3
XFILLER_12_298 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__412__B _416_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
+ _366_/Y vgnd vpwr scs8hd_diode_2
XFILLER_79_232 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_416 vpwr vgnd scs8hd_fill_2
XFILLER_62_121 vgnd vpwr scs8hd_decap_3
XFILLER_62_110 vgnd vpwr scs8hd_decap_8
XFILLER_47_184 vgnd vpwr scs8hd_fill_1
XFILLER_62_165 vgnd vpwr scs8hd_fill_1
XFILLER_62_187 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ _156_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _155_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_280 vpwr vgnd scs8hd_fill_2
XANTENNA__322__B _325_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _137_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/Y _145_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_66_471 vgnd vpwr scs8hd_decap_12
XFILLER_26_302 vgnd vpwr scs8hd_decap_4
XFILLER_53_132 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_81_452 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch_SLEEPB _356_/Y vgnd vpwr scs8hd_diode_2
XFILLER_41_327 vgnd vpwr scs8hd_decap_3
XFILLER_34_390 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_56 vgnd vpwr scs8hd_decap_12
XFILLER_5_217 vpwr vgnd scs8hd_fill_2
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XANTENNA__232__B _231_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ _155_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_76_202 vgnd vpwr scs8hd_decap_12
XFILLER_49_416 vgnd vpwr scs8hd_fill_1
XFILLER_1_489 vgnd vpwr scs8hd_decap_12
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XFILLER_17_302 vgnd vpwr scs8hd_decap_3
XFILLER_57_482 vgnd vpwr scs8hd_decap_6
XFILLER_29_195 vpwr vgnd scs8hd_fill_2
XFILLER_55_74 vgnd vpwr scs8hd_decap_12
XFILLER_44_154 vpwr vgnd scs8hd_fill_2
XFILLER_44_187 vgnd vpwr scs8hd_decap_3
XFILLER_9_501 vgnd vpwr scs8hd_decap_12
XANTENNA__407__B _406_/X vgnd vpwr scs8hd_diode_2
XFILLER_71_62 vgnd vpwr scs8hd_decap_12
XFILLER_71_51 vgnd vpwr scs8hd_decap_8
XANTENNA__423__A _210_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_250 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_67_202 vpwr vgnd scs8hd_fill_2
XFILLER_82_249 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_143 vgnd vpwr scs8hd_decap_4
XFILLER_63_485 vgnd vpwr scs8hd_decap_3
XFILLER_50_102 vpwr vgnd scs8hd_fill_2
XANTENNA__317__B address[7] vgnd vpwr scs8hd_diode_2
XFILLER_31_382 vpwr vgnd scs8hd_fill_2
XANTENNA__333__A _279_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_227 vpwr vgnd scs8hd_fill_2
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_81_293 vgnd vpwr scs8hd_decap_12
XFILLER_14_349 vgnd vpwr scs8hd_decap_8
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_decap_3
XFILLER_41_157 vpwr vgnd scs8hd_fill_2
XPHY_88 vgnd vpwr scs8hd_decap_3
XANTENNA__227__B _231_/B vgnd vpwr scs8hd_diode_2
XPHY_99 vgnd vpwr scs8hd_decap_3
XFILLER_41_179 vpwr vgnd scs8hd_fill_2
X_260_ _287_/A _262_/B _260_/Y vgnd vpwr scs8hd_nor2_4
X_191_ _122_/Y _280_/A _371_/A vgnd vpwr scs8hd_or2_4
XFILLER_22_393 vgnd vpwr scs8hd_decap_4
XFILLER_6_515 vgnd vpwr scs8hd_fill_1
XANTENNA__243__A _280_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q
+ _341_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_297 vpwr vgnd scs8hd_fill_2
XFILLER_49_257 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _133_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q
+ _306_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_132 vpwr vgnd scs8hd_fill_2
XFILLER_45_441 vpwr vgnd scs8hd_fill_2
XFILLER_45_463 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_72_260 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__418__A _200_/B vgnd vpwr scs8hd_diode_2
XFILLER_17_165 vpwr vgnd scs8hd_fill_2
XFILLER_17_176 vgnd vpwr scs8hd_decap_4
XFILLER_60_433 vpwr vgnd scs8hd_fill_2
XFILLER_82_94 vgnd vpwr scs8hd_decap_12
XFILLER_32_179 vgnd vpwr scs8hd_decap_4
X_389_ _367_/A _391_/B _389_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_382 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q
+ _271_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__153__A _153_/A vgnd vpwr scs8hd_diode_2
XFILLER_56_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ _367_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_408 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_430 vgnd vpwr scs8hd_decap_8
XFILLER_63_271 vpwr vgnd scs8hd_fill_2
XFILLER_63_260 vpwr vgnd scs8hd_fill_2
XANTENNA__328__A _274_/A vgnd vpwr scs8hd_diode_2
XPHY_609 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_455 vpwr vgnd scs8hd_fill_2
XFILLER_51_444 vgnd vpwr scs8hd_decap_3
XFILLER_23_179 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_419 vpwr vgnd scs8hd_fill_2
XFILLER_27_441 vpwr vgnd scs8hd_fill_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XANTENNA__238__A _247_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_113 vgnd vpwr scs8hd_decap_4
XFILLER_14_124 vpwr vgnd scs8hd_fill_2
X_312_ _276_/A _314_/B _312_/Y vgnd vpwr scs8hd_nor2_4
X_243_ _280_/A _243_/B _243_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_301 vgnd vpwr scs8hd_decap_4
X_174_ _181_/C address[1] _187_/B vgnd vpwr scs8hd_or2_4
XFILLER_6_323 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__420__B _416_/B vgnd vpwr scs8hd_diode_2
XFILLER_77_330 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_227 vpwr vgnd scs8hd_fill_2
XANTENNA__148__A _148_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ _131_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch/Q ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_60_263 vpwr vgnd scs8hd_fill_2
XFILLER_60_241 vgnd vpwr scs8hd_decap_4
XFILLER_9_150 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _151_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__330__B _326_/X vgnd vpwr scs8hd_diode_2
XFILLER_28_238 vgnd vpwr scs8hd_fill_1
XFILLER_24_444 vgnd vpwr scs8hd_decap_3
XPHY_406 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_417 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_252 vpwr vgnd scs8hd_fill_2
XPHY_428 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_439 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch/Q ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_56 vgnd vpwr scs8hd_decap_12
XFILLER_3_315 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/Y _147_/A vgnd vpwr scs8hd_buf_1
XFILLER_3_359 vgnd vpwr scs8hd_decap_4
XFILLER_78_105 vgnd vpwr scs8hd_decap_12
XANTENNA__240__B _243_/B vgnd vpwr scs8hd_diode_2
XFILLER_59_352 vpwr vgnd scs8hd_fill_2
XFILLER_74_300 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_47_86 vgnd vpwr scs8hd_decap_4
XFILLER_42_230 vgnd vpwr scs8hd_decap_8
XFILLER_63_74 vgnd vpwr scs8hd_decap_12
XFILLER_30_447 vgnd vpwr scs8hd_decap_8
X_226_ address[8] _235_/B _215_/X _263_/D _231_/B vgnd vpwr scs8hd_or4_4
XANTENNA__415__B _416_/B vgnd vpwr scs8hd_diode_2
X_157_ _157_/A _157_/Y vgnd vpwr scs8hd_inv_8
XFILLER_69_127 vgnd vpwr scs8hd_fill_1
XFILLER_77_171 vgnd vpwr scs8hd_decap_12
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_377 vpwr vgnd scs8hd_fill_2
XFILLER_21_414 vpwr vgnd scs8hd_fill_2
XANTENNA__325__B _325_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__341__A _287_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_68_160 vgnd vpwr scs8hd_decap_4
XFILLER_56_333 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_377 vgnd vpwr scs8hd_decap_3
XFILLER_56_366 vgnd vpwr scs8hd_fill_1
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_274 vgnd vpwr scs8hd_fill_1
XFILLER_24_285 vgnd vpwr scs8hd_decap_3
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_407 vgnd vpwr scs8hd_decap_12
XANTENNA__235__B _235_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
+ _202_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__251__A _279_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_134 vpwr vgnd scs8hd_fill_2
XFILLER_79_403 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_182 vgnd vpwr scs8hd_fill_1
XFILLER_74_141 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _147_/Y vgnd vpwr scs8hd_diode_2
XFILLER_47_333 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch/Q ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_47_388 vgnd vpwr scs8hd_decap_3
XFILLER_62_369 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XPHY_781 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_770 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__426__A _187_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_244 vgnd vpwr scs8hd_fill_1
XPHY_792 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_440 vgnd vpwr scs8hd_decap_12
X_209_ address[3] _280_/A _210_/B vgnd vpwr scs8hd_or2_4
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ _142_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_57_119 vgnd vpwr scs8hd_decap_3
XFILLER_38_300 vgnd vpwr scs8hd_decap_6
XFILLER_80_166 vgnd vpwr scs8hd_decap_12
XFILLER_53_358 vpwr vgnd scs8hd_fill_2
XFILLER_21_222 vpwr vgnd scs8hd_fill_2
XANTENNA__336__A _273_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_44 vgnd vpwr scs8hd_decap_12
XFILLER_29_355 vpwr vgnd scs8hd_fill_2
XFILLER_44_314 vgnd vpwr scs8hd_decap_8
XFILLER_56_185 vpwr vgnd scs8hd_fill_2
XFILLER_44_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__246__A _274_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_222 vpwr vgnd scs8hd_fill_2
XFILLER_8_215 vpwr vgnd scs8hd_fill_2
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_59 vpwr vgnd scs8hd_fill_2
XFILLER_69_62 vgnd vpwr scs8hd_decap_12
XFILLER_69_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_119 vgnd vpwr scs8hd_fill_1
XFILLER_62_133 vpwr vgnd scs8hd_fill_2
XFILLER_47_196 vpwr vgnd scs8hd_fill_2
XFILLER_62_177 vgnd vpwr scs8hd_decap_8
XANTENNA__156__A _156_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ _413_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
+ set vgnd vpwr scs8hd_diode_2
XFILLER_58_439 vpwr vgnd scs8hd_fill_2
XFILLER_38_130 vgnd vpwr scs8hd_decap_12
XFILLER_38_163 vgnd vpwr scs8hd_decap_8
XFILLER_66_483 vgnd vpwr scs8hd_decap_12
XFILLER_26_325 vgnd vpwr scs8hd_fill_1
XFILLER_81_464 vgnd vpwr scs8hd_decap_12
XFILLER_53_144 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _138_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_68 vgnd vpwr scs8hd_decap_12
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
+ _428_/HI vgnd vpwr scs8hd_diode_2
XFILLER_1_424 vgnd vpwr scs8hd_decap_3
XFILLER_39_98 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch/Q ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_57_450 vpwr vgnd scs8hd_fill_2
XFILLER_29_141 vpwr vgnd scs8hd_fill_2
XFILLER_29_163 vgnd vpwr scs8hd_fill_1
XFILLER_17_325 vgnd vpwr scs8hd_decap_4
XFILLER_44_122 vgnd vpwr scs8hd_decap_8
XFILLER_55_86 vgnd vpwr scs8hd_decap_8
XFILLER_17_358 vpwr vgnd scs8hd_fill_2
XFILLER_44_133 vgnd vpwr scs8hd_decap_8
XFILLER_44_144 vgnd vpwr scs8hd_decap_6
XFILLER_32_328 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_391 vpwr vgnd scs8hd_fill_2
XFILLER_71_74 vgnd vpwr scs8hd_decap_12
XFILLER_9_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _156_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_383 vgnd vpwr scs8hd_fill_1
XFILLER_40_394 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__423__B _416_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_258 vpwr vgnd scs8hd_fill_2
XFILLER_67_236 vpwr vgnd scs8hd_fill_2
XFILLER_0_490 vgnd vpwr scs8hd_decap_6
XFILLER_48_450 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_166 vpwr vgnd scs8hd_fill_2
XFILLER_35_177 vpwr vgnd scs8hd_fill_2
XFILLER_35_188 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_50_125 vgnd vpwr scs8hd_decap_4
XANTENNA__317__C _272_/C vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__333__B _326_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_80 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_236 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_461 vpwr vgnd scs8hd_fill_2
XFILLER_46_409 vpwr vgnd scs8hd_fill_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_133 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_23 vgnd vpwr scs8hd_decap_3
XFILLER_14_328 vgnd vpwr scs8hd_decap_8
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_41_114 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_decap_3
XFILLER_41_136 vpwr vgnd scs8hd_fill_2
XPHY_89 vgnd vpwr scs8hd_decap_3
X_190_ address[2] _178_/B _280_/A vgnd vpwr scs8hd_or2_4
XANTENNA__243__B _243_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_210 vpwr vgnd scs8hd_fill_2
XFILLER_1_243 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_501 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_265 vpwr vgnd scs8hd_fill_2
XFILLER_49_203 vpwr vgnd scs8hd_fill_2
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_64_206 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_37_409 vpwr vgnd scs8hd_fill_2
XFILLER_17_111 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__418__B _416_/B vgnd vpwr scs8hd_diode_2
XFILLER_17_199 vgnd vpwr scs8hd_decap_4
XFILLER_9_310 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_388_ _176_/B _391_/B _388_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_40_180 vgnd vpwr scs8hd_decap_3
XFILLER_9_365 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_49_3 vgnd vpwr scs8hd_decap_12
XFILLER_55_228 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__328__B _326_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_136 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _160_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__344__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_59_501 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_74_515 vgnd vpwr scs8hd_fill_1
XFILLER_46_206 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XFILLER_61_209 vgnd vpwr scs8hd_decap_6
XFILLER_27_464 vpwr vgnd scs8hd_fill_2
XFILLER_42_401 vpwr vgnd scs8hd_fill_2
XANTENNA__238__B _243_/B vgnd vpwr scs8hd_diode_2
XFILLER_54_283 vgnd vpwr scs8hd_decap_4
XFILLER_52_32 vgnd vpwr scs8hd_decap_12
X_311_ _247_/A _314_/B _311_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_42_456 vpwr vgnd scs8hd_fill_2
X_242_ _279_/A _243_/B _242_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_331 vgnd vpwr scs8hd_decap_4
X_173_ _202_/A _173_/B _173_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__254__A _263_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_346 vpwr vgnd scs8hd_fill_2
XFILLER_77_62 vgnd vpwr scs8hd_decap_12
XFILLER_77_51 vgnd vpwr scs8hd_decap_8
XFILLER_77_342 vgnd vpwr scs8hd_decap_12
XFILLER_37_217 vgnd vpwr scs8hd_fill_1
XFILLER_37_239 vpwr vgnd scs8hd_fill_2
XFILLER_80_507 vgnd vpwr scs8hd_decap_8
XFILLER_18_442 vgnd vpwr scs8hd_decap_12
XFILLER_45_272 vpwr vgnd scs8hd_fill_2
XFILLER_33_445 vpwr vgnd scs8hd_fill_2
XFILLER_33_456 vpwr vgnd scs8hd_fill_2
XFILLER_33_467 vpwr vgnd scs8hd_fill_2
XFILLER_33_489 vgnd vpwr scs8hd_decap_12
XANTENNA__164__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_13_191 vpwr vgnd scs8hd_fill_2
XFILLER_9_184 vgnd vpwr scs8hd_decap_8
XFILLER_68_320 vgnd vpwr scs8hd_decap_3
XFILLER_68_364 vgnd vpwr scs8hd_decap_12
XFILLER_68_353 vgnd vpwr scs8hd_decap_8
XFILLER_68_342 vpwr vgnd scs8hd_fill_2
XFILLER_28_206 vpwr vgnd scs8hd_fill_2
XANTENNA__339__A _276_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_261 vgnd vpwr scs8hd_decap_12
XPHY_407 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_418 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_429 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_297 vpwr vgnd scs8hd_fill_2
XFILLER_51_286 vpwr vgnd scs8hd_fill_2
XFILLER_11_128 vpwr vgnd scs8hd_fill_2
XFILLER_11_106 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
+ _176_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_68 vgnd vpwr scs8hd_decap_12
XFILLER_3_349 vpwr vgnd scs8hd_fill_2
XFILLER_78_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ _140_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_74_312 vgnd vpwr scs8hd_decap_12
XANTENNA__249__A _231_/A vgnd vpwr scs8hd_diode_2
XFILLER_62_507 vgnd vpwr scs8hd_decap_8
XFILLER_47_98 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_283 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_253 vgnd vpwr scs8hd_decap_3
XFILLER_63_86 vgnd vpwr scs8hd_decap_12
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
XFILLER_15_489 vgnd vpwr scs8hd_decap_12
XFILLER_30_415 vgnd vpwr scs8hd_decap_8
XFILLER_30_426 vgnd vpwr scs8hd_fill_1
X_225_ _280_/A _225_/B _225_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_194 vgnd vpwr scs8hd_decap_4
XFILLER_6_121 vpwr vgnd scs8hd_fill_2
X_156_ _156_/A _156_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_154 vgnd vpwr scs8hd_decap_3
XFILLER_6_187 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _152_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_393 vgnd vpwr scs8hd_decap_4
XFILLER_65_323 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ _139_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_515 vgnd vpwr scs8hd_fill_1
XFILLER_65_356 vgnd vpwr scs8hd_fill_1
XANTENNA__159__A _159_/A vgnd vpwr scs8hd_diode_2
XFILLER_65_367 vgnd vpwr scs8hd_decap_3
XFILLER_80_337 vgnd vpwr scs8hd_decap_12
XFILLER_33_220 vpwr vgnd scs8hd_fill_2
XFILLER_33_231 vpwr vgnd scs8hd_fill_2
XFILLER_21_437 vpwr vgnd scs8hd_fill_2
XFILLER_33_297 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__341__B _343_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_71_304 vgnd vpwr scs8hd_fill_1
XFILLER_56_389 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch_SLEEPB _257_/Y vgnd vpwr scs8hd_diode_2
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_459 vgnd vpwr scs8hd_decap_12
XFILLER_8_419 vgnd vpwr scs8hd_decap_12
XANTENNA__235__C _235_/C vgnd vpwr scs8hd_diode_2
XFILLER_3_102 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/Y _156_/A vgnd vpwr scs8hd_inv_1
XFILLER_79_415 vgnd vpwr scs8hd_decap_12
XANTENNA__251__B _252_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_168 vpwr vgnd scs8hd_fill_2
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XFILLER_59_172 vgnd vpwr scs8hd_decap_4
XFILLER_47_356 vgnd vpwr scs8hd_decap_4
XFILLER_62_337 vpwr vgnd scs8hd_fill_2
XFILLER_15_231 vpwr vgnd scs8hd_fill_2
XPHY_771 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_760 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_392 vgnd vpwr scs8hd_decap_4
XANTENNA__426__B _424_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_223 vgnd vpwr scs8hd_decap_4
XPHY_793 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_782 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_208_ _202_/A _208_/B _208_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_452 vgnd vpwr scs8hd_decap_12
X_139_ _139_/A _139_/Y vgnd vpwr scs8hd_inv_8
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_323 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_378 vgnd vpwr scs8hd_decap_4
XFILLER_53_348 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XFILLER_80_178 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ _135_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_245 vgnd vpwr scs8hd_decap_3
XANTENNA__336__B _343_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_289 vpwr vgnd scs8hd_fill_2
XANTENNA__352__A _280_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch_SLEEPB _229_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_0_105 vpwr vgnd scs8hd_fill_2
XFILLER_29_301 vgnd vpwr scs8hd_fill_1
XFILLER_48_109 vpwr vgnd scs8hd_fill_2
XFILLER_56_120 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _148_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_56 vgnd vpwr scs8hd_decap_12
XFILLER_29_345 vgnd vpwr scs8hd_fill_1
XFILLER_56_142 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
+ _394_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_378 vgnd vpwr scs8hd_decap_4
XFILLER_71_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_44_44 vgnd vpwr scs8hd_decap_12
XFILLER_71_189 vpwr vgnd scs8hd_fill_2
XANTENNA__246__B _252_/B vgnd vpwr scs8hd_diode_2
XFILLER_44_99 vgnd vpwr scs8hd_decap_3
XFILLER_60_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ _387_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__262__A _280_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_79_245 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch_SLEEPB _328_/Y vgnd vpwr scs8hd_diode_2
XFILLER_75_440 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_120 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_164 vpwr vgnd scs8hd_fill_2
XFILLER_35_315 vgnd vpwr scs8hd_decap_6
XFILLER_47_175 vpwr vgnd scs8hd_fill_2
XFILLER_62_145 vgnd vpwr scs8hd_decap_8
XFILLER_35_359 vgnd vpwr scs8hd_decap_4
XFILLER_50_329 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_79_3 vgnd vpwr scs8hd_decap_12
XPHY_590 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__172__A _122_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_66_451 vgnd vpwr scs8hd_decap_6
XFILLER_66_440 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_66_495 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_337 vgnd vpwr scs8hd_decap_4
XFILLER_53_156 vpwr vgnd scs8hd_fill_2
XFILLER_26_348 vgnd vpwr scs8hd_fill_1
XFILLER_81_476 vgnd vpwr scs8hd_decap_12
XANTENNA__347__A _247_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_215 vgnd vpwr scs8hd_decap_12
XFILLER_29_120 vpwr vgnd scs8hd_fill_2
XFILLER_29_153 vgnd vpwr scs8hd_decap_4
XFILLER_72_410 vgnd vpwr scs8hd_decap_12
XFILLER_29_175 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__257__A _247_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_340 vpwr vgnd scs8hd_fill_2
XFILLER_40_362 vpwr vgnd scs8hd_fill_2
XFILLER_71_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch_SLEEPB _301_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_230 vpwr vgnd scs8hd_fill_2
XFILLER_4_285 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_296 vgnd vpwr scs8hd_decap_6
XFILLER_67_226 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
+ _429_/HI vgnd vpwr scs8hd_diode_2
XFILLER_48_462 vpwr vgnd scs8hd_fill_2
XFILLER_82_218 vgnd vpwr scs8hd_decap_12
XFILLER_75_281 vgnd vpwr scs8hd_decap_12
XFILLER_63_421 vpwr vgnd scs8hd_fill_2
XFILLER_63_410 vpwr vgnd scs8hd_fill_2
XFILLER_48_473 vgnd vpwr scs8hd_decap_12
XFILLER_35_123 vgnd vpwr scs8hd_decap_3
XANTENNA__167__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_23_318 vpwr vgnd scs8hd_fill_2
XFILLER_50_148 vgnd vpwr scs8hd_decap_3
XFILLER_31_362 vpwr vgnd scs8hd_fill_2
XANTENNA__317__D _263_/D vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch/Q ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_31_395 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ _157_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_58_215 vpwr vgnd scs8hd_fill_2
XFILLER_58_204 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_451 vpwr vgnd scs8hd_fill_2
XFILLER_54_443 vgnd vpwr scs8hd_decap_4
XPHY_13 vgnd vpwr scs8hd_decap_3
XFILLER_26_123 vgnd vpwr scs8hd_fill_1
XFILLER_26_145 vgnd vpwr scs8hd_decap_6
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XFILLER_77_513 vgnd vpwr scs8hd_decap_3
XFILLER_49_237 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch_SLEEPB _274_/Y vgnd vpwr scs8hd_diode_2
XFILLER_45_454 vgnd vpwr scs8hd_decap_3
XFILLER_72_273 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _447_/HI ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_32_104 vpwr vgnd scs8hd_fill_2
XFILLER_45_476 vgnd vpwr scs8hd_decap_4
XFILLER_45_487 vgnd vpwr scs8hd_fill_1
XFILLER_82_63 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_446 vgnd vpwr scs8hd_decap_12
XFILLER_32_115 vgnd vpwr scs8hd_decap_12
XFILLER_13_351 vpwr vgnd scs8hd_fill_2
XFILLER_13_362 vpwr vgnd scs8hd_fill_2
X_387_ _173_/B _391_/B _387_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
+ _411_/Y vgnd vpwr scs8hd_diode_2
XFILLER_51_424 vgnd vpwr scs8hd_fill_1
XFILLER_23_115 vgnd vpwr scs8hd_decap_6
XANTENNA__344__B _272_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_59 vpwr vgnd scs8hd_fill_2
XANTENNA__360__A _279_/A vgnd vpwr scs8hd_diode_2
XFILLER_59_513 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_39_270 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch/Q ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_281 vpwr vgnd scs8hd_fill_2
XFILLER_54_262 vpwr vgnd scs8hd_fill_2
XFILLER_54_251 vpwr vgnd scs8hd_fill_2
XFILLER_27_487 vgnd vpwr scs8hd_fill_1
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
X_310_ _274_/A _314_/B _310_/Y vgnd vpwr scs8hd_nor2_4
X_241_ _287_/A _243_/B _241_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_52_44 vgnd vpwr scs8hd_decap_12
XFILLER_22_170 vgnd vpwr scs8hd_decap_6
X_172_ _122_/Y _178_/A address[0] _181_/B _173_/B vgnd vpwr scs8hd_or4_4
XANTENNA__254__B _272_/B vgnd vpwr scs8hd_diode_2
XFILLER_10_376 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch_SLEEPB _246_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__270__A _279_/A vgnd vpwr scs8hd_diode_2
XFILLER_77_354 vgnd vpwr scs8hd_decap_12
XFILLER_77_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_454 vgnd vpwr scs8hd_decap_4
XFILLER_45_240 vpwr vgnd scs8hd_fill_2
XFILLER_45_251 vpwr vgnd scs8hd_fill_2
XFILLER_33_413 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch/Q ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_60_276 vgnd vpwr scs8hd_decap_6
XFILLER_20_107 vgnd vpwr scs8hd_decap_4
XFILLER_20_129 vpwr vgnd scs8hd_fill_2
X_439_ _439_/HI _439_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__164__B address[7] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _423_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_163 vpwr vgnd scs8hd_fill_2
XFILLER_61_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_391 vgnd vpwr scs8hd_decap_4
XANTENNA__180__A _202_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch_SLEEPB _345_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_56_505 vgnd vpwr scs8hd_decap_8
XFILLER_68_398 vgnd vpwr scs8hd_decap_8
XFILLER_68_376 vpwr vgnd scs8hd_fill_2
XANTENNA__339__B _343_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_51_221 vpwr vgnd scs8hd_fill_2
XFILLER_24_413 vgnd vpwr scs8hd_decap_12
XPHY_408 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_36_273 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_457 vgnd vpwr scs8hd_fill_1
XPHY_419 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_265 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__355__A _274_/A vgnd vpwr scs8hd_diode_2
XFILLER_78_129 vgnd vpwr scs8hd_decap_12
XFILLER_74_324 vgnd vpwr scs8hd_decap_12
XFILLER_19_207 vpwr vgnd scs8hd_fill_2
XANTENNA__249__B _252_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_402 vpwr vgnd scs8hd_fill_2
XFILLER_27_240 vpwr vgnd scs8hd_fill_2
XFILLER_27_262 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ _180_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_63_98 vgnd vpwr scs8hd_decap_8
XANTENNA__265__A _274_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_276 vpwr vgnd scs8hd_fill_2
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
X_224_ _279_/A _225_/B _224_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_100 vpwr vgnd scs8hd_fill_2
X_155_ _155_/A _155_/Y vgnd vpwr scs8hd_inv_8
Xltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_12_80 vgnd vpwr scs8hd_fill_1
XFILLER_6_166 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch/Q
+ _356_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _147_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_350 vgnd vpwr scs8hd_decap_4
XFILLER_2_383 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_184 vgnd vpwr scs8hd_decap_12
XFILLER_65_335 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch/Q
+ _321_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_80_349 vgnd vpwr scs8hd_decap_12
XFILLER_33_254 vpwr vgnd scs8hd_fill_2
XANTENNA__175__A _122_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch_SLEEPB _318_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _140_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q
+ _286_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch/Q ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_56_302 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_346 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q
+ _250_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_64_390 vgnd vpwr scs8hd_decap_6
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_232 vpwr vgnd scs8hd_fill_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_265 vgnd vpwr scs8hd_decap_3
XANTENNA__235__D _272_/D vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ _148_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_471 vgnd vpwr scs8hd_decap_12
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_302 vgnd vpwr scs8hd_fill_1
XFILLER_74_154 vgnd vpwr scs8hd_decap_12
XFILLER_62_305 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_70_371 vgnd vpwr scs8hd_decap_12
XFILLER_70_360 vgnd vpwr scs8hd_decap_8
XFILLER_15_254 vpwr vgnd scs8hd_fill_2
XPHY_772 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_761 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_750 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_794 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_783 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_257 vpwr vgnd scs8hd_fill_2
X_207_ _181_/C address[1] address[3] address[2] _208_/B vgnd vpwr scs8hd_or4_4
XFILLER_7_464 vgnd vpwr scs8hd_decap_12
X_138_ _138_/A _138_/Y vgnd vpwr scs8hd_inv_8
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch/Q
+ _300_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ _147_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_78_471 vgnd vpwr scs8hd_decap_12
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
XFILLER_65_132 vpwr vgnd scs8hd_fill_2
XFILLER_38_335 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch/Q
+ _265_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_94 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_371 vgnd vpwr scs8hd_fill_1
XFILLER_61_360 vgnd vpwr scs8hd_fill_1
XFILLER_61_393 vgnd vpwr scs8hd_fill_1
XFILLER_21_257 vpwr vgnd scs8hd_fill_2
XFILLER_21_268 vpwr vgnd scs8hd_fill_2
XFILLER_9_92 vpwr vgnd scs8hd_fill_2
XANTENNA__352__B _352_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch/Q
+ _229_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_29_313 vpwr vgnd scs8hd_fill_2
XFILLER_28_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_71_135 vgnd vpwr scs8hd_decap_8
XFILLER_71_179 vgnd vpwr scs8hd_decap_4
XFILLER_44_56 vgnd vpwr scs8hd_decap_12
XFILLER_60_44 vgnd vpwr scs8hd_decap_12
XFILLER_8_239 vgnd vpwr scs8hd_decap_4
XANTENNA__262__B _262_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
XFILLER_79_257 vgnd vpwr scs8hd_decap_12
XFILLER_69_86 vgnd vpwr scs8hd_decap_12
XFILLER_75_452 vgnd vpwr scs8hd_decap_12
XFILLER_35_327 vpwr vgnd scs8hd_fill_2
XFILLER_35_338 vpwr vgnd scs8hd_fill_2
XFILLER_62_157 vgnd vpwr scs8hd_decap_8
XFILLER_50_308 vgnd vpwr scs8hd_decap_6
XFILLER_43_382 vpwr vgnd scs8hd_fill_2
XPHY_580 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_591 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__172__B _178_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch_SLEEPB _298_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_408 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_53_179 vpwr vgnd scs8hd_fill_2
XFILLER_41_319 vgnd vpwr scs8hd_decap_8
XANTENNA__347__B _352_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
XANTENNA__363__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_1_404 vgnd vpwr scs8hd_decap_12
XFILLER_49_419 vpwr vgnd scs8hd_fill_2
XFILLER_76_227 vgnd vpwr scs8hd_decap_12
XFILLER_72_422 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
+ _390_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_187 vpwr vgnd scs8hd_fill_2
XFILLER_17_338 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_55_99 vpwr vgnd scs8hd_fill_2
XANTENNA__257__B _262_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_190 vpwr vgnd scs8hd_fill_2
XFILLER_40_352 vgnd vpwr scs8hd_fill_1
XFILLER_71_98 vgnd vpwr scs8hd_decap_12
XANTENNA__273__A _273_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_400 vgnd vpwr scs8hd_fill_1
XFILLER_48_485 vgnd vpwr scs8hd_decap_12
XFILLER_75_293 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__167__B _166_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch_SLEEPB _271_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_341 vpwr vgnd scs8hd_fill_2
XANTENNA__183__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_374 vpwr vgnd scs8hd_fill_2
XFILLER_6_93 vgnd vpwr scs8hd_decap_4
XFILLER_73_208 vgnd vpwr scs8hd_decap_12
XFILLER_39_485 vgnd vpwr scs8hd_decap_3
XANTENNA__358__A _231_/A vgnd vpwr scs8hd_diode_2
XFILLER_54_422 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_69 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
+ _430_/HI vgnd vpwr scs8hd_diode_2
XFILLER_6_507 vgnd vpwr scs8hd_decap_8
XFILLER_49_216 vpwr vgnd scs8hd_fill_2
XFILLER_66_32 vgnd vpwr scs8hd_decap_12
XFILLER_45_400 vgnd vpwr scs8hd_decap_3
XFILLER_57_293 vpwr vgnd scs8hd_fill_2
XFILLER_57_282 vpwr vgnd scs8hd_fill_2
XANTENNA__268__A _231_/A vgnd vpwr scs8hd_diode_2
XFILLER_82_75 vgnd vpwr scs8hd_decap_12
XFILLER_32_127 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
X_386_ _170_/B _391_/B _386_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_356 vgnd vpwr scs8hd_decap_3
XFILLER_9_345 vpwr vgnd scs8hd_fill_2
XFILLER_9_378 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch_SLEEPB _243_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_411 vgnd vpwr scs8hd_decap_8
XFILLER_63_230 vpwr vgnd scs8hd_fill_2
XANTENNA__178__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_48_293 vgnd vpwr scs8hd_fill_1
XFILLER_63_252 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_296 vgnd vpwr scs8hd_fill_1
XFILLER_23_127 vpwr vgnd scs8hd_fill_2
XFILLER_31_193 vpwr vgnd scs8hd_fill_2
XANTENNA__344__C _163_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_27 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q
+ _351_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__360__B _359_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/Y _137_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch_SLEEPB _342_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_477 vpwr vgnd scs8hd_fill_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _139_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q
+ _316_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_240_ _231_/A _243_/B _240_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_52_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_171_ address[0] _181_/B _171_/X vgnd vpwr scs8hd_or2_4
XANTENNA__254__C _272_/C vgnd vpwr scs8hd_diode_2
XANTENNA__270__B _269_/B vgnd vpwr scs8hd_diode_2
XFILLER_77_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_285 vpwr vgnd scs8hd_fill_2
XFILLER_45_296 vgnd vpwr scs8hd_decap_4
X_438_ _438_/HI _438_/LO vgnd vpwr scs8hd_conb_1
XFILLER_9_142 vpwr vgnd scs8hd_fill_2
XFILLER_13_171 vpwr vgnd scs8hd_fill_2
X_369_ _391_/A _367_/B _369_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XFILLER_54_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_370 vgnd vpwr scs8hd_decap_4
XANTENNA__180__B _367_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_94 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_51_211 vgnd vpwr scs8hd_fill_1
XFILLER_24_425 vgnd vpwr scs8hd_fill_1
XFILLER_36_285 vgnd vpwr scs8hd_decap_3
XPHY_409 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch/Q
+ _330_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_119 vgnd vpwr scs8hd_decap_3
XANTENNA__355__B _359_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XFILLER_32_491 vgnd vpwr scs8hd_decap_12
XANTENNA__371__A _371_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _161_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch_SLEEPB _315_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q
+ _295_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_59_300 vpwr vgnd scs8hd_fill_2
XFILLER_59_333 vgnd vpwr scs8hd_decap_4
XFILLER_59_377 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_414 vgnd vpwr scs8hd_fill_1
XFILLER_27_274 vgnd vpwr scs8hd_decap_6
XFILLER_27_296 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q
+ _260_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__265__B _269_/B vgnd vpwr scs8hd_diode_2
XFILLER_42_288 vgnd vpwr scs8hd_decap_4
X_223_ _287_/A _225_/B _223_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_174 vgnd vpwr scs8hd_decap_3
X_154_ _154_/A _154_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__281__A address[6] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q
+ _224_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_373 vgnd vpwr scs8hd_fill_1
XFILLER_77_196 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
+ _376_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_230 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _157_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_391 vgnd vpwr scs8hd_decap_12
XANTENNA__175__B _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_277 vgnd vpwr scs8hd_fill_1
XANTENNA__191__A _122_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_152 vgnd vpwr scs8hd_fill_1
XFILLER_68_141 vgnd vpwr scs8hd_decap_4
XFILLER_56_314 vpwr vgnd scs8hd_fill_2
XFILLER_56_325 vpwr vgnd scs8hd_fill_2
XFILLER_71_306 vgnd vpwr scs8hd_decap_4
XFILLER_56_369 vgnd vpwr scs8hd_decap_8
XFILLER_56_358 vgnd vpwr scs8hd_fill_1
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XFILLER_44_509 vgnd vpwr scs8hd_decap_6
XFILLER_71_317 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch_SLEEPB _288_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_59 vpwr vgnd scs8hd_fill_2
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__366__A _176_/B vgnd vpwr scs8hd_diode_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_483 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _148_/Y vgnd vpwr scs8hd_diode_2
XFILLER_79_428 vgnd vpwr scs8hd_decap_12
XFILLER_58_44 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _141_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_47_325 vgnd vpwr scs8hd_fill_1
XFILLER_74_166 vgnd vpwr scs8hd_decap_12
XFILLER_74_32 vgnd vpwr scs8hd_decap_12
XFILLER_15_211 vgnd vpwr scs8hd_fill_1
XANTENNA__276__A _276_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_762 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_751 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_740 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_383 vgnd vpwr scs8hd_decap_6
XFILLER_15_288 vgnd vpwr scs8hd_decap_4
XPHY_795 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_784 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_773 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch/Q ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_247 vgnd vpwr scs8hd_fill_1
XFILLER_30_269 vgnd vpwr scs8hd_decap_6
X_206_ _202_/A _377_/A _206_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_476 vgnd vpwr scs8hd_decap_12
X_137_ _137_/A _137_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_192 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_78_483 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XFILLER_65_177 vgnd vpwr scs8hd_decap_4
XFILLER_65_166 vpwr vgnd scs8hd_fill_2
XFILLER_53_328 vgnd vpwr scs8hd_decap_3
XFILLER_53_317 vpwr vgnd scs8hd_fill_2
XANTENNA__186__A _202_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
+ _369_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_236 vpwr vgnd scs8hd_fill_2
XFILLER_0_129 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_336 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _446_/HI ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_44_328 vgnd vpwr scs8hd_decap_8
XFILLER_71_147 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ _156_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_44_68 vgnd vpwr scs8hd_decap_12
XFILLER_52_383 vgnd vpwr scs8hd_decap_4
XFILLER_52_372 vpwr vgnd scs8hd_fill_2
XFILLER_60_56 vgnd vpwr scs8hd_decap_12
XFILLER_20_291 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _135_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/Y _139_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_4_457 vgnd vpwr scs8hd_fill_1
XFILLER_69_98 vgnd vpwr scs8hd_decap_12
XFILLER_79_269 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch_SLEEPB _359_/Y vgnd vpwr scs8hd_diode_2
XFILLER_75_464 vgnd vpwr scs8hd_decap_12
XFILLER_47_144 vgnd vpwr scs8hd_decap_4
XFILLER_18_80 vgnd vpwr scs8hd_decap_12
XFILLER_31_501 vgnd vpwr scs8hd_decap_12
XFILLER_43_350 vpwr vgnd scs8hd_fill_2
XPHY_570 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_592 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_581 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_240 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_284 vpwr vgnd scs8hd_fill_2
XANTENNA__172__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_66_420 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_114 vpwr vgnd scs8hd_fill_2
XFILLER_53_103 vpwr vgnd scs8hd_fill_2
XFILLER_26_328 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_136 vpwr vgnd scs8hd_fill_2
XFILLER_81_489 vgnd vpwr scs8hd_decap_12
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_394 vgnd vpwr scs8hd_decap_3
XANTENNA__363__B _362_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
+ _415_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_416 vgnd vpwr scs8hd_decap_8
XFILLER_76_239 vgnd vpwr scs8hd_decap_12
XFILLER_17_306 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_72_434 vgnd vpwr scs8hd_decap_12
XFILLER_29_199 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch/Q ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_501 vgnd vpwr scs8hd_decap_12
XFILLER_44_158 vpwr vgnd scs8hd_fill_2
XFILLER_44_169 vgnd vpwr scs8hd_decap_4
XFILLER_25_372 vpwr vgnd scs8hd_fill_2
XANTENNA__273__B _280_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_40_386 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ _152_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_210 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_254 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_67_206 vpwr vgnd scs8hd_fill_2
XFILLER_29_90 vpwr vgnd scs8hd_fill_2
XFILLER_63_445 vpwr vgnd scs8hd_fill_2
XFILLER_63_434 vpwr vgnd scs8hd_fill_2
XFILLER_35_114 vpwr vgnd scs8hd_fill_2
XFILLER_48_497 vgnd vpwr scs8hd_decap_12
XFILLER_63_489 vgnd vpwr scs8hd_decap_12
XFILLER_23_309 vgnd vpwr scs8hd_decap_3
XFILLER_50_117 vgnd vpwr scs8hd_decap_6
XFILLER_16_372 vpwr vgnd scs8hd_fill_2
XFILLER_31_331 vgnd vpwr scs8hd_decap_6
XFILLER_43_180 vgnd vpwr scs8hd_decap_3
XANTENNA__183__B _183_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _153_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _131_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _443_/HI ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_66_250 vpwr vgnd scs8hd_fill_2
XFILLER_81_220 vgnd vpwr scs8hd_decap_12
XANTENNA__358__B _359_/B vgnd vpwr scs8hd_diode_2
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XFILLER_14_309 vgnd vpwr scs8hd_decap_8
XPHY_37 vgnd vpwr scs8hd_decap_3
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_25_59 vpwr vgnd scs8hd_fill_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XANTENNA__374__A _200_/B vgnd vpwr scs8hd_diode_2
XFILLER_10_515 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_202 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_235 vpwr vgnd scs8hd_fill_2
XFILLER_66_44 vgnd vpwr scs8hd_decap_12
XFILLER_57_250 vpwr vgnd scs8hd_fill_2
XFILLER_45_412 vgnd vpwr scs8hd_decap_4
XFILLER_72_231 vgnd vpwr scs8hd_decap_12
XANTENNA__268__B _269_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_136 vpwr vgnd scs8hd_fill_2
XFILLER_45_423 vpwr vgnd scs8hd_fill_2
XFILLER_82_32 vgnd vpwr scs8hd_decap_12
XFILLER_45_489 vgnd vpwr scs8hd_decap_12
XFILLER_82_87 vgnd vpwr scs8hd_decap_6
XFILLER_60_459 vgnd vpwr scs8hd_decap_12
XANTENNA__284__A _247_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_139 vpwr vgnd scs8hd_fill_2
X_385_ address[4] _384_/X _391_/B vgnd vpwr scs8hd_or2_4
XFILLER_9_324 vgnd vpwr scs8hd_decap_4
XFILLER_9_302 vgnd vpwr scs8hd_fill_1
XFILLER_13_386 vgnd vpwr scs8hd_decap_4
XFILLER_40_161 vpwr vgnd scs8hd_fill_2
XFILLER_40_172 vgnd vpwr scs8hd_decap_8
XFILLER_40_194 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
+ _431_/HI vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ _132_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_515 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch/Q ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__178__B _178_/B vgnd vpwr scs8hd_diode_2
XFILLER_63_264 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch_SLEEPB _218_/Y vgnd vpwr scs8hd_diode_2
XFILLER_63_275 vpwr vgnd scs8hd_fill_2
XFILLER_51_459 vpwr vgnd scs8hd_fill_2
XFILLER_16_191 vpwr vgnd scs8hd_fill_2
XANTENNA__194__A _202_/A vgnd vpwr scs8hd_diode_2
XANTENNA__344__D _272_/D vgnd vpwr scs8hd_diode_2
XFILLER_11_39 vgnd vpwr scs8hd_decap_12
XANTENNA__369__A _391_/A vgnd vpwr scs8hd_diode_2
XFILLER_74_507 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ _131_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_401 vgnd vpwr scs8hd_decap_3
XFILLER_54_220 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch/Q ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_423 vpwr vgnd scs8hd_fill_2
XFILLER_39_294 vgnd vpwr scs8hd_decap_6
XFILLER_27_445 vpwr vgnd scs8hd_fill_2
XFILLER_14_128 vpwr vgnd scs8hd_fill_2
XFILLER_27_489 vgnd vpwr scs8hd_decap_12
XFILLER_42_426 vpwr vgnd scs8hd_fill_2
XFILLER_42_448 vgnd vpwr scs8hd_decap_8
XFILLER_42_459 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_50_470 vgnd vpwr scs8hd_decap_8
XFILLER_52_68 vgnd vpwr scs8hd_decap_12
XFILLER_50_481 vgnd vpwr scs8hd_decap_12
XFILLER_10_323 vgnd vpwr scs8hd_fill_1
X_170_ _202_/A _170_/B _170_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__254__D _272_/D vgnd vpwr scs8hd_diode_2
XFILLER_6_305 vgnd vpwr scs8hd_fill_1
XFILLER_10_389 vgnd vpwr scs8hd_decap_8
XFILLER_6_327 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _149_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__279__A _279_/A vgnd vpwr scs8hd_diode_2
XFILLER_77_367 vgnd vpwr scs8hd_decap_12
XFILLER_77_98 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_209 vpwr vgnd scs8hd_fill_2
XFILLER_18_423 vgnd vpwr scs8hd_decap_8
XFILLER_60_245 vgnd vpwr scs8hd_fill_1
XFILLER_26_80 vgnd vpwr scs8hd_decap_12
XFILLER_60_267 vgnd vpwr scs8hd_decap_4
XFILLER_13_150 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_437_ _437_/HI _437_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_368_ _183_/B _367_/B _368_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_470 vpwr vgnd scs8hd_fill_2
X_299_ _263_/A address[7] _272_/C _263_/D _304_/B vgnd vpwr scs8hd_or4_4
XFILLER_5_360 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_3 vgnd vpwr scs8hd_decap_12
XFILLER_68_301 vgnd vpwr scs8hd_decap_4
XFILLER_3_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XFILLER_68_389 vgnd vpwr scs8hd_decap_8
XANTENNA__189__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_253 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_437 vgnd vpwr scs8hd_decap_4
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XANTENNA__371__B _367_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_319 vpwr vgnd scs8hd_fill_2
XFILLER_59_367 vgnd vpwr scs8hd_fill_1
XFILLER_59_356 vgnd vpwr scs8hd_decap_4
XFILLER_74_337 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_42_212 vpwr vgnd scs8hd_fill_2
XFILLER_42_267 vpwr vgnd scs8hd_fill_2
X_222_ _231_/A _225_/B _222_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_131 vgnd vpwr scs8hd_fill_1
XFILLER_10_186 vgnd vpwr scs8hd_decap_6
XFILLER_6_113 vgnd vpwr scs8hd_decap_8
X_153_ _153_/A _153_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__281__B _272_/B vgnd vpwr scs8hd_diode_2
XFILLER_12_93 vpwr vgnd scs8hd_fill_2
XFILLER_2_363 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_507 vgnd vpwr scs8hd_decap_8
XFILLER_65_359 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
+ _208_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_253 vgnd vpwr scs8hd_decap_4
XFILLER_33_201 vpwr vgnd scs8hd_fill_2
XFILLER_18_297 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__175__C _181_/C vgnd vpwr scs8hd_diode_2
XFILLER_21_418 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__191__B _280_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ _381_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_212 vpwr vgnd scs8hd_fill_2
XANTENNA__366__B _367_/B vgnd vpwr scs8hd_diode_2
XFILLER_12_407 vgnd vpwr scs8hd_decap_12
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XANTENNA__382__A _187_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_495 vgnd vpwr scs8hd_decap_12
XFILLER_58_56 vgnd vpwr scs8hd_decap_12
XFILLER_59_142 vpwr vgnd scs8hd_fill_2
XFILLER_59_131 vpwr vgnd scs8hd_fill_2
XFILLER_59_197 vpwr vgnd scs8hd_fill_2
XFILLER_47_348 vpwr vgnd scs8hd_fill_2
XFILLER_74_178 vgnd vpwr scs8hd_decap_12
XFILLER_74_44 vgnd vpwr scs8hd_decap_12
XANTENNA__276__B _280_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_223 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_763 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_752 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_741 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_730 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_215 vpwr vgnd scs8hd_fill_2
XPHY_796 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_785 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_774 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_440 vgnd vpwr scs8hd_decap_12
XANTENNA__292__A _274_/A vgnd vpwr scs8hd_diode_2
X_205_ address[0] _181_/B address[3] address[2] _377_/A vgnd vpwr scs8hd_or4_4
XFILLER_23_92 vpwr vgnd scs8hd_fill_2
X_136_ _136_/A _136_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_495 vgnd vpwr scs8hd_decap_12
XFILLER_65_145 vpwr vgnd scs8hd_fill_2
XFILLER_38_348 vgnd vpwr scs8hd_decap_12
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XANTENNA__186__B _391_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_226 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ _200_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_69_440 vgnd vpwr scs8hd_decap_12
XFILLER_56_101 vpwr vgnd scs8hd_fill_2
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_304 vgnd vpwr scs8hd_fill_1
XFILLER_29_359 vgnd vpwr scs8hd_decap_4
XFILLER_56_189 vgnd vpwr scs8hd_decap_3
XANTENNA__377__A _377_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_259 vgnd vpwr scs8hd_decap_12
XFILLER_12_237 vgnd vpwr scs8hd_decap_12
XFILLER_8_219 vgnd vpwr scs8hd_decap_3
XFILLER_60_68 vgnd vpwr scs8hd_decap_12
XFILLER_4_403 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2/Z
+ _149_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_47_123 vgnd vpwr scs8hd_decap_4
XFILLER_75_476 vgnd vpwr scs8hd_decap_12
XANTENNA__287__A _287_/A vgnd vpwr scs8hd_diode_2
XFILLER_62_137 vpwr vgnd scs8hd_fill_2
XFILLER_28_392 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_31_513 vgnd vpwr scs8hd_decap_3
XFILLER_43_395 vpwr vgnd scs8hd_fill_2
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
XPHY_560 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_571 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_593 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_582 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_281 vgnd vpwr scs8hd_decap_4
XANTENNA__172__D _181_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_263 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_145 vgnd vpwr scs8hd_decap_6
XANTENNA__197__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_53_148 vpwr vgnd scs8hd_fill_2
XFILLER_38_189 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_373 vgnd vpwr scs8hd_decap_3
XFILLER_61_192 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_428 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_57_454 vgnd vpwr scs8hd_decap_4
XFILLER_57_443 vpwr vgnd scs8hd_fill_2
XFILLER_29_123 vgnd vpwr scs8hd_decap_3
XFILLER_29_145 vgnd vpwr scs8hd_fill_1
XFILLER_72_446 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_513 vgnd vpwr scs8hd_decap_3
XFILLER_25_362 vpwr vgnd scs8hd_fill_2
XFILLER_25_395 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_398 vpwr vgnd scs8hd_fill_2
XFILLER_20_93 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_340 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ _418_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_362 vgnd vpwr scs8hd_fill_1
XFILLER_45_90 vgnd vpwr scs8hd_fill_1
XFILLER_77_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_390 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_465 vgnd vpwr scs8hd_decap_12
XFILLER_54_413 vgnd vpwr scs8hd_decap_6
XFILLER_26_115 vgnd vpwr scs8hd_decap_8
XFILLER_81_232 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_25_27 vgnd vpwr scs8hd_decap_12
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_41_118 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__374__B _367_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_365 vpwr vgnd scs8hd_fill_2
XFILLER_22_398 vgnd vpwr scs8hd_decap_6
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XANTENNA__390__A _183_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_214 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ _425_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_269 vpwr vgnd scs8hd_fill_2
XFILLER_66_56 vgnd vpwr scs8hd_decap_12
XFILLER_72_221 vgnd vpwr scs8hd_fill_1
XFILLER_17_115 vgnd vpwr scs8hd_fill_1
XFILLER_72_254 vgnd vpwr scs8hd_decap_4
XFILLER_72_243 vgnd vpwr scs8hd_decap_8
XFILLER_82_44 vgnd vpwr scs8hd_decap_12
XFILLER_72_276 vgnd vpwr scs8hd_fill_1
XFILLER_72_265 vgnd vpwr scs8hd_decap_8
XANTENNA__284__B _286_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_321 vpwr vgnd scs8hd_fill_2
XFILLER_13_376 vgnd vpwr scs8hd_decap_4
XFILLER_15_82 vgnd vpwr scs8hd_decap_3
X_384_ _263_/A address[7] _163_/X _263_/D _384_/X vgnd vpwr scs8hd_or4_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _132_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_457 vgnd vpwr scs8hd_fill_1
XFILLER_36_468 vgnd vpwr scs8hd_decap_12
XFILLER_51_416 vpwr vgnd scs8hd_fill_2
XFILLER_51_405 vpwr vgnd scs8hd_fill_2
XFILLER_23_107 vpwr vgnd scs8hd_fill_2
XFILLER_51_449 vgnd vpwr scs8hd_decap_3
XFILLER_16_170 vgnd vpwr scs8hd_decap_8
XANTENNA__194__B _194_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_162 vpwr vgnd scs8hd_fill_2
XFILLER_8_391 vgnd vpwr scs8hd_decap_6
XFILLER_8_380 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__369__B _367_/B vgnd vpwr scs8hd_diode_2
XFILLER_54_210 vgnd vpwr scs8hd_decap_4
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_54_243 vpwr vgnd scs8hd_fill_2
XANTENNA__385__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_42_405 vgnd vpwr scs8hd_decap_4
XFILLER_54_298 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch/Q ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_50_493 vgnd vpwr scs8hd_decap_12
XFILLER_10_335 vgnd vpwr scs8hd_fill_1
XFILLER_10_368 vgnd vpwr scs8hd_decap_6
XFILLER_10_346 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ _396_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_77_379 vgnd vpwr scs8hd_decap_12
XANTENNA__279__B _280_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
+ _186_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_402 vgnd vpwr scs8hd_decap_4
XANTENNA__295__A _231_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_60_224 vpwr vgnd scs8hd_fill_2
XFILLER_33_449 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_436_ _436_/HI _436_/LO vgnd vpwr scs8hd_conb_1
XFILLER_41_460 vgnd vpwr scs8hd_fill_1
XFILLER_9_111 vgnd vpwr scs8hd_decap_4
X_367_ _367_/A _367_/B _367_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_195 vgnd vpwr scs8hd_decap_4
XFILLER_42_80 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ _140_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_298_ _280_/A _295_/B _298_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_3_74 vgnd vpwr scs8hd_decap_12
XANTENNA__189__B _189_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _445_/HI ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_36_243 vpwr vgnd scs8hd_fill_2
XFILLER_24_449 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _150_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_313 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ _139_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_74_349 vgnd vpwr scs8hd_decap_12
XFILLER_27_221 vpwr vgnd scs8hd_fill_2
XFILLER_27_254 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_221_ _276_/A _225_/B _221_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_110 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_152_ _152_/A _152_/Y vgnd vpwr scs8hd_inv_8
XFILLER_10_154 vpwr vgnd scs8hd_fill_2
XFILLER_6_125 vpwr vgnd scs8hd_fill_2
XANTENNA__281__C _272_/C vgnd vpwr scs8hd_diode_2
XFILLER_10_198 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch_SLEEPB _260_/Y vgnd vpwr scs8hd_diode_2
XFILLER_77_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_65_327 vgnd vpwr scs8hd_decap_3
XFILLER_18_276 vpwr vgnd scs8hd_fill_2
XFILLER_33_224 vpwr vgnd scs8hd_fill_2
XFILLER_33_235 vpwr vgnd scs8hd_fill_2
XANTENNA__175__D address[1] vgnd vpwr scs8hd_diode_2
X_419_ _202_/B _416_/B _419_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_471 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_180 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _136_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_154 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_39 vgnd vpwr scs8hd_decap_12
XFILLER_64_382 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch/Q ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_419 vgnd vpwr scs8hd_decap_12
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_290 vgnd vpwr scs8hd_decap_3
XANTENNA__382__B _380_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ _374_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_58_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_187 vpwr vgnd scs8hd_fill_2
XFILLER_74_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_55_382 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XPHY_720 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_753 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_742 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_396 vgnd vpwr scs8hd_fill_1
XPHY_731 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch_SLEEPB _232_/Y vgnd vpwr scs8hd_diode_2
XPHY_786 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_775 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_764 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_204_ _202_/A _204_/B _204_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_797 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_452 vgnd vpwr scs8hd_decap_12
XANTENNA__292__B _295_/B vgnd vpwr scs8hd_diode_2
X_135_ _135_/A _135_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_489 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
+ _397_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _442_/HI ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_65_102 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_80_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XFILLER_46_371 vgnd vpwr scs8hd_decap_8
XFILLER_61_363 vgnd vpwr scs8hd_decap_3
XFILLER_61_341 vpwr vgnd scs8hd_fill_2
XFILLER_61_396 vpwr vgnd scs8hd_fill_2
XFILLER_61_385 vpwr vgnd scs8hd_fill_2
XFILLER_9_62 vgnd vpwr scs8hd_decap_12
XFILLER_9_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch_SLEEPB _331_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_109 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_452 vgnd vpwr scs8hd_decap_12
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XFILLER_56_146 vgnd vpwr scs8hd_fill_1
XFILLER_56_157 vgnd vpwr scs8hd_decap_12
XANTENNA__377__B _367_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_15 vgnd vpwr scs8hd_decap_12
XFILLER_52_341 vpwr vgnd scs8hd_fill_2
XFILLER_52_396 vgnd vpwr scs8hd_fill_1
XANTENNA__393__A _371_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_249 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch/Q
+ _345_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_260 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_415 vgnd vpwr scs8hd_decap_12
XFILLER_4_459 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch/Q
+ _310_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_47_113 vgnd vpwr scs8hd_decap_4
XANTENNA__287__B _286_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_360 vgnd vpwr scs8hd_decap_8
XFILLER_47_168 vpwr vgnd scs8hd_fill_2
XFILLER_47_179 vpwr vgnd scs8hd_fill_2
XFILLER_18_93 vpwr vgnd scs8hd_fill_2
XFILLER_43_363 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch/Q
+ _275_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_550 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_561 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_594 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_583 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_572 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_50_80 vgnd vpwr scs8hd_decap_12
XFILLER_7_297 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch/Q
+ _239_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch/Q ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_81_403 vgnd vpwr scs8hd_decap_12
XANTENNA__197__B _197_/B vgnd vpwr scs8hd_diode_2
XFILLER_26_308 vpwr vgnd scs8hd_fill_2
XFILLER_26_319 vgnd vpwr scs8hd_decap_6
XFILLER_19_382 vpwr vgnd scs8hd_fill_2
XFILLER_19_393 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch_SLEEPB _304_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _158_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_352 vpwr vgnd scs8hd_fill_2
XFILLER_34_385 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _131_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XFILLER_69_293 vgnd vpwr scs8hd_decap_8
XANTENNA__388__A _176_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_179 vpwr vgnd scs8hd_fill_2
XFILLER_44_105 vgnd vpwr scs8hd_decap_8
XFILLER_40_344 vgnd vpwr scs8hd_decap_8
XFILLER_40_366 vpwr vgnd scs8hd_fill_2
XFILLER_4_267 vgnd vpwr scs8hd_decap_8
XFILLER_4_234 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _439_/HI ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_289 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__298__A _280_/A vgnd vpwr scs8hd_diode_2
XFILLER_48_466 vpwr vgnd scs8hd_fill_2
XFILLER_63_425 vpwr vgnd scs8hd_fill_2
XFILLER_35_149 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch/Q
+ _218_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_380 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_391 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_399 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch_SLEEPB _277_/Y vgnd vpwr scs8hd_diode_2
XFILLER_58_219 vpwr vgnd scs8hd_fill_2
XFILLER_58_208 vgnd vpwr scs8hd_decap_6
XFILLER_39_400 vpwr vgnd scs8hd_fill_2
XFILLER_39_455 vgnd vpwr scs8hd_decap_4
XFILLER_39_477 vgnd vpwr scs8hd_decap_8
XFILLER_54_469 vpwr vgnd scs8hd_fill_2
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_25_39 vgnd vpwr scs8hd_decap_12
XFILLER_34_193 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
+ _189_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_377 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XANTENNA__390__B _391_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_248 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_68 vgnd vpwr scs8hd_decap_12
XFILLER_57_263 vpwr vgnd scs8hd_fill_2
XFILLER_72_200 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_82_56 vgnd vpwr scs8hd_decap_6
XFILLER_60_417 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_383_ _178_/B _380_/X _383_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_193 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_152 vgnd vpwr scs8hd_fill_1
XFILLER_15_94 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2/A
+ ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch/Q ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_48_285 vgnd vpwr scs8hd_decap_8
XFILLER_36_447 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch_SLEEPB _249_/Y vgnd vpwr scs8hd_diode_2
XFILLER_63_288 vpwr vgnd scs8hd_fill_2
XFILLER_51_428 vgnd vpwr scs8hd_decap_4
XFILLER_16_160 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_63_299 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XFILLER_39_274 vgnd vpwr scs8hd_fill_1
XFILLER_54_266 vpwr vgnd scs8hd_fill_2
XANTENNA__385__B _384_/X vgnd vpwr scs8hd_diode_2
XFILLER_52_15 vgnd vpwr scs8hd_decap_12
XFILLER_22_196 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch_SLEEPB _348_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_200 vpwr vgnd scs8hd_fill_2
XANTENNA__295__B _295_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_428 vpwr vgnd scs8hd_fill_2
XFILLER_33_417 vpwr vgnd scs8hd_fill_2
XFILLER_45_255 vpwr vgnd scs8hd_fill_2
XFILLER_26_93 vgnd vpwr scs8hd_decap_3
XFILLER_26_480 vgnd vpwr scs8hd_decap_12
X_435_ _435_/HI _435_/LO vgnd vpwr scs8hd_conb_1
XFILLER_9_134 vpwr vgnd scs8hd_fill_2
X_366_ _176_/B _367_/B _366_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_167 vpwr vgnd scs8hd_fill_2
X_297_ _279_/A _295_/B _297_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_86 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ _133_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q
+ _361_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_51_203 vpwr vgnd scs8hd_fill_2
XFILLER_51_236 vpwr vgnd scs8hd_fill_2
XFILLER_51_269 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch_SLEEPB _321_/Y vgnd vpwr scs8hd_diode_2
XFILLER_47_59 vpwr vgnd scs8hd_fill_2
XANTENNA__396__A _200_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_406 vgnd vpwr scs8hd_decap_8
XFILLER_15_417 vpwr vgnd scs8hd_fill_2
XFILLER_42_203 vgnd vpwr scs8hd_decap_3
XFILLER_15_428 vgnd vpwr scs8hd_decap_12
XFILLER_42_225 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_461 vgnd vpwr scs8hd_decap_12
X_220_ _247_/A _225_/B _220_/Y vgnd vpwr scs8hd_nor2_4
X_151_ _151_/A _151_/Y vgnd vpwr scs8hd_inv_8
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/Y _159_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__281__D _263_/D vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_12_84 vgnd vpwr scs8hd_decap_8
XFILLER_2_387 vgnd vpwr scs8hd_decap_4
XFILLER_65_339 vpwr vgnd scs8hd_fill_2
XFILLER_65_306 vpwr vgnd scs8hd_fill_2
XFILLER_61_501 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ _148_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_258 vgnd vpwr scs8hd_decap_4
X_418_ _200_/B _416_/B _418_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_483 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q
+ _340_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_349_ _231_/A _352_/B _349_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_52_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_68_177 vgnd vpwr scs8hd_decap_12
XFILLER_68_166 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q
+ _305_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_380 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q
+ _270_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ _366_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_59_155 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q
+ _234_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_47_317 vpwr vgnd scs8hd_fill_2
XFILLER_74_68 vgnd vpwr scs8hd_decap_12
XFILLER_55_361 vgnd vpwr scs8hd_decap_3
XFILLER_43_501 vgnd vpwr scs8hd_decap_12
XFILLER_82_180 vgnd vpwr scs8hd_decap_6
XFILLER_15_203 vpwr vgnd scs8hd_fill_2
XPHY_710 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_236 vpwr vgnd scs8hd_fill_2
XFILLER_15_269 vpwr vgnd scs8hd_fill_2
XPHY_754 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_743 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_732 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_721 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_30_206 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_787 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_776 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_765 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_203_ address[3] _231_/A _204_/B vgnd vpwr scs8hd_or2_4
XPHY_798 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_464 vgnd vpwr scs8hd_decap_12
XFILLER_7_402 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_134_ _134_/A _134_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_151 vpwr vgnd scs8hd_fill_2
XFILLER_65_114 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_136 vpwr vgnd scs8hd_fill_2
XFILLER_48_80 vgnd vpwr scs8hd_decap_12
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _156_/Y vgnd vpwr scs8hd_diode_2
XFILLER_80_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_87 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ _155_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_280 vgnd vpwr scs8hd_decap_3
XFILLER_9_74 vgnd vpwr scs8hd_decap_4
XFILLER_69_464 vgnd vpwr scs8hd_decap_12
XFILLER_29_317 vpwr vgnd scs8hd_fill_2
XFILLER_56_125 vgnd vpwr scs8hd_decap_8
XFILLER_29_339 vgnd vpwr scs8hd_decap_6
XFILLER_56_169 vgnd vpwr scs8hd_fill_1
XFILLER_25_501 vgnd vpwr scs8hd_decap_12
XFILLER_44_27 vgnd vpwr scs8hd_decap_4
XFILLER_12_206 vpwr vgnd scs8hd_fill_2
XANTENNA__393__B _391_/B vgnd vpwr scs8hd_diode_2
XFILLER_40_504 vgnd vpwr scs8hd_decap_12
XFILLER_60_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_250 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_427 vgnd vpwr scs8hd_decap_12
XFILLER_75_489 vgnd vpwr scs8hd_decap_12
XPHY_540 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_551 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_562 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_595 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_584 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_573 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_34_93 vgnd vpwr scs8hd_decap_8
XFILLER_7_221 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
XFILLER_81_415 vgnd vpwr scs8hd_decap_12
XFILLER_22_515 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_27 vgnd vpwr scs8hd_decap_12
XFILLER_57_412 vpwr vgnd scs8hd_fill_2
XFILLER_29_103 vpwr vgnd scs8hd_fill_2
XFILLER_69_272 vpwr vgnd scs8hd_fill_2
XFILLER_57_423 vpwr vgnd scs8hd_fill_2
XANTENNA__388__B _391_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_114 vgnd vpwr scs8hd_decap_4
XFILLER_55_15 vgnd vpwr scs8hd_decap_12
XFILLER_57_489 vgnd vpwr scs8hd_decap_12
XFILLER_55_59 vpwr vgnd scs8hd_fill_2
XFILLER_72_459 vgnd vpwr scs8hd_decap_12
XFILLER_37_180 vgnd vpwr scs8hd_decap_3
XFILLER_52_172 vgnd vpwr scs8hd_fill_1
XFILLER_40_334 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_220 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__298__B _295_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _444_/HI ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_106 vgnd vpwr scs8hd_decap_3
XFILLER_28_180 vgnd vpwr scs8hd_decap_4
XFILLER_35_139 vpwr vgnd scs8hd_fill_2
XFILLER_31_301 vpwr vgnd scs8hd_fill_2
XFILLER_31_323 vpwr vgnd scs8hd_fill_2
XPHY_370 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_345 vpwr vgnd scs8hd_fill_2
XFILLER_31_378 vpwr vgnd scs8hd_fill_2
XPHY_381 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_392 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_97 vgnd vpwr scs8hd_fill_1
XFILLER_3_290 vgnd vpwr scs8hd_decap_3
XFILLER_39_434 vpwr vgnd scs8hd_fill_2
XFILLER_39_489 vgnd vpwr scs8hd_decap_12
XFILLER_81_245 vgnd vpwr scs8hd_decap_12
XFILLER_54_459 vgnd vpwr scs8hd_fill_1
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_507 vgnd vpwr scs8hd_decap_8
XFILLER_22_389 vpwr vgnd scs8hd_fill_2
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__399__A _377_/A vgnd vpwr scs8hd_diode_2
XFILLER_72_212 vpwr vgnd scs8hd_fill_2
XFILLER_57_286 vpwr vgnd scs8hd_fill_2
XFILLER_57_297 vpwr vgnd scs8hd_fill_2
XFILLER_45_437 vpwr vgnd scs8hd_fill_2
XFILLER_45_459 vpwr vgnd scs8hd_fill_2
XFILLER_60_429 vpwr vgnd scs8hd_fill_2
XFILLER_53_470 vpwr vgnd scs8hd_fill_2
X_382_ _187_/B _380_/X _382_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_334 vpwr vgnd scs8hd_fill_2
XFILLER_15_51 vgnd vpwr scs8hd_decap_8
XFILLER_15_62 vgnd vpwr scs8hd_decap_12
XFILLER_40_120 vgnd vpwr scs8hd_decap_3
XFILLER_9_349 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/Y _131_/A vgnd vpwr scs8hd_buf_1
XFILLER_31_94 vgnd vpwr scs8hd_fill_1
XFILLER_68_507 vgnd vpwr scs8hd_decap_8
XFILLER_63_234 vpwr vgnd scs8hd_fill_2
XFILLER_63_223 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch/Q ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_56_80 vgnd vpwr scs8hd_decap_12
XFILLER_63_256 vgnd vpwr scs8hd_fill_1
XFILLER_82_3 vgnd vpwr scs8hd_decap_12
XFILLER_31_175 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_231 vpwr vgnd scs8hd_fill_2
XFILLER_27_415 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_437 vpwr vgnd scs8hd_fill_2
XFILLER_14_109 vpwr vgnd scs8hd_fill_2
XFILLER_42_418 vgnd vpwr scs8hd_decap_8
XFILLER_52_27 vgnd vpwr scs8hd_decap_4
XFILLER_22_142 vgnd vpwr scs8hd_decap_4
XFILLER_10_315 vpwr vgnd scs8hd_fill_2
XFILLER_10_304 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ _412_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_319 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _441_/HI ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
+ clk ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff/QN
+ reset set vgnd vpwr scs8hd_dfbbp_1
XFILLER_18_459 vgnd vpwr scs8hd_decap_12
XFILLER_45_245 vgnd vpwr scs8hd_decap_3
X_434_ _434_/HI _434_/LO vgnd vpwr scs8hd_conb_1
XFILLER_26_492 vgnd vpwr scs8hd_decap_12
XFILLER_45_289 vpwr vgnd scs8hd_fill_2
XFILLER_60_248 vgnd vpwr scs8hd_decap_4
XFILLER_13_142 vpwr vgnd scs8hd_fill_2
XFILLER_13_175 vpwr vgnd scs8hd_fill_2
X_365_ _173_/B _367_/B _365_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_146 vpwr vgnd scs8hd_fill_2
X_296_ _287_/A _295_/B _296_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_93 vgnd vpwr scs8hd_decap_4
XFILLER_5_374 vgnd vpwr scs8hd_fill_1
XFILLER_5_352 vpwr vgnd scs8hd_fill_2
XFILLER_68_337 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_98 vpwr vgnd scs8hd_fill_2
XFILLER_36_212 vpwr vgnd scs8hd_fill_2
XFILLER_51_248 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _379_/Y vgnd vpwr scs8hd_diode_2
XFILLER_59_304 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _155_/Y vgnd vpwr scs8hd_diode_2
XFILLER_59_348 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_47_27 vgnd vpwr scs8hd_decap_12
XANTENNA__396__B _391_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_234 vgnd vpwr scs8hd_decap_4
XFILLER_63_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_82_373 vgnd vpwr scs8hd_decap_12
XFILLER_42_215 vgnd vpwr scs8hd_decap_8
XFILLER_63_59 vpwr vgnd scs8hd_fill_2
XFILLER_23_451 vpwr vgnd scs8hd_fill_2
XFILLER_23_473 vgnd vpwr scs8hd_decap_12
XFILLER_10_134 vpwr vgnd scs8hd_fill_2
X_150_ _150_/A _150_/Y vgnd vpwr scs8hd_inv_8
XFILLER_10_145 vgnd vpwr scs8hd_decap_8
XFILLER_6_138 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_123 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch/Q ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_58_370 vgnd vpwr scs8hd_decap_4
XFILLER_18_267 vgnd vpwr scs8hd_decap_8
XFILLER_61_513 vgnd vpwr scs8hd_decap_3
X_417_ _197_/B _416_/B _417_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_495 vgnd vpwr scs8hd_decap_12
X_348_ _276_/A _352_/B _348_/Y vgnd vpwr scs8hd_nor2_4
X_279_ _279_/A _280_/B _279_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ _141_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_45_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_68_145 vgnd vpwr scs8hd_fill_1
XFILLER_56_329 vpwr vgnd scs8hd_fill_2
XFILLER_24_204 vgnd vpwr scs8hd_decap_8
XFILLER_24_226 vgnd vpwr scs8hd_decap_4
XFILLER_24_237 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _438_/HI ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_112 vpwr vgnd scs8hd_fill_2
XFILLER_58_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_123 vgnd vpwr scs8hd_fill_1
XFILLER_59_178 vpwr vgnd scs8hd_fill_2
XFILLER_47_329 vpwr vgnd scs8hd_fill_2
XANTENNA__200__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_43_513 vgnd vpwr scs8hd_decap_3
XPHY_711 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_700 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_248 vgnd vpwr scs8hd_decap_4
XPHY_744 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_733 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_722 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_777 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_766 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_755 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_398 vgnd vpwr scs8hd_decap_6
XFILLER_23_281 vpwr vgnd scs8hd_fill_2
XFILLER_23_292 vgnd vpwr scs8hd_decap_3
X_202_ _202_/A _202_/B _202_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_229 vpwr vgnd scs8hd_fill_2
XPHY_799 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_788 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_51 vgnd vpwr scs8hd_decap_8
XFILLER_23_62 vgnd vpwr scs8hd_decap_12
XFILLER_11_476 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
X_133_ _133_/A _133_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_410 vgnd vpwr scs8hd_decap_12
XFILLER_2_196 vgnd vpwr scs8hd_decap_4
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ _156_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_80_129 vgnd vpwr scs8hd_decap_12
XFILLER_64_80 vgnd vpwr scs8hd_decap_12
XFILLER_61_354 vgnd vpwr scs8hd_decap_6
XFILLER_21_218 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _133_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_14_292 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_476 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _137_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_340 vpwr vgnd scs8hd_fill_2
XFILLER_52_310 vgnd vpwr scs8hd_fill_1
XFILLER_25_513 vgnd vpwr scs8hd_decap_3
XFILLER_37_362 vgnd vpwr scs8hd_fill_1
XFILLER_37_384 vgnd vpwr scs8hd_decap_3
XFILLER_64_181 vgnd vpwr scs8hd_decap_4
XFILLER_52_387 vgnd vpwr scs8hd_fill_1
XFILLER_52_376 vpwr vgnd scs8hd_fill_2
XFILLER_12_218 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_398 vpwr vgnd scs8hd_fill_2
XFILLER_60_27 vgnd vpwr scs8hd_decap_4
XFILLER_4_439 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch/Q ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_340 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_148 vgnd vpwr scs8hd_fill_1
XFILLER_62_118 vgnd vpwr scs8hd_fill_1
XFILLER_70_162 vgnd vpwr scs8hd_decap_3
XFILLER_43_354 vgnd vpwr scs8hd_decap_3
XFILLER_70_195 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
+ _418_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_530 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_541 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_552 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_596 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_585 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_574 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_563 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_50_93 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_251 vgnd vpwr scs8hd_decap_12
XFILLER_66_413 vgnd vpwr scs8hd_decap_4
XFILLER_38_126 vpwr vgnd scs8hd_fill_2
XFILLER_66_457 vgnd vpwr scs8hd_fill_1
XFILLER_19_340 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_53_118 vpwr vgnd scs8hd_fill_2
XFILLER_53_107 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_162 vpwr vgnd scs8hd_fill_2
XFILLER_34_365 vpwr vgnd scs8hd_fill_2
XFILLER_61_184 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_398 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _435_/HI ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_39 vgnd vpwr scs8hd_decap_12
XFILLER_69_251 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_137 vpwr vgnd scs8hd_fill_2
XFILLER_29_159 vgnd vpwr scs8hd_decap_4
XFILLER_55_27 vgnd vpwr scs8hd_decap_12
XFILLER_25_343 vpwr vgnd scs8hd_fill_2
XFILLER_80_471 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _151_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_354 vpwr vgnd scs8hd_fill_2
XFILLER_25_376 vpwr vgnd scs8hd_fill_2
XFILLER_71_15 vgnd vpwr scs8hd_decap_12
XFILLER_40_313 vpwr vgnd scs8hd_fill_2
XFILLER_71_59 vpwr vgnd scs8hd_fill_2
XFILLER_40_379 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_497 vgnd vpwr scs8hd_decap_12
XFILLER_48_435 vpwr vgnd scs8hd_fill_2
XFILLER_75_232 vgnd vpwr scs8hd_decap_12
XFILLER_48_446 vpwr vgnd scs8hd_fill_2
XFILLER_35_118 vpwr vgnd scs8hd_fill_2
XFILLER_63_449 vgnd vpwr scs8hd_decap_12
XFILLER_63_438 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_376 vgnd vpwr scs8hd_decap_4
XFILLER_43_140 vpwr vgnd scs8hd_fill_2
XFILLER_43_162 vgnd vpwr scs8hd_decap_3
XFILLER_43_184 vpwr vgnd scs8hd_fill_2
XFILLER_45_93 vpwr vgnd scs8hd_fill_2
XPHY_360 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_371 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_382 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_393 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_66_254 vgnd vpwr scs8hd_decap_4
XFILLER_66_276 vgnd vpwr scs8hd_decap_4
XFILLER_26_107 vgnd vpwr scs8hd_decap_6
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_81_257 vgnd vpwr scs8hd_decap_12
XFILLER_34_151 vpwr vgnd scs8hd_fill_2
XFILLER_62_471 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _159_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ _132_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_206 vpwr vgnd scs8hd_fill_2
XFILLER_1_239 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch_SLEEPB _221_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__399__B _391_/B vgnd vpwr scs8hd_diode_2
XFILLER_66_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_243 vgnd vpwr scs8hd_fill_1
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_416 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_25_140 vpwr vgnd scs8hd_fill_2
XFILLER_25_151 vpwr vgnd scs8hd_fill_2
X_381_ _171_/X _380_/X _381_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_302 vgnd vpwr scs8hd_decap_3
XFILLER_25_162 vpwr vgnd scs8hd_fill_2
XFILLER_9_306 vpwr vgnd scs8hd_fill_2
XFILLER_15_74 vgnd vpwr scs8hd_decap_8
XFILLER_40_143 vgnd vpwr scs8hd_fill_1
XFILLER_40_154 vpwr vgnd scs8hd_fill_2
XFILLER_40_165 vgnd vpwr scs8hd_decap_4
XFILLER_21_390 vpwr vgnd scs8hd_fill_2
XFILLER_40_198 vgnd vpwr scs8hd_decap_4
XFILLER_5_501 vgnd vpwr scs8hd_decap_12
XFILLER_31_51 vgnd vpwr scs8hd_decap_8
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_272 vgnd vpwr scs8hd_fill_1
XFILLER_48_210 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_63_202 vpwr vgnd scs8hd_fill_2
XFILLER_48_254 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_72_80 vgnd vpwr scs8hd_decap_12
XFILLER_16_195 vgnd vpwr scs8hd_decap_4
XFILLER_31_132 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _147_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ _386_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_75_3 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_187 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_8_383 vgnd vpwr scs8hd_fill_1
XFILLER_39_254 vpwr vgnd scs8hd_fill_2
XFILLER_54_224 vgnd vpwr scs8hd_decap_4
XFILLER_54_279 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_290 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_22_154 vgnd vpwr scs8hd_decap_3
XFILLER_10_327 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ _139_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_515 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__203__A address[3] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_45_213 vgnd vpwr scs8hd_decap_4
XFILLER_45_268 vpwr vgnd scs8hd_fill_2
X_433_ _433_/HI _433_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_154 vpwr vgnd scs8hd_fill_2
X_364_ _170_/B _367_/B _364_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_452 vpwr vgnd scs8hd_fill_2
XFILLER_41_474 vgnd vpwr scs8hd_decap_12
X_295_ _231_/A _295_/B _295_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch_SLEEPB _293_/Y vgnd vpwr scs8hd_diode_2
XFILLER_68_316 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_39 vgnd vpwr scs8hd_decap_12
XFILLER_67_393 vgnd vpwr scs8hd_decap_4
XFILLER_82_385 vgnd vpwr scs8hd_decap_12
XFILLER_63_27 vgnd vpwr scs8hd_decap_12
XFILLER_42_238 vpwr vgnd scs8hd_fill_2
XFILLER_42_249 vpwr vgnd scs8hd_fill_2
XFILLER_23_485 vgnd vpwr scs8hd_decap_3
XFILLER_2_301 vgnd vpwr scs8hd_decap_4
XFILLER_2_312 vgnd vpwr scs8hd_decap_6
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_367 vgnd vpwr scs8hd_decap_6
XFILLER_77_135 vgnd vpwr scs8hd_decap_12
XFILLER_58_393 vgnd vpwr scs8hd_decap_4
XFILLER_18_202 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_330 vgnd vpwr scs8hd_decap_12
XFILLER_18_257 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch_SLEEPB _266_/Y vgnd vpwr scs8hd_diode_2
XFILLER_33_205 vgnd vpwr scs8hd_decap_4
X_416_ _194_/B _416_/B _416_/Y vgnd vpwr scs8hd_nor2_4
X_347_ _247_/A _352_/B _347_/Y vgnd vpwr scs8hd_nor2_4
X_278_ _287_/A _280_/B _278_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_172 vpwr vgnd scs8hd_fill_2
XFILLER_5_150 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _156_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_68_124 vgnd vpwr scs8hd_decap_8
XFILLER_56_308 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_190 vgnd vpwr scs8hd_decap_12
XFILLER_64_352 vpwr vgnd scs8hd_fill_2
XFILLER_64_396 vgnd vpwr scs8hd_fill_1
XFILLER_24_249 vgnd vpwr scs8hd_fill_1
XFILLER_20_411 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_74_105 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ _210_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_74_15 vgnd vpwr scs8hd_decap_12
XANTENNA__200__B _200_/B vgnd vpwr scs8hd_diode_2
XPHY_701 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ _150_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_227 vpwr vgnd scs8hd_fill_2
XPHY_745 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_734 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_723 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_712 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_219 vgnd vpwr scs8hd_fill_1
XPHY_778 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_767 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_756 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_400 vgnd vpwr scs8hd_fill_1
X_201_ address[3] _276_/A _202_/B vgnd vpwr scs8hd_or2_4
XPHY_789 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_132_ _132_/A _132_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_426 vgnd vpwr scs8hd_fill_1
XFILLER_23_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch_SLEEPB _238_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_422 vgnd vpwr scs8hd_decap_12
XFILLER_2_175 vgnd vpwr scs8hd_decap_6
XFILLER_38_319 vpwr vgnd scs8hd_fill_2
XFILLER_48_93 vpwr vgnd scs8hd_fill_2
XFILLER_65_149 vpwr vgnd scs8hd_fill_2
XFILLER_73_171 vgnd vpwr scs8hd_decap_12
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_61_333 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_80_80 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/Y _136_/A vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__301__A _274_/A vgnd vpwr scs8hd_diode_2
XFILLER_56_105 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch_SLEEPB _337_/Y vgnd vpwr scs8hd_diode_2
XFILLER_56_149 vgnd vpwr scs8hd_decap_4
XFILLER_37_352 vgnd vpwr scs8hd_fill_1
XFILLER_52_355 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_69_15 vgnd vpwr scs8hd_decap_12
XFILLER_79_208 vgnd vpwr scs8hd_decap_12
XFILLER_69_59 vpwr vgnd scs8hd_fill_2
XFILLER_75_403 vgnd vpwr scs8hd_decap_12
XANTENNA__211__A _380_/A vgnd vpwr scs8hd_diode_2
XFILLER_47_127 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_55_160 vgnd vpwr scs8hd_decap_4
XFILLER_55_193 vpwr vgnd scs8hd_fill_2
XFILLER_28_396 vgnd vpwr scs8hd_fill_1
XFILLER_43_333 vpwr vgnd scs8hd_fill_2
XFILLER_70_141 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _134_/Y vgnd vpwr scs8hd_diode_2
XPHY_520 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_399 vpwr vgnd scs8hd_fill_2
XPHY_531 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_542 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_553 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XPHY_586 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_575 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_241 vgnd vpwr scs8hd_fill_1
XPHY_564 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_597 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_263 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_285 vgnd vpwr scs8hd_fill_1
XFILLER_7_245 vpwr vgnd scs8hd_fill_2
XFILLER_7_267 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_440 vgnd vpwr scs8hd_decap_12
XFILLER_78_263 vgnd vpwr scs8hd_decap_12
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XFILLER_81_428 vgnd vpwr scs8hd_decap_12
XFILLER_19_363 vgnd vpwr scs8hd_fill_1
XFILLER_34_311 vgnd vpwr scs8hd_decap_8
XFILLER_46_171 vpwr vgnd scs8hd_fill_2
XFILLER_46_182 vpwr vgnd scs8hd_fill_2
XFILLER_61_152 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ _176_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_61_196 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch_SLEEPB _310_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ _423_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch/Q
+ _355_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _440_/HI ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_458 vgnd vpwr scs8hd_fill_1
XFILLER_29_149 vpwr vgnd scs8hd_fill_2
XFILLER_55_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch/Q
+ _320_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_160 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/Y _154_/A vgnd vpwr scs8hd_inv_1
XFILLER_25_311 vpwr vgnd scs8hd_fill_2
XFILLER_80_483 vgnd vpwr scs8hd_decap_12
XFILLER_71_27 vgnd vpwr scs8hd_decap_12
XFILLER_52_163 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__206__A _202_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch/Q
+ _285_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_215 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _139_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
+ _371_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_51 vgnd vpwr scs8hd_decap_8
XFILLER_29_62 vgnd vpwr scs8hd_decap_12
XFILLER_48_403 vpwr vgnd scs8hd_fill_2
XFILLER_48_414 vgnd vpwr scs8hd_decap_3
XFILLER_48_425 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q
+ _249_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_63_428 vgnd vpwr scs8hd_decap_3
XFILLER_63_417 vpwr vgnd scs8hd_fill_2
XFILLER_63_406 vpwr vgnd scs8hd_fill_2
XFILLER_16_322 vpwr vgnd scs8hd_fill_2
XFILLER_16_344 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_174 vgnd vpwr scs8hd_decap_4
XPHY_350 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_361 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_358 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_372 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_383 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_394 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_66_233 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch_SLEEPB _283_/Y vgnd vpwr scs8hd_diode_2
XFILLER_54_439 vpwr vgnd scs8hd_fill_2
XFILLER_81_269 vgnd vpwr scs8hd_decap_12
XFILLER_62_483 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_369 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_229 vgnd vpwr scs8hd_decap_4
XFILLER_66_27 vgnd vpwr scs8hd_decap_4
XFILLER_57_211 vpwr vgnd scs8hd_fill_2
XFILLER_57_200 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch/Q ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch/Q
+ _264_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_82_15 vgnd vpwr scs8hd_decap_12
XFILLER_60_409 vgnd vpwr scs8hd_decap_8
X_380_ _380_/A _362_/X _380_/X vgnd vpwr scs8hd_or2_4
XFILLER_13_325 vpwr vgnd scs8hd_fill_2
XFILLER_13_347 vpwr vgnd scs8hd_fill_2
XFILLER_13_358 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch/Q
+ _228_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_513 vgnd vpwr scs8hd_decap_3
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_48_233 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_93 vgnd vpwr scs8hd_decap_4
XFILLER_29_480 vgnd vpwr scs8hd_decap_8
XFILLER_51_409 vpwr vgnd scs8hd_fill_2
XFILLER_44_450 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ _401_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_152 vgnd vpwr scs8hd_fill_1
XFILLER_71_280 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
+ _364_/Y vgnd vpwr scs8hd_diode_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_68_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _437_/HI ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
.ends

