magic
tech sky130A
magscale 1 2
timestamp 1606423406
<< locali >>
rect 19073 20927 19107 21029
rect 14841 20247 14875 20349
rect 7849 19907 7883 20009
rect 3801 18615 3835 18921
rect 2237 18071 2271 18173
rect 9781 18071 9815 18241
rect 9413 16507 9447 16677
rect 17693 16575 17727 16745
rect 21281 16575 21315 16677
rect 6101 16031 6135 16133
rect 6653 15895 6687 16133
rect 8861 16031 8895 16201
rect 9505 15351 9539 15657
rect 13001 15419 13035 15657
rect 16681 14467 16715 14569
rect 3893 14331 3927 14433
rect 9413 14263 9447 14365
rect 18981 14263 19015 14433
rect 3985 13719 4019 14025
rect 19533 13855 19567 14025
rect 8309 13175 8343 13413
rect 14105 12767 14139 12869
rect 17601 12835 17635 12937
rect 17509 12631 17543 12801
rect 10793 12291 10827 12393
rect 4905 12087 4939 12189
rect 11253 12087 11287 12257
rect 11345 12155 11379 12257
rect 12633 11067 12667 11305
rect 12633 9911 12667 10149
rect 14749 9911 14783 10217
rect 20361 9979 20395 10217
rect 7481 9367 7515 9605
rect 8401 8891 8435 9061
rect 3801 8415 3835 8585
rect 9597 8347 9631 8585
rect 15393 8347 15427 8517
rect 13001 7871 13035 8041
rect 9413 7735 9447 7837
rect 13461 6783 13495 6953
rect 17141 6647 17175 6749
rect 17693 6647 17727 6749
rect 17141 6613 17233 6647
rect 20361 6647 20395 6749
rect 14657 6239 14691 6341
rect 21281 5559 21315 5661
rect 11805 4471 11839 4573
rect 14473 3927 14507 4165
rect 16221 3927 16255 4097
rect 15945 3383 15979 3689
rect 16037 3451 16071 3553
rect 16129 2839 16163 3145
<< viali >>
rect 1593 21641 1627 21675
rect 9965 21641 9999 21675
rect 15485 21641 15519 21675
rect 18521 21641 18555 21675
rect 13645 21573 13679 21607
rect 21189 21573 21223 21607
rect 2605 21505 2639 21539
rect 3617 21505 3651 21539
rect 4629 21505 4663 21539
rect 6377 21505 6411 21539
rect 7481 21505 7515 21539
rect 8953 21505 8987 21539
rect 13277 21505 13311 21539
rect 14197 21505 14231 21539
rect 16129 21505 16163 21539
rect 17049 21505 17083 21539
rect 21833 21505 21867 21539
rect 1409 21437 1443 21471
rect 5089 21437 5123 21471
rect 9781 21437 9815 21471
rect 10701 21437 10735 21471
rect 13093 21437 13127 21471
rect 14841 21437 14875 21471
rect 15945 21437 15979 21471
rect 17693 21437 17727 21471
rect 18337 21437 18371 21471
rect 18889 21437 18923 21471
rect 20545 21437 20579 21471
rect 22201 21437 22235 21471
rect 2329 21369 2363 21403
rect 6193 21369 6227 21403
rect 7941 21369 7975 21403
rect 8861 21369 8895 21403
rect 10968 21369 11002 21403
rect 13001 21369 13035 21403
rect 14013 21369 14047 21403
rect 19156 21369 19190 21403
rect 1961 21301 1995 21335
rect 2421 21301 2455 21335
rect 2973 21301 3007 21335
rect 3341 21301 3375 21335
rect 3433 21301 3467 21335
rect 4077 21301 4111 21335
rect 4445 21301 4479 21335
rect 4537 21301 4571 21335
rect 5273 21301 5307 21335
rect 5825 21301 5859 21335
rect 6285 21301 6319 21335
rect 6929 21301 6963 21335
rect 7297 21301 7331 21335
rect 7389 21301 7423 21335
rect 8401 21301 8435 21335
rect 8769 21301 8803 21335
rect 12081 21301 12115 21335
rect 12633 21301 12667 21335
rect 14105 21301 14139 21335
rect 15025 21301 15059 21335
rect 15853 21301 15887 21335
rect 16497 21301 16531 21335
rect 16865 21301 16899 21335
rect 16957 21301 16991 21335
rect 17877 21301 17911 21335
rect 20269 21301 20303 21335
rect 20729 21301 20763 21335
rect 21557 21301 21591 21335
rect 21649 21301 21683 21335
rect 22385 21301 22419 21335
rect 1593 21097 1627 21131
rect 4445 21097 4479 21131
rect 7205 21097 7239 21131
rect 8953 21097 8987 21131
rect 17141 21097 17175 21131
rect 20545 21097 20579 21131
rect 4537 21029 4571 21063
rect 7818 21029 7852 21063
rect 10149 21029 10183 21063
rect 11336 21029 11370 21063
rect 13360 21029 13394 21063
rect 19073 21029 19107 21063
rect 19432 21029 19466 21063
rect 21180 21029 21214 21063
rect 1409 20961 1443 20995
rect 2228 20961 2262 20995
rect 5089 20961 5123 20995
rect 6092 20961 6126 20995
rect 10057 20961 10091 20995
rect 13093 20961 13127 20995
rect 15557 20961 15591 20995
rect 16957 20961 16991 20995
rect 17509 20961 17543 20995
rect 17776 20961 17810 20995
rect 1961 20893 1995 20927
rect 4721 20893 4755 20927
rect 5825 20893 5859 20927
rect 7573 20893 7607 20927
rect 10241 20893 10275 20927
rect 11069 20893 11103 20927
rect 15301 20893 15335 20927
rect 19073 20893 19107 20927
rect 19165 20893 19199 20927
rect 20913 20893 20947 20927
rect 5273 20825 5307 20859
rect 3341 20757 3375 20791
rect 4077 20757 4111 20791
rect 9689 20757 9723 20791
rect 12449 20757 12483 20791
rect 14473 20757 14507 20791
rect 16681 20757 16715 20791
rect 18889 20757 18923 20791
rect 22293 20757 22327 20791
rect 3065 20553 3099 20587
rect 4813 20553 4847 20587
rect 6469 20553 6503 20587
rect 8217 20553 8251 20587
rect 9873 20553 9907 20587
rect 11805 20553 11839 20587
rect 12909 20553 12943 20587
rect 14657 20553 14691 20587
rect 19441 20553 19475 20587
rect 5089 20417 5123 20451
rect 6837 20417 6871 20451
rect 17049 20417 17083 20451
rect 17141 20417 17175 20451
rect 20177 20417 20211 20451
rect 20361 20417 20395 20451
rect 1685 20349 1719 20383
rect 3433 20349 3467 20383
rect 3700 20349 3734 20383
rect 5356 20349 5390 20383
rect 7104 20349 7138 20383
rect 8493 20349 8527 20383
rect 10425 20349 10459 20383
rect 10692 20349 10726 20383
rect 12725 20349 12759 20383
rect 13277 20349 13311 20383
rect 13544 20349 13578 20383
rect 14841 20349 14875 20383
rect 14933 20349 14967 20383
rect 15200 20349 15234 20383
rect 18061 20349 18095 20383
rect 20821 20349 20855 20383
rect 21088 20349 21122 20383
rect 22477 20349 22511 20383
rect 1952 20281 1986 20315
rect 8760 20281 8794 20315
rect 16957 20281 16991 20315
rect 18328 20281 18362 20315
rect 20085 20281 20119 20315
rect 14841 20213 14875 20247
rect 16313 20213 16347 20247
rect 16589 20213 16623 20247
rect 19717 20213 19751 20247
rect 22201 20213 22235 20247
rect 22661 20213 22695 20247
rect 3249 20009 3283 20043
rect 6561 20009 6595 20043
rect 7849 20009 7883 20043
rect 11805 20009 11839 20043
rect 13461 20009 13495 20043
rect 14013 20009 14047 20043
rect 19165 20009 19199 20043
rect 19901 20009 19935 20043
rect 4690 19941 4724 19975
rect 6653 19941 6687 19975
rect 9689 19941 9723 19975
rect 15660 19941 15694 19975
rect 17233 19941 17267 19975
rect 19809 19941 19843 19975
rect 1676 19873 1710 19907
rect 3065 19873 3099 19907
rect 7389 19873 7423 19907
rect 7849 19873 7883 19907
rect 7941 19873 7975 19907
rect 8208 19873 8242 19907
rect 9873 19873 9907 19907
rect 10692 19873 10726 19907
rect 12081 19873 12115 19907
rect 12348 19873 12382 19907
rect 13921 19873 13955 19907
rect 17049 19873 17083 19907
rect 17785 19873 17819 19907
rect 18052 19873 18086 19907
rect 21649 19873 21683 19907
rect 22293 19873 22327 19907
rect 22477 19873 22511 19907
rect 1409 19805 1443 19839
rect 4445 19805 4479 19839
rect 6837 19805 6871 19839
rect 10425 19805 10459 19839
rect 14197 19805 14231 19839
rect 14657 19805 14691 19839
rect 14749 19805 14783 19839
rect 15393 19805 15427 19839
rect 20085 19805 20119 19839
rect 21741 19805 21775 19839
rect 21833 19805 21867 19839
rect 5825 19737 5859 19771
rect 2789 19669 2823 19703
rect 6193 19669 6227 19703
rect 7573 19669 7607 19703
rect 9321 19669 9355 19703
rect 10057 19669 10091 19703
rect 13553 19669 13587 19703
rect 16773 19669 16807 19703
rect 17417 19669 17451 19703
rect 19441 19669 19475 19703
rect 21281 19669 21315 19703
rect 22661 19669 22695 19703
rect 4445 19465 4479 19499
rect 14289 19465 14323 19499
rect 13921 19397 13955 19431
rect 19441 19397 19475 19431
rect 3065 19329 3099 19363
rect 5365 19329 5399 19363
rect 6285 19329 6319 19363
rect 8125 19329 8159 19363
rect 10885 19329 10919 19363
rect 11897 19329 11931 19363
rect 13093 19329 13127 19363
rect 14749 19329 14783 19363
rect 14933 19329 14967 19363
rect 15853 19329 15887 19363
rect 16865 19329 16899 19363
rect 20269 19329 20303 19363
rect 1409 19261 1443 19295
rect 3332 19261 3366 19295
rect 5089 19261 5123 19295
rect 6193 19261 6227 19295
rect 7021 19261 7055 19295
rect 7941 19261 7975 19295
rect 8585 19261 8619 19295
rect 12817 19261 12851 19295
rect 13737 19261 13771 19295
rect 15669 19261 15703 19295
rect 16681 19261 16715 19295
rect 17417 19261 17451 19295
rect 18061 19261 18095 19295
rect 20177 19261 20211 19295
rect 21005 19261 21039 19295
rect 21272 19261 21306 19295
rect 1676 19193 1710 19227
rect 5181 19193 5215 19227
rect 6101 19193 6135 19227
rect 8830 19193 8864 19227
rect 12909 19193 12943 19227
rect 15761 19193 15795 19227
rect 18328 19193 18362 19227
rect 20085 19193 20119 19227
rect 2789 19125 2823 19159
rect 4721 19125 4755 19159
rect 5733 19125 5767 19159
rect 7205 19125 7239 19159
rect 7573 19125 7607 19159
rect 8033 19125 8067 19159
rect 9965 19125 9999 19159
rect 10333 19125 10367 19159
rect 10701 19125 10735 19159
rect 10793 19125 10827 19159
rect 11345 19125 11379 19159
rect 11713 19125 11747 19159
rect 11805 19125 11839 19159
rect 12449 19125 12483 19159
rect 14657 19125 14691 19159
rect 15301 19125 15335 19159
rect 16313 19125 16347 19159
rect 16773 19125 16807 19159
rect 17601 19125 17635 19159
rect 19717 19125 19751 19159
rect 22385 19125 22419 19159
rect 3801 18921 3835 18955
rect 4077 18921 4111 18955
rect 4445 18921 4479 18955
rect 9321 18921 9355 18955
rect 11621 18921 11655 18955
rect 16773 18921 16807 18955
rect 17049 18921 17083 18955
rect 18889 18921 18923 18955
rect 19533 18921 19567 18955
rect 22661 18921 22695 18955
rect 1777 18785 1811 18819
rect 2596 18785 2630 18819
rect 2329 18717 2363 18751
rect 4537 18853 4571 18887
rect 8208 18853 8242 18887
rect 14013 18853 14047 18887
rect 15660 18853 15694 18887
rect 17776 18853 17810 18887
rect 19625 18853 19659 18887
rect 21548 18853 21582 18887
rect 5457 18785 5491 18819
rect 6285 18785 6319 18819
rect 7205 18785 7239 18819
rect 9689 18785 9723 18819
rect 10508 18785 10542 18819
rect 11897 18785 11931 18819
rect 12164 18785 12198 18819
rect 13921 18785 13955 18819
rect 14657 18785 14691 18819
rect 15393 18785 15427 18819
rect 20177 18785 20211 18819
rect 4629 18717 4663 18751
rect 5549 18717 5583 18751
rect 5733 18717 5767 18751
rect 7297 18717 7331 18751
rect 7481 18717 7515 18751
rect 7941 18717 7975 18751
rect 10241 18717 10275 18751
rect 14197 18717 14231 18751
rect 17509 18717 17543 18751
rect 19809 18717 19843 18751
rect 21281 18717 21315 18751
rect 14841 18649 14875 18683
rect 1961 18581 1995 18615
rect 3709 18581 3743 18615
rect 3801 18581 3835 18615
rect 5089 18581 5123 18615
rect 6469 18581 6503 18615
rect 6837 18581 6871 18615
rect 9873 18581 9907 18615
rect 13277 18581 13311 18615
rect 13553 18581 13587 18615
rect 19165 18581 19199 18615
rect 20361 18581 20395 18615
rect 1961 18377 1995 18411
rect 4169 18377 4203 18411
rect 9965 18377 9999 18411
rect 11621 18377 11655 18411
rect 14381 18377 14415 18411
rect 16681 18377 16715 18411
rect 19441 18377 19475 18411
rect 3709 18309 3743 18343
rect 7297 18309 7331 18343
rect 17693 18309 17727 18343
rect 4537 18241 4571 18275
rect 7757 18241 7791 18275
rect 7941 18241 7975 18275
rect 9781 18241 9815 18275
rect 10241 18241 10275 18275
rect 15209 18241 15243 18275
rect 16221 18241 16255 18275
rect 17233 18241 17267 18275
rect 18061 18241 18095 18275
rect 20913 18241 20947 18275
rect 1777 18173 1811 18207
rect 2237 18173 2271 18207
rect 2329 18173 2363 18207
rect 3985 18173 4019 18207
rect 6193 18173 6227 18207
rect 8309 18173 8343 18207
rect 2596 18105 2630 18139
rect 4804 18105 4838 18139
rect 7665 18105 7699 18139
rect 8576 18105 8610 18139
rect 10149 18173 10183 18207
rect 12449 18173 12483 18207
rect 13001 18173 13035 18207
rect 16037 18173 16071 18207
rect 17141 18173 17175 18207
rect 17877 18173 17911 18207
rect 19809 18173 19843 18207
rect 21373 18173 21407 18207
rect 21640 18173 21674 18207
rect 10508 18105 10542 18139
rect 13268 18105 13302 18139
rect 15025 18105 15059 18139
rect 16129 18105 16163 18139
rect 18328 18105 18362 18139
rect 20729 18105 20763 18139
rect 2237 18037 2271 18071
rect 5917 18037 5951 18071
rect 6377 18037 6411 18071
rect 6837 18037 6871 18071
rect 9689 18037 9723 18071
rect 9781 18037 9815 18071
rect 11897 18037 11931 18071
rect 12633 18037 12667 18071
rect 14657 18037 14691 18071
rect 15117 18037 15151 18071
rect 15669 18037 15703 18071
rect 17049 18037 17083 18071
rect 19993 18037 20027 18071
rect 20361 18037 20395 18071
rect 20821 18037 20855 18071
rect 22753 18037 22787 18071
rect 14289 17833 14323 17867
rect 14841 17833 14875 17867
rect 18797 17833 18831 17867
rect 19533 17833 19567 17867
rect 10600 17765 10634 17799
rect 15546 17765 15580 17799
rect 16957 17765 16991 17799
rect 19441 17765 19475 17799
rect 21180 17765 21214 17799
rect 1685 17697 1719 17731
rect 2237 17697 2271 17731
rect 2504 17697 2538 17731
rect 4261 17697 4295 17731
rect 5069 17697 5103 17731
rect 6725 17697 6759 17731
rect 8493 17697 8527 17731
rect 9689 17697 9723 17731
rect 12357 17697 12391 17731
rect 12916 17697 12950 17731
rect 13176 17697 13210 17731
rect 14657 17697 14691 17731
rect 17417 17697 17451 17731
rect 17684 17697 17718 17731
rect 20269 17697 20303 17731
rect 22569 17697 22603 17731
rect 4813 17629 4847 17663
rect 6469 17629 6503 17663
rect 8585 17629 8619 17663
rect 8677 17629 8711 17663
rect 9137 17629 9171 17663
rect 10333 17629 10367 17663
rect 15301 17629 15335 17663
rect 19717 17629 19751 17663
rect 20913 17629 20947 17663
rect 3617 17561 3651 17595
rect 9873 17561 9907 17595
rect 11713 17561 11747 17595
rect 12541 17561 12575 17595
rect 1869 17493 1903 17527
rect 4445 17493 4479 17527
rect 6193 17493 6227 17527
rect 7849 17493 7883 17527
rect 8125 17493 8159 17527
rect 16681 17493 16715 17527
rect 19073 17493 19107 17527
rect 20453 17493 20487 17527
rect 22293 17493 22327 17527
rect 3525 17289 3559 17323
rect 11713 17289 11747 17323
rect 14013 17289 14047 17323
rect 16497 17289 16531 17323
rect 16957 17289 16991 17323
rect 3801 17221 3835 17255
rect 4813 17221 4847 17255
rect 9873 17221 9907 17255
rect 14841 17221 14875 17255
rect 22201 17221 22235 17255
rect 4445 17153 4479 17187
rect 5365 17153 5399 17187
rect 12633 17153 12667 17187
rect 17601 17153 17635 17187
rect 19257 17153 19291 17187
rect 20269 17153 20303 17187
rect 20453 17153 20487 17187
rect 1593 17085 1627 17119
rect 2145 17085 2179 17119
rect 4169 17085 4203 17119
rect 5181 17085 5215 17119
rect 6101 17085 6135 17119
rect 6193 17085 6227 17119
rect 6837 17085 6871 17119
rect 7104 17085 7138 17119
rect 8493 17085 8527 17119
rect 10333 17085 10367 17119
rect 12900 17085 12934 17119
rect 14289 17085 14323 17119
rect 15025 17085 15059 17119
rect 15117 17085 15151 17119
rect 17325 17085 17359 17119
rect 18061 17085 18095 17119
rect 18981 17085 19015 17119
rect 19073 17085 19107 17119
rect 20177 17085 20211 17119
rect 20821 17085 20855 17119
rect 21088 17085 21122 17119
rect 22477 17085 22511 17119
rect 2412 17017 2446 17051
rect 8738 17017 8772 17051
rect 10600 17017 10634 17051
rect 15384 17017 15418 17051
rect 1777 16949 1811 16983
rect 4261 16949 4295 16983
rect 5273 16949 5307 16983
rect 5917 16949 5951 16983
rect 6377 16949 6411 16983
rect 8217 16949 8251 16983
rect 14473 16949 14507 16983
rect 17417 16949 17451 16983
rect 18245 16949 18279 16983
rect 18613 16949 18647 16983
rect 19809 16949 19843 16983
rect 22661 16949 22695 16983
rect 1593 16745 1627 16779
rect 3341 16745 3375 16779
rect 4077 16745 4111 16779
rect 5089 16745 5123 16779
rect 11345 16745 11379 16779
rect 13093 16745 13127 16779
rect 13369 16745 13403 16779
rect 13829 16745 13863 16779
rect 14841 16745 14875 16779
rect 16681 16745 16715 16779
rect 16957 16745 16991 16779
rect 17693 16745 17727 16779
rect 19165 16745 19199 16779
rect 22753 16745 22787 16779
rect 4537 16677 4571 16711
rect 8208 16677 8242 16711
rect 9413 16677 9447 16711
rect 9956 16677 9990 16711
rect 11958 16677 11992 16711
rect 13737 16677 13771 16711
rect 1409 16609 1443 16643
rect 1961 16609 1995 16643
rect 2228 16609 2262 16643
rect 4445 16609 4479 16643
rect 5457 16609 5491 16643
rect 6541 16609 6575 16643
rect 4629 16541 4663 16575
rect 5549 16541 5583 16575
rect 5641 16541 5675 16575
rect 6285 16541 6319 16575
rect 7941 16541 7975 16575
rect 11529 16609 11563 16643
rect 14565 16609 14599 16643
rect 14657 16609 14691 16643
rect 15568 16609 15602 16643
rect 17141 16609 17175 16643
rect 17233 16609 17267 16643
rect 18052 16677 18086 16711
rect 21281 16677 21315 16711
rect 21640 16677 21674 16711
rect 19809 16609 19843 16643
rect 9689 16541 9723 16575
rect 11713 16541 11747 16575
rect 13921 16541 13955 16575
rect 15301 16541 15335 16575
rect 17693 16541 17727 16575
rect 17785 16541 17819 16575
rect 19901 16541 19935 16575
rect 19993 16541 20027 16575
rect 20913 16541 20947 16575
rect 21281 16541 21315 16575
rect 21373 16541 21407 16575
rect 9321 16473 9355 16507
rect 9413 16473 9447 16507
rect 11069 16473 11103 16507
rect 17417 16473 17451 16507
rect 7665 16405 7699 16439
rect 14381 16405 14415 16439
rect 19441 16405 19475 16439
rect 1685 16201 1719 16235
rect 3433 16201 3467 16235
rect 8861 16201 8895 16235
rect 16957 16201 16991 16235
rect 17509 16201 17543 16235
rect 19441 16201 19475 16235
rect 21557 16201 21591 16235
rect 6101 16133 6135 16167
rect 4077 16065 4111 16099
rect 4540 16065 4574 16099
rect 4813 16065 4847 16099
rect 6653 16133 6687 16167
rect 1501 15997 1535 16031
rect 2053 15997 2087 16031
rect 3985 15997 4019 16031
rect 6101 15997 6135 16031
rect 6193 15997 6227 16031
rect 2320 15929 2354 15963
rect 7300 16065 7334 16099
rect 10793 16133 10827 16167
rect 9276 16065 9310 16099
rect 9459 16065 9493 16099
rect 11621 16065 11655 16099
rect 13001 16065 13035 16099
rect 13369 16065 13403 16099
rect 13832 16065 13866 16099
rect 15577 16065 15611 16099
rect 22109 16065 22143 16099
rect 22569 16065 22603 16099
rect 6837 15997 6871 16031
rect 7573 15997 7607 16031
rect 8861 15997 8895 16031
rect 8953 15997 8987 16031
rect 9689 15997 9723 16031
rect 11437 15997 11471 16031
rect 11529 15997 11563 16031
rect 11989 15997 12023 16031
rect 13692 15997 13726 16031
rect 14105 15997 14139 16031
rect 17325 15997 17359 16031
rect 18061 15997 18095 16031
rect 19901 15997 19935 16031
rect 20168 15997 20202 16031
rect 21925 15997 21959 16031
rect 12909 15929 12943 15963
rect 15822 15929 15856 15963
rect 18328 15929 18362 15963
rect 22017 15929 22051 15963
rect 3801 15861 3835 15895
rect 4543 15861 4577 15895
rect 5917 15861 5951 15895
rect 6377 15861 6411 15895
rect 6653 15861 6687 15895
rect 7303 15861 7337 15895
rect 8677 15861 8711 15895
rect 11069 15861 11103 15895
rect 12173 15861 12207 15895
rect 12449 15861 12483 15895
rect 12817 15861 12851 15895
rect 15209 15861 15243 15895
rect 21281 15861 21315 15895
rect 8769 15657 8803 15691
rect 9229 15657 9263 15691
rect 9505 15657 9539 15691
rect 9689 15657 9723 15691
rect 13001 15657 13035 15691
rect 14933 15657 14967 15691
rect 19349 15657 19383 15691
rect 20269 15657 20303 15691
rect 7380 15589 7414 15623
rect 1501 15521 1535 15555
rect 1768 15521 1802 15555
rect 3157 15521 3191 15555
rect 4445 15521 4479 15555
rect 4997 15521 5031 15555
rect 5733 15521 5767 15555
rect 8953 15521 8987 15555
rect 9045 15521 9079 15555
rect 3341 15453 3375 15487
rect 5320 15453 5354 15487
rect 5460 15453 5494 15487
rect 7113 15453 7147 15487
rect 10057 15521 10091 15555
rect 10977 15521 11011 15555
rect 11392 15521 11426 15555
rect 11805 15521 11839 15555
rect 10149 15453 10183 15487
rect 10241 15453 10275 15487
rect 11069 15453 11103 15487
rect 11575 15453 11609 15487
rect 18236 15589 18270 15623
rect 21180 15589 21214 15623
rect 13441 15521 13475 15555
rect 15117 15521 15151 15555
rect 15301 15521 15335 15555
rect 15624 15521 15658 15555
rect 16037 15521 16071 15555
rect 17417 15521 17451 15555
rect 20177 15521 20211 15555
rect 22569 15521 22603 15555
rect 13185 15453 13219 15487
rect 15764 15453 15798 15487
rect 17969 15453 18003 15487
rect 20453 15453 20487 15487
rect 20913 15453 20947 15487
rect 13001 15385 13035 15419
rect 17141 15385 17175 15419
rect 2881 15317 2915 15351
rect 4629 15317 4663 15351
rect 6837 15317 6871 15351
rect 8493 15317 8527 15351
rect 9505 15317 9539 15351
rect 10793 15317 10827 15351
rect 12909 15317 12943 15351
rect 14565 15317 14599 15351
rect 17601 15317 17635 15351
rect 19809 15317 19843 15351
rect 22293 15317 22327 15351
rect 10333 15113 10367 15147
rect 12081 15113 12115 15147
rect 17693 15113 17727 15147
rect 21189 15113 21223 15147
rect 3801 15045 3835 15079
rect 12541 15045 12575 15079
rect 22661 15045 22695 15079
rect 1869 14977 1903 15011
rect 4675 14977 4709 15011
rect 13093 14977 13127 15011
rect 15853 14977 15887 15011
rect 18429 14977 18463 15011
rect 19855 14977 19889 15011
rect 22017 14977 22051 15011
rect 3617 14909 3651 14943
rect 4169 14909 4203 14943
rect 4905 14909 4939 14943
rect 6837 14909 6871 14943
rect 8953 14909 8987 14943
rect 9220 14909 9254 14943
rect 10701 14909 10735 14943
rect 12909 14909 12943 14943
rect 13461 14909 13495 14943
rect 16313 14909 16347 14943
rect 18245 14909 18279 14943
rect 19349 14909 19383 14943
rect 19672 14909 19706 14943
rect 20085 14909 20119 14943
rect 22477 14909 22511 14943
rect 2136 14841 2170 14875
rect 7104 14841 7138 14875
rect 10968 14841 11002 14875
rect 13706 14841 13740 14875
rect 16580 14841 16614 14875
rect 21925 14841 21959 14875
rect 1409 14773 1443 14807
rect 3249 14773 3283 14807
rect 4635 14773 4669 14807
rect 6009 14773 6043 14807
rect 6285 14773 6319 14807
rect 8217 14773 8251 14807
rect 8493 14773 8527 14807
rect 13001 14773 13035 14807
rect 14841 14773 14875 14807
rect 15301 14773 15335 14807
rect 15669 14773 15703 14807
rect 15761 14773 15795 14807
rect 21465 14773 21499 14807
rect 21833 14773 21867 14807
rect 3065 14569 3099 14603
rect 3617 14569 3651 14603
rect 4077 14569 4111 14603
rect 4537 14569 4571 14603
rect 5089 14569 5123 14603
rect 6285 14569 6319 14603
rect 9045 14569 9079 14603
rect 11529 14569 11563 14603
rect 14381 14569 14415 14603
rect 14933 14569 14967 14603
rect 16681 14569 16715 14603
rect 20269 14569 20303 14603
rect 1952 14501 1986 14535
rect 5549 14501 5583 14535
rect 8953 14501 8987 14535
rect 10118 14501 10152 14535
rect 12716 14501 12750 14535
rect 14289 14501 14323 14535
rect 20177 14501 20211 14535
rect 21456 14501 21490 14535
rect 1685 14433 1719 14467
rect 3433 14433 3467 14467
rect 3893 14433 3927 14467
rect 4445 14433 4479 14467
rect 5457 14433 5491 14467
rect 6101 14433 6135 14467
rect 6909 14433 6943 14467
rect 8493 14433 8527 14467
rect 11897 14433 11931 14467
rect 14749 14433 14783 14467
rect 16129 14433 16163 14467
rect 16681 14433 16715 14467
rect 16773 14433 16807 14467
rect 17509 14433 17543 14467
rect 17776 14433 17810 14467
rect 18981 14433 19015 14467
rect 19183 14433 19217 14467
rect 19347 14433 19381 14467
rect 4629 14365 4663 14399
rect 5641 14365 5675 14399
rect 6653 14365 6687 14399
rect 9229 14365 9263 14399
rect 9413 14365 9447 14399
rect 9873 14365 9907 14399
rect 11989 14365 12023 14399
rect 12081 14365 12115 14399
rect 12449 14365 12483 14399
rect 14473 14365 14507 14399
rect 15301 14365 15335 14399
rect 16221 14365 16255 14399
rect 16405 14365 16439 14399
rect 3893 14297 3927 14331
rect 8585 14297 8619 14331
rect 11253 14297 11287 14331
rect 20453 14365 20487 14399
rect 21189 14365 21223 14399
rect 19533 14297 19567 14331
rect 19809 14297 19843 14331
rect 8033 14229 8067 14263
rect 8309 14229 8343 14263
rect 9413 14229 9447 14263
rect 13829 14229 13863 14263
rect 13921 14229 13955 14263
rect 15761 14229 15795 14263
rect 16957 14229 16991 14263
rect 18889 14229 18923 14263
rect 18981 14229 19015 14263
rect 22569 14229 22603 14263
rect 2881 14025 2915 14059
rect 3985 14025 4019 14059
rect 4353 14025 4387 14059
rect 9689 14025 9723 14059
rect 10977 14025 11011 14059
rect 17693 14025 17727 14059
rect 19533 14025 19567 14059
rect 21465 14025 21499 14059
rect 1501 13889 1535 13923
rect 3709 13889 3743 13923
rect 1768 13821 1802 13855
rect 3525 13753 3559 13787
rect 6837 13957 6871 13991
rect 9965 13957 9999 13991
rect 11989 13957 12023 13991
rect 18245 13957 18279 13991
rect 7389 13889 7423 13923
rect 7849 13889 7883 13923
rect 10609 13889 10643 13923
rect 11621 13889 11655 13923
rect 18889 13889 18923 13923
rect 21741 13957 21775 13991
rect 19948 13889 19982 13923
rect 20131 13889 20165 13923
rect 22385 13889 22419 13923
rect 4169 13821 4203 13855
rect 4905 13821 4939 13855
rect 5172 13821 5206 13855
rect 8309 13821 8343 13855
rect 8576 13821 8610 13855
rect 10425 13821 10459 13855
rect 11345 13821 11379 13855
rect 12173 13821 12207 13855
rect 12817 13821 12851 13855
rect 13084 13821 13118 13855
rect 14565 13821 14599 13855
rect 16313 13821 16347 13855
rect 18705 13821 18739 13855
rect 19441 13821 19475 13855
rect 19533 13821 19567 13855
rect 19625 13821 19659 13855
rect 20361 13821 20395 13855
rect 22201 13821 22235 13855
rect 14810 13753 14844 13787
rect 16580 13753 16614 13787
rect 3157 13685 3191 13719
rect 3617 13685 3651 13719
rect 3985 13685 4019 13719
rect 6285 13685 6319 13719
rect 7205 13685 7239 13719
rect 7297 13685 7331 13719
rect 10333 13685 10367 13719
rect 11437 13685 11471 13719
rect 14197 13685 14231 13719
rect 15945 13685 15979 13719
rect 18613 13685 18647 13719
rect 19257 13685 19291 13719
rect 22109 13685 22143 13719
rect 2605 13481 2639 13515
rect 2697 13481 2731 13515
rect 3617 13481 3651 13515
rect 5825 13481 5859 13515
rect 8769 13481 8803 13515
rect 9321 13481 9355 13515
rect 9873 13481 9907 13515
rect 20085 13481 20119 13515
rect 20913 13481 20947 13515
rect 4712 13413 4746 13447
rect 6101 13413 6135 13447
rect 6285 13413 6319 13447
rect 7012 13413 7046 13447
rect 8309 13413 8343 13447
rect 12418 13413 12452 13447
rect 13890 13413 13924 13447
rect 18236 13413 18270 13447
rect 21640 13413 21674 13447
rect 1685 13345 1719 13379
rect 3433 13345 3467 13379
rect 2789 13277 2823 13311
rect 4445 13277 4479 13311
rect 6745 13277 6779 13311
rect 1869 13209 1903 13243
rect 6469 13209 6503 13243
rect 10241 13345 10275 13379
rect 10968 13345 11002 13379
rect 12173 13345 12207 13379
rect 13645 13345 13679 13379
rect 15301 13345 15335 13379
rect 16028 13345 16062 13379
rect 17417 13345 17451 13379
rect 19993 13345 20027 13379
rect 8861 13277 8895 13311
rect 8953 13277 8987 13311
rect 10333 13277 10367 13311
rect 10425 13277 10459 13311
rect 10701 13277 10735 13311
rect 15761 13277 15795 13311
rect 17969 13277 18003 13311
rect 20177 13277 20211 13311
rect 21373 13277 21407 13311
rect 12081 13209 12115 13243
rect 19349 13209 19383 13243
rect 2237 13141 2271 13175
rect 8125 13141 8159 13175
rect 8309 13141 8343 13175
rect 8401 13141 8435 13175
rect 13553 13141 13587 13175
rect 15025 13141 15059 13175
rect 17141 13141 17175 13175
rect 17601 13141 17635 13175
rect 19625 13141 19659 13175
rect 22753 13141 22787 13175
rect 1593 12937 1627 12971
rect 4997 12937 5031 12971
rect 8493 12937 8527 12971
rect 11713 12937 11747 12971
rect 14197 12937 14231 12971
rect 17601 12937 17635 12971
rect 20453 12937 20487 12971
rect 22385 12937 22419 12971
rect 14013 12869 14047 12903
rect 14105 12869 14139 12903
rect 16589 12869 16623 12903
rect 5733 12801 5767 12835
rect 5825 12801 5859 12835
rect 9045 12801 9079 12835
rect 10057 12801 10091 12835
rect 17693 12869 17727 12903
rect 18245 12869 18279 12903
rect 21189 12869 21223 12903
rect 14657 12801 14691 12835
rect 14749 12801 14783 12835
rect 17325 12801 17359 12835
rect 17509 12801 17543 12835
rect 17601 12801 17635 12835
rect 21649 12801 21683 12835
rect 21833 12801 21867 12835
rect 1409 12733 1443 12767
rect 1961 12733 1995 12767
rect 3617 12733 3651 12767
rect 5641 12733 5675 12767
rect 6285 12733 6319 12767
rect 6837 12733 6871 12767
rect 9873 12733 9907 12767
rect 10333 12733 10367 12767
rect 10600 12733 10634 12767
rect 11897 12733 11931 12767
rect 12081 12733 12115 12767
rect 12633 12733 12667 12767
rect 14105 12733 14139 12767
rect 15209 12733 15243 12767
rect 2228 12665 2262 12699
rect 3862 12665 3896 12699
rect 7104 12665 7138 12699
rect 12900 12665 12934 12699
rect 14565 12665 14599 12699
rect 15454 12665 15488 12699
rect 17049 12665 17083 12699
rect 17141 12665 17175 12699
rect 17877 12733 17911 12767
rect 18061 12733 18095 12767
rect 18613 12733 18647 12767
rect 18880 12733 18914 12767
rect 20269 12733 20303 12767
rect 22201 12733 22235 12767
rect 3341 12597 3375 12631
rect 5273 12597 5307 12631
rect 8217 12597 8251 12631
rect 8861 12597 8895 12631
rect 8953 12597 8987 12631
rect 9505 12597 9539 12631
rect 9965 12597 9999 12631
rect 12265 12597 12299 12631
rect 16681 12597 16715 12631
rect 17509 12597 17543 12631
rect 19993 12597 20027 12631
rect 21557 12597 21591 12631
rect 2973 12393 3007 12427
rect 3617 12393 3651 12427
rect 4445 12393 4479 12427
rect 5733 12393 5767 12427
rect 8677 12393 8711 12427
rect 9229 12393 9263 12427
rect 9965 12393 9999 12427
rect 10517 12393 10551 12427
rect 10793 12393 10827 12427
rect 14657 12393 14691 12427
rect 14933 12393 14967 12427
rect 15669 12393 15703 12427
rect 16405 12393 16439 12427
rect 17049 12393 17083 12427
rect 5825 12325 5859 12359
rect 7288 12325 7322 12359
rect 16497 12325 16531 12359
rect 1593 12257 1627 12291
rect 1860 12257 1894 12291
rect 3433 12257 3467 12291
rect 5273 12257 5307 12291
rect 6469 12257 6503 12291
rect 7021 12257 7055 12291
rect 8861 12257 8895 12291
rect 9045 12257 9079 12291
rect 9781 12257 9815 12291
rect 10701 12257 10735 12291
rect 10793 12257 10827 12291
rect 11161 12257 11195 12291
rect 11253 12257 11287 12291
rect 4537 12189 4571 12223
rect 4721 12189 4755 12223
rect 4905 12189 4939 12223
rect 5917 12189 5951 12223
rect 5089 12121 5123 12155
rect 11345 12257 11379 12291
rect 11437 12257 11471 12291
rect 13533 12257 13567 12291
rect 15117 12257 15151 12291
rect 15485 12257 15519 12291
rect 17509 12257 17543 12291
rect 17776 12257 17810 12291
rect 19809 12257 19843 12291
rect 20913 12257 20947 12291
rect 21180 12257 21214 12291
rect 13277 12189 13311 12223
rect 16589 12189 16623 12223
rect 19901 12189 19935 12223
rect 19993 12189 20027 12223
rect 22569 12189 22603 12223
rect 11345 12121 11379 12155
rect 18889 12121 18923 12155
rect 4077 12053 4111 12087
rect 4905 12053 4939 12087
rect 5365 12053 5399 12087
rect 6653 12053 6687 12087
rect 8401 12053 8435 12087
rect 10977 12053 11011 12087
rect 11253 12053 11287 12087
rect 12725 12053 12759 12087
rect 16037 12053 16071 12087
rect 19441 12053 19475 12087
rect 22293 12053 22327 12087
rect 6469 11849 6503 11883
rect 8861 11849 8895 11883
rect 9321 11849 9355 11883
rect 11713 11849 11747 11883
rect 13921 11849 13955 11883
rect 15485 11849 15519 11883
rect 20913 11849 20947 11883
rect 22753 11849 22787 11883
rect 12173 11781 12207 11815
rect 15945 11781 15979 11815
rect 3525 11713 3559 11747
rect 3709 11713 3743 11747
rect 4721 11713 4755 11747
rect 7205 11713 7239 11747
rect 9873 11713 9907 11747
rect 10333 11713 10367 11747
rect 15117 11713 15151 11747
rect 16497 11713 16531 11747
rect 17509 11713 17543 11747
rect 18705 11713 18739 11747
rect 19536 11713 19570 11747
rect 1409 11645 1443 11679
rect 1676 11645 1710 11679
rect 4537 11645 4571 11679
rect 5089 11645 5123 11679
rect 9045 11645 9079 11679
rect 11989 11645 12023 11679
rect 14841 11645 14875 11679
rect 15301 11645 15335 11679
rect 17417 11645 17451 11679
rect 18429 11645 18463 11679
rect 19073 11645 19107 11679
rect 19809 11645 19843 11679
rect 21373 11645 21407 11679
rect 4445 11577 4479 11611
rect 5356 11577 5390 11611
rect 7472 11577 7506 11611
rect 9689 11577 9723 11611
rect 10600 11577 10634 11611
rect 12633 11577 12667 11611
rect 14933 11577 14967 11611
rect 17325 11577 17359 11611
rect 21640 11577 21674 11611
rect 2789 11509 2823 11543
rect 3065 11509 3099 11543
rect 3433 11509 3467 11543
rect 4077 11509 4111 11543
rect 8585 11509 8619 11543
rect 9781 11509 9815 11543
rect 14473 11509 14507 11543
rect 16313 11509 16347 11543
rect 16405 11509 16439 11543
rect 16957 11509 16991 11543
rect 18061 11509 18095 11543
rect 18521 11509 18555 11543
rect 19539 11509 19573 11543
rect 2789 11305 2823 11339
rect 6561 11305 6595 11339
rect 8677 11305 8711 11339
rect 9229 11305 9263 11339
rect 10057 11305 10091 11339
rect 11805 11305 11839 11339
rect 12633 11305 12667 11339
rect 14841 11305 14875 11339
rect 17141 11305 17175 11339
rect 18435 11305 18469 11339
rect 19809 11305 19843 11339
rect 22661 11305 22695 11339
rect 1676 11169 1710 11203
rect 3341 11169 3375 11203
rect 3433 11169 3467 11203
rect 4445 11169 4479 11203
rect 5181 11169 5215 11203
rect 5448 11169 5482 11203
rect 7297 11169 7331 11203
rect 7564 11169 7598 11203
rect 9045 11169 9079 11203
rect 9873 11169 9907 11203
rect 10425 11169 10459 11203
rect 10692 11169 10726 11203
rect 12265 11169 12299 11203
rect 1409 11101 1443 11135
rect 4537 11101 4571 11135
rect 4721 11101 4755 11135
rect 6837 11101 6871 11135
rect 21548 11237 21582 11271
rect 12817 11169 12851 11203
rect 13084 11169 13118 11203
rect 14657 11169 14691 11203
rect 15925 11169 15959 11203
rect 17509 11169 17543 11203
rect 17601 11169 17635 11203
rect 17969 11169 18003 11203
rect 20269 11169 20303 11203
rect 15669 11101 15703 11135
rect 17693 11101 17727 11135
rect 18432 11101 18466 11135
rect 18705 11101 18739 11135
rect 21281 11101 21315 11135
rect 4077 11033 4111 11067
rect 12449 11033 12483 11067
rect 12633 11033 12667 11067
rect 20453 11033 20487 11067
rect 3157 10965 3191 10999
rect 3617 10965 3651 10999
rect 14197 10965 14231 10999
rect 17049 10965 17083 10999
rect 3157 10761 3191 10795
rect 4813 10761 4847 10795
rect 6469 10761 6503 10795
rect 7021 10761 7055 10795
rect 9321 10761 9355 10795
rect 17509 10761 17543 10795
rect 18245 10761 18279 10795
rect 21097 10761 21131 10795
rect 9689 10693 9723 10727
rect 11989 10693 12023 10727
rect 9965 10625 9999 10659
rect 12541 10625 12575 10659
rect 15853 10625 15887 10659
rect 18705 10625 18739 10659
rect 18889 10625 18923 10659
rect 21925 10625 21959 10659
rect 1777 10557 1811 10591
rect 2044 10557 2078 10591
rect 3433 10557 3467 10591
rect 3700 10557 3734 10591
rect 5089 10557 5123 10591
rect 6837 10557 6871 10591
rect 7481 10557 7515 10591
rect 9137 10557 9171 10591
rect 9873 10557 9907 10591
rect 11805 10557 11839 10591
rect 12797 10557 12831 10591
rect 14197 10557 14231 10591
rect 17325 10557 17359 10591
rect 19717 10557 19751 10591
rect 19984 10557 20018 10591
rect 21833 10557 21867 10591
rect 22385 10557 22419 10591
rect 5356 10489 5390 10523
rect 7748 10489 7782 10523
rect 10232 10489 10266 10523
rect 14442 10489 14476 10523
rect 16120 10489 16154 10523
rect 18613 10489 18647 10523
rect 19257 10489 19291 10523
rect 21741 10489 21775 10523
rect 8861 10421 8895 10455
rect 11345 10421 11379 10455
rect 13921 10421 13955 10455
rect 15577 10421 15611 10455
rect 17233 10421 17267 10455
rect 17693 10421 17727 10455
rect 21373 10421 21407 10455
rect 22569 10421 22603 10455
rect 1685 10217 1719 10251
rect 1961 10217 1995 10251
rect 5549 10217 5583 10251
rect 7205 10217 7239 10251
rect 11069 10217 11103 10251
rect 14105 10217 14139 10251
rect 14565 10217 14599 10251
rect 14749 10217 14783 10251
rect 16865 10217 16899 10251
rect 20085 10217 20119 10251
rect 20361 10217 20395 10251
rect 22293 10217 22327 10251
rect 4436 10149 4470 10183
rect 6070 10149 6104 10183
rect 12173 10149 12207 10183
rect 12633 10149 12667 10183
rect 12970 10149 13004 10183
rect 1501 10081 1535 10115
rect 2053 10081 2087 10115
rect 2320 10081 2354 10115
rect 4169 10081 4203 10115
rect 8197 10081 8231 10115
rect 9956 10081 9990 10115
rect 12081 10081 12115 10115
rect 5825 10013 5859 10047
rect 7941 10013 7975 10047
rect 9689 10013 9723 10047
rect 12357 10013 12391 10047
rect 12725 10081 12759 10115
rect 14381 10081 14415 10115
rect 3433 9877 3467 9911
rect 9321 9877 9355 9911
rect 11713 9877 11747 9911
rect 12633 9877 12667 9911
rect 15752 10149 15786 10183
rect 15117 10081 15151 10115
rect 17601 10081 17635 10115
rect 17693 10081 17727 10115
rect 18245 10081 18279 10115
rect 18512 10081 18546 10115
rect 19901 10081 19935 10115
rect 15485 10013 15519 10047
rect 17785 10013 17819 10047
rect 22201 10149 22235 10183
rect 20637 10081 20671 10115
rect 21281 10081 21315 10115
rect 22477 10013 22511 10047
rect 20361 9945 20395 9979
rect 20453 9945 20487 9979
rect 14749 9877 14783 9911
rect 14933 9877 14967 9911
rect 17233 9877 17267 9911
rect 19625 9877 19659 9911
rect 21465 9877 21499 9911
rect 21833 9877 21867 9911
rect 7665 9673 7699 9707
rect 14381 9673 14415 9707
rect 2789 9605 2823 9639
rect 4445 9605 4479 9639
rect 7297 9605 7331 9639
rect 7481 9605 7515 9639
rect 10057 9605 10091 9639
rect 11713 9605 11747 9639
rect 12081 9605 12115 9639
rect 14105 9605 14139 9639
rect 16681 9605 16715 9639
rect 21005 9605 21039 9639
rect 1409 9537 1443 9571
rect 4721 9537 4755 9571
rect 5641 9537 5675 9571
rect 5733 9537 5767 9571
rect 3065 9469 3099 9503
rect 3332 9469 3366 9503
rect 6193 9469 6227 9503
rect 7113 9469 7147 9503
rect 1654 9401 1688 9435
rect 5549 9401 5583 9435
rect 8309 9537 8343 9571
rect 12725 9537 12759 9571
rect 15301 9537 15335 9571
rect 17417 9537 17451 9571
rect 17601 9537 17635 9571
rect 18797 9537 18831 9571
rect 19165 9537 19199 9571
rect 19671 9537 19705 9571
rect 19901 9537 19935 9571
rect 21373 9537 21407 9571
rect 8125 9469 8159 9503
rect 8677 9469 8711 9503
rect 8944 9469 8978 9503
rect 10333 9469 10367 9503
rect 12265 9469 12299 9503
rect 14565 9469 14599 9503
rect 14657 9469 14691 9503
rect 15568 9469 15602 9503
rect 19488 9469 19522 9503
rect 10578 9401 10612 9435
rect 12992 9401 13026 9435
rect 14841 9401 14875 9435
rect 21640 9401 21674 9435
rect 5181 9333 5215 9367
rect 6377 9333 6411 9367
rect 7481 9333 7515 9367
rect 8033 9333 8067 9367
rect 15025 9333 15059 9367
rect 16957 9333 16991 9367
rect 17325 9333 17359 9367
rect 18153 9333 18187 9367
rect 18521 9333 18555 9367
rect 18613 9333 18647 9367
rect 22753 9333 22787 9367
rect 2329 9129 2363 9163
rect 3249 9129 3283 9163
rect 4077 9129 4111 9163
rect 4445 9129 4479 9163
rect 5089 9129 5123 9163
rect 5457 9129 5491 9163
rect 7941 9129 7975 9163
rect 8033 9129 8067 9163
rect 8585 9129 8619 9163
rect 8953 9129 8987 9163
rect 10241 9129 10275 9163
rect 11621 9129 11655 9163
rect 13185 9129 13219 9163
rect 15853 9129 15887 9163
rect 22661 9129 22695 9163
rect 2237 9061 2271 9095
rect 5549 9061 5583 9095
rect 8401 9061 8435 9095
rect 9045 9061 9079 9095
rect 11989 9061 12023 9095
rect 15945 9061 15979 9095
rect 3341 8993 3375 9027
rect 6929 8993 6963 9027
rect 2513 8925 2547 8959
rect 3525 8925 3559 8959
rect 4537 8925 4571 8959
rect 4721 8925 4755 8959
rect 5733 8925 5767 8959
rect 7021 8925 7055 8959
rect 7205 8925 7239 8959
rect 8125 8925 8159 8959
rect 10057 8993 10091 9027
rect 10977 8993 11011 9027
rect 12081 8993 12115 9027
rect 12909 8993 12943 9027
rect 13001 8993 13035 9027
rect 13820 8993 13854 9027
rect 16497 8993 16531 9027
rect 16764 8993 16798 9027
rect 18660 8993 18694 9027
rect 21537 8993 21571 9027
rect 9229 8925 9263 8959
rect 11069 8925 11103 8959
rect 11253 8925 11287 8959
rect 12265 8925 12299 8959
rect 13553 8925 13587 8959
rect 16129 8925 16163 8959
rect 18337 8925 18371 8959
rect 18843 8925 18877 8959
rect 19073 8925 19107 8959
rect 21281 8925 21315 8959
rect 2881 8857 2915 8891
rect 7573 8857 7607 8891
rect 8401 8857 8435 8891
rect 20177 8857 20211 8891
rect 1869 8789 1903 8823
rect 6561 8789 6595 8823
rect 10609 8789 10643 8823
rect 12725 8789 12759 8823
rect 14933 8789 14967 8823
rect 15485 8789 15519 8823
rect 17877 8789 17911 8823
rect 2973 8585 3007 8619
rect 3801 8585 3835 8619
rect 4169 8585 4203 8619
rect 4721 8585 4755 8619
rect 7021 8585 7055 8619
rect 7757 8585 7791 8619
rect 9597 8585 9631 8619
rect 11989 8585 12023 8619
rect 13093 8585 13127 8619
rect 14749 8585 14783 8619
rect 15209 8585 15243 8619
rect 16957 8585 16991 8619
rect 18153 8585 18187 8619
rect 20545 8585 20579 8619
rect 22201 8585 22235 8619
rect 1961 8517 1995 8551
rect 2605 8449 2639 8483
rect 3433 8449 3467 8483
rect 3617 8449 3651 8483
rect 5733 8517 5767 8551
rect 5181 8449 5215 8483
rect 5273 8449 5307 8483
rect 6377 8449 6411 8483
rect 8401 8449 8435 8483
rect 9321 8449 9355 8483
rect 2329 8381 2363 8415
rect 3341 8381 3375 8415
rect 3801 8381 3835 8415
rect 3985 8381 4019 8415
rect 5089 8381 5123 8415
rect 6837 8381 6871 8415
rect 11161 8517 11195 8551
rect 12633 8517 12667 8551
rect 15393 8517 15427 8551
rect 22661 8517 22695 8551
rect 9781 8449 9815 8483
rect 13369 8449 13403 8483
rect 11437 8381 11471 8415
rect 12173 8381 12207 8415
rect 12449 8381 12483 8415
rect 13277 8381 13311 8415
rect 13636 8381 13670 8415
rect 15025 8381 15059 8415
rect 17417 8449 17451 8483
rect 18797 8449 18831 8483
rect 15577 8381 15611 8415
rect 17233 8381 17267 8415
rect 18521 8381 18555 8415
rect 19165 8381 19199 8415
rect 19432 8381 19466 8415
rect 20821 8381 20855 8415
rect 21077 8381 21111 8415
rect 22477 8381 22511 8415
rect 2421 8313 2455 8347
rect 6101 8313 6135 8347
rect 8125 8313 8159 8347
rect 9137 8313 9171 8347
rect 9597 8313 9631 8347
rect 10048 8313 10082 8347
rect 15393 8313 15427 8347
rect 15822 8313 15856 8347
rect 18613 8313 18647 8347
rect 6193 8245 6227 8279
rect 8217 8245 8251 8279
rect 8769 8245 8803 8279
rect 9229 8245 9263 8279
rect 11621 8245 11655 8279
rect 5917 8041 5951 8075
rect 6929 8041 6963 8075
rect 8953 8041 8987 8075
rect 9045 8041 9079 8075
rect 12817 8041 12851 8075
rect 13001 8041 13035 8075
rect 14473 8041 14507 8075
rect 14749 8041 14783 8075
rect 17509 8041 17543 8075
rect 19349 8041 19383 8075
rect 19625 8041 19659 8075
rect 22201 8041 22235 8075
rect 7941 7973 7975 8007
rect 8033 7973 8067 8007
rect 10048 7973 10082 8007
rect 2513 7905 2547 7939
rect 3157 7905 3191 7939
rect 4445 7905 4479 7939
rect 5733 7905 5767 7939
rect 9781 7905 9815 7939
rect 11693 7905 11727 7939
rect 21281 7973 21315 8007
rect 22109 7973 22143 8007
rect 13360 7905 13394 7939
rect 15936 7905 15970 7939
rect 17325 7905 17359 7939
rect 18225 7905 18259 7939
rect 19993 7905 20027 7939
rect 21005 7905 21039 7939
rect 4997 7837 5031 7871
rect 7021 7837 7055 7871
rect 7205 7837 7239 7871
rect 8125 7837 8159 7871
rect 9229 7837 9263 7871
rect 9413 7837 9447 7871
rect 11437 7837 11471 7871
rect 13001 7837 13035 7871
rect 13093 7837 13127 7871
rect 15669 7837 15703 7871
rect 17969 7837 18003 7871
rect 20085 7837 20119 7871
rect 20177 7837 20211 7871
rect 22385 7837 22419 7871
rect 7573 7769 7607 7803
rect 11161 7769 11195 7803
rect 21741 7769 21775 7803
rect 6561 7701 6595 7735
rect 8585 7701 8619 7735
rect 9413 7701 9447 7735
rect 17049 7701 17083 7735
rect 4721 7497 4755 7531
rect 5733 7497 5767 7531
rect 7573 7497 7607 7531
rect 17693 7497 17727 7531
rect 20269 7497 20303 7531
rect 3709 7429 3743 7463
rect 9965 7429 9999 7463
rect 14933 7429 14967 7463
rect 4353 7361 4387 7395
rect 5365 7361 5399 7395
rect 6285 7361 6319 7395
rect 8217 7361 8251 7395
rect 8585 7361 8619 7395
rect 10241 7361 10275 7395
rect 13185 7361 13219 7395
rect 15853 7361 15887 7395
rect 16316 7361 16350 7395
rect 18429 7361 18463 7395
rect 18892 7361 18926 7395
rect 19165 7361 19199 7395
rect 4169 7293 4203 7327
rect 8033 7293 8067 7327
rect 10508 7293 10542 7327
rect 13553 7293 13587 7327
rect 15301 7293 15335 7327
rect 16589 7293 16623 7327
rect 20545 7293 20579 7327
rect 22201 7293 22235 7327
rect 5181 7225 5215 7259
rect 6193 7225 6227 7259
rect 7941 7225 7975 7259
rect 8852 7225 8886 7259
rect 13820 7225 13854 7259
rect 20790 7225 20824 7259
rect 22477 7225 22511 7259
rect 4077 7157 4111 7191
rect 5089 7157 5123 7191
rect 6101 7157 6135 7191
rect 11621 7157 11655 7191
rect 12541 7157 12575 7191
rect 12909 7157 12943 7191
rect 13001 7157 13035 7191
rect 15485 7157 15519 7191
rect 16319 7157 16353 7191
rect 18895 7157 18929 7191
rect 21925 7157 21959 7191
rect 5917 6953 5951 6987
rect 6561 6953 6595 6987
rect 6929 6953 6963 6987
rect 7941 6953 7975 6987
rect 8033 6953 8067 6987
rect 8953 6953 8987 6987
rect 13461 6953 13495 6987
rect 14933 6953 14967 6987
rect 19441 6953 19475 6987
rect 4905 6885 4939 6919
rect 12909 6885 12943 6919
rect 4997 6817 5031 6851
rect 7021 6817 7055 6851
rect 9873 6817 9907 6851
rect 10692 6817 10726 6851
rect 19809 6885 19843 6919
rect 21158 6885 21192 6919
rect 13820 6817 13854 6851
rect 15669 6817 15703 6851
rect 15936 6817 15970 6851
rect 18052 6817 18086 6851
rect 20637 6817 20671 6851
rect 22569 6817 22603 6851
rect 5181 6749 5215 6783
rect 6009 6749 6043 6783
rect 6193 6749 6227 6783
rect 7113 6749 7147 6783
rect 8217 6749 8251 6783
rect 9045 6749 9079 6783
rect 9137 6749 9171 6783
rect 10425 6749 10459 6783
rect 13001 6749 13035 6783
rect 13185 6749 13219 6783
rect 13461 6749 13495 6783
rect 13553 6749 13587 6783
rect 17141 6749 17175 6783
rect 17325 6749 17359 6783
rect 17693 6749 17727 6783
rect 17785 6749 17819 6783
rect 19901 6749 19935 6783
rect 19993 6749 20027 6783
rect 20361 6749 20395 6783
rect 20913 6749 20947 6783
rect 4537 6681 4571 6715
rect 5549 6681 5583 6715
rect 8585 6681 8619 6715
rect 10057 6681 10091 6715
rect 19165 6681 19199 6715
rect 7573 6613 7607 6647
rect 11805 6613 11839 6647
rect 12541 6613 12575 6647
rect 17049 6613 17083 6647
rect 17233 6613 17267 6647
rect 17693 6613 17727 6647
rect 20361 6613 20395 6647
rect 20453 6613 20487 6647
rect 22293 6613 22327 6647
rect 5641 6409 5675 6443
rect 7665 6409 7699 6443
rect 9689 6409 9723 6443
rect 21097 6409 21131 6443
rect 8677 6341 8711 6375
rect 14657 6341 14691 6375
rect 20177 6341 20211 6375
rect 6101 6273 6135 6307
rect 6285 6273 6319 6307
rect 8217 6273 8251 6307
rect 9137 6273 9171 6307
rect 9321 6273 9355 6307
rect 10333 6273 10367 6307
rect 13093 6273 13127 6307
rect 17417 6273 17451 6307
rect 17601 6273 17635 6307
rect 6009 6205 6043 6239
rect 8033 6205 8067 6239
rect 9045 6205 9079 6239
rect 10701 6205 10735 6239
rect 12541 6205 12575 6239
rect 14657 6205 14691 6239
rect 14749 6205 14783 6239
rect 16405 6205 16439 6239
rect 17325 6205 17359 6239
rect 18245 6205 18279 6239
rect 18797 6205 18831 6239
rect 20729 6205 20763 6239
rect 21373 6205 21407 6239
rect 8125 6137 8159 6171
rect 10057 6137 10091 6171
rect 10968 6137 11002 6171
rect 13360 6137 13394 6171
rect 14994 6137 15028 6171
rect 19064 6137 19098 6171
rect 20913 6137 20947 6171
rect 21640 6137 21674 6171
rect 10149 6069 10183 6103
rect 12081 6069 12115 6103
rect 12725 6069 12759 6103
rect 14473 6069 14507 6103
rect 16129 6069 16163 6103
rect 16589 6069 16623 6103
rect 16957 6069 16991 6103
rect 18429 6069 18463 6103
rect 22753 6069 22787 6103
rect 5549 5865 5583 5899
rect 6561 5865 6595 5899
rect 7021 5865 7055 5899
rect 7573 5865 7607 5899
rect 7941 5865 7975 5899
rect 9045 5865 9079 5899
rect 11989 5865 12023 5899
rect 13645 5865 13679 5899
rect 14289 5865 14323 5899
rect 14933 5865 14967 5899
rect 15761 5865 15795 5899
rect 18521 5865 18555 5899
rect 19165 5865 19199 5899
rect 20269 5865 20303 5899
rect 22661 5865 22695 5899
rect 5917 5797 5951 5831
rect 6009 5797 6043 5831
rect 8033 5797 8067 5831
rect 8953 5797 8987 5831
rect 12532 5797 12566 5831
rect 14381 5797 14415 5831
rect 16497 5797 16531 5831
rect 20177 5797 20211 5831
rect 6929 5729 6963 5763
rect 10609 5729 10643 5763
rect 10876 5729 10910 5763
rect 15117 5729 15151 5763
rect 15577 5729 15611 5763
rect 17141 5729 17175 5763
rect 17408 5729 17442 5763
rect 19257 5729 19291 5763
rect 20913 5729 20947 5763
rect 21833 5729 21867 5763
rect 21925 5729 21959 5763
rect 22477 5729 22511 5763
rect 6101 5661 6135 5695
rect 7113 5661 7147 5695
rect 8217 5661 8251 5695
rect 9229 5661 9263 5695
rect 12265 5661 12299 5695
rect 14565 5661 14599 5695
rect 16589 5661 16623 5695
rect 16773 5661 16807 5695
rect 19441 5661 19475 5695
rect 20361 5661 20395 5695
rect 21281 5661 21315 5695
rect 22109 5661 22143 5695
rect 8585 5593 8619 5627
rect 18797 5593 18831 5627
rect 13921 5525 13955 5559
rect 16129 5525 16163 5559
rect 19809 5525 19843 5559
rect 21097 5525 21131 5559
rect 21281 5525 21315 5559
rect 21465 5525 21499 5559
rect 7665 5321 7699 5355
rect 9137 5321 9171 5355
rect 10149 5321 10183 5355
rect 11161 5321 11195 5355
rect 12449 5321 12483 5355
rect 16589 5321 16623 5355
rect 16865 5321 16899 5355
rect 18521 5321 18555 5355
rect 20821 5321 20855 5355
rect 22569 5321 22603 5355
rect 19625 5253 19659 5287
rect 8217 5185 8251 5219
rect 9781 5185 9815 5219
rect 10701 5185 10735 5219
rect 11621 5185 11655 5219
rect 11805 5185 11839 5219
rect 12909 5185 12943 5219
rect 13093 5185 13127 5219
rect 15209 5185 15243 5219
rect 17509 5185 17543 5219
rect 18061 5185 18095 5219
rect 18981 5185 19015 5219
rect 19165 5185 19199 5219
rect 20269 5185 20303 5219
rect 8033 5117 8067 5151
rect 10517 5117 10551 5151
rect 10609 5117 10643 5151
rect 11529 5117 11563 5151
rect 13553 5117 13587 5151
rect 13820 5117 13854 5151
rect 20637 5117 20671 5151
rect 21189 5117 21223 5151
rect 8125 5049 8159 5083
rect 9505 5049 9539 5083
rect 15454 5049 15488 5083
rect 17325 5049 17359 5083
rect 19993 5049 20027 5083
rect 21456 5049 21490 5083
rect 9597 4981 9631 5015
rect 12817 4981 12851 5015
rect 14933 4981 14967 5015
rect 17233 4981 17267 5015
rect 18889 4981 18923 5015
rect 20085 4981 20119 5015
rect 9873 4777 9907 4811
rect 10241 4777 10275 4811
rect 11345 4777 11379 4811
rect 11897 4777 11931 4811
rect 12357 4777 12391 4811
rect 12909 4777 12943 4811
rect 13277 4777 13311 4811
rect 13921 4777 13955 4811
rect 14289 4777 14323 4811
rect 15485 4777 15519 4811
rect 17785 4777 17819 4811
rect 18245 4777 18279 4811
rect 19165 4777 19199 4811
rect 19809 4777 19843 4811
rect 20177 4777 20211 4811
rect 22477 4777 22511 4811
rect 10333 4709 10367 4743
rect 13369 4709 13403 4743
rect 14381 4709 14415 4743
rect 19257 4709 19291 4743
rect 11253 4641 11287 4675
rect 12265 4641 12299 4675
rect 15301 4641 15335 4675
rect 16109 4641 16143 4675
rect 18153 4641 18187 4675
rect 20269 4641 20303 4675
rect 21097 4641 21131 4675
rect 21364 4641 21398 4675
rect 10517 4573 10551 4607
rect 11529 4573 11563 4607
rect 11805 4573 11839 4607
rect 12449 4573 12483 4607
rect 13461 4573 13495 4607
rect 14473 4573 14507 4607
rect 15853 4573 15887 4607
rect 18337 4573 18371 4607
rect 19441 4573 19475 4607
rect 20361 4573 20395 4607
rect 10885 4505 10919 4539
rect 18797 4505 18831 4539
rect 11805 4437 11839 4471
rect 17233 4437 17267 4471
rect 13645 4233 13679 4267
rect 18061 4233 18095 4267
rect 14473 4165 14507 4199
rect 16037 4165 16071 4199
rect 11805 4097 11839 4131
rect 11897 4097 11931 4131
rect 13185 4097 13219 4131
rect 14289 4097 14323 4131
rect 14013 4029 14047 4063
rect 16221 4097 16255 4131
rect 16313 4097 16347 4131
rect 18705 4097 18739 4131
rect 19073 4097 19107 4131
rect 14657 4029 14691 4063
rect 14924 4029 14958 4063
rect 11345 3893 11379 3927
rect 11713 3893 11747 3927
rect 12633 3893 12667 3927
rect 13001 3893 13035 3927
rect 13093 3893 13127 3927
rect 14105 3893 14139 3927
rect 14473 3893 14507 3927
rect 18429 4029 18463 4063
rect 19533 4029 19567 4063
rect 21373 4029 21407 4063
rect 21640 4029 21674 4063
rect 16580 3961 16614 3995
rect 19778 3961 19812 3995
rect 16221 3893 16255 3927
rect 17693 3893 17727 3927
rect 18521 3893 18555 3927
rect 20913 3893 20947 3927
rect 22753 3893 22787 3927
rect 11161 3689 11195 3723
rect 11621 3689 11655 3723
rect 13553 3689 13587 3723
rect 13645 3689 13679 3723
rect 14197 3689 14231 3723
rect 14565 3689 14599 3723
rect 15945 3689 15979 3723
rect 16129 3689 16163 3723
rect 16497 3689 16531 3723
rect 18521 3689 18555 3723
rect 20913 3689 20947 3723
rect 22753 3689 22787 3723
rect 11529 3621 11563 3655
rect 12633 3621 12667 3655
rect 12541 3553 12575 3587
rect 14657 3553 14691 3587
rect 15577 3553 15611 3587
rect 11713 3485 11747 3519
rect 12817 3485 12851 3519
rect 13829 3485 13863 3519
rect 14841 3485 14875 3519
rect 12173 3417 12207 3451
rect 17408 3621 17442 3655
rect 16037 3553 16071 3587
rect 19248 3553 19282 3587
rect 21373 3553 21407 3587
rect 21640 3553 21674 3587
rect 16589 3485 16623 3519
rect 16681 3485 16715 3519
rect 17141 3485 17175 3519
rect 18981 3485 19015 3519
rect 16037 3417 16071 3451
rect 13185 3349 13219 3383
rect 15761 3349 15795 3383
rect 15945 3349 15979 3383
rect 20361 3349 20395 3383
rect 13277 3145 13311 3179
rect 14105 3145 14139 3179
rect 15301 3145 15335 3179
rect 16129 3145 16163 3179
rect 19625 3145 19659 3179
rect 22109 3145 22143 3179
rect 1961 3009 1995 3043
rect 13921 3009 13955 3043
rect 14749 3009 14783 3043
rect 15761 3009 15795 3043
rect 15853 3009 15887 3043
rect 1777 2941 1811 2975
rect 2513 2941 2547 2975
rect 5089 2941 5123 2975
rect 13737 2941 13771 2975
rect 13645 2873 13679 2907
rect 22569 3077 22603 3111
rect 20729 3009 20763 3043
rect 16313 2941 16347 2975
rect 16580 2941 16614 2975
rect 18245 2941 18279 2975
rect 19993 2941 20027 2975
rect 22385 2941 22419 2975
rect 18490 2873 18524 2907
rect 20269 2873 20303 2907
rect 20974 2873 21008 2907
rect 2697 2805 2731 2839
rect 14473 2805 14507 2839
rect 14565 2805 14599 2839
rect 15209 2805 15243 2839
rect 15669 2805 15703 2839
rect 16129 2805 16163 2839
rect 17693 2805 17727 2839
rect 13737 2601 13771 2635
rect 14841 2601 14875 2635
rect 16589 2601 16623 2635
rect 19717 2601 19751 2635
rect 20453 2601 20487 2635
rect 20545 2601 20579 2635
rect 22569 2601 22603 2635
rect 14749 2533 14783 2567
rect 16681 2533 16715 2567
rect 17601 2533 17635 2567
rect 18604 2533 18638 2567
rect 18337 2465 18371 2499
rect 21189 2465 21223 2499
rect 21445 2465 21479 2499
rect 13829 2397 13863 2431
rect 13921 2397 13955 2431
rect 15025 2397 15059 2431
rect 16865 2397 16899 2431
rect 17693 2397 17727 2431
rect 17877 2397 17911 2431
rect 20637 2397 20671 2431
rect 14381 2329 14415 2363
rect 13369 2261 13403 2295
rect 16221 2261 16255 2295
rect 17233 2261 17267 2295
rect 20085 2261 20119 2295
<< metal1 >>
rect 7558 21972 7564 22024
rect 7616 22012 7622 22024
rect 16666 22012 16672 22024
rect 7616 21984 16672 22012
rect 7616 21972 7622 21984
rect 16666 21972 16672 21984
rect 16724 21972 16730 22024
rect 9950 21904 9956 21956
rect 10008 21944 10014 21956
rect 16942 21944 16948 21956
rect 10008 21916 16948 21944
rect 10008 21904 10014 21916
rect 16942 21904 16948 21916
rect 17000 21904 17006 21956
rect 18690 21904 18696 21956
rect 18748 21944 18754 21956
rect 19518 21944 19524 21956
rect 18748 21916 19524 21944
rect 18748 21904 18754 21916
rect 19518 21904 19524 21916
rect 19576 21904 19582 21956
rect 18322 21836 18328 21888
rect 18380 21876 18386 21888
rect 20070 21876 20076 21888
rect 18380 21848 20076 21876
rect 18380 21836 18386 21848
rect 20070 21836 20076 21848
rect 20128 21836 20134 21888
rect 1104 21786 23276 21808
rect 1104 21734 4680 21786
rect 4732 21734 4744 21786
rect 4796 21734 4808 21786
rect 4860 21734 4872 21786
rect 4924 21734 12078 21786
rect 12130 21734 12142 21786
rect 12194 21734 12206 21786
rect 12258 21734 12270 21786
rect 12322 21734 19475 21786
rect 19527 21734 19539 21786
rect 19591 21734 19603 21786
rect 19655 21734 19667 21786
rect 19719 21734 23276 21786
rect 1104 21712 23276 21734
rect 1486 21632 1492 21684
rect 1544 21672 1550 21684
rect 1581 21675 1639 21681
rect 1581 21672 1593 21675
rect 1544 21644 1593 21672
rect 1544 21632 1550 21644
rect 1581 21641 1593 21644
rect 1627 21641 1639 21675
rect 1581 21635 1639 21641
rect 8110 21632 8116 21684
rect 8168 21672 8174 21684
rect 8570 21672 8576 21684
rect 8168 21644 8576 21672
rect 8168 21632 8174 21644
rect 8570 21632 8576 21644
rect 8628 21632 8634 21684
rect 9950 21672 9956 21684
rect 9911 21644 9956 21672
rect 9950 21632 9956 21644
rect 10008 21632 10014 21684
rect 14734 21632 14740 21684
rect 14792 21672 14798 21684
rect 15473 21675 15531 21681
rect 15473 21672 15485 21675
rect 14792 21644 15485 21672
rect 14792 21632 14798 21644
rect 15473 21641 15485 21644
rect 15519 21641 15531 21675
rect 15473 21635 15531 21641
rect 18509 21675 18567 21681
rect 18509 21641 18521 21675
rect 18555 21672 18567 21675
rect 19794 21672 19800 21684
rect 18555 21644 19800 21672
rect 18555 21641 18567 21644
rect 18509 21635 18567 21641
rect 19794 21632 19800 21644
rect 19852 21632 19858 21684
rect 7558 21604 7564 21616
rect 2608 21576 7564 21604
rect 2608 21545 2636 21576
rect 7558 21564 7564 21576
rect 7616 21564 7622 21616
rect 13633 21607 13691 21613
rect 13633 21573 13645 21607
rect 13679 21604 13691 21607
rect 16758 21604 16764 21616
rect 13679 21576 16764 21604
rect 13679 21573 13691 21576
rect 13633 21567 13691 21573
rect 16758 21564 16764 21576
rect 16816 21564 16822 21616
rect 17678 21604 17684 21616
rect 17604 21576 17684 21604
rect 2593 21539 2651 21545
rect 2593 21505 2605 21539
rect 2639 21505 2651 21539
rect 2593 21499 2651 21505
rect 3605 21539 3663 21545
rect 3605 21505 3617 21539
rect 3651 21536 3663 21539
rect 4617 21539 4675 21545
rect 4617 21536 4629 21539
rect 3651 21508 4629 21536
rect 3651 21505 3663 21508
rect 3605 21499 3663 21505
rect 4617 21505 4629 21508
rect 4663 21536 4675 21539
rect 5534 21536 5540 21548
rect 4663 21508 5540 21536
rect 4663 21505 4675 21508
rect 4617 21499 4675 21505
rect 5534 21496 5540 21508
rect 5592 21536 5598 21548
rect 6365 21539 6423 21545
rect 6365 21536 6377 21539
rect 5592 21508 6377 21536
rect 5592 21496 5598 21508
rect 6365 21505 6377 21508
rect 6411 21536 6423 21539
rect 7469 21539 7527 21545
rect 7469 21536 7481 21539
rect 6411 21508 7481 21536
rect 6411 21505 6423 21508
rect 6365 21499 6423 21505
rect 7469 21505 7481 21508
rect 7515 21536 7527 21539
rect 8941 21539 8999 21545
rect 8941 21536 8953 21539
rect 7515 21508 8953 21536
rect 7515 21505 7527 21508
rect 7469 21499 7527 21505
rect 8941 21505 8953 21508
rect 8987 21505 8999 21539
rect 8941 21499 8999 21505
rect 13265 21539 13323 21545
rect 13265 21505 13277 21539
rect 13311 21536 13323 21539
rect 14182 21536 14188 21548
rect 13311 21508 14188 21536
rect 13311 21505 13323 21508
rect 13265 21499 13323 21505
rect 14182 21496 14188 21508
rect 14240 21496 14246 21548
rect 14844 21508 16068 21536
rect 1397 21471 1455 21477
rect 1397 21437 1409 21471
rect 1443 21468 1455 21471
rect 1443 21440 4108 21468
rect 1443 21437 1455 21440
rect 1397 21431 1455 21437
rect 2317 21403 2375 21409
rect 2317 21369 2329 21403
rect 2363 21400 2375 21403
rect 2682 21400 2688 21412
rect 2363 21372 2688 21400
rect 2363 21369 2375 21372
rect 2317 21363 2375 21369
rect 2682 21360 2688 21372
rect 2740 21360 2746 21412
rect 4080 21400 4108 21440
rect 4154 21428 4160 21480
rect 4212 21468 4218 21480
rect 5077 21471 5135 21477
rect 5077 21468 5089 21471
rect 4212 21440 5089 21468
rect 4212 21428 4218 21440
rect 5077 21437 5089 21440
rect 5123 21437 5135 21471
rect 5077 21431 5135 21437
rect 9122 21428 9128 21480
rect 9180 21468 9186 21480
rect 9769 21471 9827 21477
rect 9769 21468 9781 21471
rect 9180 21440 9781 21468
rect 9180 21428 9186 21440
rect 9769 21437 9781 21440
rect 9815 21437 9827 21471
rect 9769 21431 9827 21437
rect 10410 21428 10416 21480
rect 10468 21468 10474 21480
rect 10689 21471 10747 21477
rect 10689 21468 10701 21471
rect 10468 21440 10701 21468
rect 10468 21428 10474 21440
rect 10689 21437 10701 21440
rect 10735 21437 10747 21471
rect 10689 21431 10747 21437
rect 12158 21428 12164 21480
rect 12216 21468 12222 21480
rect 14844 21477 14872 21508
rect 13081 21471 13139 21477
rect 13081 21468 13093 21471
rect 12216 21440 13093 21468
rect 12216 21428 12222 21440
rect 13081 21437 13093 21440
rect 13127 21437 13139 21471
rect 13081 21431 13139 21437
rect 14829 21471 14887 21477
rect 14829 21437 14841 21471
rect 14875 21437 14887 21471
rect 14829 21431 14887 21437
rect 15562 21428 15568 21480
rect 15620 21468 15626 21480
rect 15933 21471 15991 21477
rect 15933 21468 15945 21471
rect 15620 21440 15945 21468
rect 15620 21428 15626 21440
rect 15933 21437 15945 21440
rect 15979 21437 15991 21471
rect 16040 21468 16068 21508
rect 16114 21496 16120 21548
rect 16172 21536 16178 21548
rect 16172 21508 16217 21536
rect 16172 21496 16178 21508
rect 16482 21496 16488 21548
rect 16540 21536 16546 21548
rect 17037 21539 17095 21545
rect 17037 21536 17049 21539
rect 16540 21508 17049 21536
rect 16540 21496 16546 21508
rect 17037 21505 17049 21508
rect 17083 21505 17095 21539
rect 17037 21499 17095 21505
rect 17604 21468 17632 21576
rect 17678 21564 17684 21576
rect 17736 21564 17742 21616
rect 21177 21607 21235 21613
rect 21177 21573 21189 21607
rect 21223 21604 21235 21607
rect 21910 21604 21916 21616
rect 21223 21576 21916 21604
rect 21223 21573 21235 21576
rect 21177 21567 21235 21573
rect 21910 21564 21916 21576
rect 21968 21564 21974 21616
rect 18598 21536 18604 21548
rect 17696 21508 18604 21536
rect 17696 21477 17724 21508
rect 18598 21496 18604 21508
rect 18656 21496 18662 21548
rect 21818 21536 21824 21548
rect 21779 21508 21824 21536
rect 21818 21496 21824 21508
rect 21876 21496 21882 21548
rect 16040 21440 17632 21468
rect 17681 21471 17739 21477
rect 15933 21431 15991 21437
rect 17681 21437 17693 21471
rect 17727 21437 17739 21471
rect 18322 21468 18328 21480
rect 18283 21440 18328 21468
rect 17681 21431 17739 21437
rect 18322 21428 18328 21440
rect 18380 21428 18386 21480
rect 18874 21468 18880 21480
rect 18835 21440 18880 21468
rect 18874 21428 18880 21440
rect 18932 21428 18938 21480
rect 19886 21468 19892 21480
rect 18984 21440 19892 21468
rect 6086 21400 6092 21412
rect 4080 21372 6092 21400
rect 6086 21360 6092 21372
rect 6144 21360 6150 21412
rect 6181 21403 6239 21409
rect 6181 21369 6193 21403
rect 6227 21400 6239 21403
rect 6454 21400 6460 21412
rect 6227 21372 6460 21400
rect 6227 21369 6239 21372
rect 6181 21363 6239 21369
rect 6454 21360 6460 21372
rect 6512 21360 6518 21412
rect 7006 21360 7012 21412
rect 7064 21400 7070 21412
rect 7929 21403 7987 21409
rect 7929 21400 7941 21403
rect 7064 21372 7941 21400
rect 7064 21360 7070 21372
rect 7929 21369 7941 21372
rect 7975 21369 7987 21403
rect 8846 21400 8852 21412
rect 8807 21372 8852 21400
rect 7929 21363 7987 21369
rect 8846 21360 8852 21372
rect 8904 21360 8910 21412
rect 10956 21403 11014 21409
rect 10956 21369 10968 21403
rect 11002 21400 11014 21403
rect 11790 21400 11796 21412
rect 11002 21372 11796 21400
rect 11002 21369 11014 21372
rect 10956 21363 11014 21369
rect 11790 21360 11796 21372
rect 11848 21400 11854 21412
rect 12989 21403 13047 21409
rect 12989 21400 13001 21403
rect 11848 21372 13001 21400
rect 11848 21360 11854 21372
rect 12989 21369 13001 21372
rect 13035 21369 13047 21403
rect 12989 21363 13047 21369
rect 14001 21403 14059 21409
rect 14001 21369 14013 21403
rect 14047 21400 14059 21403
rect 14458 21400 14464 21412
rect 14047 21372 14464 21400
rect 14047 21369 14059 21372
rect 14001 21363 14059 21369
rect 14458 21360 14464 21372
rect 14516 21360 14522 21412
rect 18984 21400 19012 21440
rect 19886 21428 19892 21440
rect 19944 21428 19950 21480
rect 20530 21468 20536 21480
rect 20491 21440 20536 21468
rect 20530 21428 20536 21440
rect 20588 21428 20594 21480
rect 22186 21468 22192 21480
rect 22147 21440 22192 21468
rect 22186 21428 22192 21440
rect 22244 21428 22250 21480
rect 15028 21372 19012 21400
rect 19144 21403 19202 21409
rect 1946 21332 1952 21344
rect 1907 21304 1952 21332
rect 1946 21292 1952 21304
rect 2004 21292 2010 21344
rect 2406 21292 2412 21344
rect 2464 21332 2470 21344
rect 2958 21332 2964 21344
rect 2464 21304 2509 21332
rect 2919 21304 2964 21332
rect 2464 21292 2470 21304
rect 2958 21292 2964 21304
rect 3016 21292 3022 21344
rect 3326 21332 3332 21344
rect 3287 21304 3332 21332
rect 3326 21292 3332 21304
rect 3384 21292 3390 21344
rect 3418 21292 3424 21344
rect 3476 21332 3482 21344
rect 4062 21332 4068 21344
rect 3476 21304 3521 21332
rect 4023 21304 4068 21332
rect 3476 21292 3482 21304
rect 4062 21292 4068 21304
rect 4120 21292 4126 21344
rect 4430 21332 4436 21344
rect 4391 21304 4436 21332
rect 4430 21292 4436 21304
rect 4488 21292 4494 21344
rect 4522 21292 4528 21344
rect 4580 21332 4586 21344
rect 5258 21332 5264 21344
rect 4580 21304 4625 21332
rect 5219 21304 5264 21332
rect 4580 21292 4586 21304
rect 5258 21292 5264 21304
rect 5316 21292 5322 21344
rect 5810 21332 5816 21344
rect 5771 21304 5816 21332
rect 5810 21292 5816 21304
rect 5868 21292 5874 21344
rect 6270 21332 6276 21344
rect 6231 21304 6276 21332
rect 6270 21292 6276 21304
rect 6328 21292 6334 21344
rect 6914 21332 6920 21344
rect 6875 21304 6920 21332
rect 6914 21292 6920 21304
rect 6972 21292 6978 21344
rect 7282 21332 7288 21344
rect 7243 21304 7288 21332
rect 7282 21292 7288 21304
rect 7340 21292 7346 21344
rect 7374 21292 7380 21344
rect 7432 21332 7438 21344
rect 8389 21335 8447 21341
rect 7432 21304 7477 21332
rect 7432 21292 7438 21304
rect 8389 21301 8401 21335
rect 8435 21332 8447 21335
rect 8662 21332 8668 21344
rect 8435 21304 8668 21332
rect 8435 21301 8447 21304
rect 8389 21295 8447 21301
rect 8662 21292 8668 21304
rect 8720 21292 8726 21344
rect 8754 21292 8760 21344
rect 8812 21332 8818 21344
rect 12066 21332 12072 21344
rect 8812 21304 8857 21332
rect 12027 21304 12072 21332
rect 8812 21292 8818 21304
rect 12066 21292 12072 21304
rect 12124 21292 12130 21344
rect 12621 21335 12679 21341
rect 12621 21301 12633 21335
rect 12667 21332 12679 21335
rect 12894 21332 12900 21344
rect 12667 21304 12900 21332
rect 12667 21301 12679 21304
rect 12621 21295 12679 21301
rect 12894 21292 12900 21304
rect 12952 21292 12958 21344
rect 13722 21292 13728 21344
rect 13780 21332 13786 21344
rect 15028 21341 15056 21372
rect 19144 21369 19156 21403
rect 19190 21400 19202 21403
rect 19334 21400 19340 21412
rect 19190 21372 19340 21400
rect 19190 21369 19202 21372
rect 19144 21363 19202 21369
rect 19334 21360 19340 21372
rect 19392 21360 19398 21412
rect 14093 21335 14151 21341
rect 14093 21332 14105 21335
rect 13780 21304 14105 21332
rect 13780 21292 13786 21304
rect 14093 21301 14105 21304
rect 14139 21301 14151 21335
rect 14093 21295 14151 21301
rect 15013 21335 15071 21341
rect 15013 21301 15025 21335
rect 15059 21301 15071 21335
rect 15013 21295 15071 21301
rect 15102 21292 15108 21344
rect 15160 21332 15166 21344
rect 15841 21335 15899 21341
rect 15841 21332 15853 21335
rect 15160 21304 15853 21332
rect 15160 21292 15166 21304
rect 15841 21301 15853 21304
rect 15887 21301 15899 21335
rect 15841 21295 15899 21301
rect 16298 21292 16304 21344
rect 16356 21332 16362 21344
rect 16485 21335 16543 21341
rect 16485 21332 16497 21335
rect 16356 21304 16497 21332
rect 16356 21292 16362 21304
rect 16485 21301 16497 21304
rect 16531 21301 16543 21335
rect 16850 21332 16856 21344
rect 16811 21304 16856 21332
rect 16485 21295 16543 21301
rect 16850 21292 16856 21304
rect 16908 21292 16914 21344
rect 16942 21292 16948 21344
rect 17000 21332 17006 21344
rect 17865 21335 17923 21341
rect 17000 21304 17045 21332
rect 17000 21292 17006 21304
rect 17865 21301 17877 21335
rect 17911 21332 17923 21335
rect 19242 21332 19248 21344
rect 17911 21304 19248 21332
rect 17911 21301 17923 21304
rect 17865 21295 17923 21301
rect 19242 21292 19248 21304
rect 19300 21292 19306 21344
rect 20254 21332 20260 21344
rect 20215 21304 20260 21332
rect 20254 21292 20260 21304
rect 20312 21292 20318 21344
rect 20717 21335 20775 21341
rect 20717 21301 20729 21335
rect 20763 21332 20775 21335
rect 21082 21332 21088 21344
rect 20763 21304 21088 21332
rect 20763 21301 20775 21304
rect 20717 21295 20775 21301
rect 21082 21292 21088 21304
rect 21140 21292 21146 21344
rect 21542 21332 21548 21344
rect 21503 21304 21548 21332
rect 21542 21292 21548 21304
rect 21600 21292 21606 21344
rect 21634 21292 21640 21344
rect 21692 21332 21698 21344
rect 21692 21304 21737 21332
rect 21692 21292 21698 21304
rect 22278 21292 22284 21344
rect 22336 21332 22342 21344
rect 22373 21335 22431 21341
rect 22373 21332 22385 21335
rect 22336 21304 22385 21332
rect 22336 21292 22342 21304
rect 22373 21301 22385 21304
rect 22419 21301 22431 21335
rect 22373 21295 22431 21301
rect 1104 21242 23276 21264
rect 1104 21190 8379 21242
rect 8431 21190 8443 21242
rect 8495 21190 8507 21242
rect 8559 21190 8571 21242
rect 8623 21190 15776 21242
rect 15828 21190 15840 21242
rect 15892 21190 15904 21242
rect 15956 21190 15968 21242
rect 16020 21190 23276 21242
rect 1104 21168 23276 21190
rect 290 21088 296 21140
rect 348 21128 354 21140
rect 1581 21131 1639 21137
rect 1581 21128 1593 21131
rect 348 21100 1593 21128
rect 348 21088 354 21100
rect 1581 21097 1593 21100
rect 1627 21097 1639 21131
rect 1581 21091 1639 21097
rect 4062 21088 4068 21140
rect 4120 21128 4126 21140
rect 4433 21131 4491 21137
rect 4433 21128 4445 21131
rect 4120 21100 4445 21128
rect 4120 21088 4126 21100
rect 4433 21097 4445 21100
rect 4479 21097 4491 21131
rect 4433 21091 4491 21097
rect 7193 21131 7251 21137
rect 7193 21097 7205 21131
rect 7239 21128 7251 21131
rect 7374 21128 7380 21140
rect 7239 21100 7380 21128
rect 7239 21097 7251 21100
rect 7193 21091 7251 21097
rect 7374 21088 7380 21100
rect 7432 21088 7438 21140
rect 8846 21088 8852 21140
rect 8904 21128 8910 21140
rect 8941 21131 8999 21137
rect 8941 21128 8953 21131
rect 8904 21100 8953 21128
rect 8904 21088 8910 21100
rect 8941 21097 8953 21100
rect 8987 21097 8999 21131
rect 8941 21091 8999 21097
rect 11514 21088 11520 21140
rect 11572 21128 11578 21140
rect 16942 21128 16948 21140
rect 11572 21100 16948 21128
rect 11572 21088 11578 21100
rect 16942 21088 16948 21100
rect 17000 21088 17006 21140
rect 17129 21131 17187 21137
rect 17129 21097 17141 21131
rect 17175 21128 17187 21131
rect 19150 21128 19156 21140
rect 17175 21100 19156 21128
rect 17175 21097 17187 21100
rect 17129 21091 17187 21097
rect 19150 21088 19156 21100
rect 19208 21088 19214 21140
rect 20533 21131 20591 21137
rect 19260 21100 20392 21128
rect 2958 21020 2964 21072
rect 3016 21060 3022 21072
rect 4525 21063 4583 21069
rect 4525 21060 4537 21063
rect 3016 21032 4537 21060
rect 3016 21020 3022 21032
rect 4525 21029 4537 21032
rect 4571 21029 4583 21063
rect 5442 21060 5448 21072
rect 4525 21023 4583 21029
rect 4632 21032 5448 21060
rect 1397 20995 1455 21001
rect 1397 20961 1409 20995
rect 1443 20961 1455 20995
rect 1397 20955 1455 20961
rect 2216 20995 2274 21001
rect 2216 20961 2228 20995
rect 2262 20992 2274 20995
rect 3418 20992 3424 21004
rect 2262 20964 3424 20992
rect 2262 20961 2274 20964
rect 2216 20955 2274 20961
rect 1412 20788 1440 20955
rect 3418 20952 3424 20964
rect 3476 20952 3482 21004
rect 1762 20884 1768 20936
rect 1820 20924 1826 20936
rect 1949 20927 2007 20933
rect 1949 20924 1961 20927
rect 1820 20896 1961 20924
rect 1820 20884 1826 20896
rect 1949 20893 1961 20896
rect 1995 20893 2007 20927
rect 4338 20924 4344 20936
rect 1949 20887 2007 20893
rect 3160 20896 4344 20924
rect 3160 20788 3188 20896
rect 4338 20884 4344 20896
rect 4396 20924 4402 20936
rect 4632 20924 4660 21032
rect 5442 21020 5448 21032
rect 5500 21020 5506 21072
rect 5736 21032 6868 21060
rect 5077 20995 5135 21001
rect 5077 20961 5089 20995
rect 5123 20992 5135 20995
rect 5166 20992 5172 21004
rect 5123 20964 5172 20992
rect 5123 20961 5135 20964
rect 5077 20955 5135 20961
rect 5166 20952 5172 20964
rect 5224 20952 5230 21004
rect 4396 20896 4660 20924
rect 4709 20927 4767 20933
rect 4396 20884 4402 20896
rect 4709 20893 4721 20927
rect 4755 20924 4767 20927
rect 5736 20924 5764 21032
rect 6840 21004 6868 21032
rect 7282 21020 7288 21072
rect 7340 21060 7346 21072
rect 7806 21063 7864 21069
rect 7806 21060 7818 21063
rect 7340 21032 7818 21060
rect 7340 21020 7346 21032
rect 7806 21029 7818 21032
rect 7852 21060 7864 21063
rect 8202 21060 8208 21072
rect 7852 21032 8208 21060
rect 7852 21029 7864 21032
rect 7806 21023 7864 21029
rect 8202 21020 8208 21032
rect 8260 21020 8266 21072
rect 8662 21020 8668 21072
rect 8720 21060 8726 21072
rect 10137 21063 10195 21069
rect 10137 21060 10149 21063
rect 8720 21032 10149 21060
rect 8720 21020 8726 21032
rect 10137 21029 10149 21032
rect 10183 21029 10195 21063
rect 10137 21023 10195 21029
rect 11324 21063 11382 21069
rect 11324 21029 11336 21063
rect 11370 21060 11382 21063
rect 12066 21060 12072 21072
rect 11370 21032 12072 21060
rect 11370 21029 11382 21032
rect 11324 21023 11382 21029
rect 12066 21020 12072 21032
rect 12124 21060 12130 21072
rect 13348 21063 13406 21069
rect 12124 21032 13308 21060
rect 12124 21020 12130 21032
rect 6080 20995 6138 21001
rect 6080 20961 6092 20995
rect 6126 20992 6138 20995
rect 6454 20992 6460 21004
rect 6126 20964 6460 20992
rect 6126 20961 6138 20964
rect 6080 20955 6138 20961
rect 6454 20952 6460 20964
rect 6512 20952 6518 21004
rect 6822 20952 6828 21004
rect 6880 20992 6886 21004
rect 10042 20992 10048 21004
rect 6880 20964 8616 20992
rect 10003 20964 10048 20992
rect 6880 20952 6886 20964
rect 4755 20896 5764 20924
rect 5813 20927 5871 20933
rect 4755 20893 4767 20896
rect 4709 20887 4767 20893
rect 5813 20893 5825 20927
rect 5859 20893 5871 20927
rect 7558 20924 7564 20936
rect 7519 20896 7564 20924
rect 5813 20887 5871 20893
rect 3878 20816 3884 20868
rect 3936 20856 3942 20868
rect 5261 20859 5319 20865
rect 5261 20856 5273 20859
rect 3936 20828 5273 20856
rect 3936 20816 3942 20828
rect 5261 20825 5273 20828
rect 5307 20825 5319 20859
rect 5261 20819 5319 20825
rect 3326 20788 3332 20800
rect 1412 20760 3188 20788
rect 3287 20760 3332 20788
rect 3326 20748 3332 20760
rect 3384 20748 3390 20800
rect 3970 20748 3976 20800
rect 4028 20788 4034 20800
rect 4065 20791 4123 20797
rect 4065 20788 4077 20791
rect 4028 20760 4077 20788
rect 4028 20748 4034 20760
rect 4065 20757 4077 20760
rect 4111 20757 4123 20791
rect 4065 20751 4123 20757
rect 5074 20748 5080 20800
rect 5132 20788 5138 20800
rect 5828 20788 5856 20887
rect 7558 20884 7564 20896
rect 7616 20884 7622 20936
rect 8588 20924 8616 20964
rect 10042 20952 10048 20964
rect 10100 20952 10106 21004
rect 13081 20995 13139 21001
rect 13081 20961 13093 20995
rect 13127 20992 13139 20995
rect 13170 20992 13176 21004
rect 13127 20964 13176 20992
rect 13127 20961 13139 20964
rect 13081 20955 13139 20961
rect 13170 20952 13176 20964
rect 13228 20952 13234 21004
rect 13280 20992 13308 21032
rect 13348 21029 13360 21063
rect 13394 21060 13406 21063
rect 13722 21060 13728 21072
rect 13394 21032 13728 21060
rect 13394 21029 13406 21032
rect 13348 21023 13406 21029
rect 13722 21020 13728 21032
rect 13780 21020 13786 21072
rect 18046 21060 18052 21072
rect 17512 21032 18052 21060
rect 13814 20992 13820 21004
rect 13280 20964 13820 20992
rect 13814 20952 13820 20964
rect 13872 20952 13878 21004
rect 14642 20952 14648 21004
rect 14700 20992 14706 21004
rect 17512 21001 17540 21032
rect 18046 21020 18052 21032
rect 18104 21060 18110 21072
rect 18874 21060 18880 21072
rect 18104 21032 18880 21060
rect 18104 21020 18110 21032
rect 18874 21020 18880 21032
rect 18932 21060 18938 21072
rect 19061 21063 19119 21069
rect 19061 21060 19073 21063
rect 18932 21032 19073 21060
rect 18932 21020 18938 21032
rect 19061 21029 19073 21032
rect 19107 21060 19119 21063
rect 19260 21060 19288 21100
rect 19107 21032 19288 21060
rect 19420 21063 19478 21069
rect 19107 21029 19119 21032
rect 19061 21023 19119 21029
rect 19420 21029 19432 21063
rect 19466 21060 19478 21063
rect 20254 21060 20260 21072
rect 19466 21032 20260 21060
rect 19466 21029 19478 21032
rect 19420 21023 19478 21029
rect 20254 21020 20260 21032
rect 20312 21020 20318 21072
rect 15545 20995 15603 21001
rect 15545 20992 15557 20995
rect 14700 20964 15557 20992
rect 14700 20952 14706 20964
rect 15545 20961 15557 20964
rect 15591 20961 15603 20995
rect 15545 20955 15603 20961
rect 16945 20995 17003 21001
rect 16945 20961 16957 20995
rect 16991 20961 17003 20995
rect 16945 20955 17003 20961
rect 17497 20995 17555 21001
rect 17497 20961 17509 20995
rect 17543 20961 17555 20995
rect 17497 20955 17555 20961
rect 17764 20995 17822 21001
rect 17764 20961 17776 20995
rect 17810 20992 17822 20995
rect 19794 20992 19800 21004
rect 17810 20964 19800 20992
rect 17810 20961 17822 20964
rect 17764 20955 17822 20961
rect 10229 20927 10287 20933
rect 10229 20924 10241 20927
rect 8588 20896 10241 20924
rect 10229 20893 10241 20896
rect 10275 20893 10287 20927
rect 10229 20887 10287 20893
rect 10410 20884 10416 20936
rect 10468 20924 10474 20936
rect 11057 20927 11115 20933
rect 11057 20924 11069 20927
rect 10468 20896 11069 20924
rect 10468 20884 10474 20896
rect 11057 20893 11069 20896
rect 11103 20893 11115 20927
rect 15286 20924 15292 20936
rect 15247 20896 15292 20924
rect 11057 20887 11115 20893
rect 15286 20884 15292 20896
rect 15344 20884 15350 20936
rect 6546 20788 6552 20800
rect 5132 20760 6552 20788
rect 5132 20748 5138 20760
rect 6546 20748 6552 20760
rect 6604 20748 6610 20800
rect 9677 20791 9735 20797
rect 9677 20757 9689 20791
rect 9723 20788 9735 20791
rect 9766 20788 9772 20800
rect 9723 20760 9772 20788
rect 9723 20757 9735 20760
rect 9677 20751 9735 20757
rect 9766 20748 9772 20760
rect 9824 20748 9830 20800
rect 12434 20748 12440 20800
rect 12492 20788 12498 20800
rect 14458 20788 14464 20800
rect 12492 20760 12537 20788
rect 14419 20760 14464 20788
rect 12492 20748 12498 20760
rect 14458 20748 14464 20760
rect 14516 20748 14522 20800
rect 14550 20748 14556 20800
rect 14608 20788 14614 20800
rect 15102 20788 15108 20800
rect 14608 20760 15108 20788
rect 14608 20748 14614 20760
rect 15102 20748 15108 20760
rect 15160 20748 15166 20800
rect 15194 20748 15200 20800
rect 15252 20788 15258 20800
rect 16669 20791 16727 20797
rect 16669 20788 16681 20791
rect 15252 20760 16681 20788
rect 15252 20748 15258 20760
rect 16669 20757 16681 20760
rect 16715 20757 16727 20791
rect 16960 20788 16988 20955
rect 19794 20952 19800 20964
rect 19852 20952 19858 21004
rect 20364 20992 20392 21100
rect 20533 21097 20545 21131
rect 20579 21097 20591 21131
rect 20533 21091 20591 21097
rect 20548 21060 20576 21091
rect 21168 21063 21226 21069
rect 21168 21060 21180 21063
rect 20548 21032 21180 21060
rect 21168 21029 21180 21032
rect 21214 21060 21226 21063
rect 21634 21060 21640 21072
rect 21214 21032 21640 21060
rect 21214 21029 21226 21032
rect 21168 21023 21226 21029
rect 21634 21020 21640 21032
rect 21692 21020 21698 21072
rect 20364 20964 20944 20992
rect 20916 20936 20944 20964
rect 19061 20927 19119 20933
rect 19061 20893 19073 20927
rect 19107 20924 19119 20927
rect 19153 20927 19211 20933
rect 19153 20924 19165 20927
rect 19107 20896 19165 20924
rect 19107 20893 19119 20896
rect 19061 20887 19119 20893
rect 19153 20893 19165 20896
rect 19199 20893 19211 20927
rect 20898 20924 20904 20936
rect 20859 20896 20904 20924
rect 19153 20887 19211 20893
rect 20898 20884 20904 20896
rect 20956 20884 20962 20936
rect 17770 20788 17776 20800
rect 16960 20760 17776 20788
rect 16669 20751 16727 20757
rect 17770 20748 17776 20760
rect 17828 20748 17834 20800
rect 18877 20791 18935 20797
rect 18877 20757 18889 20791
rect 18923 20788 18935 20791
rect 19334 20788 19340 20800
rect 18923 20760 19340 20788
rect 18923 20757 18935 20760
rect 18877 20751 18935 20757
rect 19334 20748 19340 20760
rect 19392 20788 19398 20800
rect 20162 20788 20168 20800
rect 19392 20760 20168 20788
rect 19392 20748 19398 20760
rect 20162 20748 20168 20760
rect 20220 20748 20226 20800
rect 21542 20748 21548 20800
rect 21600 20788 21606 20800
rect 22281 20791 22339 20797
rect 22281 20788 22293 20791
rect 21600 20760 22293 20788
rect 21600 20748 21606 20760
rect 22281 20757 22293 20760
rect 22327 20757 22339 20791
rect 22281 20751 22339 20757
rect 1104 20698 23276 20720
rect 1104 20646 4680 20698
rect 4732 20646 4744 20698
rect 4796 20646 4808 20698
rect 4860 20646 4872 20698
rect 4924 20646 12078 20698
rect 12130 20646 12142 20698
rect 12194 20646 12206 20698
rect 12258 20646 12270 20698
rect 12322 20646 19475 20698
rect 19527 20646 19539 20698
rect 19591 20646 19603 20698
rect 19655 20646 19667 20698
rect 19719 20646 23276 20698
rect 1104 20624 23276 20646
rect 3053 20587 3111 20593
rect 3053 20553 3065 20587
rect 3099 20584 3111 20587
rect 3418 20584 3424 20596
rect 3099 20556 3424 20584
rect 3099 20553 3111 20556
rect 3053 20547 3111 20553
rect 3418 20544 3424 20556
rect 3476 20544 3482 20596
rect 4430 20544 4436 20596
rect 4488 20584 4494 20596
rect 4801 20587 4859 20593
rect 4801 20584 4813 20587
rect 4488 20556 4813 20584
rect 4488 20544 4494 20556
rect 4801 20553 4813 20556
rect 4847 20553 4859 20587
rect 6454 20584 6460 20596
rect 6415 20556 6460 20584
rect 4801 20547 4859 20553
rect 6454 20544 6460 20556
rect 6512 20544 6518 20596
rect 6546 20544 6552 20596
rect 6604 20584 6610 20596
rect 7558 20584 7564 20596
rect 6604 20556 7564 20584
rect 6604 20544 6610 20556
rect 5074 20448 5080 20460
rect 5035 20420 5080 20448
rect 5074 20408 5080 20420
rect 5132 20408 5138 20460
rect 6840 20457 6868 20556
rect 7558 20544 7564 20556
rect 7616 20544 7622 20596
rect 8202 20584 8208 20596
rect 8163 20556 8208 20584
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 8754 20544 8760 20596
rect 8812 20584 8818 20596
rect 9861 20587 9919 20593
rect 9861 20584 9873 20587
rect 8812 20556 9873 20584
rect 8812 20544 8818 20556
rect 9861 20553 9873 20556
rect 9907 20553 9919 20587
rect 11790 20584 11796 20596
rect 9861 20547 9919 20553
rect 10428 20556 11376 20584
rect 11751 20556 11796 20584
rect 9490 20476 9496 20528
rect 9548 20516 9554 20528
rect 10428 20516 10456 20556
rect 9548 20488 10456 20516
rect 11348 20516 11376 20556
rect 11790 20544 11796 20556
rect 11848 20544 11854 20596
rect 12897 20587 12955 20593
rect 12897 20553 12909 20587
rect 12943 20584 12955 20587
rect 14642 20584 14648 20596
rect 12943 20556 14504 20584
rect 14603 20556 14648 20584
rect 12943 20553 12955 20556
rect 12897 20547 12955 20553
rect 13078 20516 13084 20528
rect 11348 20488 13084 20516
rect 9548 20476 9554 20488
rect 13078 20476 13084 20488
rect 13136 20476 13142 20528
rect 14476 20516 14504 20556
rect 14642 20544 14648 20556
rect 14700 20544 14706 20596
rect 19058 20584 19064 20596
rect 14936 20556 19064 20584
rect 14936 20516 14964 20556
rect 19058 20544 19064 20556
rect 19116 20544 19122 20596
rect 19429 20587 19487 20593
rect 19429 20553 19441 20587
rect 19475 20584 19487 20587
rect 19794 20584 19800 20596
rect 19475 20556 19800 20584
rect 19475 20553 19487 20556
rect 19429 20547 19487 20553
rect 19794 20544 19800 20556
rect 19852 20544 19858 20596
rect 21818 20584 21824 20596
rect 20364 20556 21824 20584
rect 14476 20488 14964 20516
rect 16206 20476 16212 20528
rect 16264 20516 16270 20528
rect 16264 20488 17172 20516
rect 16264 20476 16270 20488
rect 6825 20451 6883 20457
rect 6825 20417 6837 20451
rect 6871 20417 6883 20451
rect 6825 20411 6883 20417
rect 11422 20408 11428 20460
rect 11480 20448 11486 20460
rect 11480 20420 13400 20448
rect 11480 20408 11486 20420
rect 1673 20383 1731 20389
rect 1673 20349 1685 20383
rect 1719 20380 1731 20383
rect 1762 20380 1768 20392
rect 1719 20352 1768 20380
rect 1719 20349 1731 20352
rect 1673 20343 1731 20349
rect 1762 20340 1768 20352
rect 1820 20380 1826 20392
rect 3418 20380 3424 20392
rect 1820 20352 3424 20380
rect 1820 20340 1826 20352
rect 3418 20340 3424 20352
rect 3476 20340 3482 20392
rect 3688 20383 3746 20389
rect 3688 20349 3700 20383
rect 3734 20380 3746 20383
rect 4522 20380 4528 20392
rect 3734 20352 4528 20380
rect 3734 20349 3746 20352
rect 3688 20343 3746 20349
rect 4522 20340 4528 20352
rect 4580 20340 4586 20392
rect 5344 20383 5402 20389
rect 5344 20349 5356 20383
rect 5390 20380 5402 20383
rect 6270 20380 6276 20392
rect 5390 20352 6276 20380
rect 5390 20349 5402 20352
rect 5344 20343 5402 20349
rect 6270 20340 6276 20352
rect 6328 20340 6334 20392
rect 7092 20383 7150 20389
rect 7092 20349 7104 20383
rect 7138 20380 7150 20383
rect 7374 20380 7380 20392
rect 7138 20352 7380 20380
rect 7138 20349 7150 20352
rect 7092 20343 7150 20349
rect 7374 20340 7380 20352
rect 7432 20340 7438 20392
rect 8018 20340 8024 20392
rect 8076 20380 8082 20392
rect 8481 20383 8539 20389
rect 8481 20380 8493 20383
rect 8076 20352 8493 20380
rect 8076 20340 8082 20352
rect 8481 20349 8493 20352
rect 8527 20380 8539 20383
rect 10410 20380 10416 20392
rect 8527 20352 10416 20380
rect 8527 20349 8539 20352
rect 8481 20343 8539 20349
rect 10410 20340 10416 20352
rect 10468 20340 10474 20392
rect 10680 20383 10738 20389
rect 10680 20349 10692 20383
rect 10726 20380 10738 20383
rect 11974 20380 11980 20392
rect 10726 20352 11980 20380
rect 10726 20349 10738 20352
rect 10680 20343 10738 20349
rect 11974 20340 11980 20352
rect 12032 20340 12038 20392
rect 12713 20383 12771 20389
rect 12713 20349 12725 20383
rect 12759 20349 12771 20383
rect 12713 20343 12771 20349
rect 1940 20315 1998 20321
rect 1940 20281 1952 20315
rect 1986 20312 1998 20315
rect 2038 20312 2044 20324
rect 1986 20284 2044 20312
rect 1986 20281 1998 20284
rect 1940 20275 1998 20281
rect 2038 20272 2044 20284
rect 2096 20272 2102 20324
rect 4246 20272 4252 20324
rect 4304 20312 4310 20324
rect 6638 20312 6644 20324
rect 4304 20284 6644 20312
rect 4304 20272 4310 20284
rect 6638 20272 6644 20284
rect 6696 20272 6702 20324
rect 8748 20315 8806 20321
rect 8748 20281 8760 20315
rect 8794 20312 8806 20315
rect 8846 20312 8852 20324
rect 8794 20284 8852 20312
rect 8794 20281 8806 20284
rect 8748 20275 8806 20281
rect 8846 20272 8852 20284
rect 8904 20272 8910 20324
rect 9030 20272 9036 20324
rect 9088 20312 9094 20324
rect 11330 20312 11336 20324
rect 9088 20284 11336 20312
rect 9088 20272 9094 20284
rect 11330 20272 11336 20284
rect 11388 20272 11394 20324
rect 11422 20272 11428 20324
rect 11480 20312 11486 20324
rect 12526 20312 12532 20324
rect 11480 20284 12532 20312
rect 11480 20272 11486 20284
rect 12526 20272 12532 20284
rect 12584 20272 12590 20324
rect 12728 20312 12756 20343
rect 13170 20340 13176 20392
rect 13228 20380 13234 20392
rect 13265 20383 13323 20389
rect 13265 20380 13277 20383
rect 13228 20352 13277 20380
rect 13228 20340 13234 20352
rect 13265 20349 13277 20352
rect 13311 20349 13323 20383
rect 13372 20380 13400 20420
rect 16114 20408 16120 20460
rect 16172 20448 16178 20460
rect 16574 20448 16580 20460
rect 16172 20420 16580 20448
rect 16172 20408 16178 20420
rect 16574 20408 16580 20420
rect 16632 20408 16638 20460
rect 16758 20408 16764 20460
rect 16816 20448 16822 20460
rect 17144 20457 17172 20488
rect 20364 20460 20392 20556
rect 21818 20544 21824 20556
rect 21876 20544 21882 20596
rect 17037 20451 17095 20457
rect 17037 20448 17049 20451
rect 16816 20420 17049 20448
rect 16816 20408 16822 20420
rect 17037 20417 17049 20420
rect 17083 20417 17095 20451
rect 17037 20411 17095 20417
rect 17129 20451 17187 20457
rect 17129 20417 17141 20451
rect 17175 20417 17187 20451
rect 20162 20448 20168 20460
rect 20123 20420 20168 20448
rect 17129 20411 17187 20417
rect 20162 20408 20168 20420
rect 20220 20408 20226 20460
rect 20346 20448 20352 20460
rect 20259 20420 20352 20448
rect 20346 20408 20352 20420
rect 20404 20408 20410 20460
rect 13532 20383 13590 20389
rect 13372 20352 13492 20380
rect 13265 20343 13323 20349
rect 13354 20312 13360 20324
rect 12728 20284 13360 20312
rect 13354 20272 13360 20284
rect 13412 20272 13418 20324
rect 13464 20312 13492 20352
rect 13532 20349 13544 20383
rect 13578 20380 13590 20383
rect 14458 20380 14464 20392
rect 13578 20352 14464 20380
rect 13578 20349 13590 20352
rect 13532 20343 13590 20349
rect 14458 20340 14464 20352
rect 14516 20340 14522 20392
rect 15194 20389 15200 20392
rect 14829 20383 14887 20389
rect 14829 20349 14841 20383
rect 14875 20380 14887 20383
rect 14921 20383 14979 20389
rect 14921 20380 14933 20383
rect 14875 20352 14933 20380
rect 14875 20349 14887 20352
rect 14829 20343 14887 20349
rect 14921 20349 14933 20352
rect 14967 20349 14979 20383
rect 15188 20380 15200 20389
rect 15155 20352 15200 20380
rect 14921 20343 14979 20349
rect 15188 20343 15200 20352
rect 15194 20340 15200 20343
rect 15252 20340 15258 20392
rect 18046 20380 18052 20392
rect 15304 20352 17080 20380
rect 18007 20352 18052 20380
rect 15304 20312 15332 20352
rect 13464 20284 15332 20312
rect 15470 20272 15476 20324
rect 15528 20312 15534 20324
rect 16945 20315 17003 20321
rect 16945 20312 16957 20315
rect 15528 20284 16957 20312
rect 15528 20272 15534 20284
rect 16945 20281 16957 20284
rect 16991 20281 17003 20315
rect 17052 20312 17080 20352
rect 18046 20340 18052 20352
rect 18104 20340 18110 20392
rect 20809 20383 20867 20389
rect 18156 20352 20392 20380
rect 18156 20312 18184 20352
rect 17052 20284 18184 20312
rect 18316 20315 18374 20321
rect 16945 20275 17003 20281
rect 18316 20281 18328 20315
rect 18362 20312 18374 20315
rect 19150 20312 19156 20324
rect 18362 20284 19156 20312
rect 18362 20281 18374 20284
rect 18316 20275 18374 20281
rect 19150 20272 19156 20284
rect 19208 20272 19214 20324
rect 19978 20312 19984 20324
rect 19260 20284 19984 20312
rect 842 20204 848 20256
rect 900 20244 906 20256
rect 5258 20244 5264 20256
rect 900 20216 5264 20244
rect 900 20204 906 20216
rect 5258 20204 5264 20216
rect 5316 20204 5322 20256
rect 5442 20204 5448 20256
rect 5500 20244 5506 20256
rect 12158 20244 12164 20256
rect 5500 20216 12164 20244
rect 5500 20204 5506 20216
rect 12158 20204 12164 20216
rect 12216 20204 12222 20256
rect 12250 20204 12256 20256
rect 12308 20244 12314 20256
rect 12710 20244 12716 20256
rect 12308 20216 12716 20244
rect 12308 20204 12314 20216
rect 12710 20204 12716 20216
rect 12768 20204 12774 20256
rect 12802 20204 12808 20256
rect 12860 20244 12866 20256
rect 13170 20244 13176 20256
rect 12860 20216 13176 20244
rect 12860 20204 12866 20216
rect 13170 20204 13176 20216
rect 13228 20244 13234 20256
rect 14829 20247 14887 20253
rect 14829 20244 14841 20247
rect 13228 20216 14841 20244
rect 13228 20204 13234 20216
rect 14829 20213 14841 20216
rect 14875 20244 14887 20247
rect 15286 20244 15292 20256
rect 14875 20216 15292 20244
rect 14875 20213 14887 20216
rect 14829 20207 14887 20213
rect 15286 20204 15292 20216
rect 15344 20204 15350 20256
rect 16298 20244 16304 20256
rect 16259 20216 16304 20244
rect 16298 20204 16304 20216
rect 16356 20204 16362 20256
rect 16577 20247 16635 20253
rect 16577 20213 16589 20247
rect 16623 20244 16635 20247
rect 17034 20244 17040 20256
rect 16623 20216 17040 20244
rect 16623 20213 16635 20216
rect 16577 20207 16635 20213
rect 17034 20204 17040 20216
rect 17092 20204 17098 20256
rect 17218 20204 17224 20256
rect 17276 20244 17282 20256
rect 19260 20244 19288 20284
rect 19978 20272 19984 20284
rect 20036 20272 20042 20324
rect 20073 20315 20131 20321
rect 20073 20281 20085 20315
rect 20119 20312 20131 20315
rect 20254 20312 20260 20324
rect 20119 20284 20260 20312
rect 20119 20281 20131 20284
rect 20073 20275 20131 20281
rect 20254 20272 20260 20284
rect 20312 20272 20318 20324
rect 20364 20312 20392 20352
rect 20809 20349 20821 20383
rect 20855 20380 20867 20383
rect 20898 20380 20904 20392
rect 20855 20352 20904 20380
rect 20855 20349 20867 20352
rect 20809 20343 20867 20349
rect 20898 20340 20904 20352
rect 20956 20340 20962 20392
rect 21076 20383 21134 20389
rect 21076 20349 21088 20383
rect 21122 20380 21134 20383
rect 21542 20380 21548 20392
rect 21122 20352 21548 20380
rect 21122 20349 21134 20352
rect 21076 20343 21134 20349
rect 21542 20340 21548 20352
rect 21600 20340 21606 20392
rect 22465 20383 22523 20389
rect 22465 20349 22477 20383
rect 22511 20380 22523 20383
rect 22554 20380 22560 20392
rect 22511 20352 22560 20380
rect 22511 20349 22523 20352
rect 22465 20343 22523 20349
rect 22554 20340 22560 20352
rect 22612 20340 22618 20392
rect 21450 20312 21456 20324
rect 20364 20284 21456 20312
rect 21450 20272 21456 20284
rect 21508 20272 21514 20324
rect 24026 20312 24032 20324
rect 21560 20284 24032 20312
rect 17276 20216 19288 20244
rect 19705 20247 19763 20253
rect 17276 20204 17282 20216
rect 19705 20213 19717 20247
rect 19751 20244 19763 20247
rect 20162 20244 20168 20256
rect 19751 20216 20168 20244
rect 19751 20213 19763 20216
rect 19705 20207 19763 20213
rect 20162 20204 20168 20216
rect 20220 20204 20226 20256
rect 20438 20204 20444 20256
rect 20496 20244 20502 20256
rect 21560 20244 21588 20284
rect 24026 20272 24032 20284
rect 24084 20272 24090 20324
rect 20496 20216 21588 20244
rect 20496 20204 20502 20216
rect 21726 20204 21732 20256
rect 21784 20244 21790 20256
rect 22189 20247 22247 20253
rect 22189 20244 22201 20247
rect 21784 20216 22201 20244
rect 21784 20204 21790 20216
rect 22189 20213 22201 20216
rect 22235 20213 22247 20247
rect 22189 20207 22247 20213
rect 22649 20247 22707 20253
rect 22649 20213 22661 20247
rect 22695 20244 22707 20247
rect 22922 20244 22928 20256
rect 22695 20216 22928 20244
rect 22695 20213 22707 20216
rect 22649 20207 22707 20213
rect 22922 20204 22928 20216
rect 22980 20204 22986 20256
rect 1104 20154 23276 20176
rect 1104 20102 8379 20154
rect 8431 20102 8443 20154
rect 8495 20102 8507 20154
rect 8559 20102 8571 20154
rect 8623 20102 15776 20154
rect 15828 20102 15840 20154
rect 15892 20102 15904 20154
rect 15956 20102 15968 20154
rect 16020 20102 23276 20154
rect 1104 20080 23276 20102
rect 2130 20000 2136 20052
rect 2188 20040 2194 20052
rect 3237 20043 3295 20049
rect 3237 20040 3249 20043
rect 2188 20012 3249 20040
rect 2188 20000 2194 20012
rect 3237 20009 3249 20012
rect 3283 20009 3295 20043
rect 3237 20003 3295 20009
rect 4154 20000 4160 20052
rect 4212 20040 4218 20052
rect 4212 20012 4936 20040
rect 4212 20000 4218 20012
rect 1762 19932 1768 19984
rect 1820 19972 1826 19984
rect 3786 19972 3792 19984
rect 1820 19944 3792 19972
rect 1820 19932 1826 19944
rect 3786 19932 3792 19944
rect 3844 19932 3850 19984
rect 4430 19932 4436 19984
rect 4488 19972 4494 19984
rect 4678 19975 4736 19981
rect 4678 19972 4690 19975
rect 4488 19944 4690 19972
rect 4488 19932 4494 19944
rect 4678 19941 4690 19944
rect 4724 19941 4736 19975
rect 4908 19972 4936 20012
rect 4982 20000 4988 20052
rect 5040 20040 5046 20052
rect 5442 20040 5448 20052
rect 5040 20012 5448 20040
rect 5040 20000 5046 20012
rect 5442 20000 5448 20012
rect 5500 20000 5506 20052
rect 6549 20043 6607 20049
rect 6549 20009 6561 20043
rect 6595 20040 6607 20043
rect 6914 20040 6920 20052
rect 6595 20012 6920 20040
rect 6595 20009 6607 20012
rect 6549 20003 6607 20009
rect 6914 20000 6920 20012
rect 6972 20000 6978 20052
rect 7837 20043 7895 20049
rect 7837 20009 7849 20043
rect 7883 20040 7895 20043
rect 9214 20040 9220 20052
rect 7883 20012 9220 20040
rect 7883 20009 7895 20012
rect 7837 20003 7895 20009
rect 9214 20000 9220 20012
rect 9272 20000 9278 20052
rect 9858 20000 9864 20052
rect 9916 20000 9922 20052
rect 11793 20043 11851 20049
rect 11793 20009 11805 20043
rect 11839 20040 11851 20043
rect 11974 20040 11980 20052
rect 11839 20012 11980 20040
rect 11839 20009 11851 20012
rect 11793 20003 11851 20009
rect 11974 20000 11980 20012
rect 12032 20000 12038 20052
rect 13449 20043 13507 20049
rect 13449 20009 13461 20043
rect 13495 20040 13507 20043
rect 13722 20040 13728 20052
rect 13495 20012 13728 20040
rect 13495 20009 13507 20012
rect 13449 20003 13507 20009
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 13814 20000 13820 20052
rect 13872 20040 13878 20052
rect 14001 20043 14059 20049
rect 14001 20040 14013 20043
rect 13872 20012 14013 20040
rect 13872 20000 13878 20012
rect 14001 20009 14013 20012
rect 14047 20009 14059 20043
rect 14001 20003 14059 20009
rect 15580 20012 17356 20040
rect 4908 19944 5764 19972
rect 4678 19935 4736 19941
rect 1664 19907 1722 19913
rect 1664 19873 1676 19907
rect 1710 19904 1722 19907
rect 2774 19904 2780 19916
rect 1710 19876 2780 19904
rect 1710 19873 1722 19876
rect 1664 19867 1722 19873
rect 2774 19864 2780 19876
rect 2832 19864 2838 19916
rect 3053 19907 3111 19913
rect 3053 19873 3065 19907
rect 3099 19873 3111 19907
rect 3053 19867 3111 19873
rect 1394 19836 1400 19848
rect 1355 19808 1400 19836
rect 1394 19796 1400 19808
rect 1452 19796 1458 19848
rect 3068 19836 3096 19867
rect 3418 19864 3424 19916
rect 3476 19904 3482 19916
rect 5074 19904 5080 19916
rect 3476 19876 5080 19904
rect 3476 19864 3482 19876
rect 4062 19836 4068 19848
rect 3068 19808 4068 19836
rect 4062 19796 4068 19808
rect 4120 19796 4126 19848
rect 4448 19845 4476 19876
rect 5074 19864 5080 19876
rect 5132 19864 5138 19916
rect 5736 19904 5764 19944
rect 5810 19932 5816 19984
rect 5868 19972 5874 19984
rect 6641 19975 6699 19981
rect 6641 19972 6653 19975
rect 5868 19944 6653 19972
rect 5868 19932 5874 19944
rect 6641 19941 6653 19944
rect 6687 19941 6699 19975
rect 9677 19975 9735 19981
rect 6641 19935 6699 19941
rect 7300 19944 9536 19972
rect 7300 19904 7328 19944
rect 5736 19876 7328 19904
rect 7377 19907 7435 19913
rect 7377 19873 7389 19907
rect 7423 19904 7435 19907
rect 7837 19907 7895 19913
rect 7837 19904 7849 19907
rect 7423 19876 7849 19904
rect 7423 19873 7435 19876
rect 7377 19867 7435 19873
rect 7837 19873 7849 19876
rect 7883 19873 7895 19907
rect 7837 19867 7895 19873
rect 7929 19907 7987 19913
rect 7929 19873 7941 19907
rect 7975 19904 7987 19907
rect 8018 19904 8024 19916
rect 7975 19876 8024 19904
rect 7975 19873 7987 19876
rect 7929 19867 7987 19873
rect 8018 19864 8024 19876
rect 8076 19864 8082 19916
rect 8202 19913 8208 19916
rect 8196 19867 8208 19913
rect 8260 19904 8266 19916
rect 8260 19876 8296 19904
rect 8202 19864 8208 19867
rect 8260 19864 8266 19876
rect 4433 19839 4491 19845
rect 4433 19805 4445 19839
rect 4479 19805 4491 19839
rect 4433 19799 4491 19805
rect 5442 19796 5448 19848
rect 5500 19836 5506 19848
rect 6822 19836 6828 19848
rect 5500 19808 6408 19836
rect 6783 19808 6828 19836
rect 5500 19796 5506 19808
rect 5813 19771 5871 19777
rect 5813 19737 5825 19771
rect 5859 19768 5871 19771
rect 6270 19768 6276 19780
rect 5859 19740 6276 19768
rect 5859 19737 5871 19740
rect 5813 19731 5871 19737
rect 6270 19728 6276 19740
rect 6328 19728 6334 19780
rect 6380 19768 6408 19808
rect 6822 19796 6828 19808
rect 6880 19796 6886 19848
rect 7650 19768 7656 19780
rect 6380 19740 7656 19768
rect 7650 19728 7656 19740
rect 7708 19728 7714 19780
rect 9508 19768 9536 19944
rect 9677 19941 9689 19975
rect 9723 19972 9735 19975
rect 9876 19972 9904 20000
rect 9723 19944 9904 19972
rect 10511 19944 12020 19972
rect 9723 19941 9735 19944
rect 9677 19935 9735 19941
rect 9858 19904 9864 19916
rect 9819 19876 9864 19904
rect 9858 19864 9864 19876
rect 9916 19864 9922 19916
rect 10410 19836 10416 19848
rect 10323 19808 10416 19836
rect 10410 19796 10416 19808
rect 10468 19836 10474 19848
rect 10511 19836 10539 19944
rect 11992 19916 12020 19944
rect 12158 19932 12164 19984
rect 12216 19972 12222 19984
rect 15580 19972 15608 20012
rect 12216 19944 15608 19972
rect 15648 19975 15706 19981
rect 12216 19932 12222 19944
rect 15648 19941 15660 19975
rect 15694 19972 15706 19975
rect 16298 19972 16304 19984
rect 15694 19944 16304 19972
rect 15694 19941 15706 19944
rect 15648 19935 15706 19941
rect 16298 19932 16304 19944
rect 16356 19972 16362 19984
rect 17221 19975 17279 19981
rect 17221 19972 17233 19975
rect 16356 19944 17233 19972
rect 16356 19932 16362 19944
rect 17221 19941 17233 19944
rect 17267 19941 17279 19975
rect 17328 19972 17356 20012
rect 17402 20000 17408 20052
rect 17460 20040 17466 20052
rect 18782 20040 18788 20052
rect 17460 20012 18788 20040
rect 17460 20000 17466 20012
rect 18782 20000 18788 20012
rect 18840 20000 18846 20052
rect 19150 20040 19156 20052
rect 19111 20012 19156 20040
rect 19150 20000 19156 20012
rect 19208 20040 19214 20052
rect 19889 20043 19947 20049
rect 19889 20040 19901 20043
rect 19208 20012 19901 20040
rect 19208 20000 19214 20012
rect 19889 20009 19901 20012
rect 19935 20009 19947 20043
rect 19889 20003 19947 20009
rect 18690 19972 18696 19984
rect 17328 19944 18696 19972
rect 17221 19935 17279 19941
rect 18690 19932 18696 19944
rect 18748 19932 18754 19984
rect 19794 19972 19800 19984
rect 19755 19944 19800 19972
rect 19794 19932 19800 19944
rect 19852 19932 19858 19984
rect 10686 19913 10692 19916
rect 10680 19904 10692 19913
rect 10647 19876 10692 19904
rect 10680 19867 10692 19876
rect 10686 19864 10692 19867
rect 10744 19864 10750 19916
rect 11974 19864 11980 19916
rect 12032 19904 12038 19916
rect 12342 19913 12348 19916
rect 12069 19907 12127 19913
rect 12069 19904 12081 19907
rect 12032 19876 12081 19904
rect 12032 19864 12038 19876
rect 12069 19873 12081 19876
rect 12115 19873 12127 19907
rect 12336 19904 12348 19913
rect 12255 19876 12348 19904
rect 12069 19867 12127 19873
rect 12336 19867 12348 19876
rect 12400 19904 12406 19916
rect 13909 19907 13967 19913
rect 13909 19904 13921 19907
rect 12400 19876 13921 19904
rect 12342 19864 12348 19867
rect 12400 19864 12406 19876
rect 13909 19873 13921 19876
rect 13955 19873 13967 19907
rect 13909 19867 13967 19873
rect 15010 19864 15016 19916
rect 15068 19904 15074 19916
rect 17037 19907 17095 19913
rect 17037 19904 17049 19907
rect 15068 19876 17049 19904
rect 15068 19864 15074 19876
rect 17037 19873 17049 19876
rect 17083 19873 17095 19907
rect 17037 19867 17095 19873
rect 17773 19907 17831 19913
rect 17773 19873 17785 19907
rect 17819 19904 17831 19907
rect 17862 19904 17868 19916
rect 17819 19876 17868 19904
rect 17819 19873 17831 19876
rect 17773 19867 17831 19873
rect 17862 19864 17868 19876
rect 17920 19864 17926 19916
rect 18040 19907 18098 19913
rect 18040 19873 18052 19907
rect 18086 19904 18098 19907
rect 18874 19904 18880 19916
rect 18086 19876 18880 19904
rect 18086 19873 18098 19876
rect 18040 19867 18098 19873
rect 18874 19864 18880 19876
rect 18932 19864 18938 19916
rect 20806 19904 20812 19916
rect 18984 19876 20812 19904
rect 14182 19836 14188 19848
rect 10468 19808 10539 19836
rect 14095 19808 14188 19836
rect 10468 19796 10474 19808
rect 14182 19796 14188 19808
rect 14240 19796 14246 19848
rect 14645 19839 14703 19845
rect 14645 19805 14657 19839
rect 14691 19836 14703 19839
rect 14737 19839 14795 19845
rect 14737 19836 14749 19839
rect 14691 19808 14749 19836
rect 14691 19805 14703 19808
rect 14645 19799 14703 19805
rect 14737 19805 14749 19808
rect 14783 19836 14795 19839
rect 14826 19836 14832 19848
rect 14783 19808 14832 19836
rect 14783 19805 14795 19808
rect 14737 19799 14795 19805
rect 14826 19796 14832 19808
rect 14884 19796 14890 19848
rect 15286 19796 15292 19848
rect 15344 19836 15350 19848
rect 15381 19839 15439 19845
rect 15381 19836 15393 19839
rect 15344 19808 15393 19836
rect 15344 19796 15350 19808
rect 15381 19805 15393 19808
rect 15427 19805 15439 19839
rect 15381 19799 15439 19805
rect 18782 19796 18788 19848
rect 18840 19836 18846 19848
rect 18984 19836 19012 19876
rect 20806 19864 20812 19876
rect 20864 19864 20870 19916
rect 21634 19904 21640 19916
rect 21595 19876 21640 19904
rect 21634 19864 21640 19876
rect 21692 19864 21698 19916
rect 22002 19864 22008 19916
rect 22060 19904 22066 19916
rect 22281 19907 22339 19913
rect 22281 19904 22293 19907
rect 22060 19876 22293 19904
rect 22060 19864 22066 19876
rect 22281 19873 22293 19876
rect 22327 19873 22339 19907
rect 22462 19904 22468 19916
rect 22423 19876 22468 19904
rect 22281 19867 22339 19873
rect 22462 19864 22468 19876
rect 22520 19864 22526 19916
rect 18840 19808 19012 19836
rect 18840 19796 18846 19808
rect 19794 19796 19800 19848
rect 19852 19836 19858 19848
rect 20073 19839 20131 19845
rect 20073 19836 20085 19839
rect 19852 19808 20085 19836
rect 19852 19796 19858 19808
rect 20073 19805 20085 19808
rect 20119 19836 20131 19839
rect 20346 19836 20352 19848
rect 20119 19808 20352 19836
rect 20119 19805 20131 19808
rect 20073 19799 20131 19805
rect 20346 19796 20352 19808
rect 20404 19796 20410 19848
rect 21726 19836 21732 19848
rect 21687 19808 21732 19836
rect 21726 19796 21732 19808
rect 21784 19796 21790 19848
rect 21818 19796 21824 19848
rect 21876 19836 21882 19848
rect 21876 19808 21921 19836
rect 21876 19796 21882 19808
rect 12066 19768 12072 19780
rect 9508 19740 10456 19768
rect 2038 19660 2044 19712
rect 2096 19700 2102 19712
rect 2777 19703 2835 19709
rect 2777 19700 2789 19703
rect 2096 19672 2789 19700
rect 2096 19660 2102 19672
rect 2777 19669 2789 19672
rect 2823 19700 2835 19703
rect 5074 19700 5080 19712
rect 2823 19672 5080 19700
rect 2823 19669 2835 19672
rect 2777 19663 2835 19669
rect 5074 19660 5080 19672
rect 5132 19660 5138 19712
rect 5994 19660 6000 19712
rect 6052 19700 6058 19712
rect 6181 19703 6239 19709
rect 6181 19700 6193 19703
rect 6052 19672 6193 19700
rect 6052 19660 6058 19672
rect 6181 19669 6193 19672
rect 6227 19669 6239 19703
rect 7558 19700 7564 19712
rect 7519 19672 7564 19700
rect 6181 19663 6239 19669
rect 7558 19660 7564 19672
rect 7616 19660 7622 19712
rect 8294 19660 8300 19712
rect 8352 19700 8358 19712
rect 9309 19703 9367 19709
rect 9309 19700 9321 19703
rect 8352 19672 9321 19700
rect 8352 19660 8358 19672
rect 9309 19669 9321 19672
rect 9355 19669 9367 19703
rect 9309 19663 9367 19669
rect 9674 19660 9680 19712
rect 9732 19700 9738 19712
rect 10045 19703 10103 19709
rect 10045 19700 10057 19703
rect 9732 19672 10057 19700
rect 9732 19660 9738 19672
rect 10045 19669 10057 19672
rect 10091 19669 10103 19703
rect 10428 19700 10456 19740
rect 11808 19740 12072 19768
rect 11808 19700 11836 19740
rect 12066 19728 12072 19740
rect 12124 19728 12130 19780
rect 14200 19768 14228 19796
rect 14918 19768 14924 19780
rect 13004 19740 13768 19768
rect 14200 19740 14924 19768
rect 10428 19672 11836 19700
rect 10045 19663 10103 19669
rect 11882 19660 11888 19712
rect 11940 19700 11946 19712
rect 12434 19700 12440 19712
rect 11940 19672 12440 19700
rect 11940 19660 11946 19672
rect 12434 19660 12440 19672
rect 12492 19660 12498 19712
rect 12710 19660 12716 19712
rect 12768 19700 12774 19712
rect 13004 19700 13032 19740
rect 12768 19672 13032 19700
rect 12768 19660 12774 19672
rect 13538 19660 13544 19712
rect 13596 19700 13602 19712
rect 13740 19700 13768 19740
rect 14918 19728 14924 19740
rect 14976 19728 14982 19780
rect 17218 19768 17224 19780
rect 16316 19740 17224 19768
rect 16316 19700 16344 19740
rect 17218 19728 17224 19740
rect 17276 19728 17282 19780
rect 19886 19768 19892 19780
rect 18708 19740 19892 19768
rect 13596 19672 13641 19700
rect 13740 19672 16344 19700
rect 13596 19660 13602 19672
rect 16390 19660 16396 19712
rect 16448 19700 16454 19712
rect 16666 19700 16672 19712
rect 16448 19672 16672 19700
rect 16448 19660 16454 19672
rect 16666 19660 16672 19672
rect 16724 19700 16730 19712
rect 16761 19703 16819 19709
rect 16761 19700 16773 19703
rect 16724 19672 16773 19700
rect 16724 19660 16730 19672
rect 16761 19669 16773 19672
rect 16807 19669 16819 19703
rect 16761 19663 16819 19669
rect 17126 19660 17132 19712
rect 17184 19700 17190 19712
rect 17405 19703 17463 19709
rect 17405 19700 17417 19703
rect 17184 19672 17417 19700
rect 17184 19660 17190 19672
rect 17405 19669 17417 19672
rect 17451 19669 17463 19703
rect 17405 19663 17463 19669
rect 17954 19660 17960 19712
rect 18012 19700 18018 19712
rect 18708 19700 18736 19740
rect 19886 19728 19892 19740
rect 19944 19728 19950 19780
rect 18012 19672 18736 19700
rect 18012 19660 18018 19672
rect 19242 19660 19248 19712
rect 19300 19700 19306 19712
rect 19429 19703 19487 19709
rect 19429 19700 19441 19703
rect 19300 19672 19441 19700
rect 19300 19660 19306 19672
rect 19429 19669 19441 19672
rect 19475 19669 19487 19703
rect 19429 19663 19487 19669
rect 21269 19703 21327 19709
rect 21269 19669 21281 19703
rect 21315 19700 21327 19703
rect 21358 19700 21364 19712
rect 21315 19672 21364 19700
rect 21315 19669 21327 19672
rect 21269 19663 21327 19669
rect 21358 19660 21364 19672
rect 21416 19660 21422 19712
rect 22646 19700 22652 19712
rect 22607 19672 22652 19700
rect 22646 19660 22652 19672
rect 22704 19660 22710 19712
rect 1104 19610 23276 19632
rect 1104 19558 4680 19610
rect 4732 19558 4744 19610
rect 4796 19558 4808 19610
rect 4860 19558 4872 19610
rect 4924 19558 12078 19610
rect 12130 19558 12142 19610
rect 12194 19558 12206 19610
rect 12258 19558 12270 19610
rect 12322 19558 19475 19610
rect 19527 19558 19539 19610
rect 19591 19558 19603 19610
rect 19655 19558 19667 19610
rect 19719 19558 23276 19610
rect 1104 19536 23276 19558
rect 3418 19496 3424 19508
rect 3068 19468 3424 19496
rect 3068 19369 3096 19468
rect 3418 19456 3424 19468
rect 3476 19456 3482 19508
rect 3786 19456 3792 19508
rect 3844 19496 3850 19508
rect 4433 19499 4491 19505
rect 3844 19468 4016 19496
rect 3844 19456 3850 19468
rect 3988 19428 4016 19468
rect 4433 19465 4445 19499
rect 4479 19496 4491 19499
rect 4522 19496 4528 19508
rect 4479 19468 4528 19496
rect 4479 19465 4491 19468
rect 4433 19459 4491 19465
rect 4522 19456 4528 19468
rect 4580 19456 4586 19508
rect 5350 19456 5356 19508
rect 5408 19456 5414 19508
rect 5442 19456 5448 19508
rect 5500 19496 5506 19508
rect 5500 19468 9996 19496
rect 5500 19456 5506 19468
rect 5368 19428 5396 19456
rect 3988 19400 5396 19428
rect 7834 19388 7840 19440
rect 7892 19428 7898 19440
rect 7892 19400 8340 19428
rect 7892 19388 7898 19400
rect 3053 19363 3111 19369
rect 3053 19329 3065 19363
rect 3099 19329 3111 19363
rect 5353 19363 5411 19369
rect 3053 19323 3111 19329
rect 4908 19332 5212 19360
rect 1394 19292 1400 19304
rect 1307 19264 1400 19292
rect 1394 19252 1400 19264
rect 1452 19292 1458 19304
rect 3326 19301 3332 19304
rect 1452 19264 2360 19292
rect 1452 19252 1458 19264
rect 2332 19236 2360 19264
rect 3320 19255 3332 19301
rect 3384 19292 3390 19304
rect 3384 19264 3420 19292
rect 3326 19252 3332 19255
rect 3384 19252 3390 19264
rect 3694 19252 3700 19304
rect 3752 19292 3758 19304
rect 4908 19292 4936 19332
rect 5074 19292 5080 19304
rect 3752 19264 4936 19292
rect 5035 19264 5080 19292
rect 3752 19252 3758 19264
rect 5074 19252 5080 19264
rect 5132 19252 5138 19304
rect 5184 19292 5212 19332
rect 5353 19329 5365 19363
rect 5399 19360 5411 19363
rect 5534 19360 5540 19372
rect 5399 19332 5540 19360
rect 5399 19329 5411 19332
rect 5353 19323 5411 19329
rect 5534 19320 5540 19332
rect 5592 19360 5598 19372
rect 6273 19363 6331 19369
rect 6273 19360 6285 19363
rect 5592 19332 6285 19360
rect 5592 19320 5598 19332
rect 6273 19329 6285 19332
rect 6319 19360 6331 19363
rect 6454 19360 6460 19372
rect 6319 19332 6460 19360
rect 6319 19329 6331 19332
rect 6273 19323 6331 19329
rect 6454 19320 6460 19332
rect 6512 19360 6518 19372
rect 8113 19363 8171 19369
rect 8113 19360 8125 19363
rect 6512 19332 8125 19360
rect 6512 19320 6518 19332
rect 8113 19329 8125 19332
rect 8159 19329 8171 19363
rect 8312 19360 8340 19400
rect 9968 19360 9996 19468
rect 10134 19456 10140 19508
rect 10192 19496 10198 19508
rect 12526 19496 12532 19508
rect 10192 19468 12532 19496
rect 10192 19456 10198 19468
rect 12526 19456 12532 19468
rect 12584 19456 12590 19508
rect 14182 19496 14188 19508
rect 12636 19468 14188 19496
rect 10873 19363 10931 19369
rect 10873 19360 10885 19363
rect 8312 19332 8708 19360
rect 9968 19332 10885 19360
rect 8113 19323 8171 19329
rect 6181 19295 6239 19301
rect 6181 19292 6193 19295
rect 5184 19264 6193 19292
rect 6181 19261 6193 19264
rect 6227 19261 6239 19295
rect 6181 19255 6239 19261
rect 7009 19295 7067 19301
rect 7009 19261 7021 19295
rect 7055 19261 7067 19295
rect 7009 19255 7067 19261
rect 7929 19295 7987 19301
rect 7929 19261 7941 19295
rect 7975 19292 7987 19295
rect 8294 19292 8300 19304
rect 7975 19264 8300 19292
rect 7975 19261 7987 19264
rect 7929 19255 7987 19261
rect 1670 19233 1676 19236
rect 1664 19224 1676 19233
rect 1631 19196 1676 19224
rect 1664 19187 1676 19196
rect 1670 19184 1676 19187
rect 1728 19184 1734 19236
rect 2314 19184 2320 19236
rect 2372 19184 2378 19236
rect 2958 19184 2964 19236
rect 3016 19224 3022 19236
rect 5169 19227 5227 19233
rect 5169 19224 5181 19227
rect 3016 19196 5181 19224
rect 3016 19184 3022 19196
rect 5169 19193 5181 19196
rect 5215 19193 5227 19227
rect 5169 19187 5227 19193
rect 5258 19184 5264 19236
rect 5316 19224 5322 19236
rect 6089 19227 6147 19233
rect 6089 19224 6101 19227
rect 5316 19196 6101 19224
rect 5316 19184 5322 19196
rect 6089 19193 6101 19196
rect 6135 19193 6147 19227
rect 7024 19224 7052 19255
rect 8294 19252 8300 19264
rect 8352 19252 8358 19304
rect 8573 19295 8631 19301
rect 8573 19261 8585 19295
rect 8619 19261 8631 19295
rect 8680 19292 8708 19332
rect 10873 19329 10885 19332
rect 10919 19360 10931 19363
rect 11885 19363 11943 19369
rect 11885 19360 11897 19363
rect 10919 19332 11897 19360
rect 10919 19329 10931 19332
rect 10873 19323 10931 19329
rect 11885 19329 11897 19332
rect 11931 19360 11943 19363
rect 12636 19360 12664 19468
rect 14182 19456 14188 19468
rect 14240 19456 14246 19508
rect 14277 19499 14335 19505
rect 14277 19465 14289 19499
rect 14323 19496 14335 19499
rect 15470 19496 15476 19508
rect 14323 19468 15476 19496
rect 14323 19465 14335 19468
rect 14277 19459 14335 19465
rect 15470 19456 15476 19468
rect 15528 19456 15534 19508
rect 19334 19496 19340 19508
rect 15764 19468 15976 19496
rect 13909 19431 13967 19437
rect 11931 19332 12664 19360
rect 12728 19400 13860 19428
rect 11931 19329 11943 19332
rect 11885 19323 11943 19329
rect 10042 19292 10048 19304
rect 8680 19264 10048 19292
rect 8573 19255 8631 19261
rect 8478 19224 8484 19236
rect 7024 19196 8484 19224
rect 6089 19187 6147 19193
rect 8478 19184 8484 19196
rect 8536 19184 8542 19236
rect 8588 19224 8616 19255
rect 10042 19252 10048 19264
rect 10100 19252 10106 19304
rect 12728 19292 12756 19400
rect 13078 19360 13084 19372
rect 13039 19332 13084 19360
rect 13078 19320 13084 19332
rect 13136 19320 13142 19372
rect 10336 19264 12756 19292
rect 12805 19295 12863 19301
rect 8662 19224 8668 19236
rect 8588 19196 8668 19224
rect 8662 19184 8668 19196
rect 8720 19184 8726 19236
rect 8754 19184 8760 19236
rect 8812 19233 8818 19236
rect 8812 19227 8876 19233
rect 8812 19193 8830 19227
rect 8864 19193 8876 19227
rect 8812 19187 8876 19193
rect 8812 19184 8818 19187
rect 9766 19184 9772 19236
rect 9824 19224 9830 19236
rect 10226 19224 10232 19236
rect 9824 19196 10232 19224
rect 9824 19184 9830 19196
rect 10226 19184 10232 19196
rect 10284 19184 10290 19236
rect 2774 19156 2780 19168
rect 2735 19128 2780 19156
rect 2774 19116 2780 19128
rect 2832 19116 2838 19168
rect 3234 19116 3240 19168
rect 3292 19156 3298 19168
rect 4154 19156 4160 19168
rect 3292 19128 4160 19156
rect 3292 19116 3298 19128
rect 4154 19116 4160 19128
rect 4212 19116 4218 19168
rect 4706 19156 4712 19168
rect 4667 19128 4712 19156
rect 4706 19116 4712 19128
rect 4764 19116 4770 19168
rect 5718 19156 5724 19168
rect 5679 19128 5724 19156
rect 5718 19116 5724 19128
rect 5776 19116 5782 19168
rect 6822 19116 6828 19168
rect 6880 19156 6886 19168
rect 7193 19159 7251 19165
rect 7193 19156 7205 19159
rect 6880 19128 7205 19156
rect 6880 19116 6886 19128
rect 7193 19125 7205 19128
rect 7239 19125 7251 19159
rect 7193 19119 7251 19125
rect 7561 19159 7619 19165
rect 7561 19125 7573 19159
rect 7607 19156 7619 19159
rect 7834 19156 7840 19168
rect 7607 19128 7840 19156
rect 7607 19125 7619 19128
rect 7561 19119 7619 19125
rect 7834 19116 7840 19128
rect 7892 19116 7898 19168
rect 8021 19159 8079 19165
rect 8021 19125 8033 19159
rect 8067 19156 8079 19159
rect 8110 19156 8116 19168
rect 8067 19128 8116 19156
rect 8067 19125 8079 19128
rect 8021 19119 8079 19125
rect 8110 19116 8116 19128
rect 8168 19156 8174 19168
rect 10336 19165 10364 19264
rect 12805 19261 12817 19295
rect 12851 19292 12863 19295
rect 13538 19292 13544 19304
rect 12851 19264 13544 19292
rect 12851 19261 12863 19264
rect 12805 19255 12863 19261
rect 13538 19252 13544 19264
rect 13596 19252 13602 19304
rect 13630 19252 13636 19304
rect 13688 19292 13694 19304
rect 13725 19295 13783 19301
rect 13725 19292 13737 19295
rect 13688 19264 13737 19292
rect 13688 19252 13694 19264
rect 13725 19261 13737 19264
rect 13771 19261 13783 19295
rect 13832 19292 13860 19400
rect 13909 19397 13921 19431
rect 13955 19428 13967 19431
rect 15764 19428 15792 19468
rect 13955 19400 15792 19428
rect 15948 19428 15976 19468
rect 17420 19468 19340 19496
rect 17420 19428 17448 19468
rect 19334 19456 19340 19468
rect 19392 19456 19398 19508
rect 19426 19428 19432 19440
rect 15948 19400 17448 19428
rect 19387 19400 19432 19428
rect 13955 19397 13967 19400
rect 13909 19391 13967 19397
rect 19426 19388 19432 19400
rect 19484 19388 19490 19440
rect 14642 19320 14648 19372
rect 14700 19360 14706 19372
rect 14737 19363 14795 19369
rect 14737 19360 14749 19363
rect 14700 19332 14749 19360
rect 14700 19320 14706 19332
rect 14737 19329 14749 19332
rect 14783 19329 14795 19363
rect 14918 19360 14924 19372
rect 14879 19332 14924 19360
rect 14737 19323 14795 19329
rect 14918 19320 14924 19332
rect 14976 19320 14982 19372
rect 15841 19363 15899 19369
rect 15841 19329 15853 19363
rect 15887 19329 15899 19363
rect 15841 19323 15899 19329
rect 15657 19295 15715 19301
rect 15657 19292 15669 19295
rect 13832 19264 15669 19292
rect 13725 19255 13783 19261
rect 15657 19261 15669 19264
rect 15703 19261 15715 19295
rect 15856 19292 15884 19323
rect 15930 19320 15936 19372
rect 15988 19360 15994 19372
rect 16574 19360 16580 19372
rect 15988 19332 16580 19360
rect 15988 19320 15994 19332
rect 16574 19320 16580 19332
rect 16632 19360 16638 19372
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 16632 19332 16865 19360
rect 16632 19320 16638 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 19886 19320 19892 19372
rect 19944 19360 19950 19372
rect 20257 19363 20315 19369
rect 20257 19360 20269 19363
rect 19944 19332 20269 19360
rect 19944 19320 19950 19332
rect 20257 19329 20269 19332
rect 20303 19329 20315 19363
rect 20257 19323 20315 19329
rect 16114 19292 16120 19304
rect 15856 19264 16120 19292
rect 15657 19255 15715 19261
rect 16114 19252 16120 19264
rect 16172 19252 16178 19304
rect 16666 19292 16672 19304
rect 16627 19264 16672 19292
rect 16666 19252 16672 19264
rect 16724 19252 16730 19304
rect 17402 19292 17408 19304
rect 17363 19264 17408 19292
rect 17402 19252 17408 19264
rect 17460 19252 17466 19304
rect 18046 19292 18052 19304
rect 18007 19264 18052 19292
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 18690 19252 18696 19304
rect 18748 19292 18754 19304
rect 20165 19295 20223 19301
rect 20165 19292 20177 19295
rect 18748 19264 20177 19292
rect 18748 19252 18754 19264
rect 20165 19261 20177 19264
rect 20211 19261 20223 19295
rect 20165 19255 20223 19261
rect 20898 19252 20904 19304
rect 20956 19292 20962 19304
rect 20993 19295 21051 19301
rect 20993 19292 21005 19295
rect 20956 19264 21005 19292
rect 20956 19252 20962 19264
rect 20993 19261 21005 19264
rect 21039 19261 21051 19295
rect 20993 19255 21051 19261
rect 21260 19295 21318 19301
rect 21260 19261 21272 19295
rect 21306 19292 21318 19295
rect 21726 19292 21732 19304
rect 21306 19264 21732 19292
rect 21306 19261 21318 19264
rect 21260 19255 21318 19261
rect 12894 19224 12900 19236
rect 11348 19196 12756 19224
rect 12855 19196 12900 19224
rect 9953 19159 10011 19165
rect 9953 19156 9965 19159
rect 8168 19128 9965 19156
rect 8168 19116 8174 19128
rect 9953 19125 9965 19128
rect 9999 19125 10011 19159
rect 9953 19119 10011 19125
rect 10321 19159 10379 19165
rect 10321 19125 10333 19159
rect 10367 19125 10379 19159
rect 10686 19156 10692 19168
rect 10647 19128 10692 19156
rect 10321 19119 10379 19125
rect 10686 19116 10692 19128
rect 10744 19116 10750 19168
rect 10778 19116 10784 19168
rect 10836 19156 10842 19168
rect 11348 19165 11376 19196
rect 11333 19159 11391 19165
rect 10836 19128 10881 19156
rect 10836 19116 10842 19128
rect 11333 19125 11345 19159
rect 11379 19125 11391 19159
rect 11698 19156 11704 19168
rect 11659 19128 11704 19156
rect 11333 19119 11391 19125
rect 11698 19116 11704 19128
rect 11756 19116 11762 19168
rect 11790 19116 11796 19168
rect 11848 19156 11854 19168
rect 11848 19128 11893 19156
rect 11848 19116 11854 19128
rect 12342 19116 12348 19168
rect 12400 19156 12406 19168
rect 12437 19159 12495 19165
rect 12437 19156 12449 19159
rect 12400 19128 12449 19156
rect 12400 19116 12406 19128
rect 12437 19125 12449 19128
rect 12483 19125 12495 19159
rect 12728 19156 12756 19196
rect 12894 19184 12900 19196
rect 12952 19184 12958 19236
rect 15749 19227 15807 19233
rect 15749 19224 15761 19227
rect 13004 19196 15761 19224
rect 13004 19156 13032 19196
rect 15749 19193 15761 19196
rect 15795 19193 15807 19227
rect 15749 19187 15807 19193
rect 18316 19227 18374 19233
rect 18316 19193 18328 19227
rect 18362 19224 18374 19227
rect 19242 19224 19248 19236
rect 18362 19196 19248 19224
rect 18362 19193 18374 19196
rect 18316 19187 18374 19193
rect 19242 19184 19248 19196
rect 19300 19184 19306 19236
rect 20073 19227 20131 19233
rect 20073 19224 20085 19227
rect 19352 19196 20085 19224
rect 12728 19128 13032 19156
rect 14645 19159 14703 19165
rect 12437 19119 12495 19125
rect 14645 19125 14657 19159
rect 14691 19156 14703 19159
rect 15194 19156 15200 19168
rect 14691 19128 15200 19156
rect 14691 19125 14703 19128
rect 14645 19119 14703 19125
rect 15194 19116 15200 19128
rect 15252 19116 15258 19168
rect 15286 19116 15292 19168
rect 15344 19156 15350 19168
rect 16298 19156 16304 19168
rect 15344 19128 15389 19156
rect 16259 19128 16304 19156
rect 15344 19116 15350 19128
rect 16298 19116 16304 19128
rect 16356 19116 16362 19168
rect 16758 19156 16764 19168
rect 16719 19128 16764 19156
rect 16758 19116 16764 19128
rect 16816 19116 16822 19168
rect 17310 19116 17316 19168
rect 17368 19156 17374 19168
rect 17589 19159 17647 19165
rect 17589 19156 17601 19159
rect 17368 19128 17601 19156
rect 17368 19116 17374 19128
rect 17589 19125 17601 19128
rect 17635 19125 17647 19159
rect 17589 19119 17647 19125
rect 17954 19116 17960 19168
rect 18012 19156 18018 19168
rect 19352 19156 19380 19196
rect 20073 19193 20085 19196
rect 20119 19193 20131 19227
rect 20073 19187 20131 19193
rect 18012 19128 19380 19156
rect 19705 19159 19763 19165
rect 18012 19116 18018 19128
rect 19705 19125 19717 19159
rect 19751 19156 19763 19159
rect 20254 19156 20260 19168
rect 19751 19128 20260 19156
rect 19751 19125 19763 19128
rect 19705 19119 19763 19125
rect 20254 19116 20260 19128
rect 20312 19116 20318 19168
rect 21008 19156 21036 19255
rect 21726 19252 21732 19264
rect 21784 19252 21790 19304
rect 21266 19156 21272 19168
rect 21008 19128 21272 19156
rect 21266 19116 21272 19128
rect 21324 19116 21330 19168
rect 21634 19116 21640 19168
rect 21692 19156 21698 19168
rect 22373 19159 22431 19165
rect 22373 19156 22385 19159
rect 21692 19128 22385 19156
rect 21692 19116 21698 19128
rect 22373 19125 22385 19128
rect 22419 19125 22431 19159
rect 22373 19119 22431 19125
rect 1104 19066 23276 19088
rect 1104 19014 8379 19066
rect 8431 19014 8443 19066
rect 8495 19014 8507 19066
rect 8559 19014 8571 19066
rect 8623 19014 15776 19066
rect 15828 19014 15840 19066
rect 15892 19014 15904 19066
rect 15956 19014 15968 19066
rect 16020 19014 23276 19066
rect 1104 18992 23276 19014
rect 1670 18912 1676 18964
rect 1728 18952 1734 18964
rect 3789 18955 3847 18961
rect 3789 18952 3801 18955
rect 1728 18924 3801 18952
rect 1728 18912 1734 18924
rect 3789 18921 3801 18924
rect 3835 18921 3847 18955
rect 3789 18915 3847 18921
rect 4065 18955 4123 18961
rect 4065 18921 4077 18955
rect 4111 18921 4123 18955
rect 4065 18915 4123 18921
rect 4433 18955 4491 18961
rect 4433 18921 4445 18955
rect 4479 18952 4491 18955
rect 4706 18952 4712 18964
rect 4479 18924 4712 18952
rect 4479 18921 4491 18924
rect 4433 18915 4491 18921
rect 4080 18884 4108 18915
rect 4706 18912 4712 18924
rect 4764 18912 4770 18964
rect 4798 18912 4804 18964
rect 4856 18952 4862 18964
rect 6822 18952 6828 18964
rect 4856 18924 6828 18952
rect 4856 18912 4862 18924
rect 6822 18912 6828 18924
rect 6880 18912 6886 18964
rect 9309 18955 9367 18961
rect 9309 18921 9321 18955
rect 9355 18952 9367 18955
rect 9858 18952 9864 18964
rect 9355 18924 9864 18952
rect 9355 18921 9367 18924
rect 9309 18915 9367 18921
rect 9858 18912 9864 18924
rect 9916 18912 9922 18964
rect 10686 18912 10692 18964
rect 10744 18952 10750 18964
rect 11609 18955 11667 18961
rect 11609 18952 11621 18955
rect 10744 18924 11621 18952
rect 10744 18912 10750 18924
rect 11609 18921 11621 18924
rect 11655 18921 11667 18955
rect 12526 18952 12532 18964
rect 11609 18915 11667 18921
rect 11716 18924 12532 18952
rect 1780 18856 4108 18884
rect 4525 18887 4583 18893
rect 1780 18825 1808 18856
rect 4525 18853 4537 18887
rect 4571 18884 4583 18887
rect 5718 18884 5724 18896
rect 4571 18856 5724 18884
rect 4571 18853 4583 18856
rect 4525 18847 4583 18853
rect 5718 18844 5724 18856
rect 5776 18844 5782 18896
rect 7926 18884 7932 18896
rect 6288 18856 7932 18884
rect 1765 18819 1823 18825
rect 1765 18785 1777 18819
rect 1811 18785 1823 18819
rect 1765 18779 1823 18785
rect 2584 18819 2642 18825
rect 2584 18785 2596 18819
rect 2630 18816 2642 18819
rect 3694 18816 3700 18828
rect 2630 18788 3700 18816
rect 2630 18785 2642 18788
rect 2584 18779 2642 18785
rect 3694 18776 3700 18788
rect 3752 18776 3758 18828
rect 4154 18776 4160 18828
rect 4212 18816 4218 18828
rect 6288 18825 6316 18856
rect 7926 18844 7932 18856
rect 7984 18844 7990 18896
rect 8202 18893 8208 18896
rect 8196 18884 8208 18893
rect 8163 18856 8208 18884
rect 8196 18847 8208 18856
rect 8202 18844 8208 18847
rect 8260 18844 8266 18896
rect 8294 18844 8300 18896
rect 8352 18884 8358 18896
rect 11716 18884 11744 18924
rect 12526 18912 12532 18924
rect 12584 18912 12590 18964
rect 16114 18912 16120 18964
rect 16172 18952 16178 18964
rect 16761 18955 16819 18961
rect 16761 18952 16773 18955
rect 16172 18924 16773 18952
rect 16172 18912 16178 18924
rect 16761 18921 16773 18924
rect 16807 18921 16819 18955
rect 16761 18915 16819 18921
rect 16850 18912 16856 18964
rect 16908 18952 16914 18964
rect 17037 18955 17095 18961
rect 17037 18952 17049 18955
rect 16908 18924 17049 18952
rect 16908 18912 16914 18924
rect 17037 18921 17049 18924
rect 17083 18921 17095 18955
rect 18874 18952 18880 18964
rect 18835 18924 18880 18952
rect 17037 18915 17095 18921
rect 18874 18912 18880 18924
rect 18932 18952 18938 18964
rect 19521 18955 19579 18961
rect 19521 18952 19533 18955
rect 18932 18924 19533 18952
rect 18932 18912 18938 18924
rect 19521 18921 19533 18924
rect 19567 18921 19579 18955
rect 19521 18915 19579 18921
rect 22462 18912 22468 18964
rect 22520 18952 22526 18964
rect 22649 18955 22707 18961
rect 22649 18952 22661 18955
rect 22520 18924 22661 18952
rect 22520 18912 22526 18924
rect 22649 18921 22661 18924
rect 22695 18921 22707 18955
rect 22649 18915 22707 18921
rect 14001 18887 14059 18893
rect 14001 18884 14013 18887
rect 8352 18856 11744 18884
rect 12167 18856 14013 18884
rect 8352 18844 8358 18856
rect 12167 18828 12195 18856
rect 14001 18853 14013 18856
rect 14047 18853 14059 18887
rect 14001 18847 14059 18853
rect 15648 18887 15706 18893
rect 15648 18853 15660 18887
rect 15694 18884 15706 18887
rect 16206 18884 16212 18896
rect 15694 18856 16212 18884
rect 15694 18853 15706 18856
rect 15648 18847 15706 18853
rect 16206 18844 16212 18856
rect 16264 18844 16270 18896
rect 17764 18887 17822 18893
rect 17764 18853 17776 18887
rect 17810 18884 17822 18887
rect 19426 18884 19432 18896
rect 17810 18856 19432 18884
rect 17810 18853 17822 18856
rect 17764 18847 17822 18853
rect 19426 18844 19432 18856
rect 19484 18884 19490 18896
rect 19613 18887 19671 18893
rect 19613 18884 19625 18887
rect 19484 18856 19625 18884
rect 19484 18844 19490 18856
rect 19613 18853 19625 18856
rect 19659 18853 19671 18887
rect 19613 18847 19671 18853
rect 21536 18887 21594 18893
rect 21536 18853 21548 18887
rect 21582 18884 21594 18887
rect 21634 18884 21640 18896
rect 21582 18856 21640 18884
rect 21582 18853 21594 18856
rect 21536 18847 21594 18853
rect 21634 18844 21640 18856
rect 21692 18844 21698 18896
rect 5445 18819 5503 18825
rect 5445 18816 5457 18819
rect 4212 18788 5457 18816
rect 4212 18776 4218 18788
rect 5445 18785 5457 18788
rect 5491 18785 5503 18819
rect 5445 18779 5503 18785
rect 6273 18819 6331 18825
rect 6273 18785 6285 18819
rect 6319 18785 6331 18819
rect 6273 18779 6331 18785
rect 7193 18819 7251 18825
rect 7193 18785 7205 18819
rect 7239 18816 7251 18819
rect 9490 18816 9496 18828
rect 7239 18788 9496 18816
rect 7239 18785 7251 18788
rect 7193 18779 7251 18785
rect 9490 18776 9496 18788
rect 9548 18776 9554 18828
rect 9674 18816 9680 18828
rect 9635 18788 9680 18816
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 10496 18819 10554 18825
rect 10496 18785 10508 18819
rect 10542 18816 10554 18819
rect 10778 18816 10784 18828
rect 10542 18788 10784 18816
rect 10542 18785 10554 18788
rect 10496 18779 10554 18785
rect 10778 18776 10784 18788
rect 10836 18816 10842 18828
rect 11606 18816 11612 18828
rect 10836 18788 11612 18816
rect 10836 18776 10842 18788
rect 11606 18776 11612 18788
rect 11664 18776 11670 18828
rect 11885 18819 11943 18825
rect 11885 18785 11897 18819
rect 11931 18816 11943 18819
rect 11974 18816 11980 18828
rect 11931 18788 11980 18816
rect 11931 18785 11943 18788
rect 11885 18779 11943 18785
rect 11974 18776 11980 18788
rect 12032 18776 12038 18828
rect 12158 18825 12164 18828
rect 12152 18779 12164 18825
rect 12216 18816 12222 18828
rect 12216 18788 12300 18816
rect 12158 18776 12164 18779
rect 12216 18776 12222 18788
rect 12618 18776 12624 18828
rect 12676 18816 12682 18828
rect 12676 18788 12940 18816
rect 12676 18776 12682 18788
rect 2314 18748 2320 18760
rect 2275 18720 2320 18748
rect 2314 18708 2320 18720
rect 2372 18708 2378 18760
rect 4614 18748 4620 18760
rect 4575 18720 4620 18748
rect 4614 18708 4620 18720
rect 4672 18708 4678 18760
rect 5537 18751 5595 18757
rect 5537 18748 5549 18751
rect 4724 18720 5549 18748
rect 4724 18680 4752 18720
rect 5537 18717 5549 18720
rect 5583 18717 5595 18751
rect 5537 18711 5595 18717
rect 5721 18751 5779 18757
rect 5721 18717 5733 18751
rect 5767 18717 5779 18751
rect 7282 18748 7288 18760
rect 7243 18720 7288 18748
rect 5721 18711 5779 18717
rect 5258 18680 5264 18692
rect 3620 18652 4752 18680
rect 4816 18652 5264 18680
rect 1949 18615 2007 18621
rect 1949 18581 1961 18615
rect 1995 18612 2007 18615
rect 3620 18612 3648 18652
rect 1995 18584 3648 18612
rect 3697 18615 3755 18621
rect 1995 18581 2007 18584
rect 1949 18575 2007 18581
rect 3697 18581 3709 18615
rect 3743 18612 3755 18615
rect 3789 18615 3847 18621
rect 3789 18612 3801 18615
rect 3743 18584 3801 18612
rect 3743 18581 3755 18584
rect 3697 18575 3755 18581
rect 3789 18581 3801 18584
rect 3835 18612 3847 18615
rect 4816 18612 4844 18652
rect 5258 18640 5264 18652
rect 5316 18640 5322 18692
rect 5736 18680 5764 18711
rect 7282 18708 7288 18720
rect 7340 18708 7346 18760
rect 7469 18751 7527 18757
rect 7469 18717 7481 18751
rect 7515 18748 7527 18751
rect 7558 18748 7564 18760
rect 7515 18720 7564 18748
rect 7515 18717 7527 18720
rect 7469 18711 7527 18717
rect 7484 18680 7512 18711
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 7926 18748 7932 18760
rect 7887 18720 7932 18748
rect 7926 18708 7932 18720
rect 7984 18708 7990 18760
rect 9766 18708 9772 18760
rect 9824 18748 9830 18760
rect 10229 18751 10287 18757
rect 10229 18748 10241 18751
rect 9824 18720 10241 18748
rect 9824 18708 9830 18720
rect 10229 18717 10241 18720
rect 10275 18717 10287 18751
rect 10229 18711 10287 18717
rect 12912 18680 12940 18788
rect 13262 18776 13268 18828
rect 13320 18816 13326 18828
rect 13909 18819 13967 18825
rect 13909 18816 13921 18819
rect 13320 18788 13921 18816
rect 13320 18776 13326 18788
rect 13909 18785 13921 18788
rect 13955 18785 13967 18819
rect 13909 18779 13967 18785
rect 14645 18819 14703 18825
rect 14645 18785 14657 18819
rect 14691 18816 14703 18819
rect 15102 18816 15108 18828
rect 14691 18788 15108 18816
rect 14691 18785 14703 18788
rect 14645 18779 14703 18785
rect 15102 18776 15108 18788
rect 15160 18776 15166 18828
rect 15194 18776 15200 18828
rect 15252 18816 15258 18828
rect 15378 18816 15384 18828
rect 15252 18788 15384 18816
rect 15252 18776 15258 18788
rect 15378 18776 15384 18788
rect 15436 18776 15442 18828
rect 15470 18776 15476 18828
rect 15528 18816 15534 18828
rect 20165 18819 20223 18825
rect 20165 18816 20177 18819
rect 15528 18788 20177 18816
rect 15528 18776 15534 18788
rect 20165 18785 20177 18788
rect 20211 18785 20223 18819
rect 22094 18816 22100 18828
rect 20165 18779 20223 18785
rect 20272 18788 22100 18816
rect 14185 18751 14243 18757
rect 14185 18717 14197 18751
rect 14231 18748 14243 18751
rect 14918 18748 14924 18760
rect 14231 18720 14924 18748
rect 14231 18717 14243 18720
rect 14185 18711 14243 18717
rect 14918 18708 14924 18720
rect 14976 18708 14982 18760
rect 17494 18748 17500 18760
rect 17455 18720 17500 18748
rect 17494 18708 17500 18720
rect 17552 18708 17558 18760
rect 19794 18748 19800 18760
rect 19755 18720 19800 18748
rect 19794 18708 19800 18720
rect 19852 18708 19858 18760
rect 14829 18683 14887 18689
rect 5736 18652 7512 18680
rect 8864 18652 10180 18680
rect 12912 18652 13676 18680
rect 5074 18612 5080 18624
rect 3835 18584 4844 18612
rect 5035 18584 5080 18612
rect 3835 18581 3847 18584
rect 3789 18575 3847 18581
rect 5074 18572 5080 18584
rect 5132 18572 5138 18624
rect 6454 18612 6460 18624
rect 6415 18584 6460 18612
rect 6454 18572 6460 18584
rect 6512 18572 6518 18624
rect 6822 18612 6828 18624
rect 6783 18584 6828 18612
rect 6822 18572 6828 18584
rect 6880 18572 6886 18624
rect 7558 18572 7564 18624
rect 7616 18612 7622 18624
rect 8864 18612 8892 18652
rect 7616 18584 8892 18612
rect 9861 18615 9919 18621
rect 7616 18572 7622 18584
rect 9861 18581 9873 18615
rect 9907 18612 9919 18615
rect 10042 18612 10048 18624
rect 9907 18584 10048 18612
rect 9907 18581 9919 18584
rect 9861 18575 9919 18581
rect 10042 18572 10048 18584
rect 10100 18572 10106 18624
rect 10152 18612 10180 18652
rect 13078 18612 13084 18624
rect 10152 18584 13084 18612
rect 13078 18572 13084 18584
rect 13136 18572 13142 18624
rect 13262 18612 13268 18624
rect 13223 18584 13268 18612
rect 13262 18572 13268 18584
rect 13320 18572 13326 18624
rect 13538 18612 13544 18624
rect 13499 18584 13544 18612
rect 13538 18572 13544 18584
rect 13596 18572 13602 18624
rect 13648 18612 13676 18652
rect 14829 18649 14841 18683
rect 14875 18680 14887 18683
rect 15010 18680 15016 18692
rect 14875 18652 15016 18680
rect 14875 18649 14887 18652
rect 14829 18643 14887 18649
rect 15010 18640 15016 18652
rect 15068 18640 15074 18692
rect 20272 18680 20300 18788
rect 22094 18776 22100 18788
rect 22152 18776 22158 18828
rect 21266 18748 21272 18760
rect 21227 18720 21272 18748
rect 21266 18708 21272 18720
rect 21324 18708 21330 18760
rect 18432 18652 20300 18680
rect 18432 18612 18460 18652
rect 13648 18584 18460 18612
rect 18506 18572 18512 18624
rect 18564 18612 18570 18624
rect 19153 18615 19211 18621
rect 19153 18612 19165 18615
rect 18564 18584 19165 18612
rect 18564 18572 18570 18584
rect 19153 18581 19165 18584
rect 19199 18581 19211 18615
rect 20346 18612 20352 18624
rect 20307 18584 20352 18612
rect 19153 18575 19211 18581
rect 20346 18572 20352 18584
rect 20404 18572 20410 18624
rect 1104 18522 23276 18544
rect 1104 18470 4680 18522
rect 4732 18470 4744 18522
rect 4796 18470 4808 18522
rect 4860 18470 4872 18522
rect 4924 18470 12078 18522
rect 12130 18470 12142 18522
rect 12194 18470 12206 18522
rect 12258 18470 12270 18522
rect 12322 18470 19475 18522
rect 19527 18470 19539 18522
rect 19591 18470 19603 18522
rect 19655 18470 19667 18522
rect 19719 18470 23276 18522
rect 1104 18448 23276 18470
rect 1949 18411 2007 18417
rect 1949 18377 1961 18411
rect 1995 18408 2007 18411
rect 4154 18408 4160 18420
rect 1995 18380 4016 18408
rect 4115 18380 4160 18408
rect 1995 18377 2007 18380
rect 1949 18371 2007 18377
rect 3694 18340 3700 18352
rect 3655 18312 3700 18340
rect 3694 18300 3700 18312
rect 3752 18300 3758 18352
rect 3988 18340 4016 18380
rect 4154 18368 4160 18380
rect 4212 18368 4218 18420
rect 9582 18408 9588 18420
rect 4543 18380 9588 18408
rect 4543 18340 4571 18380
rect 9582 18368 9588 18380
rect 9640 18368 9646 18420
rect 9766 18368 9772 18420
rect 9824 18408 9830 18420
rect 9953 18411 10011 18417
rect 9953 18408 9965 18411
rect 9824 18380 9965 18408
rect 9824 18368 9830 18380
rect 9953 18377 9965 18380
rect 9999 18377 10011 18411
rect 11606 18408 11612 18420
rect 11567 18380 11612 18408
rect 9953 18371 10011 18377
rect 11606 18368 11612 18380
rect 11664 18368 11670 18420
rect 14369 18411 14427 18417
rect 14369 18408 14381 18411
rect 13004 18380 14381 18408
rect 3988 18312 4571 18340
rect 7190 18300 7196 18352
rect 7248 18340 7254 18352
rect 7285 18343 7343 18349
rect 7285 18340 7297 18343
rect 7248 18312 7297 18340
rect 7248 18300 7254 18312
rect 7285 18309 7297 18312
rect 7331 18309 7343 18343
rect 8294 18340 8300 18352
rect 7285 18303 7343 18309
rect 7760 18312 8300 18340
rect 3418 18232 3424 18284
rect 3476 18272 3482 18284
rect 4525 18275 4583 18281
rect 4525 18272 4537 18275
rect 3476 18244 4537 18272
rect 3476 18232 3482 18244
rect 4525 18241 4537 18244
rect 4571 18241 4583 18275
rect 7558 18272 7564 18284
rect 4525 18235 4583 18241
rect 6104 18244 7564 18272
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18173 1823 18207
rect 1765 18167 1823 18173
rect 2225 18207 2283 18213
rect 2225 18173 2237 18207
rect 2271 18204 2283 18207
rect 2317 18207 2375 18213
rect 2317 18204 2329 18207
rect 2271 18176 2329 18204
rect 2271 18173 2283 18176
rect 2225 18167 2283 18173
rect 2317 18173 2329 18176
rect 2363 18173 2375 18207
rect 3970 18204 3976 18216
rect 2317 18167 2375 18173
rect 2516 18176 3832 18204
rect 3931 18176 3976 18204
rect 1780 18136 1808 18167
rect 2516 18136 2544 18176
rect 1780 18108 2544 18136
rect 2584 18139 2642 18145
rect 2584 18105 2596 18139
rect 2630 18136 2642 18139
rect 3602 18136 3608 18148
rect 2630 18108 3608 18136
rect 2630 18105 2642 18108
rect 2584 18099 2642 18105
rect 3602 18096 3608 18108
rect 3660 18096 3666 18148
rect 3804 18136 3832 18176
rect 3970 18164 3976 18176
rect 4028 18164 4034 18216
rect 6104 18204 6132 18244
rect 7558 18232 7564 18244
rect 7616 18232 7622 18284
rect 7760 18281 7788 18312
rect 8294 18300 8300 18312
rect 8352 18300 8358 18352
rect 10134 18300 10140 18352
rect 10192 18300 10198 18352
rect 7745 18275 7803 18281
rect 7745 18241 7757 18275
rect 7791 18241 7803 18275
rect 7926 18272 7932 18284
rect 7887 18244 7932 18272
rect 7745 18235 7803 18241
rect 7926 18232 7932 18244
rect 7984 18232 7990 18284
rect 9769 18275 9827 18281
rect 9769 18272 9781 18275
rect 9324 18244 9781 18272
rect 4632 18176 6132 18204
rect 6181 18207 6239 18213
rect 4632 18136 4660 18176
rect 6181 18173 6193 18207
rect 6227 18204 6239 18207
rect 6822 18204 6828 18216
rect 6227 18176 6828 18204
rect 6227 18173 6239 18176
rect 6181 18167 6239 18173
rect 3804 18108 4660 18136
rect 4792 18139 4850 18145
rect 4792 18105 4804 18139
rect 4838 18105 4850 18139
rect 4792 18099 4850 18105
rect 2225 18071 2283 18077
rect 2225 18037 2237 18071
rect 2271 18068 2283 18071
rect 2314 18068 2320 18080
rect 2271 18040 2320 18068
rect 2271 18037 2283 18040
rect 2225 18031 2283 18037
rect 2314 18028 2320 18040
rect 2372 18068 2378 18080
rect 3418 18068 3424 18080
rect 2372 18040 3424 18068
rect 2372 18028 2378 18040
rect 3418 18028 3424 18040
rect 3476 18028 3482 18080
rect 4807 18068 4835 18099
rect 5626 18096 5632 18148
rect 5684 18136 5690 18148
rect 6196 18136 6224 18167
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 8202 18164 8208 18216
rect 8260 18204 8266 18216
rect 8297 18207 8355 18213
rect 8297 18204 8309 18207
rect 8260 18176 8309 18204
rect 8260 18164 8266 18176
rect 8297 18173 8309 18176
rect 8343 18204 8355 18207
rect 8386 18204 8392 18216
rect 8343 18176 8392 18204
rect 8343 18173 8355 18176
rect 8297 18167 8355 18173
rect 8386 18164 8392 18176
rect 8444 18164 8450 18216
rect 9324 18204 9352 18244
rect 9769 18241 9781 18244
rect 9815 18241 9827 18275
rect 9769 18235 9827 18241
rect 9858 18204 9864 18216
rect 8496 18176 9352 18204
rect 9600 18176 9864 18204
rect 5684 18108 6224 18136
rect 7653 18139 7711 18145
rect 5684 18096 5690 18108
rect 7653 18105 7665 18139
rect 7699 18136 7711 18139
rect 8496 18136 8524 18176
rect 7699 18108 8524 18136
rect 8564 18139 8622 18145
rect 7699 18105 7711 18108
rect 7653 18099 7711 18105
rect 8564 18105 8576 18139
rect 8610 18136 8622 18139
rect 9600 18136 9628 18176
rect 9858 18164 9864 18176
rect 9916 18164 9922 18216
rect 10152 18213 10180 18300
rect 10229 18275 10287 18281
rect 10229 18241 10241 18275
rect 10275 18272 10287 18275
rect 10275 18244 10364 18272
rect 10275 18241 10287 18244
rect 10229 18235 10287 18241
rect 10336 18216 10364 18244
rect 12066 18232 12072 18284
rect 12124 18272 12130 18284
rect 13004 18272 13032 18380
rect 14369 18377 14381 18380
rect 14415 18377 14427 18411
rect 14369 18371 14427 18377
rect 14826 18368 14832 18420
rect 14884 18408 14890 18420
rect 16390 18408 16396 18420
rect 14884 18380 16396 18408
rect 14884 18368 14890 18380
rect 16390 18368 16396 18380
rect 16448 18368 16454 18420
rect 16669 18411 16727 18417
rect 16669 18377 16681 18411
rect 16715 18408 16727 18411
rect 18690 18408 18696 18420
rect 16715 18380 18696 18408
rect 16715 18377 16727 18380
rect 16669 18371 16727 18377
rect 18690 18368 18696 18380
rect 18748 18368 18754 18420
rect 19334 18368 19340 18420
rect 19392 18408 19398 18420
rect 19429 18411 19487 18417
rect 19429 18408 19441 18411
rect 19392 18380 19441 18408
rect 19392 18368 19398 18380
rect 19429 18377 19441 18380
rect 19475 18377 19487 18411
rect 19429 18371 19487 18377
rect 14090 18300 14096 18352
rect 14148 18340 14154 18352
rect 14148 18312 17264 18340
rect 14148 18300 14154 18312
rect 12124 18244 13032 18272
rect 12124 18232 12130 18244
rect 14918 18232 14924 18284
rect 14976 18272 14982 18284
rect 15197 18275 15255 18281
rect 15197 18272 15209 18275
rect 14976 18244 15209 18272
rect 14976 18232 14982 18244
rect 15197 18241 15209 18244
rect 15243 18241 15255 18275
rect 16206 18272 16212 18284
rect 16167 18244 16212 18272
rect 15197 18235 15255 18241
rect 16206 18232 16212 18244
rect 16264 18232 16270 18284
rect 17236 18281 17264 18312
rect 17494 18300 17500 18352
rect 17552 18340 17558 18352
rect 17681 18343 17739 18349
rect 17681 18340 17693 18343
rect 17552 18312 17693 18340
rect 17552 18300 17558 18312
rect 17681 18309 17693 18312
rect 17727 18309 17739 18343
rect 17681 18303 17739 18309
rect 17221 18275 17279 18281
rect 17221 18241 17233 18275
rect 17267 18241 17279 18275
rect 17696 18272 17724 18303
rect 20070 18300 20076 18352
rect 20128 18340 20134 18352
rect 20128 18312 20392 18340
rect 20128 18300 20134 18312
rect 18046 18272 18052 18284
rect 17696 18244 18052 18272
rect 17221 18235 17279 18241
rect 18046 18232 18052 18244
rect 18104 18232 18110 18284
rect 10137 18207 10195 18213
rect 10137 18173 10149 18207
rect 10183 18173 10195 18207
rect 10137 18167 10195 18173
rect 10318 18164 10324 18216
rect 10376 18164 10382 18216
rect 10778 18204 10784 18216
rect 10428 18176 10784 18204
rect 10428 18136 10456 18176
rect 10778 18164 10784 18176
rect 10836 18164 10842 18216
rect 12434 18164 12440 18216
rect 12492 18204 12498 18216
rect 12492 18176 12537 18204
rect 12492 18164 12498 18176
rect 12802 18164 12808 18216
rect 12860 18204 12866 18216
rect 12989 18207 13047 18213
rect 12989 18204 13001 18207
rect 12860 18176 13001 18204
rect 12860 18164 12866 18176
rect 12989 18173 13001 18176
rect 13035 18173 13047 18207
rect 14734 18204 14740 18216
rect 12989 18167 13047 18173
rect 13188 18176 14740 18204
rect 8610 18108 9628 18136
rect 9692 18108 10456 18136
rect 10496 18139 10554 18145
rect 8610 18105 8622 18108
rect 8564 18099 8622 18105
rect 5718 18068 5724 18080
rect 4807 18040 5724 18068
rect 5718 18028 5724 18040
rect 5776 18028 5782 18080
rect 5902 18068 5908 18080
rect 5863 18040 5908 18068
rect 5902 18028 5908 18040
rect 5960 18028 5966 18080
rect 6270 18028 6276 18080
rect 6328 18068 6334 18080
rect 6365 18071 6423 18077
rect 6365 18068 6377 18071
rect 6328 18040 6377 18068
rect 6328 18028 6334 18040
rect 6365 18037 6377 18040
rect 6411 18037 6423 18071
rect 6365 18031 6423 18037
rect 6825 18071 6883 18077
rect 6825 18037 6837 18071
rect 6871 18068 6883 18071
rect 8938 18068 8944 18080
rect 6871 18040 8944 18068
rect 6871 18037 6883 18040
rect 6825 18031 6883 18037
rect 8938 18028 8944 18040
rect 8996 18028 9002 18080
rect 9692 18077 9720 18108
rect 10496 18105 10508 18139
rect 10542 18136 10554 18139
rect 11698 18136 11704 18148
rect 10542 18108 11704 18136
rect 10542 18105 10554 18108
rect 10496 18099 10554 18105
rect 11698 18096 11704 18108
rect 11756 18096 11762 18148
rect 12342 18096 12348 18148
rect 12400 18136 12406 18148
rect 13188 18136 13216 18176
rect 14734 18164 14740 18176
rect 14792 18204 14798 18216
rect 16025 18207 16083 18213
rect 16025 18204 16037 18207
rect 14792 18176 16037 18204
rect 14792 18164 14798 18176
rect 16025 18173 16037 18176
rect 16071 18173 16083 18207
rect 16025 18167 16083 18173
rect 16850 18164 16856 18216
rect 16908 18204 16914 18216
rect 17129 18207 17187 18213
rect 17129 18204 17141 18207
rect 16908 18176 17141 18204
rect 16908 18164 16914 18176
rect 17129 18173 17141 18176
rect 17175 18173 17187 18207
rect 17862 18204 17868 18216
rect 17823 18176 17868 18204
rect 17129 18167 17187 18173
rect 17862 18164 17868 18176
rect 17920 18164 17926 18216
rect 19797 18207 19855 18213
rect 19797 18173 19809 18207
rect 19843 18204 19855 18207
rect 20070 18204 20076 18216
rect 19843 18176 20076 18204
rect 19843 18173 19855 18176
rect 19797 18167 19855 18173
rect 20070 18164 20076 18176
rect 20128 18164 20134 18216
rect 12400 18108 13216 18136
rect 13256 18139 13314 18145
rect 12400 18096 12406 18108
rect 13256 18105 13268 18139
rect 13302 18136 13314 18139
rect 14274 18136 14280 18148
rect 13302 18108 14280 18136
rect 13302 18105 13314 18108
rect 13256 18099 13314 18105
rect 14274 18096 14280 18108
rect 14332 18136 14338 18148
rect 15013 18139 15071 18145
rect 15013 18136 15025 18139
rect 14332 18108 15025 18136
rect 14332 18096 14338 18108
rect 15013 18105 15025 18108
rect 15059 18105 15071 18139
rect 15013 18099 15071 18105
rect 15378 18096 15384 18148
rect 15436 18136 15442 18148
rect 16117 18139 16175 18145
rect 16117 18136 16129 18139
rect 15436 18108 16129 18136
rect 15436 18096 15442 18108
rect 16117 18105 16129 18108
rect 16163 18136 16175 18139
rect 16298 18136 16304 18148
rect 16163 18108 16304 18136
rect 16163 18105 16175 18108
rect 16117 18099 16175 18105
rect 16298 18096 16304 18108
rect 16356 18096 16362 18148
rect 18316 18139 18374 18145
rect 18316 18105 18328 18139
rect 18362 18136 18374 18139
rect 18782 18136 18788 18148
rect 18362 18108 18788 18136
rect 18362 18105 18374 18108
rect 18316 18099 18374 18105
rect 18782 18096 18788 18108
rect 18840 18096 18846 18148
rect 20364 18080 20392 18312
rect 20714 18232 20720 18284
rect 20772 18272 20778 18284
rect 20901 18275 20959 18281
rect 20901 18272 20913 18275
rect 20772 18244 20913 18272
rect 20772 18232 20778 18244
rect 20901 18241 20913 18244
rect 20947 18241 20959 18275
rect 20901 18235 20959 18241
rect 20806 18164 20812 18216
rect 20864 18204 20870 18216
rect 21266 18204 21272 18216
rect 20864 18176 21272 18204
rect 20864 18164 20870 18176
rect 21266 18164 21272 18176
rect 21324 18204 21330 18216
rect 21361 18207 21419 18213
rect 21361 18204 21373 18207
rect 21324 18176 21373 18204
rect 21324 18164 21330 18176
rect 21361 18173 21373 18176
rect 21407 18173 21419 18207
rect 21361 18167 21419 18173
rect 21628 18207 21686 18213
rect 21628 18173 21640 18207
rect 21674 18204 21686 18207
rect 22462 18204 22468 18216
rect 21674 18176 22468 18204
rect 21674 18173 21686 18176
rect 21628 18167 21686 18173
rect 22462 18164 22468 18176
rect 22520 18164 22526 18216
rect 20717 18139 20775 18145
rect 20717 18105 20729 18139
rect 20763 18136 20775 18139
rect 22370 18136 22376 18148
rect 20763 18108 22376 18136
rect 20763 18105 20775 18108
rect 20717 18099 20775 18105
rect 22370 18096 22376 18108
rect 22428 18096 22434 18148
rect 9677 18071 9735 18077
rect 9677 18037 9689 18071
rect 9723 18037 9735 18071
rect 9677 18031 9735 18037
rect 9769 18071 9827 18077
rect 9769 18037 9781 18071
rect 9815 18068 9827 18071
rect 11885 18071 11943 18077
rect 11885 18068 11897 18071
rect 9815 18040 11897 18068
rect 9815 18037 9827 18040
rect 9769 18031 9827 18037
rect 11885 18037 11897 18040
rect 11931 18037 11943 18071
rect 11885 18031 11943 18037
rect 12526 18028 12532 18080
rect 12584 18068 12590 18080
rect 12621 18071 12679 18077
rect 12621 18068 12633 18071
rect 12584 18040 12633 18068
rect 12584 18028 12590 18040
rect 12621 18037 12633 18040
rect 12667 18037 12679 18071
rect 12621 18031 12679 18037
rect 13906 18028 13912 18080
rect 13964 18068 13970 18080
rect 14645 18071 14703 18077
rect 14645 18068 14657 18071
rect 13964 18040 14657 18068
rect 13964 18028 13970 18040
rect 14645 18037 14657 18040
rect 14691 18037 14703 18071
rect 14645 18031 14703 18037
rect 14918 18028 14924 18080
rect 14976 18068 14982 18080
rect 15105 18071 15163 18077
rect 15105 18068 15117 18071
rect 14976 18040 15117 18068
rect 14976 18028 14982 18040
rect 15105 18037 15117 18040
rect 15151 18037 15163 18071
rect 15105 18031 15163 18037
rect 15657 18071 15715 18077
rect 15657 18037 15669 18071
rect 15703 18068 15715 18071
rect 16942 18068 16948 18080
rect 15703 18040 16948 18068
rect 15703 18037 15715 18040
rect 15657 18031 15715 18037
rect 16942 18028 16948 18040
rect 17000 18028 17006 18080
rect 17037 18071 17095 18077
rect 17037 18037 17049 18071
rect 17083 18068 17095 18071
rect 17494 18068 17500 18080
rect 17083 18040 17500 18068
rect 17083 18037 17095 18040
rect 17037 18031 17095 18037
rect 17494 18028 17500 18040
rect 17552 18028 17558 18080
rect 19978 18068 19984 18080
rect 19939 18040 19984 18068
rect 19978 18028 19984 18040
rect 20036 18028 20042 18080
rect 20346 18068 20352 18080
rect 20307 18040 20352 18068
rect 20346 18028 20352 18040
rect 20404 18028 20410 18080
rect 20438 18028 20444 18080
rect 20496 18068 20502 18080
rect 20809 18071 20867 18077
rect 20809 18068 20821 18071
rect 20496 18040 20821 18068
rect 20496 18028 20502 18040
rect 20809 18037 20821 18040
rect 20855 18037 20867 18071
rect 20809 18031 20867 18037
rect 21174 18028 21180 18080
rect 21232 18068 21238 18080
rect 22741 18071 22799 18077
rect 22741 18068 22753 18071
rect 21232 18040 22753 18068
rect 21232 18028 21238 18040
rect 22741 18037 22753 18040
rect 22787 18037 22799 18071
rect 22741 18031 22799 18037
rect 1104 17978 23276 18000
rect 1104 17926 8379 17978
rect 8431 17926 8443 17978
rect 8495 17926 8507 17978
rect 8559 17926 8571 17978
rect 8623 17926 15776 17978
rect 15828 17926 15840 17978
rect 15892 17926 15904 17978
rect 15956 17926 15968 17978
rect 16020 17926 23276 17978
rect 1104 17904 23276 17926
rect 2774 17824 2780 17876
rect 2832 17864 2838 17876
rect 2832 17836 12572 17864
rect 2832 17824 2838 17836
rect 2590 17796 2596 17808
rect 1688 17768 2596 17796
rect 1688 17737 1716 17768
rect 2590 17756 2596 17768
rect 2648 17756 2654 17808
rect 10588 17799 10646 17805
rect 3988 17768 9904 17796
rect 1673 17731 1731 17737
rect 1673 17697 1685 17731
rect 1719 17697 1731 17731
rect 1673 17691 1731 17697
rect 2225 17731 2283 17737
rect 2225 17697 2237 17731
rect 2271 17728 2283 17731
rect 2314 17728 2320 17740
rect 2271 17700 2320 17728
rect 2271 17697 2283 17700
rect 2225 17691 2283 17697
rect 2314 17688 2320 17700
rect 2372 17688 2378 17740
rect 2492 17731 2550 17737
rect 2492 17697 2504 17731
rect 2538 17728 2550 17731
rect 3510 17728 3516 17740
rect 2538 17700 3516 17728
rect 2538 17697 2550 17700
rect 2492 17691 2550 17697
rect 3510 17688 3516 17700
rect 3568 17688 3574 17740
rect 3602 17592 3608 17604
rect 3563 17564 3608 17592
rect 3602 17552 3608 17564
rect 3660 17552 3666 17604
rect 1857 17527 1915 17533
rect 1857 17493 1869 17527
rect 1903 17524 1915 17527
rect 3988 17524 4016 17768
rect 4062 17688 4068 17740
rect 4120 17688 4126 17740
rect 4249 17731 4307 17737
rect 4249 17697 4261 17731
rect 4295 17728 4307 17731
rect 4430 17728 4436 17740
rect 4295 17700 4436 17728
rect 4295 17697 4307 17700
rect 4249 17691 4307 17697
rect 4430 17688 4436 17700
rect 4488 17688 4494 17740
rect 5057 17731 5115 17737
rect 5057 17728 5069 17731
rect 4540 17700 5069 17728
rect 4080 17592 4108 17688
rect 4154 17620 4160 17672
rect 4212 17660 4218 17672
rect 4540 17660 4568 17700
rect 5057 17697 5069 17700
rect 5103 17728 5115 17731
rect 5902 17728 5908 17740
rect 5103 17700 5908 17728
rect 5103 17697 5115 17700
rect 5057 17691 5115 17697
rect 5902 17688 5908 17700
rect 5960 17688 5966 17740
rect 6713 17731 6771 17737
rect 6713 17728 6725 17731
rect 6196 17700 6725 17728
rect 4798 17660 4804 17672
rect 4212 17632 4568 17660
rect 4759 17632 4804 17660
rect 4212 17620 4218 17632
rect 4798 17620 4804 17632
rect 4856 17620 4862 17672
rect 4080 17564 4568 17592
rect 1903 17496 4016 17524
rect 1903 17493 1915 17496
rect 1857 17487 1915 17493
rect 4154 17484 4160 17536
rect 4212 17524 4218 17536
rect 4433 17527 4491 17533
rect 4433 17524 4445 17527
rect 4212 17496 4445 17524
rect 4212 17484 4218 17496
rect 4433 17493 4445 17496
rect 4479 17493 4491 17527
rect 4540 17524 4568 17564
rect 5442 17524 5448 17536
rect 4540 17496 5448 17524
rect 4433 17487 4491 17493
rect 5442 17484 5448 17496
rect 5500 17484 5506 17536
rect 6086 17484 6092 17536
rect 6144 17524 6150 17536
rect 6196 17533 6224 17700
rect 6713 17697 6725 17700
rect 6759 17697 6771 17731
rect 6713 17691 6771 17697
rect 8481 17731 8539 17737
rect 8481 17697 8493 17731
rect 8527 17728 8539 17731
rect 8754 17728 8760 17740
rect 8527 17700 8760 17728
rect 8527 17697 8539 17700
rect 8481 17691 8539 17697
rect 8754 17688 8760 17700
rect 8812 17688 8818 17740
rect 9677 17731 9735 17737
rect 9677 17697 9689 17731
rect 9723 17697 9735 17731
rect 9876 17728 9904 17768
rect 10588 17765 10600 17799
rect 10634 17796 10646 17799
rect 11790 17796 11796 17808
rect 10634 17768 11796 17796
rect 10634 17765 10646 17768
rect 10588 17759 10646 17765
rect 11790 17756 11796 17768
rect 11848 17796 11854 17808
rect 12066 17796 12072 17808
rect 11848 17768 12072 17796
rect 11848 17756 11854 17768
rect 12066 17756 12072 17768
rect 12124 17756 12130 17808
rect 12434 17796 12440 17808
rect 12176 17768 12440 17796
rect 12176 17728 12204 17768
rect 12434 17756 12440 17768
rect 12492 17756 12498 17808
rect 12544 17796 12572 17836
rect 12710 17824 12716 17876
rect 12768 17864 12774 17876
rect 13722 17864 13728 17876
rect 12768 17836 13728 17864
rect 12768 17824 12774 17836
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 14274 17864 14280 17876
rect 14235 17836 14280 17864
rect 14274 17824 14280 17836
rect 14332 17824 14338 17876
rect 14829 17867 14887 17873
rect 14829 17833 14841 17867
rect 14875 17864 14887 17867
rect 16206 17864 16212 17876
rect 14875 17836 16212 17864
rect 14875 17833 14887 17836
rect 14829 17827 14887 17833
rect 16206 17824 16212 17836
rect 16264 17824 16270 17876
rect 18782 17864 18788 17876
rect 18743 17836 18788 17864
rect 18782 17824 18788 17836
rect 18840 17864 18846 17876
rect 19521 17867 19579 17873
rect 19521 17864 19533 17867
rect 18840 17836 19533 17864
rect 18840 17824 18846 17836
rect 19521 17833 19533 17836
rect 19567 17833 19579 17867
rect 22646 17864 22652 17876
rect 19521 17827 19579 17833
rect 19628 17836 22652 17864
rect 15286 17796 15292 17808
rect 12544 17768 15292 17796
rect 15286 17756 15292 17768
rect 15344 17756 15350 17808
rect 15470 17756 15476 17808
rect 15528 17805 15534 17808
rect 15528 17799 15592 17805
rect 15528 17765 15546 17799
rect 15580 17796 15592 17799
rect 16114 17796 16120 17808
rect 15580 17768 16120 17796
rect 15580 17765 15592 17768
rect 15528 17759 15592 17765
rect 15528 17756 15534 17759
rect 16114 17756 16120 17768
rect 16172 17756 16178 17808
rect 16298 17756 16304 17808
rect 16356 17796 16362 17808
rect 16945 17799 17003 17805
rect 16945 17796 16957 17799
rect 16356 17768 16957 17796
rect 16356 17756 16362 17768
rect 16945 17765 16957 17768
rect 16991 17765 17003 17799
rect 18046 17796 18052 17808
rect 16945 17759 17003 17765
rect 17420 17768 18052 17796
rect 12342 17728 12348 17740
rect 9876 17700 12204 17728
rect 12303 17700 12348 17728
rect 9677 17691 9735 17697
rect 6454 17660 6460 17672
rect 6415 17632 6460 17660
rect 6454 17620 6460 17632
rect 6512 17620 6518 17672
rect 8570 17660 8576 17672
rect 8531 17632 8576 17660
rect 8570 17620 8576 17632
rect 8628 17620 8634 17672
rect 8665 17663 8723 17669
rect 8665 17629 8677 17663
rect 8711 17660 8723 17663
rect 9030 17660 9036 17672
rect 8711 17632 9036 17660
rect 8711 17629 8723 17632
rect 8665 17623 8723 17629
rect 9030 17620 9036 17632
rect 9088 17620 9094 17672
rect 9125 17663 9183 17669
rect 9125 17629 9137 17663
rect 9171 17660 9183 17663
rect 9398 17660 9404 17672
rect 9171 17632 9404 17660
rect 9171 17629 9183 17632
rect 9125 17623 9183 17629
rect 9398 17620 9404 17632
rect 9456 17620 9462 17672
rect 9692 17660 9720 17691
rect 12342 17688 12348 17700
rect 12400 17688 12406 17740
rect 12802 17688 12808 17740
rect 12860 17728 12866 17740
rect 12904 17731 12962 17737
rect 12904 17728 12916 17731
rect 12860 17700 12916 17728
rect 12860 17688 12866 17700
rect 12904 17697 12916 17700
rect 12950 17697 12962 17731
rect 12904 17691 12962 17697
rect 13164 17731 13222 17737
rect 13164 17697 13176 17731
rect 13210 17728 13222 17731
rect 14645 17731 14703 17737
rect 13210 17700 13952 17728
rect 13210 17697 13222 17700
rect 13164 17691 13222 17697
rect 10318 17660 10324 17672
rect 9692 17632 10180 17660
rect 10279 17632 10324 17660
rect 9490 17552 9496 17604
rect 9548 17592 9554 17604
rect 9861 17595 9919 17601
rect 9861 17592 9873 17595
rect 9548 17564 9873 17592
rect 9548 17552 9554 17564
rect 9861 17561 9873 17564
rect 9907 17561 9919 17595
rect 10152 17592 10180 17632
rect 10318 17620 10324 17632
rect 10376 17620 10382 17672
rect 13924 17660 13952 17700
rect 14645 17697 14657 17731
rect 14691 17728 14703 17731
rect 17126 17728 17132 17740
rect 14691 17700 17132 17728
rect 14691 17697 14703 17700
rect 14645 17691 14703 17697
rect 17126 17688 17132 17700
rect 17184 17688 17190 17740
rect 17420 17737 17448 17768
rect 18046 17756 18052 17768
rect 18104 17756 18110 17808
rect 19334 17756 19340 17808
rect 19392 17796 19398 17808
rect 19429 17799 19487 17805
rect 19429 17796 19441 17799
rect 19392 17768 19441 17796
rect 19392 17756 19398 17768
rect 19429 17765 19441 17768
rect 19475 17765 19487 17799
rect 19628 17796 19656 17836
rect 22646 17824 22652 17836
rect 22704 17824 22710 17876
rect 21174 17805 21180 17808
rect 21168 17796 21180 17805
rect 19429 17759 19487 17765
rect 19536 17768 19656 17796
rect 21135 17768 21180 17796
rect 17405 17731 17463 17737
rect 17405 17697 17417 17731
rect 17451 17697 17463 17731
rect 17405 17691 17463 17697
rect 17672 17731 17730 17737
rect 17672 17697 17684 17731
rect 17718 17728 17730 17731
rect 18966 17728 18972 17740
rect 17718 17700 18972 17728
rect 17718 17697 17730 17700
rect 17672 17691 17730 17697
rect 18966 17688 18972 17700
rect 19024 17688 19030 17740
rect 19242 17688 19248 17740
rect 19300 17728 19306 17740
rect 19536 17728 19564 17768
rect 21168 17759 21180 17768
rect 21174 17756 21180 17759
rect 21232 17756 21238 17808
rect 19886 17728 19892 17740
rect 19300 17700 19564 17728
rect 19628 17700 19892 17728
rect 19300 17688 19306 17700
rect 13998 17660 14004 17672
rect 13924 17632 14004 17660
rect 13998 17620 14004 17632
rect 14056 17620 14062 17672
rect 15289 17663 15347 17669
rect 15289 17629 15301 17663
rect 15335 17629 15347 17663
rect 15289 17623 15347 17629
rect 10226 17592 10232 17604
rect 10152 17564 10232 17592
rect 9861 17555 9919 17561
rect 10226 17552 10232 17564
rect 10284 17552 10290 17604
rect 11698 17592 11704 17604
rect 11659 17564 11704 17592
rect 11698 17552 11704 17564
rect 11756 17552 11762 17604
rect 12529 17595 12587 17601
rect 12529 17561 12541 17595
rect 12575 17592 12587 17595
rect 12894 17592 12900 17604
rect 12575 17564 12900 17592
rect 12575 17561 12587 17564
rect 12529 17555 12587 17561
rect 12894 17552 12900 17564
rect 12952 17552 12958 17604
rect 14826 17552 14832 17604
rect 14884 17592 14890 17604
rect 15102 17592 15108 17604
rect 14884 17564 15108 17592
rect 14884 17552 14890 17564
rect 15102 17552 15108 17564
rect 15160 17592 15166 17604
rect 15304 17592 15332 17623
rect 18414 17620 18420 17672
rect 18472 17660 18478 17672
rect 19628 17660 19656 17700
rect 19886 17688 19892 17700
rect 19944 17688 19950 17740
rect 20257 17731 20315 17737
rect 20257 17697 20269 17731
rect 20303 17728 20315 17731
rect 20530 17728 20536 17740
rect 20303 17700 20536 17728
rect 20303 17697 20315 17700
rect 20257 17691 20315 17697
rect 20530 17688 20536 17700
rect 20588 17688 20594 17740
rect 22557 17731 22615 17737
rect 22557 17728 22569 17731
rect 20640 17700 22569 17728
rect 18472 17632 19656 17660
rect 19705 17663 19763 17669
rect 18472 17620 18478 17632
rect 19705 17629 19717 17663
rect 19751 17660 19763 17663
rect 19794 17660 19800 17672
rect 19751 17632 19800 17660
rect 19751 17629 19763 17632
rect 19705 17623 19763 17629
rect 19794 17620 19800 17632
rect 19852 17620 19858 17672
rect 20346 17620 20352 17672
rect 20404 17660 20410 17672
rect 20640 17660 20668 17700
rect 22557 17697 22569 17700
rect 22603 17697 22615 17731
rect 22557 17691 22615 17697
rect 20404 17632 20668 17660
rect 20404 17620 20410 17632
rect 20806 17620 20812 17672
rect 20864 17660 20870 17672
rect 20901 17663 20959 17669
rect 20901 17660 20913 17663
rect 20864 17632 20913 17660
rect 20864 17620 20870 17632
rect 20901 17629 20913 17632
rect 20947 17629 20959 17663
rect 20901 17623 20959 17629
rect 15160 17564 15332 17592
rect 18892 17564 20944 17592
rect 15160 17552 15166 17564
rect 6181 17527 6239 17533
rect 6181 17524 6193 17527
rect 6144 17496 6193 17524
rect 6144 17484 6150 17496
rect 6181 17493 6193 17496
rect 6227 17493 6239 17527
rect 7834 17524 7840 17536
rect 7795 17496 7840 17524
rect 6181 17487 6239 17493
rect 7834 17484 7840 17496
rect 7892 17484 7898 17536
rect 8018 17484 8024 17536
rect 8076 17524 8082 17536
rect 8113 17527 8171 17533
rect 8113 17524 8125 17527
rect 8076 17496 8125 17524
rect 8076 17484 8082 17496
rect 8113 17493 8125 17496
rect 8159 17493 8171 17527
rect 8113 17487 8171 17493
rect 9214 17484 9220 17536
rect 9272 17524 9278 17536
rect 11514 17524 11520 17536
rect 9272 17496 11520 17524
rect 9272 17484 9278 17496
rect 11514 17484 11520 17496
rect 11572 17484 11578 17536
rect 16666 17524 16672 17536
rect 16627 17496 16672 17524
rect 16666 17484 16672 17496
rect 16724 17484 16730 17536
rect 17402 17484 17408 17536
rect 17460 17524 17466 17536
rect 18892 17524 18920 17564
rect 19058 17524 19064 17536
rect 17460 17496 18920 17524
rect 19019 17496 19064 17524
rect 17460 17484 17466 17496
rect 19058 17484 19064 17496
rect 19116 17484 19122 17536
rect 20162 17484 20168 17536
rect 20220 17524 20226 17536
rect 20441 17527 20499 17533
rect 20441 17524 20453 17527
rect 20220 17496 20453 17524
rect 20220 17484 20226 17496
rect 20441 17493 20453 17496
rect 20487 17493 20499 17527
rect 20916 17524 20944 17564
rect 21542 17524 21548 17536
rect 20916 17496 21548 17524
rect 20441 17487 20499 17493
rect 21542 17484 21548 17496
rect 21600 17484 21606 17536
rect 22002 17484 22008 17536
rect 22060 17524 22066 17536
rect 22281 17527 22339 17533
rect 22281 17524 22293 17527
rect 22060 17496 22293 17524
rect 22060 17484 22066 17496
rect 22281 17493 22293 17496
rect 22327 17493 22339 17527
rect 22281 17487 22339 17493
rect 1104 17434 23276 17456
rect 1104 17382 4680 17434
rect 4732 17382 4744 17434
rect 4796 17382 4808 17434
rect 4860 17382 4872 17434
rect 4924 17382 12078 17434
rect 12130 17382 12142 17434
rect 12194 17382 12206 17434
rect 12258 17382 12270 17434
rect 12322 17382 19475 17434
rect 19527 17382 19539 17434
rect 19591 17382 19603 17434
rect 19655 17382 19667 17434
rect 19719 17382 23276 17434
rect 1104 17360 23276 17382
rect 1394 17280 1400 17332
rect 1452 17320 1458 17332
rect 3510 17320 3516 17332
rect 1452 17292 3372 17320
rect 3471 17292 3516 17320
rect 1452 17280 1458 17292
rect 3344 17252 3372 17292
rect 3510 17280 3516 17292
rect 3568 17320 3574 17332
rect 4338 17320 4344 17332
rect 3568 17292 4344 17320
rect 3568 17280 3574 17292
rect 4338 17280 4344 17292
rect 4396 17280 4402 17332
rect 4430 17280 4436 17332
rect 4488 17320 4494 17332
rect 5074 17320 5080 17332
rect 4488 17292 5080 17320
rect 4488 17280 4494 17292
rect 5074 17280 5080 17292
rect 5132 17280 5138 17332
rect 5166 17280 5172 17332
rect 5224 17320 5230 17332
rect 5350 17320 5356 17332
rect 5224 17292 5356 17320
rect 5224 17280 5230 17292
rect 5350 17280 5356 17292
rect 5408 17280 5414 17332
rect 5534 17280 5540 17332
rect 5592 17320 5598 17332
rect 11701 17323 11759 17329
rect 5592 17292 11284 17320
rect 5592 17280 5598 17292
rect 3694 17252 3700 17264
rect 3344 17224 3700 17252
rect 3694 17212 3700 17224
rect 3752 17212 3758 17264
rect 3789 17255 3847 17261
rect 3789 17221 3801 17255
rect 3835 17252 3847 17255
rect 4062 17252 4068 17264
rect 3835 17224 4068 17252
rect 3835 17221 3847 17224
rect 3789 17215 3847 17221
rect 4062 17212 4068 17224
rect 4120 17212 4126 17264
rect 4614 17212 4620 17264
rect 4672 17252 4678 17264
rect 4801 17255 4859 17261
rect 4801 17252 4813 17255
rect 4672 17224 4813 17252
rect 4672 17212 4678 17224
rect 4801 17221 4813 17224
rect 4847 17221 4859 17255
rect 6822 17252 6828 17264
rect 4801 17215 4859 17221
rect 5828 17224 6828 17252
rect 3602 17144 3608 17196
rect 3660 17184 3666 17196
rect 4433 17187 4491 17193
rect 4433 17184 4445 17187
rect 3660 17156 4445 17184
rect 3660 17144 3666 17156
rect 4433 17153 4445 17156
rect 4479 17153 4491 17187
rect 4433 17147 4491 17153
rect 4706 17144 4712 17196
rect 4764 17184 4770 17196
rect 5353 17187 5411 17193
rect 5353 17184 5365 17187
rect 4764 17156 5365 17184
rect 4764 17144 4770 17156
rect 5353 17153 5365 17156
rect 5399 17153 5411 17187
rect 5353 17147 5411 17153
rect 1581 17119 1639 17125
rect 1581 17085 1593 17119
rect 1627 17085 1639 17119
rect 1581 17079 1639 17085
rect 2133 17119 2191 17125
rect 2133 17085 2145 17119
rect 2179 17116 2191 17119
rect 2222 17116 2228 17128
rect 2179 17088 2228 17116
rect 2179 17085 2191 17088
rect 2133 17079 2191 17085
rect 1596 17048 1624 17079
rect 2222 17076 2228 17088
rect 2280 17076 2286 17128
rect 4062 17116 4068 17128
rect 2332 17088 4068 17116
rect 2332 17048 2360 17088
rect 4062 17076 4068 17088
rect 4120 17076 4126 17128
rect 4157 17119 4215 17125
rect 4157 17085 4169 17119
rect 4203 17116 4215 17119
rect 5169 17119 5227 17125
rect 4203 17088 4476 17116
rect 4203 17085 4215 17088
rect 4157 17079 4215 17085
rect 1596 17020 2360 17048
rect 2400 17051 2458 17057
rect 2400 17017 2412 17051
rect 2446 17048 2458 17051
rect 3326 17048 3332 17060
rect 2446 17020 3332 17048
rect 2446 17017 2458 17020
rect 2400 17011 2458 17017
rect 3326 17008 3332 17020
rect 3384 17008 3390 17060
rect 1765 16983 1823 16989
rect 1765 16949 1777 16983
rect 1811 16980 1823 16983
rect 4062 16980 4068 16992
rect 1811 16952 4068 16980
rect 1811 16949 1823 16952
rect 1765 16943 1823 16949
rect 4062 16940 4068 16952
rect 4120 16940 4126 16992
rect 4246 16940 4252 16992
rect 4304 16980 4310 16992
rect 4448 16980 4476 17088
rect 5169 17085 5181 17119
rect 5215 17116 5227 17119
rect 5828 17116 5856 17224
rect 6822 17212 6828 17224
rect 6880 17212 6886 17264
rect 9861 17255 9919 17261
rect 9861 17252 9873 17255
rect 9508 17224 9873 17252
rect 5994 17144 6000 17196
rect 6052 17184 6058 17196
rect 6052 17156 6224 17184
rect 6052 17144 6058 17156
rect 6196 17125 6224 17156
rect 5215 17088 5856 17116
rect 6089 17119 6147 17125
rect 5215 17085 5227 17088
rect 5169 17079 5227 17085
rect 6089 17085 6101 17119
rect 6135 17085 6147 17119
rect 6089 17079 6147 17085
rect 6181 17119 6239 17125
rect 6181 17085 6193 17119
rect 6227 17085 6239 17119
rect 6181 17079 6239 17085
rect 5994 17008 6000 17060
rect 6052 17048 6058 17060
rect 6104 17048 6132 17079
rect 6546 17076 6552 17128
rect 6604 17116 6610 17128
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 6604 17088 6837 17116
rect 6604 17076 6610 17088
rect 6825 17085 6837 17088
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 7092 17119 7150 17125
rect 7092 17085 7104 17119
rect 7138 17116 7150 17119
rect 7834 17116 7840 17128
rect 7138 17088 7840 17116
rect 7138 17085 7150 17088
rect 7092 17079 7150 17085
rect 7834 17076 7840 17088
rect 7892 17076 7898 17128
rect 8294 17076 8300 17128
rect 8352 17116 8358 17128
rect 8481 17119 8539 17125
rect 8481 17116 8493 17119
rect 8352 17088 8493 17116
rect 8352 17076 8358 17088
rect 8481 17085 8493 17088
rect 8527 17085 8539 17119
rect 9508 17116 9536 17224
rect 9861 17221 9873 17224
rect 9907 17221 9919 17255
rect 11256 17252 11284 17292
rect 11701 17289 11713 17323
rect 11747 17320 11759 17323
rect 11974 17320 11980 17332
rect 11747 17292 11980 17320
rect 11747 17289 11759 17292
rect 11701 17283 11759 17289
rect 11974 17280 11980 17292
rect 12032 17280 12038 17332
rect 13998 17320 14004 17332
rect 13911 17292 14004 17320
rect 13998 17280 14004 17292
rect 14056 17320 14062 17332
rect 14918 17320 14924 17332
rect 14056 17292 14924 17320
rect 14056 17280 14062 17292
rect 14918 17280 14924 17292
rect 14976 17280 14982 17332
rect 16482 17320 16488 17332
rect 16443 17292 16488 17320
rect 16482 17280 16488 17292
rect 16540 17280 16546 17332
rect 16945 17323 17003 17329
rect 16945 17289 16957 17323
rect 16991 17320 17003 17323
rect 20438 17320 20444 17332
rect 16991 17292 20444 17320
rect 16991 17289 17003 17292
rect 16945 17283 17003 17289
rect 20438 17280 20444 17292
rect 20496 17280 20502 17332
rect 21174 17320 21180 17332
rect 20824 17292 21180 17320
rect 12250 17252 12256 17264
rect 11256 17224 12256 17252
rect 9861 17215 9919 17221
rect 12250 17212 12256 17224
rect 12308 17212 12314 17264
rect 14826 17252 14832 17264
rect 14787 17224 14832 17252
rect 14826 17212 14832 17224
rect 14884 17212 14890 17264
rect 17126 17212 17132 17264
rect 17184 17252 17190 17264
rect 17184 17224 18092 17252
rect 17184 17212 17190 17224
rect 12618 17144 12624 17196
rect 12676 17184 12682 17196
rect 17589 17187 17647 17193
rect 12676 17156 12721 17184
rect 12676 17144 12682 17156
rect 17589 17153 17601 17187
rect 17635 17153 17647 17187
rect 17589 17147 17647 17153
rect 10318 17116 10324 17128
rect 8481 17079 8539 17085
rect 8956 17088 9536 17116
rect 10279 17088 10324 17116
rect 6564 17048 6592 17076
rect 8956 17060 8984 17088
rect 10318 17076 10324 17088
rect 10376 17076 10382 17128
rect 12888 17119 12946 17125
rect 12888 17085 12900 17119
rect 12934 17116 12946 17119
rect 13262 17116 13268 17128
rect 12934 17088 13268 17116
rect 12934 17085 12946 17088
rect 12888 17079 12946 17085
rect 13262 17076 13268 17088
rect 13320 17076 13326 17128
rect 14277 17119 14335 17125
rect 14277 17085 14289 17119
rect 14323 17116 14335 17119
rect 14366 17116 14372 17128
rect 14323 17088 14372 17116
rect 14323 17085 14335 17088
rect 14277 17079 14335 17085
rect 14366 17076 14372 17088
rect 14424 17076 14430 17128
rect 14458 17076 14464 17128
rect 14516 17116 14522 17128
rect 15013 17119 15071 17125
rect 15013 17116 15025 17119
rect 14516 17088 15025 17116
rect 14516 17076 14522 17088
rect 15013 17085 15025 17088
rect 15059 17085 15071 17119
rect 15013 17079 15071 17085
rect 15105 17119 15163 17125
rect 15105 17085 15117 17119
rect 15151 17116 15163 17119
rect 15194 17116 15200 17128
rect 15151 17088 15200 17116
rect 15151 17085 15163 17088
rect 15105 17079 15163 17085
rect 15194 17076 15200 17088
rect 15252 17076 15258 17128
rect 17313 17119 17371 17125
rect 17313 17085 17325 17119
rect 17359 17116 17371 17119
rect 17402 17116 17408 17128
rect 17359 17088 17408 17116
rect 17359 17085 17371 17088
rect 17313 17079 17371 17085
rect 17402 17076 17408 17088
rect 17460 17076 17466 17128
rect 8726 17051 8784 17057
rect 8726 17048 8738 17051
rect 6052 17020 6132 17048
rect 6288 17020 6592 17048
rect 8220 17020 8738 17048
rect 6052 17008 6058 17020
rect 4798 16980 4804 16992
rect 4304 16952 4349 16980
rect 4448 16952 4804 16980
rect 4304 16940 4310 16952
rect 4798 16940 4804 16952
rect 4856 16940 4862 16992
rect 5258 16940 5264 16992
rect 5316 16980 5322 16992
rect 5905 16983 5963 16989
rect 5316 16952 5361 16980
rect 5316 16940 5322 16952
rect 5905 16949 5917 16983
rect 5951 16980 5963 16983
rect 6288 16980 6316 17020
rect 5951 16952 6316 16980
rect 6365 16983 6423 16989
rect 5951 16949 5963 16952
rect 5905 16943 5963 16949
rect 6365 16949 6377 16983
rect 6411 16980 6423 16983
rect 7282 16980 7288 16992
rect 6411 16952 7288 16980
rect 6411 16949 6423 16952
rect 6365 16943 6423 16949
rect 7282 16940 7288 16952
rect 7340 16940 7346 16992
rect 7834 16940 7840 16992
rect 7892 16980 7898 16992
rect 8220 16989 8248 17020
rect 8726 17017 8738 17020
rect 8772 17017 8784 17051
rect 8726 17011 8784 17017
rect 8938 17008 8944 17060
rect 8996 17008 9002 17060
rect 10588 17051 10646 17057
rect 10588 17017 10600 17051
rect 10634 17048 10646 17051
rect 11054 17048 11060 17060
rect 10634 17020 11060 17048
rect 10634 17017 10646 17020
rect 10588 17011 10646 17017
rect 11054 17008 11060 17020
rect 11112 17008 11118 17060
rect 13814 17048 13820 17060
rect 11440 17020 13820 17048
rect 8205 16983 8263 16989
rect 8205 16980 8217 16983
rect 7892 16952 8217 16980
rect 7892 16940 7898 16952
rect 8205 16949 8217 16952
rect 8251 16949 8263 16983
rect 8205 16943 8263 16949
rect 8846 16940 8852 16992
rect 8904 16980 8910 16992
rect 11440 16980 11468 17020
rect 13814 17008 13820 17020
rect 13872 17008 13878 17060
rect 15372 17051 15430 17057
rect 15372 17017 15384 17051
rect 15418 17017 15430 17051
rect 17604 17048 17632 17147
rect 18064 17125 18092 17224
rect 19794 17212 19800 17264
rect 19852 17212 19858 17264
rect 19245 17187 19303 17193
rect 19245 17153 19257 17187
rect 19291 17184 19303 17187
rect 19812 17184 19840 17212
rect 19291 17156 19840 17184
rect 19291 17153 19303 17156
rect 19245 17147 19303 17153
rect 19978 17144 19984 17196
rect 20036 17184 20042 17196
rect 20257 17187 20315 17193
rect 20257 17184 20269 17187
rect 20036 17156 20269 17184
rect 20036 17144 20042 17156
rect 20257 17153 20269 17156
rect 20303 17153 20315 17187
rect 20257 17147 20315 17153
rect 20441 17187 20499 17193
rect 20441 17153 20453 17187
rect 20487 17184 20499 17187
rect 20824 17184 20852 17292
rect 21174 17280 21180 17292
rect 21232 17280 21238 17332
rect 22189 17255 22247 17261
rect 22189 17221 22201 17255
rect 22235 17221 22247 17255
rect 22189 17215 22247 17221
rect 20487 17156 20852 17184
rect 20487 17153 20499 17156
rect 20441 17147 20499 17153
rect 18049 17119 18107 17125
rect 18049 17085 18061 17119
rect 18095 17085 18107 17119
rect 18966 17116 18972 17128
rect 18927 17088 18972 17116
rect 18049 17079 18107 17085
rect 18966 17076 18972 17088
rect 19024 17076 19030 17128
rect 19061 17119 19119 17125
rect 19061 17085 19073 17119
rect 19107 17116 19119 17119
rect 19794 17116 19800 17128
rect 19107 17088 19800 17116
rect 19107 17085 19119 17088
rect 19061 17079 19119 17085
rect 19794 17076 19800 17088
rect 19852 17076 19858 17128
rect 20162 17116 20168 17128
rect 20123 17088 20168 17116
rect 20162 17076 20168 17088
rect 20220 17076 20226 17128
rect 20806 17116 20812 17128
rect 20767 17088 20812 17116
rect 20806 17076 20812 17088
rect 20864 17076 20870 17128
rect 21076 17119 21134 17125
rect 21076 17085 21088 17119
rect 21122 17116 21134 17119
rect 22002 17116 22008 17128
rect 21122 17088 22008 17116
rect 21122 17085 21134 17088
rect 21076 17079 21134 17085
rect 22002 17076 22008 17088
rect 22060 17076 22066 17128
rect 21634 17048 21640 17060
rect 17604 17020 21640 17048
rect 15372 17011 15430 17017
rect 8904 16952 11468 16980
rect 8904 16940 8910 16952
rect 11514 16940 11520 16992
rect 11572 16980 11578 16992
rect 13078 16980 13084 16992
rect 11572 16952 13084 16980
rect 11572 16940 11578 16952
rect 13078 16940 13084 16952
rect 13136 16940 13142 16992
rect 14461 16983 14519 16989
rect 14461 16949 14473 16983
rect 14507 16980 14519 16983
rect 14918 16980 14924 16992
rect 14507 16952 14924 16980
rect 14507 16949 14519 16952
rect 14461 16943 14519 16949
rect 14918 16940 14924 16952
rect 14976 16940 14982 16992
rect 15010 16940 15016 16992
rect 15068 16980 15074 16992
rect 15396 16980 15424 17011
rect 21634 17008 21640 17020
rect 21692 17048 21698 17060
rect 22204 17048 22232 17215
rect 22462 17116 22468 17128
rect 22423 17088 22468 17116
rect 22462 17076 22468 17088
rect 22520 17076 22526 17128
rect 21692 17020 22232 17048
rect 21692 17008 21698 17020
rect 16666 16980 16672 16992
rect 15068 16952 16672 16980
rect 15068 16940 15074 16952
rect 16666 16940 16672 16952
rect 16724 16940 16730 16992
rect 17405 16983 17463 16989
rect 17405 16949 17417 16983
rect 17451 16980 17463 16983
rect 18046 16980 18052 16992
rect 17451 16952 18052 16980
rect 17451 16949 17463 16952
rect 17405 16943 17463 16949
rect 18046 16940 18052 16952
rect 18104 16940 18110 16992
rect 18233 16983 18291 16989
rect 18233 16949 18245 16983
rect 18279 16980 18291 16983
rect 18322 16980 18328 16992
rect 18279 16952 18328 16980
rect 18279 16949 18291 16952
rect 18233 16943 18291 16949
rect 18322 16940 18328 16952
rect 18380 16940 18386 16992
rect 18601 16983 18659 16989
rect 18601 16949 18613 16983
rect 18647 16980 18659 16983
rect 18874 16980 18880 16992
rect 18647 16952 18880 16980
rect 18647 16949 18659 16952
rect 18601 16943 18659 16949
rect 18874 16940 18880 16952
rect 18932 16940 18938 16992
rect 19797 16983 19855 16989
rect 19797 16949 19809 16983
rect 19843 16980 19855 16983
rect 21818 16980 21824 16992
rect 19843 16952 21824 16980
rect 19843 16949 19855 16952
rect 19797 16943 19855 16949
rect 21818 16940 21824 16952
rect 21876 16940 21882 16992
rect 22646 16980 22652 16992
rect 22607 16952 22652 16980
rect 22646 16940 22652 16952
rect 22704 16940 22710 16992
rect 1104 16890 23276 16912
rect 1104 16838 8379 16890
rect 8431 16838 8443 16890
rect 8495 16838 8507 16890
rect 8559 16838 8571 16890
rect 8623 16838 15776 16890
rect 15828 16838 15840 16890
rect 15892 16838 15904 16890
rect 15956 16838 15968 16890
rect 16020 16838 23276 16890
rect 1104 16816 23276 16838
rect 1581 16779 1639 16785
rect 1581 16745 1593 16779
rect 1627 16776 1639 16779
rect 3142 16776 3148 16788
rect 1627 16748 3148 16776
rect 1627 16745 1639 16748
rect 1581 16739 1639 16745
rect 3142 16736 3148 16748
rect 3200 16736 3206 16788
rect 3326 16776 3332 16788
rect 3287 16748 3332 16776
rect 3326 16736 3332 16748
rect 3384 16736 3390 16788
rect 4065 16779 4123 16785
rect 4065 16745 4077 16779
rect 4111 16776 4123 16779
rect 4246 16776 4252 16788
rect 4111 16748 4252 16776
rect 4111 16745 4123 16748
rect 4065 16739 4123 16745
rect 4246 16736 4252 16748
rect 4304 16736 4310 16788
rect 5077 16779 5135 16785
rect 5077 16745 5089 16779
rect 5123 16776 5135 16779
rect 5258 16776 5264 16788
rect 5123 16748 5264 16776
rect 5123 16745 5135 16748
rect 5077 16739 5135 16745
rect 5258 16736 5264 16748
rect 5316 16736 5322 16788
rect 5442 16736 5448 16788
rect 5500 16776 5506 16788
rect 5500 16748 10180 16776
rect 5500 16736 5506 16748
rect 2314 16708 2320 16720
rect 1964 16680 2320 16708
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 1964 16649 1992 16680
rect 2314 16668 2320 16680
rect 2372 16668 2378 16720
rect 2590 16668 2596 16720
rect 2648 16708 2654 16720
rect 3970 16708 3976 16720
rect 2648 16680 3976 16708
rect 2648 16668 2654 16680
rect 3970 16668 3976 16680
rect 4028 16668 4034 16720
rect 4525 16711 4583 16717
rect 4525 16708 4537 16711
rect 4172 16680 4537 16708
rect 1949 16643 2007 16649
rect 1949 16609 1961 16643
rect 1995 16609 2007 16643
rect 1949 16603 2007 16609
rect 2216 16643 2274 16649
rect 2216 16609 2228 16643
rect 2262 16640 2274 16643
rect 2262 16612 3464 16640
rect 2262 16609 2274 16612
rect 2216 16603 2274 16609
rect 3436 16516 3464 16612
rect 4062 16600 4068 16652
rect 4120 16640 4126 16652
rect 4172 16640 4200 16680
rect 4525 16677 4537 16680
rect 4571 16677 4583 16711
rect 4525 16671 4583 16677
rect 4798 16668 4804 16720
rect 4856 16708 4862 16720
rect 7742 16708 7748 16720
rect 4856 16680 7748 16708
rect 4856 16668 4862 16680
rect 7742 16668 7748 16680
rect 7800 16668 7806 16720
rect 7926 16668 7932 16720
rect 7984 16708 7990 16720
rect 8196 16711 8254 16717
rect 8196 16708 8208 16711
rect 7984 16680 8208 16708
rect 7984 16668 7990 16680
rect 8196 16677 8208 16680
rect 8242 16708 8254 16711
rect 9214 16708 9220 16720
rect 8242 16680 9220 16708
rect 8242 16677 8254 16680
rect 8196 16671 8254 16677
rect 9214 16668 9220 16680
rect 9272 16668 9278 16720
rect 9950 16717 9956 16720
rect 9401 16711 9459 16717
rect 9401 16677 9413 16711
rect 9447 16708 9459 16711
rect 9944 16708 9956 16717
rect 9447 16680 9956 16708
rect 9447 16677 9459 16680
rect 9401 16671 9459 16677
rect 9944 16671 9956 16680
rect 9950 16668 9956 16671
rect 10008 16668 10014 16720
rect 10152 16708 10180 16748
rect 10226 16736 10232 16788
rect 10284 16776 10290 16788
rect 10962 16776 10968 16788
rect 10284 16748 10968 16776
rect 10284 16736 10290 16748
rect 10962 16736 10968 16748
rect 11020 16776 11026 16788
rect 11333 16779 11391 16785
rect 11333 16776 11345 16779
rect 11020 16748 11345 16776
rect 11020 16736 11026 16748
rect 11333 16745 11345 16748
rect 11379 16745 11391 16779
rect 13078 16776 13084 16788
rect 13039 16748 13084 16776
rect 11333 16739 11391 16745
rect 13078 16736 13084 16748
rect 13136 16736 13142 16788
rect 13170 16736 13176 16788
rect 13228 16776 13234 16788
rect 13357 16779 13415 16785
rect 13357 16776 13369 16779
rect 13228 16748 13369 16776
rect 13228 16736 13234 16748
rect 13357 16745 13369 16748
rect 13403 16745 13415 16779
rect 13357 16739 13415 16745
rect 13538 16736 13544 16788
rect 13596 16776 13602 16788
rect 13817 16779 13875 16785
rect 13817 16776 13829 16779
rect 13596 16748 13829 16776
rect 13596 16736 13602 16748
rect 13817 16745 13829 16748
rect 13863 16745 13875 16779
rect 14829 16779 14887 16785
rect 14829 16776 14841 16779
rect 13817 16739 13875 16745
rect 14016 16748 14841 16776
rect 10152 16680 11744 16708
rect 4120 16612 4200 16640
rect 4433 16643 4491 16649
rect 4120 16600 4126 16612
rect 4433 16609 4445 16643
rect 4479 16640 4491 16643
rect 4890 16640 4896 16652
rect 4479 16612 4896 16640
rect 4479 16609 4491 16612
rect 4433 16603 4491 16609
rect 4890 16600 4896 16612
rect 4948 16600 4954 16652
rect 5442 16640 5448 16652
rect 5403 16612 5448 16640
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 5994 16640 6000 16652
rect 5552 16612 6000 16640
rect 4338 16532 4344 16584
rect 4396 16572 4402 16584
rect 5552 16581 5580 16612
rect 5994 16600 6000 16612
rect 6052 16600 6058 16652
rect 6178 16600 6184 16652
rect 6236 16640 6242 16652
rect 6529 16643 6587 16649
rect 6529 16640 6541 16643
rect 6236 16612 6541 16640
rect 6236 16600 6242 16612
rect 6529 16609 6541 16612
rect 6575 16640 6587 16643
rect 8938 16640 8944 16652
rect 6575 16612 8944 16640
rect 6575 16609 6587 16612
rect 6529 16603 6587 16609
rect 8938 16600 8944 16612
rect 8996 16600 9002 16652
rect 10226 16640 10232 16652
rect 9048 16612 10232 16640
rect 4617 16575 4675 16581
rect 4617 16572 4629 16575
rect 4396 16544 4629 16572
rect 4396 16532 4402 16544
rect 4617 16541 4629 16544
rect 4663 16541 4675 16575
rect 4617 16535 4675 16541
rect 5537 16575 5595 16581
rect 5537 16541 5549 16575
rect 5583 16541 5595 16575
rect 5537 16535 5595 16541
rect 5629 16575 5687 16581
rect 5629 16541 5641 16575
rect 5675 16541 5687 16575
rect 5629 16535 5687 16541
rect 3418 16464 3424 16516
rect 3476 16504 3482 16516
rect 5644 16504 5672 16535
rect 5718 16532 5724 16584
rect 5776 16572 5782 16584
rect 6273 16575 6331 16581
rect 6273 16572 6285 16575
rect 5776 16544 6285 16572
rect 5776 16532 5782 16544
rect 6273 16541 6285 16544
rect 6319 16541 6331 16575
rect 6273 16535 6331 16541
rect 7929 16575 7987 16581
rect 7929 16541 7941 16575
rect 7975 16541 7987 16575
rect 7929 16535 7987 16541
rect 3476 16476 5672 16504
rect 3476 16464 3482 16476
rect 6288 16436 6316 16535
rect 6454 16436 6460 16448
rect 6288 16408 6460 16436
rect 6454 16396 6460 16408
rect 6512 16396 6518 16448
rect 7466 16396 7472 16448
rect 7524 16436 7530 16448
rect 7653 16439 7711 16445
rect 7653 16436 7665 16439
rect 7524 16408 7665 16436
rect 7524 16396 7530 16408
rect 7653 16405 7665 16408
rect 7699 16405 7711 16439
rect 7944 16436 7972 16535
rect 8938 16464 8944 16516
rect 8996 16504 9002 16516
rect 9048 16504 9076 16612
rect 10226 16600 10232 16612
rect 10284 16600 10290 16652
rect 11330 16600 11336 16652
rect 11388 16640 11394 16652
rect 11517 16643 11575 16649
rect 11517 16640 11529 16643
rect 11388 16612 11529 16640
rect 11388 16600 11394 16612
rect 11517 16609 11529 16612
rect 11563 16609 11575 16643
rect 11716 16640 11744 16680
rect 11882 16668 11888 16720
rect 11940 16717 11946 16720
rect 11940 16711 12004 16717
rect 11940 16677 11958 16711
rect 11992 16677 12004 16711
rect 11940 16671 12004 16677
rect 13725 16711 13783 16717
rect 13725 16677 13737 16711
rect 13771 16708 13783 16711
rect 13906 16708 13912 16720
rect 13771 16680 13912 16708
rect 13771 16677 13783 16680
rect 13725 16671 13783 16677
rect 11940 16668 11946 16671
rect 13906 16668 13912 16680
rect 13964 16668 13970 16720
rect 14016 16640 14044 16748
rect 14829 16745 14841 16748
rect 14875 16745 14887 16779
rect 14829 16739 14887 16745
rect 15654 16736 15660 16788
rect 15712 16776 15718 16788
rect 16669 16779 16727 16785
rect 16669 16776 16681 16779
rect 15712 16748 16681 16776
rect 15712 16736 15718 16748
rect 16669 16745 16681 16748
rect 16715 16745 16727 16779
rect 16669 16739 16727 16745
rect 16945 16779 17003 16785
rect 16945 16745 16957 16779
rect 16991 16776 17003 16779
rect 17681 16779 17739 16785
rect 16991 16748 17356 16776
rect 16991 16745 17003 16748
rect 16945 16739 17003 16745
rect 14918 16708 14924 16720
rect 14568 16680 14924 16708
rect 14568 16649 14596 16680
rect 14918 16668 14924 16680
rect 14976 16708 14982 16720
rect 17328 16708 17356 16748
rect 17681 16745 17693 16779
rect 17727 16776 17739 16779
rect 17954 16776 17960 16788
rect 17727 16748 17960 16776
rect 17727 16745 17739 16748
rect 17681 16739 17739 16745
rect 17954 16736 17960 16748
rect 18012 16736 18018 16788
rect 18966 16736 18972 16788
rect 19024 16776 19030 16788
rect 19153 16779 19211 16785
rect 19153 16776 19165 16779
rect 19024 16748 19165 16776
rect 19024 16736 19030 16748
rect 19153 16745 19165 16748
rect 19199 16745 19211 16779
rect 19153 16739 19211 16745
rect 19978 16736 19984 16788
rect 20036 16776 20042 16788
rect 22646 16776 22652 16788
rect 20036 16748 22652 16776
rect 20036 16736 20042 16748
rect 22646 16736 22652 16748
rect 22704 16736 22710 16788
rect 22741 16779 22799 16785
rect 22741 16745 22753 16779
rect 22787 16745 22799 16779
rect 22741 16739 22799 16745
rect 17862 16708 17868 16720
rect 14976 16680 17172 16708
rect 17328 16680 17868 16708
rect 14976 16668 14982 16680
rect 11716 16612 14044 16640
rect 14553 16643 14611 16649
rect 11517 16603 11575 16609
rect 14553 16609 14565 16643
rect 14599 16609 14611 16643
rect 14553 16603 14611 16609
rect 14645 16643 14703 16649
rect 14645 16609 14657 16643
rect 14691 16640 14703 16643
rect 15378 16640 15384 16652
rect 14691 16612 15384 16640
rect 14691 16609 14703 16612
rect 14645 16603 14703 16609
rect 15378 16600 15384 16612
rect 15436 16600 15442 16652
rect 15556 16643 15614 16649
rect 15556 16609 15568 16643
rect 15602 16640 15614 16643
rect 16482 16640 16488 16652
rect 15602 16612 16488 16640
rect 15602 16609 15614 16612
rect 15556 16603 15614 16609
rect 16482 16600 16488 16612
rect 16540 16600 16546 16652
rect 17144 16649 17172 16680
rect 17862 16668 17868 16680
rect 17920 16668 17926 16720
rect 18040 16711 18098 16717
rect 18040 16677 18052 16711
rect 18086 16708 18098 16711
rect 19702 16708 19708 16720
rect 18086 16680 19708 16708
rect 18086 16677 18098 16680
rect 18040 16671 18098 16677
rect 19702 16668 19708 16680
rect 19760 16668 19766 16720
rect 19886 16668 19892 16720
rect 19944 16708 19950 16720
rect 20254 16708 20260 16720
rect 19944 16680 20260 16708
rect 19944 16668 19950 16680
rect 20254 16668 20260 16680
rect 20312 16668 20318 16720
rect 20806 16668 20812 16720
rect 20864 16708 20870 16720
rect 21634 16717 21640 16720
rect 21269 16711 21327 16717
rect 21269 16708 21281 16711
rect 20864 16680 21281 16708
rect 20864 16668 20870 16680
rect 21269 16677 21281 16680
rect 21315 16677 21327 16711
rect 21628 16708 21640 16717
rect 21595 16680 21640 16708
rect 21269 16671 21327 16677
rect 21628 16671 21640 16680
rect 21634 16668 21640 16671
rect 21692 16668 21698 16720
rect 17129 16643 17187 16649
rect 17129 16609 17141 16643
rect 17175 16609 17187 16643
rect 17129 16603 17187 16609
rect 17221 16643 17279 16649
rect 17221 16609 17233 16643
rect 17267 16640 17279 16643
rect 19242 16640 19248 16652
rect 17267 16612 19248 16640
rect 17267 16609 17279 16612
rect 17221 16603 17279 16609
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 19334 16600 19340 16652
rect 19392 16640 19398 16652
rect 19797 16643 19855 16649
rect 19797 16640 19809 16643
rect 19392 16612 19809 16640
rect 19392 16600 19398 16612
rect 19797 16609 19809 16612
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 20714 16600 20720 16652
rect 20772 16640 20778 16652
rect 22756 16640 22784 16739
rect 20772 16612 22784 16640
rect 20772 16600 20778 16612
rect 9677 16575 9735 16581
rect 9677 16541 9689 16575
rect 9723 16541 9735 16575
rect 11701 16575 11759 16581
rect 11701 16572 11713 16575
rect 9677 16535 9735 16541
rect 10695 16544 11713 16572
rect 8996 16476 9076 16504
rect 9309 16507 9367 16513
rect 8996 16464 9002 16476
rect 9309 16473 9321 16507
rect 9355 16504 9367 16507
rect 9401 16507 9459 16513
rect 9401 16504 9413 16507
rect 9355 16476 9413 16504
rect 9355 16473 9367 16476
rect 9309 16467 9367 16473
rect 9401 16473 9413 16476
rect 9447 16473 9459 16507
rect 9401 16467 9459 16473
rect 9692 16436 9720 16535
rect 9950 16436 9956 16448
rect 7944 16408 9956 16436
rect 7653 16399 7711 16405
rect 9950 16396 9956 16408
rect 10008 16436 10014 16448
rect 10318 16436 10324 16448
rect 10008 16408 10324 16436
rect 10008 16396 10014 16408
rect 10318 16396 10324 16408
rect 10376 16436 10382 16448
rect 10695 16436 10723 16544
rect 11701 16541 11713 16544
rect 11747 16541 11759 16575
rect 11701 16535 11759 16541
rect 12894 16532 12900 16584
rect 12952 16572 12958 16584
rect 13446 16572 13452 16584
rect 12952 16544 13452 16572
rect 12952 16532 12958 16544
rect 13446 16532 13452 16544
rect 13504 16532 13510 16584
rect 13814 16532 13820 16584
rect 13872 16572 13878 16584
rect 13909 16575 13967 16581
rect 13909 16572 13921 16575
rect 13872 16544 13921 16572
rect 13872 16532 13878 16544
rect 13909 16541 13921 16544
rect 13955 16541 13967 16575
rect 13909 16535 13967 16541
rect 15194 16532 15200 16584
rect 15252 16572 15258 16584
rect 15289 16575 15347 16581
rect 15289 16572 15301 16575
rect 15252 16544 15301 16572
rect 15252 16532 15258 16544
rect 15289 16541 15301 16544
rect 15335 16541 15347 16575
rect 15289 16535 15347 16541
rect 17681 16575 17739 16581
rect 17681 16541 17693 16575
rect 17727 16572 17739 16575
rect 17773 16575 17831 16581
rect 17773 16572 17785 16575
rect 17727 16544 17785 16572
rect 17727 16541 17739 16544
rect 17681 16535 17739 16541
rect 17773 16541 17785 16544
rect 17819 16541 17831 16575
rect 17773 16535 17831 16541
rect 18782 16532 18788 16584
rect 18840 16572 18846 16584
rect 19889 16575 19947 16581
rect 19889 16572 19901 16575
rect 18840 16544 19901 16572
rect 18840 16532 18846 16544
rect 19889 16541 19901 16544
rect 19935 16541 19947 16575
rect 19889 16535 19947 16541
rect 19978 16532 19984 16584
rect 20036 16572 20042 16584
rect 20898 16572 20904 16584
rect 20036 16544 20081 16572
rect 20859 16544 20904 16572
rect 20036 16532 20042 16544
rect 20898 16532 20904 16544
rect 20956 16532 20962 16584
rect 21269 16575 21327 16581
rect 21269 16541 21281 16575
rect 21315 16572 21327 16575
rect 21361 16575 21419 16581
rect 21361 16572 21373 16575
rect 21315 16544 21373 16572
rect 21315 16541 21327 16544
rect 21269 16535 21327 16541
rect 21361 16541 21373 16544
rect 21407 16541 21419 16575
rect 21361 16535 21419 16541
rect 11054 16504 11060 16516
rect 10967 16476 11060 16504
rect 11054 16464 11060 16476
rect 11112 16504 11118 16516
rect 17405 16507 17463 16513
rect 11112 16476 11744 16504
rect 11112 16464 11118 16476
rect 10376 16408 10723 16436
rect 11716 16436 11744 16476
rect 13648 16476 14504 16504
rect 13648 16436 13676 16476
rect 11716 16408 13676 16436
rect 10376 16396 10382 16408
rect 14274 16396 14280 16448
rect 14332 16436 14338 16448
rect 14369 16439 14427 16445
rect 14369 16436 14381 16439
rect 14332 16408 14381 16436
rect 14332 16396 14338 16408
rect 14369 16405 14381 16408
rect 14415 16405 14427 16439
rect 14476 16436 14504 16476
rect 17405 16473 17417 16507
rect 17451 16504 17463 16507
rect 17494 16504 17500 16516
rect 17451 16476 17500 16504
rect 17451 16473 17463 16476
rect 17405 16467 17463 16473
rect 17494 16464 17500 16476
rect 17552 16464 17558 16516
rect 18414 16436 18420 16448
rect 14476 16408 18420 16436
rect 14369 16399 14427 16405
rect 18414 16396 18420 16408
rect 18472 16396 18478 16448
rect 19429 16439 19487 16445
rect 19429 16405 19441 16439
rect 19475 16436 19487 16439
rect 20254 16436 20260 16448
rect 19475 16408 20260 16436
rect 19475 16405 19487 16408
rect 19429 16399 19487 16405
rect 20254 16396 20260 16408
rect 20312 16396 20318 16448
rect 1104 16346 23276 16368
rect 1104 16294 4680 16346
rect 4732 16294 4744 16346
rect 4796 16294 4808 16346
rect 4860 16294 4872 16346
rect 4924 16294 12078 16346
rect 12130 16294 12142 16346
rect 12194 16294 12206 16346
rect 12258 16294 12270 16346
rect 12322 16294 19475 16346
rect 19527 16294 19539 16346
rect 19591 16294 19603 16346
rect 19655 16294 19667 16346
rect 19719 16294 23276 16346
rect 1104 16272 23276 16294
rect 1673 16235 1731 16241
rect 1673 16201 1685 16235
rect 1719 16232 1731 16235
rect 2774 16232 2780 16244
rect 1719 16204 2780 16232
rect 1719 16201 1731 16204
rect 1673 16195 1731 16201
rect 2774 16192 2780 16204
rect 2832 16192 2838 16244
rect 3418 16232 3424 16244
rect 3379 16204 3424 16232
rect 3418 16192 3424 16204
rect 3476 16192 3482 16244
rect 5902 16232 5908 16244
rect 3988 16204 5908 16232
rect 1486 16028 1492 16040
rect 1447 16000 1492 16028
rect 1486 15988 1492 16000
rect 1544 15988 1550 16040
rect 1854 15988 1860 16040
rect 1912 16028 1918 16040
rect 3988 16037 4016 16204
rect 5902 16192 5908 16204
rect 5960 16192 5966 16244
rect 6822 16192 6828 16244
rect 6880 16232 6886 16244
rect 8849 16235 8907 16241
rect 8849 16232 8861 16235
rect 6880 16204 8861 16232
rect 6880 16192 6886 16204
rect 8849 16201 8861 16204
rect 8895 16232 8907 16235
rect 10410 16232 10416 16244
rect 8895 16204 10416 16232
rect 8895 16201 8907 16204
rect 8849 16195 8907 16201
rect 10410 16192 10416 16204
rect 10468 16192 10474 16244
rect 10686 16192 10692 16244
rect 10744 16232 10750 16244
rect 10744 16204 11836 16232
rect 10744 16192 10750 16204
rect 6089 16167 6147 16173
rect 6089 16133 6101 16167
rect 6135 16164 6147 16167
rect 6641 16167 6699 16173
rect 6641 16164 6653 16167
rect 6135 16136 6653 16164
rect 6135 16133 6147 16136
rect 6089 16127 6147 16133
rect 6641 16133 6653 16136
rect 6687 16133 6699 16167
rect 6641 16127 6699 16133
rect 10781 16167 10839 16173
rect 10781 16133 10793 16167
rect 10827 16164 10839 16167
rect 10827 16136 11560 16164
rect 10827 16133 10839 16136
rect 10781 16127 10839 16133
rect 4065 16099 4123 16105
rect 4065 16065 4077 16099
rect 4111 16096 4123 16099
rect 4246 16096 4252 16108
rect 4111 16068 4252 16096
rect 4111 16065 4123 16068
rect 4065 16059 4123 16065
rect 4246 16056 4252 16068
rect 4304 16056 4310 16108
rect 4522 16056 4528 16108
rect 4580 16096 4586 16108
rect 4801 16099 4859 16105
rect 4580 16068 4625 16096
rect 4580 16056 4586 16068
rect 4801 16065 4813 16099
rect 4847 16096 4859 16099
rect 5534 16096 5540 16108
rect 4847 16068 5540 16096
rect 4847 16065 4859 16068
rect 4801 16059 4859 16065
rect 5534 16056 5540 16068
rect 5592 16056 5598 16108
rect 5718 16056 5724 16108
rect 5776 16096 5782 16108
rect 6270 16096 6276 16108
rect 5776 16068 6276 16096
rect 5776 16056 5782 16068
rect 6270 16056 6276 16068
rect 6328 16096 6334 16108
rect 7288 16099 7346 16105
rect 7288 16096 7300 16099
rect 6328 16068 7300 16096
rect 6328 16056 6334 16068
rect 7288 16065 7300 16068
rect 7334 16065 7346 16099
rect 7288 16059 7346 16065
rect 7374 16056 7380 16108
rect 7432 16096 7438 16108
rect 9306 16105 9312 16108
rect 9264 16099 9312 16105
rect 9264 16096 9276 16099
rect 7432 16068 9276 16096
rect 7432 16056 7438 16068
rect 9264 16065 9276 16068
rect 9310 16065 9312 16099
rect 9264 16059 9312 16065
rect 9306 16056 9312 16059
rect 9364 16096 9370 16108
rect 9447 16099 9505 16105
rect 9364 16068 9412 16096
rect 9364 16056 9370 16068
rect 9447 16065 9459 16099
rect 9493 16096 9505 16099
rect 10870 16096 10876 16108
rect 9493 16068 10876 16096
rect 9493 16065 9505 16068
rect 9447 16059 9505 16065
rect 10870 16056 10876 16068
rect 10928 16056 10934 16108
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1912 16000 2053 16028
rect 1912 15988 1918 16000
rect 2041 15997 2053 16000
rect 2087 16028 2099 16031
rect 3973 16031 4031 16037
rect 2087 16000 3832 16028
rect 2087 15997 2099 16000
rect 2041 15991 2099 15997
rect 2308 15963 2366 15969
rect 2308 15929 2320 15963
rect 2354 15960 2366 15963
rect 2682 15960 2688 15972
rect 2354 15932 2688 15960
rect 2354 15929 2366 15932
rect 2308 15923 2366 15929
rect 2682 15920 2688 15932
rect 2740 15920 2746 15972
rect 3804 15901 3832 16000
rect 3973 15997 3985 16031
rect 4019 15997 4031 16031
rect 3973 15991 4031 15997
rect 4890 15988 4896 16040
rect 4948 16028 4954 16040
rect 6089 16031 6147 16037
rect 6089 16028 6101 16031
rect 4948 16000 6101 16028
rect 4948 15988 4954 16000
rect 6089 15997 6101 16000
rect 6135 15997 6147 16031
rect 6089 15991 6147 15997
rect 6181 16031 6239 16037
rect 6181 15997 6193 16031
rect 6227 16028 6239 16031
rect 6638 16028 6644 16040
rect 6227 16000 6644 16028
rect 6227 15997 6239 16000
rect 6181 15991 6239 15997
rect 6638 15988 6644 16000
rect 6696 15988 6702 16040
rect 6822 16028 6828 16040
rect 6783 16000 6828 16028
rect 6822 15988 6828 16000
rect 6880 15988 6886 16040
rect 7561 16031 7619 16037
rect 7561 16028 7573 16031
rect 6932 16000 7573 16028
rect 6730 15920 6736 15972
rect 6788 15960 6794 15972
rect 6932 15960 6960 16000
rect 7561 15997 7573 16000
rect 7607 15997 7619 16031
rect 7561 15991 7619 15997
rect 8849 16031 8907 16037
rect 8849 15997 8861 16031
rect 8895 16028 8907 16031
rect 8941 16031 8999 16037
rect 8941 16028 8953 16031
rect 8895 16000 8953 16028
rect 8895 15997 8907 16000
rect 8849 15991 8907 15997
rect 8941 15997 8953 16000
rect 8987 15997 8999 16031
rect 9674 16028 9680 16040
rect 8941 15991 8999 15997
rect 9048 16000 9680 16028
rect 9048 15960 9076 16000
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 10778 15988 10784 16040
rect 10836 16028 10842 16040
rect 11238 16028 11244 16040
rect 10836 16000 11244 16028
rect 10836 15988 10842 16000
rect 11238 15988 11244 16000
rect 11296 16028 11302 16040
rect 11532 16037 11560 16136
rect 11606 16056 11612 16108
rect 11664 16096 11670 16108
rect 11808 16096 11836 16204
rect 11974 16192 11980 16244
rect 12032 16232 12038 16244
rect 12032 16204 13032 16232
rect 12032 16192 12038 16204
rect 13004 16105 13032 16204
rect 13262 16192 13268 16244
rect 13320 16232 13326 16244
rect 16945 16235 17003 16241
rect 16945 16232 16957 16235
rect 13320 16204 16957 16232
rect 13320 16192 13326 16204
rect 16945 16201 16957 16204
rect 16991 16201 17003 16235
rect 16945 16195 17003 16201
rect 17497 16235 17555 16241
rect 17497 16201 17509 16235
rect 17543 16232 17555 16235
rect 17586 16232 17592 16244
rect 17543 16204 17592 16232
rect 17543 16201 17555 16204
rect 17497 16195 17555 16201
rect 17586 16192 17592 16204
rect 17644 16192 17650 16244
rect 19429 16235 19487 16241
rect 17696 16204 19012 16232
rect 16574 16124 16580 16176
rect 16632 16164 16638 16176
rect 17696 16164 17724 16204
rect 16632 16136 17724 16164
rect 18984 16164 19012 16204
rect 19429 16201 19441 16235
rect 19475 16232 19487 16235
rect 19794 16232 19800 16244
rect 19475 16204 19800 16232
rect 19475 16201 19487 16204
rect 19429 16195 19487 16201
rect 19794 16192 19800 16204
rect 19852 16192 19858 16244
rect 21542 16232 21548 16244
rect 19904 16204 20852 16232
rect 21503 16204 21548 16232
rect 19904 16164 19932 16204
rect 18984 16136 19932 16164
rect 20824 16164 20852 16204
rect 21542 16192 21548 16204
rect 21600 16192 21606 16244
rect 22738 16164 22744 16176
rect 20824 16136 22744 16164
rect 16632 16124 16638 16136
rect 22738 16124 22744 16136
rect 22796 16124 22802 16176
rect 12989 16099 13047 16105
rect 11664 16068 11709 16096
rect 11808 16068 12388 16096
rect 11664 16056 11670 16068
rect 11425 16031 11483 16037
rect 11425 16028 11437 16031
rect 11296 16000 11437 16028
rect 11296 15988 11302 16000
rect 11425 15997 11437 16000
rect 11471 15997 11483 16031
rect 11425 15991 11483 15997
rect 11517 16031 11575 16037
rect 11517 15997 11529 16031
rect 11563 16028 11575 16031
rect 11790 16028 11796 16040
rect 11563 16000 11796 16028
rect 11563 15997 11575 16000
rect 11517 15991 11575 15997
rect 11790 15988 11796 16000
rect 11848 15988 11854 16040
rect 11974 16028 11980 16040
rect 11935 16000 11980 16028
rect 11974 15988 11980 16000
rect 12032 15988 12038 16040
rect 12360 16028 12388 16068
rect 12989 16065 13001 16099
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 13078 16056 13084 16108
rect 13136 16096 13142 16108
rect 13357 16099 13415 16105
rect 13357 16096 13369 16099
rect 13136 16068 13369 16096
rect 13136 16056 13142 16068
rect 13357 16065 13369 16068
rect 13403 16065 13415 16099
rect 13814 16096 13820 16108
rect 13778 16068 13820 16096
rect 13357 16059 13415 16065
rect 13814 16056 13820 16068
rect 13872 16056 13878 16108
rect 15194 16056 15200 16108
rect 15252 16096 15258 16108
rect 15565 16099 15623 16105
rect 15565 16096 15577 16099
rect 15252 16068 15577 16096
rect 15252 16056 15258 16068
rect 15565 16065 15577 16068
rect 15611 16065 15623 16099
rect 15565 16059 15623 16065
rect 22002 16056 22008 16108
rect 22060 16096 22066 16108
rect 22097 16099 22155 16105
rect 22097 16096 22109 16099
rect 22060 16068 22109 16096
rect 22060 16056 22066 16068
rect 22097 16065 22109 16068
rect 22143 16065 22155 16099
rect 22097 16059 22155 16065
rect 22370 16056 22376 16108
rect 22428 16096 22434 16108
rect 22557 16099 22615 16105
rect 22557 16096 22569 16099
rect 22428 16068 22569 16096
rect 22428 16056 22434 16068
rect 22557 16065 22569 16068
rect 22603 16065 22615 16099
rect 22557 16059 22615 16065
rect 13680 16031 13738 16037
rect 13680 16028 13692 16031
rect 12360 16000 13692 16028
rect 13680 15997 13692 16000
rect 13726 16028 13738 16031
rect 13998 16028 14004 16040
rect 13726 16000 14004 16028
rect 13726 15997 13738 16000
rect 13680 15991 13738 15997
rect 13998 15988 14004 16000
rect 14056 15988 14062 16040
rect 14090 15988 14096 16040
rect 14148 16028 14154 16040
rect 14148 16000 14193 16028
rect 14148 15988 14154 16000
rect 16850 15988 16856 16040
rect 16908 16028 16914 16040
rect 17313 16031 17371 16037
rect 17313 16028 17325 16031
rect 16908 16000 17325 16028
rect 16908 15988 16914 16000
rect 17313 15997 17325 16000
rect 17359 15997 17371 16031
rect 17313 15991 17371 15997
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 16028 18107 16031
rect 18690 16028 18696 16040
rect 18095 16000 18696 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 12897 15963 12955 15969
rect 12897 15960 12909 15963
rect 6788 15932 6960 15960
rect 8680 15932 9076 15960
rect 11072 15932 12909 15960
rect 6788 15920 6794 15932
rect 3789 15895 3847 15901
rect 3789 15861 3801 15895
rect 3835 15892 3847 15895
rect 4338 15892 4344 15904
rect 3835 15864 4344 15892
rect 3835 15861 3847 15864
rect 3789 15855 3847 15861
rect 4338 15852 4344 15864
rect 4396 15852 4402 15904
rect 4531 15895 4589 15901
rect 4531 15861 4543 15895
rect 4577 15892 4589 15895
rect 4890 15892 4896 15904
rect 4577 15864 4896 15892
rect 4577 15861 4589 15864
rect 4531 15855 4589 15861
rect 4890 15852 4896 15864
rect 4948 15852 4954 15904
rect 5166 15852 5172 15904
rect 5224 15892 5230 15904
rect 5905 15895 5963 15901
rect 5905 15892 5917 15895
rect 5224 15864 5917 15892
rect 5224 15852 5230 15864
rect 5905 15861 5917 15864
rect 5951 15861 5963 15895
rect 5905 15855 5963 15861
rect 6365 15895 6423 15901
rect 6365 15861 6377 15895
rect 6411 15892 6423 15895
rect 6546 15892 6552 15904
rect 6411 15864 6552 15892
rect 6411 15861 6423 15864
rect 6365 15855 6423 15861
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 6641 15895 6699 15901
rect 6641 15861 6653 15895
rect 6687 15892 6699 15895
rect 7282 15892 7288 15904
rect 7340 15901 7346 15904
rect 6687 15864 7288 15892
rect 6687 15861 6699 15864
rect 6641 15855 6699 15861
rect 7282 15852 7288 15864
rect 7340 15855 7349 15901
rect 7340 15852 7346 15855
rect 8202 15852 8208 15904
rect 8260 15892 8266 15904
rect 8680 15901 8708 15932
rect 8665 15895 8723 15901
rect 8665 15892 8677 15895
rect 8260 15864 8677 15892
rect 8260 15852 8266 15864
rect 8665 15861 8677 15864
rect 8711 15861 8723 15895
rect 8665 15855 8723 15861
rect 9306 15852 9312 15904
rect 9364 15892 9370 15904
rect 10686 15892 10692 15904
rect 9364 15864 10692 15892
rect 9364 15852 9370 15864
rect 10686 15852 10692 15864
rect 10744 15852 10750 15904
rect 11072 15901 11100 15932
rect 12897 15929 12909 15932
rect 12943 15929 12955 15963
rect 12897 15923 12955 15929
rect 15654 15920 15660 15972
rect 15712 15960 15718 15972
rect 15810 15963 15868 15969
rect 15810 15960 15822 15963
rect 15712 15932 15822 15960
rect 15712 15920 15718 15932
rect 15810 15929 15822 15932
rect 15856 15929 15868 15963
rect 15810 15923 15868 15929
rect 11057 15895 11115 15901
rect 11057 15861 11069 15895
rect 11103 15861 11115 15895
rect 11057 15855 11115 15861
rect 11238 15852 11244 15904
rect 11296 15892 11302 15904
rect 12066 15892 12072 15904
rect 11296 15864 12072 15892
rect 11296 15852 11302 15864
rect 12066 15852 12072 15864
rect 12124 15852 12130 15904
rect 12161 15895 12219 15901
rect 12161 15861 12173 15895
rect 12207 15892 12219 15895
rect 12342 15892 12348 15904
rect 12207 15864 12348 15892
rect 12207 15861 12219 15864
rect 12161 15855 12219 15861
rect 12342 15852 12348 15864
rect 12400 15852 12406 15904
rect 12437 15895 12495 15901
rect 12437 15861 12449 15895
rect 12483 15892 12495 15895
rect 12618 15892 12624 15904
rect 12483 15864 12624 15892
rect 12483 15861 12495 15864
rect 12437 15855 12495 15861
rect 12618 15852 12624 15864
rect 12676 15852 12682 15904
rect 12802 15892 12808 15904
rect 12763 15864 12808 15892
rect 12802 15852 12808 15864
rect 12860 15852 12866 15904
rect 13446 15852 13452 15904
rect 13504 15892 13510 15904
rect 13906 15892 13912 15904
rect 13504 15864 13912 15892
rect 13504 15852 13510 15864
rect 13906 15852 13912 15864
rect 13964 15852 13970 15904
rect 15194 15892 15200 15904
rect 15155 15864 15200 15892
rect 15194 15852 15200 15864
rect 15252 15892 15258 15904
rect 16114 15892 16120 15904
rect 15252 15864 16120 15892
rect 15252 15852 15258 15864
rect 16114 15852 16120 15864
rect 16172 15852 16178 15904
rect 17328 15892 17356 15991
rect 18690 15988 18696 16000
rect 18748 16028 18754 16040
rect 19889 16031 19947 16037
rect 19889 16028 19901 16031
rect 18748 16000 19901 16028
rect 18748 15988 18754 16000
rect 19889 15997 19901 16000
rect 19935 15997 19947 16031
rect 19889 15991 19947 15997
rect 20156 16031 20214 16037
rect 20156 15997 20168 16031
rect 20202 16028 20214 16031
rect 20714 16028 20720 16040
rect 20202 16000 20720 16028
rect 20202 15997 20214 16000
rect 20156 15991 20214 15997
rect 18316 15963 18374 15969
rect 18316 15929 18328 15963
rect 18362 15960 18374 15963
rect 19334 15960 19340 15972
rect 18362 15932 19340 15960
rect 18362 15929 18374 15932
rect 18316 15923 18374 15929
rect 19334 15920 19340 15932
rect 19392 15920 19398 15972
rect 19904 15960 19932 15991
rect 20714 15988 20720 16000
rect 20772 15988 20778 16040
rect 20898 15988 20904 16040
rect 20956 16028 20962 16040
rect 21913 16031 21971 16037
rect 21913 16028 21925 16031
rect 20956 16000 21925 16028
rect 20956 15988 20962 16000
rect 21913 15997 21925 16000
rect 21959 15997 21971 16031
rect 21913 15991 21971 15997
rect 19904 15932 20944 15960
rect 20916 15904 20944 15932
rect 21818 15920 21824 15972
rect 21876 15960 21882 15972
rect 22005 15963 22063 15969
rect 22005 15960 22017 15963
rect 21876 15932 22017 15960
rect 21876 15920 21882 15932
rect 22005 15929 22017 15932
rect 22051 15929 22063 15963
rect 22005 15923 22063 15929
rect 20162 15892 20168 15904
rect 17328 15864 20168 15892
rect 20162 15852 20168 15864
rect 20220 15852 20226 15904
rect 20898 15852 20904 15904
rect 20956 15852 20962 15904
rect 21266 15892 21272 15904
rect 21227 15864 21272 15892
rect 21266 15852 21272 15864
rect 21324 15852 21330 15904
rect 1104 15802 23276 15824
rect 1104 15750 8379 15802
rect 8431 15750 8443 15802
rect 8495 15750 8507 15802
rect 8559 15750 8571 15802
rect 8623 15750 15776 15802
rect 15828 15750 15840 15802
rect 15892 15750 15904 15802
rect 15956 15750 15968 15802
rect 16020 15750 23276 15802
rect 1104 15728 23276 15750
rect 7190 15648 7196 15700
rect 7248 15688 7254 15700
rect 8757 15691 8815 15697
rect 8757 15688 8769 15691
rect 7248 15660 8769 15688
rect 7248 15648 7254 15660
rect 8757 15657 8769 15660
rect 8803 15657 8815 15691
rect 8757 15651 8815 15657
rect 9217 15691 9275 15697
rect 9217 15657 9229 15691
rect 9263 15688 9275 15691
rect 9493 15691 9551 15697
rect 9493 15688 9505 15691
rect 9263 15660 9505 15688
rect 9263 15657 9275 15660
rect 9217 15651 9275 15657
rect 9493 15657 9505 15660
rect 9539 15657 9551 15691
rect 9493 15651 9551 15657
rect 9677 15691 9735 15697
rect 9677 15657 9689 15691
rect 9723 15688 9735 15691
rect 10778 15688 10784 15700
rect 9723 15660 10784 15688
rect 9723 15657 9735 15660
rect 9677 15651 9735 15657
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 10870 15648 10876 15700
rect 10928 15688 10934 15700
rect 12710 15688 12716 15700
rect 10928 15660 12716 15688
rect 10928 15648 10934 15660
rect 12710 15648 12716 15660
rect 12768 15648 12774 15700
rect 12989 15691 13047 15697
rect 12989 15657 13001 15691
rect 13035 15688 13047 15691
rect 13078 15688 13084 15700
rect 13035 15660 13084 15688
rect 13035 15657 13047 15660
rect 12989 15651 13047 15657
rect 13078 15648 13084 15660
rect 13136 15648 13142 15700
rect 14918 15688 14924 15700
rect 14879 15660 14924 15688
rect 14918 15648 14924 15660
rect 14976 15648 14982 15700
rect 15102 15648 15108 15700
rect 15160 15688 15166 15700
rect 19334 15688 19340 15700
rect 15160 15660 18920 15688
rect 19295 15660 19340 15688
rect 15160 15648 15166 15660
rect 1854 15620 1860 15632
rect 1504 15592 1860 15620
rect 1504 15561 1532 15592
rect 1854 15580 1860 15592
rect 1912 15580 1918 15632
rect 3970 15580 3976 15632
rect 4028 15620 4034 15632
rect 4246 15620 4252 15632
rect 4028 15592 4252 15620
rect 4028 15580 4034 15592
rect 4246 15580 4252 15592
rect 4304 15620 4310 15632
rect 4304 15592 5028 15620
rect 4304 15580 4310 15592
rect 1489 15555 1547 15561
rect 1489 15521 1501 15555
rect 1535 15521 1547 15555
rect 1489 15515 1547 15521
rect 1756 15555 1814 15561
rect 1756 15521 1768 15555
rect 1802 15552 1814 15555
rect 2958 15552 2964 15564
rect 1802 15524 2964 15552
rect 1802 15521 1814 15524
rect 1756 15515 1814 15521
rect 2958 15512 2964 15524
rect 3016 15512 3022 15564
rect 3142 15552 3148 15564
rect 3103 15524 3148 15552
rect 3142 15512 3148 15524
rect 3200 15512 3206 15564
rect 4430 15552 4436 15564
rect 4391 15524 4436 15552
rect 4430 15512 4436 15524
rect 4488 15512 4494 15564
rect 5000 15561 5028 15592
rect 6822 15580 6828 15632
rect 6880 15580 6886 15632
rect 7368 15623 7426 15629
rect 7368 15589 7380 15623
rect 7414 15620 7426 15623
rect 7466 15620 7472 15632
rect 7414 15592 7472 15620
rect 7414 15589 7426 15592
rect 7368 15583 7426 15589
rect 7466 15580 7472 15592
rect 7524 15580 7530 15632
rect 10502 15620 10508 15632
rect 9048 15592 10508 15620
rect 4985 15555 5043 15561
rect 4985 15521 4997 15555
rect 5031 15552 5043 15555
rect 5721 15555 5779 15561
rect 5031 15524 5672 15552
rect 5031 15521 5043 15524
rect 4985 15515 5043 15521
rect 3326 15484 3332 15496
rect 3287 15456 3332 15484
rect 3326 15444 3332 15456
rect 3384 15444 3390 15496
rect 5308 15487 5366 15493
rect 5308 15484 5320 15487
rect 5000 15456 5320 15484
rect 5000 15428 5028 15456
rect 5308 15453 5320 15456
rect 5354 15453 5366 15487
rect 5442 15484 5448 15496
rect 5406 15456 5448 15484
rect 5308 15447 5366 15453
rect 5442 15444 5448 15456
rect 5500 15444 5506 15496
rect 5644 15484 5672 15524
rect 5721 15521 5733 15555
rect 5767 15552 5779 15555
rect 5994 15552 6000 15564
rect 5767 15524 6000 15552
rect 5767 15521 5779 15524
rect 5721 15515 5779 15521
rect 5994 15512 6000 15524
rect 6052 15512 6058 15564
rect 6840 15552 6868 15580
rect 6095 15524 6868 15552
rect 6095 15484 6123 15524
rect 8662 15512 8668 15564
rect 8720 15552 8726 15564
rect 8938 15552 8944 15564
rect 8720 15524 8944 15552
rect 8720 15512 8726 15524
rect 8938 15512 8944 15524
rect 8996 15512 9002 15564
rect 9048 15561 9076 15592
rect 10502 15580 10508 15592
rect 10560 15580 10566 15632
rect 10686 15580 10692 15632
rect 10744 15620 10750 15632
rect 10744 15592 11100 15620
rect 10744 15580 10750 15592
rect 9033 15555 9091 15561
rect 9033 15521 9045 15555
rect 9079 15521 9091 15555
rect 9033 15515 9091 15521
rect 9122 15512 9128 15564
rect 9180 15552 9186 15564
rect 10045 15555 10103 15561
rect 10045 15552 10057 15555
rect 9180 15524 9260 15552
rect 9180 15512 9186 15524
rect 5644 15456 6123 15484
rect 6454 15444 6460 15496
rect 6512 15484 6518 15496
rect 6822 15484 6828 15496
rect 6512 15456 6828 15484
rect 6512 15444 6518 15456
rect 6822 15444 6828 15456
rect 6880 15484 6886 15496
rect 7101 15487 7159 15493
rect 7101 15484 7113 15487
rect 6880 15456 7113 15484
rect 6880 15444 6886 15456
rect 7101 15453 7113 15456
rect 7147 15453 7159 15487
rect 7101 15447 7159 15453
rect 4982 15376 4988 15428
rect 5040 15376 5046 15428
rect 9232 15360 9260 15524
rect 9324 15524 10057 15552
rect 9324 15360 9352 15524
rect 10045 15521 10057 15524
rect 10091 15521 10103 15555
rect 10962 15552 10968 15564
rect 10923 15524 10968 15552
rect 10045 15515 10103 15521
rect 10962 15512 10968 15524
rect 11020 15512 11026 15564
rect 11072 15552 11100 15592
rect 13998 15580 14004 15632
rect 14056 15620 14062 15632
rect 14056 15592 15415 15620
rect 14056 15580 14062 15592
rect 11380 15555 11438 15561
rect 11380 15552 11392 15555
rect 11072 15524 11392 15552
rect 11380 15521 11392 15524
rect 11426 15521 11438 15555
rect 11790 15552 11796 15564
rect 11751 15524 11796 15552
rect 11380 15515 11438 15521
rect 11790 15512 11796 15524
rect 11848 15512 11854 15564
rect 12894 15512 12900 15564
rect 12952 15552 12958 15564
rect 13262 15552 13268 15564
rect 12952 15524 13268 15552
rect 12952 15512 12958 15524
rect 13262 15512 13268 15524
rect 13320 15552 13326 15564
rect 13429 15555 13487 15561
rect 13429 15552 13441 15555
rect 13320 15524 13441 15552
rect 13320 15512 13326 15524
rect 13429 15521 13441 15524
rect 13475 15521 13487 15555
rect 13429 15515 13487 15521
rect 13906 15512 13912 15564
rect 13964 15552 13970 15564
rect 15102 15552 15108 15564
rect 13964 15524 14228 15552
rect 15063 15524 15108 15552
rect 13964 15512 13970 15524
rect 9766 15444 9772 15496
rect 9824 15484 9830 15496
rect 10137 15487 10195 15493
rect 10137 15484 10149 15487
rect 9824 15456 10149 15484
rect 9824 15444 9830 15456
rect 10137 15453 10149 15456
rect 10183 15453 10195 15487
rect 10137 15447 10195 15453
rect 10226 15444 10232 15496
rect 10284 15484 10290 15496
rect 10284 15456 10329 15484
rect 10284 15444 10290 15456
rect 10410 15444 10416 15496
rect 10468 15484 10474 15496
rect 11057 15487 11115 15493
rect 11057 15484 11069 15487
rect 10468 15456 11069 15484
rect 10468 15444 10474 15456
rect 11057 15453 11069 15456
rect 11103 15453 11115 15487
rect 11057 15447 11115 15453
rect 11563 15487 11621 15493
rect 11563 15453 11575 15487
rect 11609 15484 11621 15487
rect 12434 15484 12440 15496
rect 11609 15456 12440 15484
rect 11609 15453 11621 15456
rect 11563 15447 11621 15453
rect 2682 15308 2688 15360
rect 2740 15348 2746 15360
rect 2869 15351 2927 15357
rect 2869 15348 2881 15351
rect 2740 15320 2881 15348
rect 2740 15308 2746 15320
rect 2869 15317 2881 15320
rect 2915 15317 2927 15351
rect 2869 15311 2927 15317
rect 4617 15351 4675 15357
rect 4617 15317 4629 15351
rect 4663 15348 4675 15351
rect 5258 15348 5264 15360
rect 4663 15320 5264 15348
rect 4663 15317 4675 15320
rect 4617 15311 4675 15317
rect 5258 15308 5264 15320
rect 5316 15308 5322 15360
rect 5902 15308 5908 15360
rect 5960 15348 5966 15360
rect 6730 15348 6736 15360
rect 5960 15320 6736 15348
rect 5960 15308 5966 15320
rect 6730 15308 6736 15320
rect 6788 15348 6794 15360
rect 6825 15351 6883 15357
rect 6825 15348 6837 15351
rect 6788 15320 6837 15348
rect 6788 15308 6794 15320
rect 6825 15317 6837 15320
rect 6871 15317 6883 15351
rect 6825 15311 6883 15317
rect 7098 15308 7104 15360
rect 7156 15348 7162 15360
rect 8481 15351 8539 15357
rect 8481 15348 8493 15351
rect 7156 15320 8493 15348
rect 7156 15308 7162 15320
rect 8481 15317 8493 15320
rect 8527 15317 8539 15351
rect 8481 15311 8539 15317
rect 9214 15308 9220 15360
rect 9272 15308 9278 15360
rect 9306 15308 9312 15360
rect 9364 15308 9370 15360
rect 9493 15351 9551 15357
rect 9493 15317 9505 15351
rect 9539 15348 9551 15351
rect 10594 15348 10600 15360
rect 9539 15320 10600 15348
rect 9539 15317 9551 15320
rect 9493 15311 9551 15317
rect 10594 15308 10600 15320
rect 10652 15308 10658 15360
rect 10778 15348 10784 15360
rect 10739 15320 10784 15348
rect 10778 15308 10784 15320
rect 10836 15308 10842 15360
rect 10870 15308 10876 15360
rect 10928 15348 10934 15360
rect 11072 15348 11100 15447
rect 12434 15444 12440 15456
rect 12492 15484 12498 15496
rect 13078 15484 13084 15496
rect 12492 15456 13084 15484
rect 12492 15444 12498 15456
rect 13078 15444 13084 15456
rect 13136 15444 13142 15496
rect 13173 15487 13231 15493
rect 13173 15453 13185 15487
rect 13219 15453 13231 15487
rect 13173 15447 13231 15453
rect 12989 15419 13047 15425
rect 12989 15416 13001 15419
rect 12452 15388 13001 15416
rect 12452 15348 12480 15388
rect 12989 15385 13001 15388
rect 13035 15385 13047 15419
rect 12989 15379 13047 15385
rect 10928 15320 12480 15348
rect 10928 15308 10934 15320
rect 12618 15308 12624 15360
rect 12676 15348 12682 15360
rect 12897 15351 12955 15357
rect 12897 15348 12909 15351
rect 12676 15320 12909 15348
rect 12676 15308 12682 15320
rect 12897 15317 12909 15320
rect 12943 15317 12955 15351
rect 13188 15348 13216 15447
rect 14200 15416 14228 15524
rect 15102 15512 15108 15524
rect 15160 15512 15166 15564
rect 15289 15555 15347 15561
rect 15289 15552 15301 15555
rect 15212 15524 15301 15552
rect 14734 15444 14740 15496
rect 14792 15484 14798 15496
rect 15212 15484 15240 15524
rect 15289 15521 15301 15524
rect 15335 15521 15347 15555
rect 15387 15552 15415 15592
rect 17954 15580 17960 15632
rect 18012 15620 18018 15632
rect 18224 15623 18282 15629
rect 18224 15620 18236 15623
rect 18012 15592 18236 15620
rect 18012 15580 18018 15592
rect 18224 15589 18236 15592
rect 18270 15620 18282 15623
rect 18782 15620 18788 15632
rect 18270 15592 18788 15620
rect 18270 15589 18282 15592
rect 18224 15583 18282 15589
rect 18782 15580 18788 15592
rect 18840 15580 18846 15632
rect 18892 15620 18920 15660
rect 19334 15648 19340 15660
rect 19392 15648 19398 15700
rect 20162 15648 20168 15700
rect 20220 15688 20226 15700
rect 20257 15691 20315 15697
rect 20257 15688 20269 15691
rect 20220 15660 20269 15688
rect 20220 15648 20226 15660
rect 20257 15657 20269 15660
rect 20303 15688 20315 15691
rect 20714 15688 20720 15700
rect 20303 15660 20720 15688
rect 20303 15657 20315 15660
rect 20257 15651 20315 15657
rect 20714 15648 20720 15660
rect 20772 15648 20778 15700
rect 19886 15620 19892 15632
rect 18892 15592 19892 15620
rect 19886 15580 19892 15592
rect 19944 15580 19950 15632
rect 21168 15623 21226 15629
rect 21168 15589 21180 15623
rect 21214 15620 21226 15623
rect 21266 15620 21272 15632
rect 21214 15592 21272 15620
rect 21214 15589 21226 15592
rect 21168 15583 21226 15589
rect 15612 15555 15670 15561
rect 15612 15552 15624 15555
rect 15387 15524 15624 15552
rect 15289 15515 15347 15521
rect 15612 15521 15624 15524
rect 15658 15552 15670 15555
rect 15838 15552 15844 15564
rect 15658 15524 15844 15552
rect 15658 15521 15670 15524
rect 15612 15515 15670 15521
rect 15838 15512 15844 15524
rect 15896 15512 15902 15564
rect 16025 15555 16083 15561
rect 16025 15521 16037 15555
rect 16071 15552 16083 15555
rect 16114 15552 16120 15564
rect 16071 15524 16120 15552
rect 16071 15521 16083 15524
rect 16025 15515 16083 15521
rect 16114 15512 16120 15524
rect 16172 15512 16178 15564
rect 17405 15555 17463 15561
rect 17405 15521 17417 15555
rect 17451 15552 17463 15555
rect 18966 15552 18972 15564
rect 17451 15524 18972 15552
rect 17451 15521 17463 15524
rect 17405 15515 17463 15521
rect 18966 15512 18972 15524
rect 19024 15512 19030 15564
rect 20162 15552 20168 15564
rect 20123 15524 20168 15552
rect 20162 15512 20168 15524
rect 20220 15512 20226 15564
rect 21183 15552 21211 15583
rect 21266 15580 21272 15592
rect 21324 15580 21330 15632
rect 20456 15524 21211 15552
rect 20456 15493 20484 15524
rect 21634 15512 21640 15564
rect 21692 15552 21698 15564
rect 22557 15555 22615 15561
rect 22557 15552 22569 15555
rect 21692 15524 22569 15552
rect 21692 15512 21698 15524
rect 22557 15521 22569 15524
rect 22603 15521 22615 15555
rect 22557 15515 22615 15521
rect 15752 15487 15810 15493
rect 15752 15484 15764 15487
rect 14792 15456 15240 15484
rect 15304 15456 15764 15484
rect 14792 15444 14798 15456
rect 15304 15416 15332 15456
rect 15752 15453 15764 15456
rect 15798 15453 15810 15487
rect 15752 15447 15810 15453
rect 17957 15487 18015 15493
rect 17957 15453 17969 15487
rect 18003 15453 18015 15487
rect 17957 15447 18015 15453
rect 20441 15487 20499 15493
rect 20441 15453 20453 15487
rect 20487 15453 20499 15487
rect 20898 15484 20904 15496
rect 20859 15456 20904 15484
rect 20441 15447 20499 15453
rect 14200 15388 15332 15416
rect 17129 15419 17187 15425
rect 17129 15385 17141 15419
rect 17175 15416 17187 15419
rect 17678 15416 17684 15428
rect 17175 15388 17684 15416
rect 17175 15385 17187 15388
rect 17129 15379 17187 15385
rect 17678 15376 17684 15388
rect 17736 15376 17742 15428
rect 13538 15348 13544 15360
rect 13188 15320 13544 15348
rect 12897 15311 12955 15317
rect 13538 15308 13544 15320
rect 13596 15308 13602 15360
rect 14182 15308 14188 15360
rect 14240 15348 14246 15360
rect 14553 15351 14611 15357
rect 14553 15348 14565 15351
rect 14240 15320 14565 15348
rect 14240 15308 14246 15320
rect 14553 15317 14565 15320
rect 14599 15317 14611 15351
rect 14553 15311 14611 15317
rect 15194 15308 15200 15360
rect 15252 15348 15258 15360
rect 15470 15348 15476 15360
rect 15252 15320 15476 15348
rect 15252 15308 15258 15320
rect 15470 15308 15476 15320
rect 15528 15308 15534 15360
rect 16114 15308 16120 15360
rect 16172 15348 16178 15360
rect 17589 15351 17647 15357
rect 17589 15348 17601 15351
rect 16172 15320 17601 15348
rect 16172 15308 16178 15320
rect 17589 15317 17601 15320
rect 17635 15317 17647 15351
rect 17972 15348 18000 15447
rect 20898 15444 20904 15456
rect 20956 15444 20962 15496
rect 18690 15348 18696 15360
rect 17972 15320 18696 15348
rect 17589 15311 17647 15317
rect 18690 15308 18696 15320
rect 18748 15308 18754 15360
rect 19794 15348 19800 15360
rect 19755 15320 19800 15348
rect 19794 15308 19800 15320
rect 19852 15308 19858 15360
rect 21542 15308 21548 15360
rect 21600 15348 21606 15360
rect 22281 15351 22339 15357
rect 22281 15348 22293 15351
rect 21600 15320 22293 15348
rect 21600 15308 21606 15320
rect 22281 15317 22293 15320
rect 22327 15317 22339 15351
rect 22281 15311 22339 15317
rect 1104 15258 23276 15280
rect 1104 15206 4680 15258
rect 4732 15206 4744 15258
rect 4796 15206 4808 15258
rect 4860 15206 4872 15258
rect 4924 15206 12078 15258
rect 12130 15206 12142 15258
rect 12194 15206 12206 15258
rect 12258 15206 12270 15258
rect 12322 15206 19475 15258
rect 19527 15206 19539 15258
rect 19591 15206 19603 15258
rect 19655 15206 19667 15258
rect 19719 15206 23276 15258
rect 1104 15184 23276 15206
rect 6730 15144 6736 15156
rect 3620 15116 6736 15144
rect 1854 15008 1860 15020
rect 1815 14980 1860 15008
rect 1854 14968 1860 14980
rect 1912 14968 1918 15020
rect 3620 14949 3648 15116
rect 6730 15104 6736 15116
rect 6788 15104 6794 15156
rect 10042 15104 10048 15156
rect 10100 15144 10106 15156
rect 10321 15147 10379 15153
rect 10321 15144 10333 15147
rect 10100 15116 10333 15144
rect 10100 15104 10106 15116
rect 10321 15113 10333 15116
rect 10367 15144 10379 15147
rect 11606 15144 11612 15156
rect 10367 15116 11612 15144
rect 10367 15113 10379 15116
rect 10321 15107 10379 15113
rect 11606 15104 11612 15116
rect 11664 15104 11670 15156
rect 11882 15104 11888 15156
rect 11940 15144 11946 15156
rect 12069 15147 12127 15153
rect 12069 15144 12081 15147
rect 11940 15116 12081 15144
rect 11940 15104 11946 15116
rect 12069 15113 12081 15116
rect 12115 15113 12127 15147
rect 12069 15107 12127 15113
rect 14458 15104 14464 15156
rect 14516 15144 14522 15156
rect 15010 15144 15016 15156
rect 14516 15116 15016 15144
rect 14516 15104 14522 15116
rect 15010 15104 15016 15116
rect 15068 15104 15074 15156
rect 17681 15147 17739 15153
rect 17681 15113 17693 15147
rect 17727 15144 17739 15147
rect 17954 15144 17960 15156
rect 17727 15116 17960 15144
rect 17727 15113 17739 15116
rect 17681 15107 17739 15113
rect 17954 15104 17960 15116
rect 18012 15104 18018 15156
rect 18966 15104 18972 15156
rect 19024 15144 19030 15156
rect 20438 15144 20444 15156
rect 19024 15116 20444 15144
rect 19024 15104 19030 15116
rect 20438 15104 20444 15116
rect 20496 15104 20502 15156
rect 20714 15104 20720 15156
rect 20772 15144 20778 15156
rect 21177 15147 21235 15153
rect 21177 15144 21189 15147
rect 20772 15116 21189 15144
rect 20772 15104 20778 15116
rect 21177 15113 21189 15116
rect 21223 15113 21235 15147
rect 21177 15107 21235 15113
rect 3789 15079 3847 15085
rect 3789 15045 3801 15079
rect 3835 15045 3847 15079
rect 3789 15039 3847 15045
rect 3804 15008 3832 15039
rect 11698 15036 11704 15088
rect 11756 15076 11762 15088
rect 12529 15079 12587 15085
rect 12529 15076 12541 15079
rect 11756 15048 12541 15076
rect 11756 15036 11762 15048
rect 12529 15045 12541 15048
rect 12575 15045 12587 15079
rect 12529 15039 12587 15045
rect 12710 15036 12716 15088
rect 12768 15076 12774 15088
rect 12986 15076 12992 15088
rect 12768 15048 12992 15076
rect 12768 15036 12774 15048
rect 12986 15036 12992 15048
rect 13044 15036 13050 15088
rect 18046 15036 18052 15088
rect 18104 15076 18110 15088
rect 19334 15076 19340 15088
rect 18104 15048 19340 15076
rect 18104 15036 18110 15048
rect 19334 15036 19340 15048
rect 19392 15036 19398 15088
rect 22649 15079 22707 15085
rect 22649 15076 22661 15079
rect 20732 15048 22661 15076
rect 4663 15011 4721 15017
rect 4663 15008 4675 15011
rect 3804 14980 4675 15008
rect 4663 14977 4675 14980
rect 4709 15008 4721 15011
rect 5350 15008 5356 15020
rect 4709 14980 5356 15008
rect 4709 14977 4721 14980
rect 4663 14971 4721 14977
rect 5350 14968 5356 14980
rect 5408 14968 5414 15020
rect 9950 14968 9956 15020
rect 10008 15008 10014 15020
rect 10008 14980 10732 15008
rect 10008 14968 10014 14980
rect 3605 14943 3663 14949
rect 3605 14909 3617 14943
rect 3651 14909 3663 14943
rect 3605 14903 3663 14909
rect 3970 14900 3976 14952
rect 4028 14940 4034 14952
rect 4157 14943 4215 14949
rect 4157 14940 4169 14943
rect 4028 14912 4169 14940
rect 4028 14900 4034 14912
rect 4157 14909 4169 14912
rect 4203 14909 4215 14943
rect 4157 14903 4215 14909
rect 4246 14900 4252 14952
rect 4304 14940 4310 14952
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4304 14912 4905 14940
rect 4304 14900 4310 14912
rect 4893 14909 4905 14912
rect 4939 14940 4951 14943
rect 5166 14940 5172 14952
rect 4939 14912 5172 14940
rect 4939 14909 4951 14912
rect 4893 14903 4951 14909
rect 5166 14900 5172 14912
rect 5224 14900 5230 14952
rect 6822 14940 6828 14952
rect 6783 14912 6828 14940
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 8941 14943 8999 14949
rect 8941 14909 8953 14943
rect 8987 14909 8999 14943
rect 8941 14903 8999 14909
rect 9208 14943 9266 14949
rect 9208 14909 9220 14943
rect 9254 14940 9266 14943
rect 9674 14940 9680 14952
rect 9254 14912 9680 14940
rect 9254 14909 9266 14912
rect 9208 14903 9266 14909
rect 2124 14875 2182 14881
rect 2124 14841 2136 14875
rect 2170 14872 2182 14875
rect 3050 14872 3056 14884
rect 2170 14844 3056 14872
rect 2170 14841 2182 14844
rect 2124 14835 2182 14841
rect 3050 14832 3056 14844
rect 3108 14832 3114 14884
rect 7098 14881 7104 14884
rect 7092 14872 7104 14881
rect 7059 14844 7104 14872
rect 7092 14835 7104 14844
rect 7098 14832 7104 14835
rect 7156 14832 7162 14884
rect 8956 14872 8984 14903
rect 9674 14900 9680 14912
rect 9732 14940 9738 14952
rect 10226 14940 10232 14952
rect 9732 14912 10232 14940
rect 9732 14900 9738 14912
rect 10226 14900 10232 14912
rect 10284 14900 10290 14952
rect 10704 14949 10732 14980
rect 12066 14968 12072 15020
rect 12124 15008 12130 15020
rect 13081 15011 13139 15017
rect 13081 15008 13093 15011
rect 12124 14980 13093 15008
rect 12124 14968 12130 14980
rect 13081 14977 13093 14980
rect 13127 14977 13139 15011
rect 13081 14971 13139 14977
rect 14918 14968 14924 15020
rect 14976 15008 14982 15020
rect 15841 15011 15899 15017
rect 15841 15008 15853 15011
rect 14976 14980 15853 15008
rect 14976 14968 14982 14980
rect 15841 14977 15853 14980
rect 15887 14977 15899 15011
rect 15841 14971 15899 14977
rect 18322 14968 18328 15020
rect 18380 15008 18386 15020
rect 18417 15011 18475 15017
rect 18417 15008 18429 15011
rect 18380 14980 18429 15008
rect 18380 14968 18386 14980
rect 18417 14977 18429 14980
rect 18463 14977 18475 15011
rect 18417 14971 18475 14977
rect 19843 15011 19901 15017
rect 19843 14977 19855 15011
rect 19889 15008 19901 15011
rect 20162 15008 20168 15020
rect 19889 14980 20168 15008
rect 19889 14977 19901 14980
rect 19843 14971 19901 14977
rect 20162 14968 20168 14980
rect 20220 15008 20226 15020
rect 20732 15008 20760 15048
rect 22649 15045 22661 15048
rect 22695 15045 22707 15079
rect 22649 15039 22707 15045
rect 20220 14980 20760 15008
rect 20220 14968 20226 14980
rect 21910 14968 21916 15020
rect 21968 15008 21974 15020
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21968 14980 22017 15008
rect 21968 14968 21974 14980
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 10689 14943 10747 14949
rect 10689 14909 10701 14943
rect 10735 14940 10747 14943
rect 10778 14940 10784 14952
rect 10735 14912 10784 14940
rect 10735 14909 10747 14912
rect 10689 14903 10747 14909
rect 10778 14900 10784 14912
rect 10836 14900 10842 14952
rect 10888 14912 11100 14940
rect 9582 14872 9588 14884
rect 8956 14844 9588 14872
rect 9582 14832 9588 14844
rect 9640 14872 9646 14884
rect 9950 14872 9956 14884
rect 9640 14844 9956 14872
rect 9640 14832 9646 14844
rect 9950 14832 9956 14844
rect 10008 14832 10014 14884
rect 10888 14872 10916 14912
rect 10244 14844 10916 14872
rect 10956 14875 11014 14881
rect 1394 14804 1400 14816
rect 1355 14776 1400 14804
rect 1394 14764 1400 14776
rect 1452 14764 1458 14816
rect 2958 14764 2964 14816
rect 3016 14804 3022 14816
rect 3237 14807 3295 14813
rect 3237 14804 3249 14807
rect 3016 14776 3249 14804
rect 3016 14764 3022 14776
rect 3237 14773 3249 14776
rect 3283 14804 3295 14807
rect 3694 14804 3700 14816
rect 3283 14776 3700 14804
rect 3283 14773 3295 14776
rect 3237 14767 3295 14773
rect 3694 14764 3700 14776
rect 3752 14764 3758 14816
rect 4623 14807 4681 14813
rect 4623 14773 4635 14807
rect 4669 14804 4681 14807
rect 4982 14804 4988 14816
rect 4669 14776 4988 14804
rect 4669 14773 4681 14776
rect 4623 14767 4681 14773
rect 4982 14764 4988 14776
rect 5040 14764 5046 14816
rect 5994 14804 6000 14816
rect 5955 14776 6000 14804
rect 5994 14764 6000 14776
rect 6052 14764 6058 14816
rect 6178 14764 6184 14816
rect 6236 14804 6242 14816
rect 6273 14807 6331 14813
rect 6273 14804 6285 14807
rect 6236 14776 6285 14804
rect 6236 14764 6242 14776
rect 6273 14773 6285 14776
rect 6319 14773 6331 14807
rect 8202 14804 8208 14816
rect 8163 14776 8208 14804
rect 6273 14767 6331 14773
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 8481 14807 8539 14813
rect 8481 14773 8493 14807
rect 8527 14804 8539 14807
rect 10244 14804 10272 14844
rect 10956 14841 10968 14875
rect 11002 14841 11014 14875
rect 11072 14872 11100 14912
rect 11790 14900 11796 14952
rect 11848 14940 11854 14952
rect 12897 14943 12955 14949
rect 12897 14940 12909 14943
rect 11848 14912 12909 14940
rect 11848 14900 11854 14912
rect 12897 14909 12909 14912
rect 12943 14909 12955 14943
rect 12897 14903 12955 14909
rect 13449 14943 13507 14949
rect 13449 14909 13461 14943
rect 13495 14940 13507 14943
rect 13538 14940 13544 14952
rect 13495 14912 13544 14940
rect 13495 14909 13507 14912
rect 13449 14903 13507 14909
rect 13538 14900 13544 14912
rect 13596 14940 13602 14952
rect 16301 14943 16359 14949
rect 16301 14940 16313 14943
rect 13596 14912 16313 14940
rect 13596 14900 13602 14912
rect 16301 14909 16313 14912
rect 16347 14909 16359 14943
rect 16301 14903 16359 14909
rect 17954 14900 17960 14952
rect 18012 14940 18018 14952
rect 18230 14940 18236 14952
rect 18012 14912 18236 14940
rect 18012 14900 18018 14912
rect 18230 14900 18236 14912
rect 18288 14900 18294 14952
rect 19242 14900 19248 14952
rect 19300 14940 19306 14952
rect 19337 14943 19395 14949
rect 19337 14940 19349 14943
rect 19300 14912 19349 14940
rect 19300 14900 19306 14912
rect 19337 14909 19349 14912
rect 19383 14909 19395 14943
rect 19337 14903 19395 14909
rect 19610 14900 19616 14952
rect 19668 14949 19674 14952
rect 19668 14943 19718 14949
rect 19668 14909 19672 14943
rect 19706 14909 19718 14943
rect 19668 14903 19718 14909
rect 19668 14900 19674 14903
rect 19978 14900 19984 14952
rect 20036 14940 20042 14952
rect 20073 14943 20131 14949
rect 20073 14940 20085 14943
rect 20036 14912 20085 14940
rect 20036 14900 20042 14912
rect 20073 14909 20085 14912
rect 20119 14940 20131 14943
rect 20714 14940 20720 14952
rect 20119 14912 20720 14940
rect 20119 14909 20131 14912
rect 20073 14903 20131 14909
rect 20714 14900 20720 14912
rect 20772 14900 20778 14952
rect 21726 14900 21732 14952
rect 21784 14940 21790 14952
rect 22465 14943 22523 14949
rect 21784 14912 21956 14940
rect 21784 14900 21790 14912
rect 12802 14872 12808 14884
rect 11072 14844 12808 14872
rect 10956 14835 11014 14841
rect 8527 14776 10272 14804
rect 10980 14804 11008 14835
rect 12802 14832 12808 14844
rect 12860 14832 12866 14884
rect 13262 14832 13268 14884
rect 13320 14872 13326 14884
rect 13694 14875 13752 14881
rect 13694 14872 13706 14875
rect 13320 14844 13706 14872
rect 13320 14832 13326 14844
rect 13694 14841 13706 14844
rect 13740 14872 13752 14875
rect 14182 14872 14188 14884
rect 13740 14844 14188 14872
rect 13740 14841 13752 14844
rect 13694 14835 13752 14841
rect 14182 14832 14188 14844
rect 14240 14832 14246 14884
rect 16568 14875 16626 14881
rect 16568 14841 16580 14875
rect 16614 14872 16626 14875
rect 18782 14872 18788 14884
rect 16614 14844 18788 14872
rect 16614 14841 16626 14844
rect 16568 14835 16626 14841
rect 18782 14832 18788 14844
rect 18840 14832 18846 14884
rect 21928 14881 21956 14912
rect 22465 14909 22477 14943
rect 22511 14940 22523 14943
rect 23014 14940 23020 14952
rect 22511 14912 23020 14940
rect 22511 14909 22523 14912
rect 22465 14903 22523 14909
rect 23014 14900 23020 14912
rect 23072 14900 23078 14952
rect 21913 14875 21971 14881
rect 21913 14841 21925 14875
rect 21959 14841 21971 14875
rect 21913 14835 21971 14841
rect 11238 14804 11244 14816
rect 10980 14776 11244 14804
rect 8527 14773 8539 14776
rect 8481 14767 8539 14773
rect 11238 14764 11244 14776
rect 11296 14764 11302 14816
rect 11422 14764 11428 14816
rect 11480 14804 11486 14816
rect 11606 14804 11612 14816
rect 11480 14776 11612 14804
rect 11480 14764 11486 14776
rect 11606 14764 11612 14776
rect 11664 14764 11670 14816
rect 12986 14804 12992 14816
rect 12947 14776 12992 14804
rect 12986 14764 12992 14776
rect 13044 14764 13050 14816
rect 14826 14804 14832 14816
rect 14787 14776 14832 14804
rect 14826 14764 14832 14776
rect 14884 14764 14890 14816
rect 15289 14807 15347 14813
rect 15289 14773 15301 14807
rect 15335 14804 15347 14807
rect 15470 14804 15476 14816
rect 15335 14776 15476 14804
rect 15335 14773 15347 14776
rect 15289 14767 15347 14773
rect 15470 14764 15476 14776
rect 15528 14764 15534 14816
rect 15562 14764 15568 14816
rect 15620 14804 15626 14816
rect 15657 14807 15715 14813
rect 15657 14804 15669 14807
rect 15620 14776 15669 14804
rect 15620 14764 15626 14776
rect 15657 14773 15669 14776
rect 15703 14773 15715 14807
rect 15657 14767 15715 14773
rect 15749 14807 15807 14813
rect 15749 14773 15761 14807
rect 15795 14804 15807 14807
rect 16206 14804 16212 14816
rect 15795 14776 16212 14804
rect 15795 14773 15807 14776
rect 15749 14767 15807 14773
rect 16206 14764 16212 14776
rect 16264 14764 16270 14816
rect 18598 14764 18604 14816
rect 18656 14804 18662 14816
rect 19610 14804 19616 14816
rect 18656 14776 19616 14804
rect 18656 14764 18662 14776
rect 19610 14764 19616 14776
rect 19668 14764 19674 14816
rect 21450 14804 21456 14816
rect 21411 14776 21456 14804
rect 21450 14764 21456 14776
rect 21508 14764 21514 14816
rect 21726 14764 21732 14816
rect 21784 14804 21790 14816
rect 21821 14807 21879 14813
rect 21821 14804 21833 14807
rect 21784 14776 21833 14804
rect 21784 14764 21790 14776
rect 21821 14773 21833 14776
rect 21867 14773 21879 14807
rect 21821 14767 21879 14773
rect 1104 14714 23276 14736
rect 1104 14662 8379 14714
rect 8431 14662 8443 14714
rect 8495 14662 8507 14714
rect 8559 14662 8571 14714
rect 8623 14662 15776 14714
rect 15828 14662 15840 14714
rect 15892 14662 15904 14714
rect 15956 14662 15968 14714
rect 16020 14662 23276 14714
rect 1104 14640 23276 14662
rect 1854 14560 1860 14612
rect 1912 14560 1918 14612
rect 3050 14600 3056 14612
rect 3011 14572 3056 14600
rect 3050 14560 3056 14572
rect 3108 14560 3114 14612
rect 3605 14603 3663 14609
rect 3605 14569 3617 14603
rect 3651 14569 3663 14603
rect 4062 14600 4068 14612
rect 4023 14572 4068 14600
rect 3605 14563 3663 14569
rect 1486 14424 1492 14476
rect 1544 14464 1550 14476
rect 1673 14467 1731 14473
rect 1673 14464 1685 14467
rect 1544 14436 1685 14464
rect 1544 14424 1550 14436
rect 1673 14433 1685 14436
rect 1719 14464 1731 14467
rect 1872 14464 1900 14560
rect 1940 14535 1998 14541
rect 1940 14501 1952 14535
rect 1986 14532 1998 14535
rect 2866 14532 2872 14544
rect 1986 14504 2872 14532
rect 1986 14501 1998 14504
rect 1940 14495 1998 14501
rect 2866 14492 2872 14504
rect 2924 14492 2930 14544
rect 3620 14532 3648 14563
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 4525 14603 4583 14609
rect 4525 14569 4537 14603
rect 4571 14600 4583 14603
rect 5077 14603 5135 14609
rect 5077 14600 5089 14603
rect 4571 14572 5089 14600
rect 4571 14569 4583 14572
rect 4525 14563 4583 14569
rect 5077 14569 5089 14572
rect 5123 14569 5135 14603
rect 5077 14563 5135 14569
rect 6273 14603 6331 14609
rect 6273 14569 6285 14603
rect 6319 14600 6331 14603
rect 9033 14603 9091 14609
rect 9033 14600 9045 14603
rect 6319 14572 9045 14600
rect 6319 14569 6331 14572
rect 6273 14563 6331 14569
rect 9033 14569 9045 14572
rect 9079 14569 9091 14603
rect 9033 14563 9091 14569
rect 9950 14560 9956 14612
rect 10008 14600 10014 14612
rect 10008 14572 11192 14600
rect 10008 14560 10014 14572
rect 5537 14535 5595 14541
rect 5537 14532 5549 14535
rect 3620 14504 5549 14532
rect 5537 14501 5549 14504
rect 5583 14501 5595 14535
rect 8941 14535 8999 14541
rect 5537 14495 5595 14501
rect 6104 14504 8607 14532
rect 1719 14436 1900 14464
rect 3421 14467 3479 14473
rect 1719 14433 1731 14436
rect 1673 14427 1731 14433
rect 3421 14433 3433 14467
rect 3467 14464 3479 14467
rect 3881 14467 3939 14473
rect 3881 14464 3893 14467
rect 3467 14436 3893 14464
rect 3467 14433 3479 14436
rect 3421 14427 3479 14433
rect 3881 14433 3893 14436
rect 3927 14433 3939 14467
rect 3881 14427 3939 14433
rect 4433 14467 4491 14473
rect 4433 14433 4445 14467
rect 4479 14464 4491 14467
rect 5258 14464 5264 14476
rect 4479 14436 5264 14464
rect 4479 14433 4491 14436
rect 4433 14427 4491 14433
rect 5258 14424 5264 14436
rect 5316 14424 5322 14476
rect 5350 14424 5356 14476
rect 5408 14464 5414 14476
rect 6104 14473 6132 14504
rect 5445 14467 5503 14473
rect 5445 14464 5457 14467
rect 5408 14436 5457 14464
rect 5408 14424 5414 14436
rect 5445 14433 5457 14436
rect 5491 14433 5503 14467
rect 5445 14427 5503 14433
rect 6089 14467 6147 14473
rect 6089 14433 6101 14467
rect 6135 14433 6147 14467
rect 6089 14427 6147 14433
rect 6454 14424 6460 14476
rect 6512 14464 6518 14476
rect 6897 14467 6955 14473
rect 6897 14464 6909 14467
rect 6512 14436 6909 14464
rect 6512 14424 6518 14436
rect 6897 14433 6909 14436
rect 6943 14464 6955 14467
rect 8202 14464 8208 14476
rect 6943 14436 8208 14464
rect 6943 14433 6955 14436
rect 6897 14427 6955 14433
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 8481 14467 8539 14473
rect 8481 14433 8493 14467
rect 8527 14433 8539 14467
rect 8579 14464 8607 14504
rect 8941 14501 8953 14535
rect 8987 14532 8999 14535
rect 9858 14532 9864 14544
rect 8987 14504 9864 14532
rect 8987 14501 8999 14504
rect 8941 14495 8999 14501
rect 9858 14492 9864 14504
rect 9916 14492 9922 14544
rect 10042 14492 10048 14544
rect 10100 14541 10106 14544
rect 10100 14535 10164 14541
rect 10100 14501 10118 14535
rect 10152 14501 10164 14535
rect 10502 14532 10508 14544
rect 10100 14495 10164 14501
rect 10336 14504 10508 14532
rect 10100 14492 10106 14495
rect 10336 14464 10364 14504
rect 10502 14492 10508 14504
rect 10560 14492 10566 14544
rect 11164 14532 11192 14572
rect 11330 14560 11336 14612
rect 11388 14600 11394 14612
rect 11517 14603 11575 14609
rect 11517 14600 11529 14603
rect 11388 14572 11529 14600
rect 11388 14560 11394 14572
rect 11517 14569 11529 14572
rect 11563 14600 11575 14603
rect 11974 14600 11980 14612
rect 11563 14572 11980 14600
rect 11563 14569 11575 14572
rect 11517 14563 11575 14569
rect 11974 14560 11980 14572
rect 12032 14560 12038 14612
rect 12618 14560 12624 14612
rect 12676 14600 12682 14612
rect 14090 14600 14096 14612
rect 12676 14572 14096 14600
rect 12676 14560 12682 14572
rect 14090 14560 14096 14572
rect 14148 14600 14154 14612
rect 14369 14603 14427 14609
rect 14369 14600 14381 14603
rect 14148 14572 14381 14600
rect 14148 14560 14154 14572
rect 14369 14569 14381 14572
rect 14415 14569 14427 14603
rect 14918 14600 14924 14612
rect 14879 14572 14924 14600
rect 14369 14563 14427 14569
rect 14918 14560 14924 14572
rect 14976 14560 14982 14612
rect 16669 14603 16727 14609
rect 16669 14569 16681 14603
rect 16715 14600 16727 14603
rect 19150 14600 19156 14612
rect 16715 14572 19156 14600
rect 16715 14569 16727 14572
rect 16669 14563 16727 14569
rect 19150 14560 19156 14572
rect 19208 14560 19214 14612
rect 19794 14560 19800 14612
rect 19852 14600 19858 14612
rect 20257 14603 20315 14609
rect 20257 14600 20269 14603
rect 19852 14572 20269 14600
rect 19852 14560 19858 14572
rect 20257 14569 20269 14572
rect 20303 14569 20315 14603
rect 21634 14600 21640 14612
rect 20257 14563 20315 14569
rect 21008 14572 21640 14600
rect 11698 14532 11704 14544
rect 11164 14504 11704 14532
rect 11698 14492 11704 14504
rect 11756 14492 11762 14544
rect 12526 14532 12532 14544
rect 12084 14504 12532 14532
rect 8579 14436 10364 14464
rect 8481 14427 8539 14433
rect 3050 14356 3056 14408
rect 3108 14396 3114 14408
rect 4617 14399 4675 14405
rect 4617 14396 4629 14399
rect 3108 14368 4629 14396
rect 3108 14356 3114 14368
rect 4617 14365 4629 14368
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 4706 14356 4712 14408
rect 4764 14396 4770 14408
rect 5629 14399 5687 14405
rect 5629 14396 5641 14399
rect 4764 14368 5641 14396
rect 4764 14356 4770 14368
rect 5629 14365 5641 14368
rect 5675 14365 5687 14399
rect 5629 14359 5687 14365
rect 6641 14399 6699 14405
rect 6641 14365 6653 14399
rect 6687 14365 6699 14399
rect 8496 14396 8524 14427
rect 10410 14424 10416 14476
rect 10468 14464 10474 14476
rect 11885 14467 11943 14473
rect 11885 14464 11897 14467
rect 10468 14436 11897 14464
rect 10468 14424 10474 14436
rect 11885 14433 11897 14436
rect 11931 14433 11943 14467
rect 11885 14427 11943 14433
rect 9030 14396 9036 14408
rect 8496 14368 9036 14396
rect 6641 14359 6699 14365
rect 3881 14331 3939 14337
rect 3881 14297 3893 14331
rect 3927 14328 3939 14331
rect 6454 14328 6460 14340
rect 3927 14300 6460 14328
rect 3927 14297 3939 14300
rect 3881 14291 3939 14297
rect 6454 14288 6460 14300
rect 6512 14288 6518 14340
rect 4338 14220 4344 14272
rect 4396 14260 4402 14272
rect 4982 14260 4988 14272
rect 4396 14232 4988 14260
rect 4396 14220 4402 14232
rect 4982 14220 4988 14232
rect 5040 14260 5046 14272
rect 6656 14260 6684 14359
rect 9030 14356 9036 14368
rect 9088 14356 9094 14408
rect 9217 14399 9275 14405
rect 9217 14365 9229 14399
rect 9263 14396 9275 14399
rect 9401 14399 9459 14405
rect 9401 14396 9413 14399
rect 9263 14368 9413 14396
rect 9263 14365 9275 14368
rect 9217 14359 9275 14365
rect 9401 14365 9413 14368
rect 9447 14365 9459 14399
rect 9401 14359 9459 14365
rect 9582 14356 9588 14408
rect 9640 14396 9646 14408
rect 9861 14399 9919 14405
rect 9861 14396 9873 14399
rect 9640 14368 9873 14396
rect 9640 14356 9646 14368
rect 9861 14365 9873 14368
rect 9907 14365 9919 14399
rect 9861 14359 9919 14365
rect 10962 14356 10968 14408
rect 11020 14396 11026 14408
rect 12084 14405 12112 14504
rect 12526 14492 12532 14504
rect 12584 14492 12590 14544
rect 12704 14535 12762 14541
rect 12704 14501 12716 14535
rect 12750 14532 12762 14535
rect 12802 14532 12808 14544
rect 12750 14504 12808 14532
rect 12750 14501 12762 14504
rect 12704 14495 12762 14501
rect 12802 14492 12808 14504
rect 12860 14492 12866 14544
rect 13078 14492 13084 14544
rect 13136 14532 13142 14544
rect 14277 14535 14335 14541
rect 14277 14532 14289 14535
rect 13136 14504 14289 14532
rect 13136 14492 13142 14504
rect 14277 14501 14289 14504
rect 14323 14501 14335 14535
rect 19978 14532 19984 14544
rect 14277 14495 14335 14501
rect 14752 14504 19984 14532
rect 14752 14473 14780 14504
rect 19978 14492 19984 14504
rect 20036 14492 20042 14544
rect 20165 14535 20223 14541
rect 20165 14501 20177 14535
rect 20211 14532 20223 14535
rect 21008 14532 21036 14572
rect 21634 14560 21640 14572
rect 21692 14560 21698 14612
rect 21444 14535 21502 14541
rect 21444 14532 21456 14535
rect 20211 14504 21036 14532
rect 21100 14504 21456 14532
rect 20211 14501 20223 14504
rect 20165 14495 20223 14501
rect 14737 14467 14795 14473
rect 14737 14433 14749 14467
rect 14783 14433 14795 14467
rect 14737 14427 14795 14433
rect 15654 14424 15660 14476
rect 15712 14464 15718 14476
rect 16117 14467 16175 14473
rect 16117 14464 16129 14467
rect 15712 14436 16129 14464
rect 15712 14424 15718 14436
rect 16117 14433 16129 14436
rect 16163 14433 16175 14467
rect 16117 14427 16175 14433
rect 16669 14467 16727 14473
rect 16669 14433 16681 14467
rect 16715 14464 16727 14467
rect 16761 14467 16819 14473
rect 16761 14464 16773 14467
rect 16715 14436 16773 14464
rect 16715 14433 16727 14436
rect 16669 14427 16727 14433
rect 16761 14433 16773 14436
rect 16807 14433 16819 14467
rect 16761 14427 16819 14433
rect 17497 14467 17555 14473
rect 17497 14433 17509 14467
rect 17543 14464 17555 14467
rect 17586 14464 17592 14476
rect 17543 14436 17592 14464
rect 17543 14433 17555 14436
rect 17497 14427 17555 14433
rect 17586 14424 17592 14436
rect 17644 14424 17650 14476
rect 17770 14473 17776 14476
rect 17764 14427 17776 14473
rect 17828 14464 17834 14476
rect 18969 14467 19027 14473
rect 18969 14464 18981 14467
rect 17828 14436 18981 14464
rect 17770 14424 17776 14427
rect 17828 14424 17834 14436
rect 18969 14433 18981 14436
rect 19015 14433 19027 14467
rect 18969 14427 19027 14433
rect 19150 14424 19156 14476
rect 19208 14473 19214 14476
rect 19208 14467 19229 14473
rect 19217 14433 19229 14467
rect 19208 14427 19229 14433
rect 19208 14424 19214 14427
rect 19334 14424 19340 14476
rect 19392 14464 19398 14476
rect 19392 14436 19435 14464
rect 19392 14424 19398 14436
rect 11977 14399 12035 14405
rect 11977 14396 11989 14399
rect 11020 14368 11989 14396
rect 11020 14356 11026 14368
rect 11977 14365 11989 14368
rect 12023 14365 12035 14399
rect 11977 14359 12035 14365
rect 12069 14399 12127 14405
rect 12069 14365 12081 14399
rect 12115 14365 12127 14399
rect 12434 14396 12440 14408
rect 12395 14368 12440 14396
rect 12069 14359 12127 14365
rect 8573 14331 8631 14337
rect 8573 14297 8585 14331
rect 8619 14328 8631 14331
rect 9766 14328 9772 14340
rect 8619 14300 9772 14328
rect 8619 14297 8631 14300
rect 8573 14291 8631 14297
rect 9766 14288 9772 14300
rect 9824 14288 9830 14340
rect 11238 14328 11244 14340
rect 11199 14300 11244 14328
rect 11238 14288 11244 14300
rect 11296 14288 11302 14340
rect 11422 14288 11428 14340
rect 11480 14328 11486 14340
rect 12084 14328 12112 14359
rect 12434 14356 12440 14368
rect 12492 14356 12498 14408
rect 14461 14399 14519 14405
rect 14461 14365 14473 14399
rect 14507 14365 14519 14399
rect 14461 14359 14519 14365
rect 14476 14328 14504 14359
rect 14642 14356 14648 14408
rect 14700 14396 14706 14408
rect 15289 14399 15347 14405
rect 15289 14396 15301 14399
rect 14700 14368 15301 14396
rect 14700 14356 14706 14368
rect 15289 14365 15301 14368
rect 15335 14365 15347 14399
rect 16206 14396 16212 14408
rect 16167 14368 16212 14396
rect 15289 14359 15347 14365
rect 16206 14356 16212 14368
rect 16264 14356 16270 14408
rect 16393 14399 16451 14405
rect 16393 14365 16405 14399
rect 16439 14396 16451 14399
rect 20441 14399 20499 14405
rect 16439 14368 16988 14396
rect 16439 14365 16451 14368
rect 16393 14359 16451 14365
rect 11480 14300 12112 14328
rect 13464 14300 14504 14328
rect 11480 14288 11486 14300
rect 6822 14260 6828 14272
rect 5040 14232 6828 14260
rect 5040 14220 5046 14232
rect 6822 14220 6828 14232
rect 6880 14220 6886 14272
rect 7006 14220 7012 14272
rect 7064 14260 7070 14272
rect 8021 14263 8079 14269
rect 8021 14260 8033 14263
rect 7064 14232 8033 14260
rect 7064 14220 7070 14232
rect 8021 14229 8033 14232
rect 8067 14229 8079 14263
rect 8021 14223 8079 14229
rect 8297 14263 8355 14269
rect 8297 14229 8309 14263
rect 8343 14260 8355 14263
rect 8662 14260 8668 14272
rect 8343 14232 8668 14260
rect 8343 14229 8355 14232
rect 8297 14223 8355 14229
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 9401 14263 9459 14269
rect 9401 14229 9413 14263
rect 9447 14260 9459 14263
rect 10042 14260 10048 14272
rect 9447 14232 10048 14260
rect 9447 14229 9459 14232
rect 9401 14223 9459 14229
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 11882 14220 11888 14272
rect 11940 14260 11946 14272
rect 13464 14260 13492 14300
rect 11940 14232 13492 14260
rect 11940 14220 11946 14232
rect 13722 14220 13728 14272
rect 13780 14260 13786 14272
rect 13817 14263 13875 14269
rect 13817 14260 13829 14263
rect 13780 14232 13829 14260
rect 13780 14220 13786 14232
rect 13817 14229 13829 14232
rect 13863 14229 13875 14263
rect 13817 14223 13875 14229
rect 13906 14220 13912 14272
rect 13964 14260 13970 14272
rect 15746 14260 15752 14272
rect 13964 14232 14009 14260
rect 15707 14232 15752 14260
rect 13964 14220 13970 14232
rect 15746 14220 15752 14232
rect 15804 14220 15810 14272
rect 16960 14269 16988 14368
rect 20441 14365 20453 14399
rect 20487 14396 20499 14399
rect 21100 14396 21128 14504
rect 21444 14501 21456 14504
rect 21490 14532 21502 14535
rect 21542 14532 21548 14544
rect 21490 14504 21548 14532
rect 21490 14501 21502 14504
rect 21444 14495 21502 14501
rect 21542 14492 21548 14504
rect 21600 14492 21606 14544
rect 20487 14368 21128 14396
rect 21177 14399 21235 14405
rect 20487 14365 20499 14368
rect 20441 14359 20499 14365
rect 21177 14365 21189 14399
rect 21223 14365 21235 14399
rect 21177 14359 21235 14365
rect 18506 14288 18512 14340
rect 18564 14328 18570 14340
rect 19521 14331 19579 14337
rect 19521 14328 19533 14331
rect 18564 14300 19533 14328
rect 18564 14288 18570 14300
rect 19521 14297 19533 14300
rect 19567 14297 19579 14331
rect 19521 14291 19579 14297
rect 19610 14288 19616 14340
rect 19668 14328 19674 14340
rect 19797 14331 19855 14337
rect 19797 14328 19809 14331
rect 19668 14300 19809 14328
rect 19668 14288 19674 14300
rect 19797 14297 19809 14300
rect 19843 14328 19855 14331
rect 19978 14328 19984 14340
rect 19843 14300 19984 14328
rect 19843 14297 19855 14300
rect 19797 14291 19855 14297
rect 19978 14288 19984 14300
rect 20036 14288 20042 14340
rect 20990 14288 20996 14340
rect 21048 14328 21054 14340
rect 21192 14328 21220 14359
rect 21048 14300 21220 14328
rect 21048 14288 21054 14300
rect 16945 14263 17003 14269
rect 16945 14229 16957 14263
rect 16991 14260 17003 14263
rect 17218 14260 17224 14272
rect 16991 14232 17224 14260
rect 16991 14229 17003 14232
rect 16945 14223 17003 14229
rect 17218 14220 17224 14232
rect 17276 14220 17282 14272
rect 18874 14260 18880 14272
rect 18835 14232 18880 14260
rect 18874 14220 18880 14232
rect 18932 14220 18938 14272
rect 18969 14263 19027 14269
rect 18969 14229 18981 14263
rect 19015 14260 19027 14263
rect 19334 14260 19340 14272
rect 19015 14232 19340 14260
rect 19015 14229 19027 14232
rect 18969 14223 19027 14229
rect 19334 14220 19340 14232
rect 19392 14220 19398 14272
rect 21910 14220 21916 14272
rect 21968 14260 21974 14272
rect 22557 14263 22615 14269
rect 22557 14260 22569 14263
rect 21968 14232 22569 14260
rect 21968 14220 21974 14232
rect 22557 14229 22569 14232
rect 22603 14229 22615 14263
rect 22557 14223 22615 14229
rect 1104 14170 23276 14192
rect 1104 14118 4680 14170
rect 4732 14118 4744 14170
rect 4796 14118 4808 14170
rect 4860 14118 4872 14170
rect 4924 14118 12078 14170
rect 12130 14118 12142 14170
rect 12194 14118 12206 14170
rect 12258 14118 12270 14170
rect 12322 14118 19475 14170
rect 19527 14118 19539 14170
rect 19591 14118 19603 14170
rect 19655 14118 19667 14170
rect 19719 14118 23276 14170
rect 1104 14096 23276 14118
rect 2866 14056 2872 14068
rect 2827 14028 2872 14056
rect 2866 14016 2872 14028
rect 2924 14016 2930 14068
rect 3973 14059 4031 14065
rect 3973 14025 3985 14059
rect 4019 14056 4031 14059
rect 4246 14056 4252 14068
rect 4019 14028 4252 14056
rect 4019 14025 4031 14028
rect 3973 14019 4031 14025
rect 4246 14016 4252 14028
rect 4304 14016 4310 14068
rect 4341 14059 4399 14065
rect 4341 14025 4353 14059
rect 4387 14056 4399 14059
rect 7374 14056 7380 14068
rect 4387 14028 7380 14056
rect 4387 14025 4399 14028
rect 4341 14019 4399 14025
rect 7374 14016 7380 14028
rect 7432 14016 7438 14068
rect 8662 14016 8668 14068
rect 8720 14056 8726 14068
rect 9214 14056 9220 14068
rect 8720 14028 9220 14056
rect 8720 14016 8726 14028
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 9674 14056 9680 14068
rect 9635 14028 9680 14056
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 10502 14016 10508 14068
rect 10560 14056 10566 14068
rect 10965 14059 11023 14065
rect 10965 14056 10977 14059
rect 10560 14028 10977 14056
rect 10560 14016 10566 14028
rect 10965 14025 10977 14028
rect 11011 14025 11023 14059
rect 10965 14019 11023 14025
rect 11606 14016 11612 14068
rect 11664 14056 11670 14068
rect 11882 14056 11888 14068
rect 11664 14028 11888 14056
rect 11664 14016 11670 14028
rect 11882 14016 11888 14028
rect 11940 14016 11946 14068
rect 17681 14059 17739 14065
rect 17681 14025 17693 14059
rect 17727 14056 17739 14059
rect 17770 14056 17776 14068
rect 17727 14028 17776 14056
rect 17727 14025 17739 14028
rect 17681 14019 17739 14025
rect 17770 14016 17776 14028
rect 17828 14016 17834 14068
rect 17862 14016 17868 14068
rect 17920 14056 17926 14068
rect 19521 14059 19579 14065
rect 19521 14056 19533 14059
rect 17920 14028 19533 14056
rect 17920 14016 17926 14028
rect 19521 14025 19533 14028
rect 19567 14025 19579 14059
rect 19521 14019 19579 14025
rect 20714 14016 20720 14068
rect 20772 14056 20778 14068
rect 21453 14059 21511 14065
rect 21453 14056 21465 14059
rect 20772 14028 21465 14056
rect 20772 14016 20778 14028
rect 21453 14025 21465 14028
rect 21499 14025 21511 14059
rect 21453 14019 21511 14025
rect 6454 13948 6460 14000
rect 6512 13988 6518 14000
rect 6825 13991 6883 13997
rect 6825 13988 6837 13991
rect 6512 13960 6837 13988
rect 6512 13948 6518 13960
rect 6825 13957 6837 13960
rect 6871 13957 6883 13991
rect 6825 13951 6883 13957
rect 9953 13991 10011 13997
rect 9953 13957 9965 13991
rect 9999 13957 10011 13991
rect 9953 13951 10011 13957
rect 1486 13920 1492 13932
rect 1447 13892 1492 13920
rect 1486 13880 1492 13892
rect 1544 13880 1550 13932
rect 3694 13920 3700 13932
rect 3655 13892 3700 13920
rect 3694 13880 3700 13892
rect 3752 13880 3758 13932
rect 4080 13892 4835 13920
rect 1756 13855 1814 13861
rect 1756 13821 1768 13855
rect 1802 13852 1814 13855
rect 4080 13852 4108 13892
rect 1802 13824 4108 13852
rect 4157 13855 4215 13861
rect 1802 13821 1814 13824
rect 1756 13815 1814 13821
rect 4157 13821 4169 13855
rect 4203 13821 4215 13855
rect 4157 13815 4215 13821
rect 3513 13787 3571 13793
rect 3513 13753 3525 13787
rect 3559 13784 3571 13787
rect 4062 13784 4068 13796
rect 3559 13756 4068 13784
rect 3559 13753 3571 13756
rect 3513 13747 3571 13753
rect 4062 13744 4068 13756
rect 4120 13744 4126 13796
rect 4172 13784 4200 13815
rect 4522 13784 4528 13796
rect 4172 13756 4528 13784
rect 4522 13744 4528 13756
rect 4580 13744 4586 13796
rect 3142 13716 3148 13728
rect 3103 13688 3148 13716
rect 3142 13676 3148 13688
rect 3200 13676 3206 13728
rect 3605 13719 3663 13725
rect 3605 13685 3617 13719
rect 3651 13716 3663 13719
rect 3973 13719 4031 13725
rect 3973 13716 3985 13719
rect 3651 13688 3985 13716
rect 3651 13685 3663 13688
rect 3605 13679 3663 13685
rect 3973 13685 3985 13688
rect 4019 13685 4031 13719
rect 4807 13716 4835 13892
rect 7190 13880 7196 13932
rect 7248 13920 7254 13932
rect 7377 13923 7435 13929
rect 7377 13920 7389 13923
rect 7248 13892 7389 13920
rect 7248 13880 7254 13892
rect 7377 13889 7389 13892
rect 7423 13889 7435 13923
rect 7377 13883 7435 13889
rect 7742 13880 7748 13932
rect 7800 13920 7806 13932
rect 7837 13923 7895 13929
rect 7837 13920 7849 13923
rect 7800 13892 7849 13920
rect 7800 13880 7806 13892
rect 7837 13889 7849 13892
rect 7883 13889 7895 13923
rect 7837 13883 7895 13889
rect 9766 13880 9772 13932
rect 9824 13920 9830 13932
rect 9968 13920 9996 13951
rect 10686 13948 10692 14000
rect 10744 13988 10750 14000
rect 11977 13991 12035 13997
rect 11977 13988 11989 13991
rect 10744 13960 11989 13988
rect 10744 13948 10750 13960
rect 11977 13957 11989 13960
rect 12023 13957 12035 13991
rect 11977 13951 12035 13957
rect 18233 13991 18291 13997
rect 18233 13957 18245 13991
rect 18279 13988 18291 13991
rect 19610 13988 19616 14000
rect 18279 13960 19616 13988
rect 18279 13957 18291 13960
rect 18233 13951 18291 13957
rect 19610 13948 19616 13960
rect 19668 13948 19674 14000
rect 21729 13991 21787 13997
rect 21729 13957 21741 13991
rect 21775 13957 21787 13991
rect 21729 13951 21787 13957
rect 10597 13923 10655 13929
rect 9824 13892 10548 13920
rect 9824 13880 9830 13892
rect 4893 13855 4951 13861
rect 4893 13821 4905 13855
rect 4939 13852 4951 13855
rect 4982 13852 4988 13864
rect 4939 13824 4988 13852
rect 4939 13821 4951 13824
rect 4893 13815 4951 13821
rect 4982 13812 4988 13824
rect 5040 13812 5046 13864
rect 5160 13855 5218 13861
rect 5160 13821 5172 13855
rect 5206 13852 5218 13855
rect 5718 13852 5724 13864
rect 5206 13824 5724 13852
rect 5206 13821 5218 13824
rect 5160 13815 5218 13821
rect 5718 13812 5724 13824
rect 5776 13812 5782 13864
rect 6270 13812 6276 13864
rect 6328 13852 6334 13864
rect 6454 13852 6460 13864
rect 6328 13824 6460 13852
rect 6328 13812 6334 13824
rect 6454 13812 6460 13824
rect 6512 13812 6518 13864
rect 8202 13812 8208 13864
rect 8260 13852 8266 13864
rect 8297 13855 8355 13861
rect 8297 13852 8309 13855
rect 8260 13824 8309 13852
rect 8260 13812 8266 13824
rect 8297 13821 8309 13824
rect 8343 13821 8355 13855
rect 8297 13815 8355 13821
rect 8564 13855 8622 13861
rect 8564 13821 8576 13855
rect 8610 13852 8622 13855
rect 10413 13855 10471 13861
rect 10413 13852 10425 13855
rect 8610 13824 9168 13852
rect 8610 13821 8622 13824
rect 8564 13815 8622 13821
rect 6270 13716 6276 13728
rect 4807 13688 6276 13716
rect 3973 13679 4031 13685
rect 6270 13676 6276 13688
rect 6328 13676 6334 13728
rect 6730 13676 6736 13728
rect 6788 13716 6794 13728
rect 7190 13716 7196 13728
rect 6788 13688 7196 13716
rect 6788 13676 6794 13688
rect 7190 13676 7196 13688
rect 7248 13676 7254 13728
rect 7282 13676 7288 13728
rect 7340 13716 7346 13728
rect 9140 13716 9168 13824
rect 9232 13824 10425 13852
rect 9232 13796 9260 13824
rect 10413 13821 10425 13824
rect 10459 13821 10471 13855
rect 10520 13852 10548 13892
rect 10597 13889 10609 13923
rect 10643 13920 10655 13923
rect 11422 13920 11428 13932
rect 10643 13892 11428 13920
rect 10643 13889 10655 13892
rect 10597 13883 10655 13889
rect 11422 13880 11428 13892
rect 11480 13880 11486 13932
rect 11606 13920 11612 13932
rect 11567 13892 11612 13920
rect 11606 13880 11612 13892
rect 11664 13880 11670 13932
rect 18874 13920 18880 13932
rect 18835 13892 18880 13920
rect 18874 13880 18880 13892
rect 18932 13880 18938 13932
rect 19242 13880 19248 13932
rect 19300 13920 19306 13932
rect 19300 13892 19656 13920
rect 19300 13880 19306 13892
rect 11330 13852 11336 13864
rect 10520 13824 11008 13852
rect 11291 13824 11336 13852
rect 10413 13815 10471 13821
rect 9214 13744 9220 13796
rect 9272 13744 9278 13796
rect 10042 13784 10048 13796
rect 9324 13756 10048 13784
rect 9324 13716 9352 13756
rect 10042 13744 10048 13756
rect 10100 13744 10106 13796
rect 7340 13688 7385 13716
rect 9140 13688 9352 13716
rect 7340 13676 7346 13688
rect 9490 13676 9496 13728
rect 9548 13716 9554 13728
rect 10321 13719 10379 13725
rect 10321 13716 10333 13719
rect 9548 13688 10333 13716
rect 9548 13676 9554 13688
rect 10321 13685 10333 13688
rect 10367 13685 10379 13719
rect 10980 13716 11008 13824
rect 11330 13812 11336 13824
rect 11388 13812 11394 13864
rect 12161 13855 12219 13861
rect 12161 13852 12173 13855
rect 11440 13824 12173 13852
rect 11054 13744 11060 13796
rect 11112 13784 11118 13796
rect 11440 13784 11468 13824
rect 12161 13821 12173 13824
rect 12207 13821 12219 13855
rect 12161 13815 12219 13821
rect 12434 13812 12440 13864
rect 12492 13852 12498 13864
rect 13078 13861 13084 13864
rect 12805 13855 12863 13861
rect 12805 13852 12817 13855
rect 12492 13824 12817 13852
rect 12492 13812 12498 13824
rect 12805 13821 12817 13824
rect 12851 13821 12863 13855
rect 12805 13815 12863 13821
rect 13072 13815 13084 13861
rect 13136 13852 13142 13864
rect 14553 13855 14611 13861
rect 13136 13824 13172 13852
rect 11112 13756 11468 13784
rect 12820 13784 12848 13815
rect 13078 13812 13084 13815
rect 13136 13812 13142 13824
rect 14553 13821 14565 13855
rect 14599 13852 14611 13855
rect 16301 13855 16359 13861
rect 14599 13824 14964 13852
rect 14599 13821 14611 13824
rect 14553 13815 14611 13821
rect 13538 13784 13544 13796
rect 12820 13756 13544 13784
rect 11112 13744 11118 13756
rect 13538 13744 13544 13756
rect 13596 13784 13602 13796
rect 14568 13784 14596 13815
rect 14936 13796 14964 13824
rect 16301 13821 16313 13855
rect 16347 13852 16359 13855
rect 17586 13852 17592 13864
rect 16347 13824 17592 13852
rect 16347 13821 16359 13824
rect 16301 13815 16359 13821
rect 17586 13812 17592 13824
rect 17644 13812 17650 13864
rect 18693 13855 18751 13861
rect 18693 13821 18705 13855
rect 18739 13852 18751 13855
rect 19150 13852 19156 13864
rect 18739 13824 19156 13852
rect 18739 13821 18751 13824
rect 18693 13815 18751 13821
rect 19150 13812 19156 13824
rect 19208 13812 19214 13864
rect 19628 13861 19656 13892
rect 19794 13880 19800 13932
rect 19852 13920 19858 13932
rect 19936 13923 19994 13929
rect 19936 13920 19948 13923
rect 19852 13892 19948 13920
rect 19852 13880 19858 13892
rect 19936 13889 19948 13892
rect 19982 13889 19994 13923
rect 19936 13883 19994 13889
rect 20119 13923 20177 13929
rect 20119 13889 20131 13923
rect 20165 13920 20177 13923
rect 21744 13920 21772 13951
rect 20165 13892 21772 13920
rect 22373 13923 22431 13929
rect 20165 13889 20177 13892
rect 20119 13883 20177 13889
rect 22373 13889 22385 13923
rect 22419 13920 22431 13923
rect 22830 13920 22836 13932
rect 22419 13892 22836 13920
rect 22419 13889 22431 13892
rect 22373 13883 22431 13889
rect 22830 13880 22836 13892
rect 22888 13880 22894 13932
rect 19429 13855 19487 13861
rect 19429 13821 19441 13855
rect 19475 13852 19487 13855
rect 19521 13855 19579 13861
rect 19521 13852 19533 13855
rect 19475 13824 19533 13852
rect 19475 13821 19487 13824
rect 19429 13815 19487 13821
rect 19521 13821 19533 13824
rect 19567 13821 19579 13855
rect 19521 13815 19579 13821
rect 19613 13855 19671 13861
rect 19613 13821 19625 13855
rect 19659 13821 19671 13855
rect 19613 13815 19671 13821
rect 20349 13855 20407 13861
rect 20349 13821 20361 13855
rect 20395 13852 20407 13855
rect 20395 13824 21220 13852
rect 20395 13821 20407 13824
rect 20349 13815 20407 13821
rect 13596 13756 14596 13784
rect 13596 13744 13602 13756
rect 14642 13744 14648 13796
rect 14700 13784 14706 13796
rect 14798 13787 14856 13793
rect 14798 13784 14810 13787
rect 14700 13756 14810 13784
rect 14700 13744 14706 13756
rect 14798 13753 14810 13756
rect 14844 13753 14856 13787
rect 14798 13747 14856 13753
rect 14918 13744 14924 13796
rect 14976 13744 14982 13796
rect 15010 13744 15016 13796
rect 15068 13784 15074 13796
rect 16568 13787 16626 13793
rect 15068 13756 16068 13784
rect 15068 13744 15074 13756
rect 11425 13719 11483 13725
rect 11425 13716 11437 13719
rect 10980 13688 11437 13716
rect 10321 13679 10379 13685
rect 11425 13685 11437 13688
rect 11471 13685 11483 13719
rect 11425 13679 11483 13685
rect 13814 13676 13820 13728
rect 13872 13716 13878 13728
rect 14185 13719 14243 13725
rect 14185 13716 14197 13719
rect 13872 13688 14197 13716
rect 13872 13676 13878 13688
rect 14185 13685 14197 13688
rect 14231 13685 14243 13719
rect 14185 13679 14243 13685
rect 15378 13676 15384 13728
rect 15436 13716 15442 13728
rect 15933 13719 15991 13725
rect 15933 13716 15945 13719
rect 15436 13688 15945 13716
rect 15436 13676 15442 13688
rect 15933 13685 15945 13688
rect 15979 13685 15991 13719
rect 16040 13716 16068 13756
rect 16568 13753 16580 13787
rect 16614 13784 16626 13787
rect 17402 13784 17408 13796
rect 16614 13756 17408 13784
rect 16614 13753 16626 13756
rect 16568 13747 16626 13753
rect 17402 13744 17408 13756
rect 17460 13744 17466 13796
rect 19334 13784 19340 13796
rect 17512 13756 19340 13784
rect 17512 13716 17540 13756
rect 19334 13744 19340 13756
rect 19392 13744 19398 13796
rect 21192 13784 21220 13824
rect 21450 13812 21456 13864
rect 21508 13852 21514 13864
rect 22189 13855 22247 13861
rect 22189 13852 22201 13855
rect 21508 13824 22201 13852
rect 21508 13812 21514 13824
rect 22189 13821 22201 13824
rect 22235 13821 22247 13855
rect 22189 13815 22247 13821
rect 21726 13784 21732 13796
rect 21192 13756 21732 13784
rect 21726 13744 21732 13756
rect 21784 13744 21790 13796
rect 16040 13688 17540 13716
rect 15933 13679 15991 13685
rect 18046 13676 18052 13728
rect 18104 13716 18110 13728
rect 18601 13719 18659 13725
rect 18601 13716 18613 13719
rect 18104 13688 18613 13716
rect 18104 13676 18110 13688
rect 18601 13685 18613 13688
rect 18647 13685 18659 13719
rect 18601 13679 18659 13685
rect 19245 13719 19303 13725
rect 19245 13685 19257 13719
rect 19291 13716 19303 13719
rect 20990 13716 20996 13728
rect 19291 13688 20996 13716
rect 19291 13685 19303 13688
rect 19245 13679 19303 13685
rect 20990 13676 20996 13688
rect 21048 13676 21054 13728
rect 22094 13676 22100 13728
rect 22152 13716 22158 13728
rect 22152 13688 22197 13716
rect 22152 13676 22158 13688
rect 1104 13626 23276 13648
rect 1104 13574 8379 13626
rect 8431 13574 8443 13626
rect 8495 13574 8507 13626
rect 8559 13574 8571 13626
rect 8623 13574 15776 13626
rect 15828 13574 15840 13626
rect 15892 13574 15904 13626
rect 15956 13574 15968 13626
rect 16020 13574 23276 13626
rect 1104 13552 23276 13574
rect 1394 13472 1400 13524
rect 1452 13512 1458 13524
rect 2593 13515 2651 13521
rect 2593 13512 2605 13515
rect 1452 13484 2605 13512
rect 1452 13472 1458 13484
rect 2593 13481 2605 13484
rect 2639 13481 2651 13515
rect 2593 13475 2651 13481
rect 2685 13515 2743 13521
rect 2685 13481 2697 13515
rect 2731 13512 2743 13515
rect 3142 13512 3148 13524
rect 2731 13484 3148 13512
rect 2731 13481 2743 13484
rect 2685 13475 2743 13481
rect 3142 13472 3148 13484
rect 3200 13472 3206 13524
rect 3605 13515 3663 13521
rect 3605 13481 3617 13515
rect 3651 13512 3663 13515
rect 5350 13512 5356 13524
rect 3651 13484 5356 13512
rect 3651 13481 3663 13484
rect 3605 13475 3663 13481
rect 5350 13472 5356 13484
rect 5408 13472 5414 13524
rect 5718 13472 5724 13524
rect 5776 13512 5782 13524
rect 5813 13515 5871 13521
rect 5813 13512 5825 13515
rect 5776 13484 5825 13512
rect 5776 13472 5782 13484
rect 5813 13481 5825 13484
rect 5859 13481 5871 13515
rect 6914 13512 6920 13524
rect 5813 13475 5871 13481
rect 6104 13484 6920 13512
rect 4700 13447 4758 13453
rect 4700 13413 4712 13447
rect 4746 13444 4758 13447
rect 4982 13444 4988 13456
rect 4746 13416 4988 13444
rect 4746 13413 4758 13416
rect 4700 13407 4758 13413
rect 4982 13404 4988 13416
rect 5040 13404 5046 13456
rect 6104 13453 6132 13484
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 7374 13472 7380 13524
rect 7432 13512 7438 13524
rect 8757 13515 8815 13521
rect 8757 13512 8769 13515
rect 7432 13484 8769 13512
rect 7432 13472 7438 13484
rect 8757 13481 8769 13484
rect 8803 13481 8815 13515
rect 9306 13512 9312 13524
rect 9267 13484 9312 13512
rect 8757 13475 8815 13481
rect 9306 13472 9312 13484
rect 9364 13472 9370 13524
rect 9861 13515 9919 13521
rect 9861 13481 9873 13515
rect 9907 13512 9919 13515
rect 9907 13484 10732 13512
rect 9907 13481 9919 13484
rect 9861 13475 9919 13481
rect 6089 13447 6147 13453
rect 6089 13413 6101 13447
rect 6135 13413 6147 13447
rect 6270 13444 6276 13456
rect 6231 13416 6276 13444
rect 6089 13407 6147 13413
rect 6270 13404 6276 13416
rect 6328 13404 6334 13456
rect 7006 13453 7012 13456
rect 7000 13444 7012 13453
rect 6967 13416 7012 13444
rect 7000 13407 7012 13416
rect 7006 13404 7012 13407
rect 7064 13404 7070 13456
rect 7190 13404 7196 13456
rect 7248 13444 7254 13456
rect 8297 13447 8355 13453
rect 8297 13444 8309 13447
rect 7248 13416 8309 13444
rect 7248 13404 7254 13416
rect 8297 13413 8309 13416
rect 8343 13413 8355 13447
rect 8297 13407 8355 13413
rect 8938 13404 8944 13456
rect 8996 13404 9002 13456
rect 10704 13444 10732 13484
rect 10778 13472 10784 13524
rect 10836 13512 10842 13524
rect 10836 13484 19012 13512
rect 10836 13472 10842 13484
rect 11790 13444 11796 13456
rect 10704 13416 11796 13444
rect 11790 13404 11796 13416
rect 11848 13404 11854 13456
rect 12406 13447 12464 13453
rect 12406 13444 12418 13447
rect 12268 13416 12418 13444
rect 1670 13376 1676 13388
rect 1631 13348 1676 13376
rect 1670 13336 1676 13348
rect 1728 13336 1734 13388
rect 3421 13379 3479 13385
rect 3421 13345 3433 13379
rect 3467 13376 3479 13379
rect 7282 13376 7288 13388
rect 3467 13348 7288 13376
rect 3467 13345 3479 13348
rect 3421 13339 3479 13345
rect 7282 13336 7288 13348
rect 7340 13376 7346 13388
rect 8478 13376 8484 13388
rect 7340 13348 8484 13376
rect 7340 13336 7346 13348
rect 8478 13336 8484 13348
rect 8536 13336 8542 13388
rect 8956 13376 8984 13404
rect 9306 13376 9312 13388
rect 8956 13348 9312 13376
rect 9306 13336 9312 13348
rect 9364 13336 9370 13388
rect 10229 13379 10287 13385
rect 10229 13345 10241 13379
rect 10275 13376 10287 13379
rect 10956 13379 11014 13385
rect 10956 13376 10968 13379
rect 10275 13348 10968 13376
rect 10275 13345 10287 13348
rect 10229 13339 10287 13345
rect 10956 13345 10968 13348
rect 11002 13376 11014 13379
rect 11698 13376 11704 13388
rect 11002 13348 11704 13376
rect 11002 13345 11014 13348
rect 10956 13339 11014 13345
rect 11698 13336 11704 13348
rect 11756 13336 11762 13388
rect 12158 13376 12164 13388
rect 12119 13348 12164 13376
rect 12158 13336 12164 13348
rect 12216 13336 12222 13388
rect 2682 13268 2688 13320
rect 2740 13308 2746 13320
rect 2777 13311 2835 13317
rect 2777 13308 2789 13311
rect 2740 13280 2789 13308
rect 2740 13268 2746 13280
rect 2777 13277 2789 13280
rect 2823 13277 2835 13311
rect 2777 13271 2835 13277
rect 4338 13268 4344 13320
rect 4396 13308 4402 13320
rect 4433 13311 4491 13317
rect 4433 13308 4445 13311
rect 4396 13280 4445 13308
rect 4396 13268 4402 13280
rect 4433 13277 4445 13280
rect 4479 13277 4491 13311
rect 6730 13308 6736 13320
rect 6691 13280 6736 13308
rect 4433 13271 4491 13277
rect 6730 13268 6736 13280
rect 6788 13268 6794 13320
rect 8849 13311 8907 13317
rect 8849 13277 8861 13311
rect 8895 13277 8907 13311
rect 8849 13271 8907 13277
rect 1854 13240 1860 13252
rect 1815 13212 1860 13240
rect 1854 13200 1860 13212
rect 1912 13200 1918 13252
rect 5534 13200 5540 13252
rect 5592 13240 5598 13252
rect 6457 13243 6515 13249
rect 6457 13240 6469 13243
rect 5592 13212 6469 13240
rect 5592 13200 5598 13212
rect 6457 13209 6469 13212
rect 6503 13209 6515 13243
rect 8864 13240 8892 13271
rect 8938 13268 8944 13320
rect 8996 13308 9002 13320
rect 10321 13311 10379 13317
rect 8996 13280 9041 13308
rect 8996 13268 9002 13280
rect 10321 13277 10333 13311
rect 10367 13277 10379 13311
rect 10321 13271 10379 13277
rect 10413 13311 10471 13317
rect 10413 13277 10425 13311
rect 10459 13308 10471 13311
rect 10594 13308 10600 13320
rect 10459 13280 10600 13308
rect 10459 13277 10471 13280
rect 10413 13271 10471 13277
rect 6457 13203 6515 13209
rect 7668 13212 8892 13240
rect 10336 13240 10364 13271
rect 10594 13268 10600 13280
rect 10652 13268 10658 13320
rect 10686 13268 10692 13320
rect 10744 13308 10750 13320
rect 12268 13308 12296 13416
rect 12406 13413 12418 13416
rect 12452 13413 12464 13447
rect 13722 13444 13728 13456
rect 12406 13407 12464 13413
rect 13464 13416 13728 13444
rect 13464 13388 13492 13416
rect 13722 13404 13728 13416
rect 13780 13404 13786 13456
rect 13814 13404 13820 13456
rect 13872 13453 13878 13456
rect 13872 13447 13936 13453
rect 13872 13413 13890 13447
rect 13924 13413 13936 13447
rect 13872 13407 13936 13413
rect 18224 13447 18282 13453
rect 18224 13413 18236 13447
rect 18270 13444 18282 13447
rect 18874 13444 18880 13456
rect 18270 13416 18880 13444
rect 18270 13413 18282 13416
rect 18224 13407 18282 13413
rect 13872 13404 13878 13407
rect 18874 13404 18880 13416
rect 18932 13404 18938 13456
rect 18984 13444 19012 13484
rect 19610 13472 19616 13524
rect 19668 13512 19674 13524
rect 20073 13515 20131 13521
rect 20073 13512 20085 13515
rect 19668 13484 20085 13512
rect 19668 13472 19674 13484
rect 20073 13481 20085 13484
rect 20119 13481 20131 13515
rect 20073 13475 20131 13481
rect 20901 13515 20959 13521
rect 20901 13481 20913 13515
rect 20947 13512 20959 13515
rect 22094 13512 22100 13524
rect 20947 13484 22100 13512
rect 20947 13481 20959 13484
rect 20901 13475 20959 13481
rect 22094 13472 22100 13484
rect 22152 13472 22158 13524
rect 20162 13444 20168 13456
rect 18984 13416 20168 13444
rect 20162 13404 20168 13416
rect 20220 13404 20226 13456
rect 21628 13447 21686 13453
rect 21628 13413 21640 13447
rect 21674 13444 21686 13447
rect 21910 13444 21916 13456
rect 21674 13416 21916 13444
rect 21674 13413 21686 13416
rect 21628 13407 21686 13413
rect 21910 13404 21916 13416
rect 21968 13404 21974 13456
rect 13446 13336 13452 13388
rect 13504 13336 13510 13388
rect 13633 13379 13691 13385
rect 13633 13345 13645 13379
rect 13679 13376 13691 13379
rect 14182 13376 14188 13388
rect 13679 13348 14188 13376
rect 13679 13345 13691 13348
rect 13633 13339 13691 13345
rect 14182 13336 14188 13348
rect 14240 13376 14246 13388
rect 14918 13376 14924 13388
rect 14240 13348 14924 13376
rect 14240 13336 14246 13348
rect 14918 13336 14924 13348
rect 14976 13336 14982 13388
rect 15289 13379 15347 13385
rect 15289 13345 15301 13379
rect 15335 13376 15347 13379
rect 15838 13376 15844 13388
rect 15335 13348 15844 13376
rect 15335 13345 15347 13348
rect 15289 13339 15347 13345
rect 15838 13336 15844 13348
rect 15896 13336 15902 13388
rect 16016 13379 16074 13385
rect 16016 13345 16028 13379
rect 16062 13376 16074 13379
rect 16298 13376 16304 13388
rect 16062 13348 16304 13376
rect 16062 13345 16074 13348
rect 16016 13339 16074 13345
rect 16298 13336 16304 13348
rect 16356 13336 16362 13388
rect 17405 13379 17463 13385
rect 17405 13345 17417 13379
rect 17451 13376 17463 13379
rect 18506 13376 18512 13388
rect 17451 13348 18512 13376
rect 17451 13345 17463 13348
rect 17405 13339 17463 13345
rect 18506 13336 18512 13348
rect 18564 13336 18570 13388
rect 19981 13379 20039 13385
rect 19981 13345 19993 13379
rect 20027 13376 20039 13379
rect 20346 13376 20352 13388
rect 20027 13348 20352 13376
rect 20027 13345 20039 13348
rect 19981 13339 20039 13345
rect 20346 13336 20352 13348
rect 20404 13336 20410 13388
rect 10744 13280 10789 13308
rect 12084 13280 12296 13308
rect 15749 13311 15807 13317
rect 10744 13268 10750 13280
rect 10502 13240 10508 13252
rect 10336 13212 10508 13240
rect 2225 13175 2283 13181
rect 2225 13141 2237 13175
rect 2271 13172 2283 13175
rect 3234 13172 3240 13184
rect 2271 13144 3240 13172
rect 2271 13141 2283 13144
rect 2225 13135 2283 13141
rect 3234 13132 3240 13144
rect 3292 13132 3298 13184
rect 4338 13132 4344 13184
rect 4396 13172 4402 13184
rect 7668 13172 7696 13212
rect 10502 13200 10508 13212
rect 10560 13200 10566 13252
rect 11974 13200 11980 13252
rect 12032 13240 12038 13252
rect 12084 13249 12112 13280
rect 15749 13277 15761 13311
rect 15795 13277 15807 13311
rect 17678 13308 17684 13320
rect 15749 13271 15807 13277
rect 16776 13280 17684 13308
rect 12069 13243 12127 13249
rect 12069 13240 12081 13243
rect 12032 13212 12081 13240
rect 12032 13200 12038 13212
rect 12069 13209 12081 13212
rect 12115 13209 12127 13243
rect 12069 13203 12127 13209
rect 8110 13172 8116 13184
rect 4396 13144 7696 13172
rect 8071 13144 8116 13172
rect 4396 13132 4402 13144
rect 8110 13132 8116 13144
rect 8168 13132 8174 13184
rect 8297 13175 8355 13181
rect 8297 13141 8309 13175
rect 8343 13172 8355 13175
rect 8389 13175 8447 13181
rect 8389 13172 8401 13175
rect 8343 13144 8401 13172
rect 8343 13141 8355 13144
rect 8297 13135 8355 13141
rect 8389 13141 8401 13144
rect 8435 13141 8447 13175
rect 8389 13135 8447 13141
rect 10042 13132 10048 13184
rect 10100 13172 10106 13184
rect 13541 13175 13599 13181
rect 13541 13172 13553 13175
rect 10100 13144 13553 13172
rect 10100 13132 10106 13144
rect 13541 13141 13553 13144
rect 13587 13141 13599 13175
rect 13541 13135 13599 13141
rect 14642 13132 14648 13184
rect 14700 13172 14706 13184
rect 15013 13175 15071 13181
rect 15013 13172 15025 13175
rect 14700 13144 15025 13172
rect 14700 13132 14706 13144
rect 15013 13141 15025 13144
rect 15059 13141 15071 13175
rect 15764 13172 15792 13271
rect 16776 13172 16804 13280
rect 17678 13268 17684 13280
rect 17736 13308 17742 13320
rect 17957 13311 18015 13317
rect 17957 13308 17969 13311
rect 17736 13280 17969 13308
rect 17736 13268 17742 13280
rect 17957 13277 17969 13280
rect 18003 13277 18015 13311
rect 20165 13311 20223 13317
rect 20165 13308 20177 13311
rect 17957 13271 18015 13277
rect 19904 13280 20177 13308
rect 16942 13200 16948 13252
rect 17000 13240 17006 13252
rect 17862 13240 17868 13252
rect 17000 13212 17868 13240
rect 17000 13200 17006 13212
rect 17862 13200 17868 13212
rect 17920 13200 17926 13252
rect 15764 13144 16804 13172
rect 17129 13175 17187 13181
rect 15013 13135 15071 13141
rect 17129 13141 17141 13175
rect 17175 13172 17187 13175
rect 17402 13172 17408 13184
rect 17175 13144 17408 13172
rect 17175 13141 17187 13144
rect 17129 13135 17187 13141
rect 17402 13132 17408 13144
rect 17460 13132 17466 13184
rect 17589 13175 17647 13181
rect 17589 13141 17601 13175
rect 17635 13172 17647 13175
rect 17678 13172 17684 13184
rect 17635 13144 17684 13172
rect 17635 13141 17647 13144
rect 17589 13135 17647 13141
rect 17678 13132 17684 13144
rect 17736 13132 17742 13184
rect 17972 13172 18000 13271
rect 19334 13240 19340 13252
rect 19247 13212 19340 13240
rect 19334 13200 19340 13212
rect 19392 13240 19398 13252
rect 19904 13240 19932 13280
rect 20165 13277 20177 13280
rect 20211 13277 20223 13311
rect 20165 13271 20223 13277
rect 20990 13268 20996 13320
rect 21048 13308 21054 13320
rect 21361 13311 21419 13317
rect 21361 13308 21373 13311
rect 21048 13280 21373 13308
rect 21048 13268 21054 13280
rect 21361 13277 21373 13280
rect 21407 13277 21419 13311
rect 21361 13271 21419 13277
rect 19392 13212 19932 13240
rect 19392 13200 19398 13212
rect 18598 13172 18604 13184
rect 17972 13144 18604 13172
rect 18598 13132 18604 13144
rect 18656 13132 18662 13184
rect 19613 13175 19671 13181
rect 19613 13141 19625 13175
rect 19659 13172 19671 13175
rect 19794 13172 19800 13184
rect 19659 13144 19800 13172
rect 19659 13141 19671 13144
rect 19613 13135 19671 13141
rect 19794 13132 19800 13144
rect 19852 13132 19858 13184
rect 22741 13175 22799 13181
rect 22741 13141 22753 13175
rect 22787 13172 22799 13175
rect 22830 13172 22836 13184
rect 22787 13144 22836 13172
rect 22787 13141 22799 13144
rect 22741 13135 22799 13141
rect 22830 13132 22836 13144
rect 22888 13132 22894 13184
rect 1104 13082 23276 13104
rect 1104 13030 4680 13082
rect 4732 13030 4744 13082
rect 4796 13030 4808 13082
rect 4860 13030 4872 13082
rect 4924 13030 12078 13082
rect 12130 13030 12142 13082
rect 12194 13030 12206 13082
rect 12258 13030 12270 13082
rect 12322 13030 19475 13082
rect 19527 13030 19539 13082
rect 19591 13030 19603 13082
rect 19655 13030 19667 13082
rect 19719 13030 23276 13082
rect 1104 13008 23276 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 4338 12968 4344 12980
rect 1627 12940 4344 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 4982 12968 4988 12980
rect 4943 12940 4988 12968
rect 4982 12928 4988 12940
rect 5040 12928 5046 12980
rect 8481 12971 8539 12977
rect 8481 12937 8493 12971
rect 8527 12937 8539 12971
rect 8481 12931 8539 12937
rect 5000 12832 5028 12928
rect 5350 12860 5356 12912
rect 5408 12900 5414 12912
rect 5408 12872 5856 12900
rect 5408 12860 5414 12872
rect 5828 12841 5856 12872
rect 8496 12844 8524 12931
rect 9122 12928 9128 12980
rect 9180 12968 9186 12980
rect 10318 12968 10324 12980
rect 9180 12940 10324 12968
rect 9180 12928 9186 12940
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 11698 12968 11704 12980
rect 11659 12940 11704 12968
rect 11698 12928 11704 12940
rect 11756 12928 11762 12980
rect 14185 12971 14243 12977
rect 11808 12940 13667 12968
rect 11330 12860 11336 12912
rect 11388 12900 11394 12912
rect 11808 12900 11836 12940
rect 11388 12872 11836 12900
rect 11388 12860 11394 12872
rect 5721 12835 5779 12841
rect 5721 12832 5733 12835
rect 5000 12804 5733 12832
rect 5721 12801 5733 12804
rect 5767 12801 5779 12835
rect 5721 12795 5779 12801
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12801 5871 12835
rect 5813 12795 5871 12801
rect 8478 12792 8484 12844
rect 8536 12792 8542 12844
rect 8938 12792 8944 12844
rect 8996 12832 9002 12844
rect 9033 12835 9091 12841
rect 9033 12832 9045 12835
rect 8996 12804 9045 12832
rect 8996 12792 9002 12804
rect 9033 12801 9045 12804
rect 9079 12801 9091 12835
rect 9033 12795 9091 12801
rect 9674 12792 9680 12844
rect 9732 12832 9738 12844
rect 10045 12835 10103 12841
rect 10045 12832 10057 12835
rect 9732 12804 10057 12832
rect 9732 12792 9738 12804
rect 10045 12801 10057 12804
rect 10091 12801 10103 12835
rect 13639 12832 13667 12940
rect 14185 12937 14197 12971
rect 14231 12968 14243 12971
rect 16390 12968 16396 12980
rect 14231 12940 16396 12968
rect 14231 12937 14243 12940
rect 14185 12931 14243 12937
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 17589 12971 17647 12977
rect 17589 12937 17601 12971
rect 17635 12968 17647 12971
rect 20441 12971 20499 12977
rect 20441 12968 20453 12971
rect 17635 12940 20453 12968
rect 17635 12937 17647 12940
rect 17589 12931 17647 12937
rect 20441 12937 20453 12940
rect 20487 12937 20499 12971
rect 20441 12931 20499 12937
rect 20622 12928 20628 12980
rect 20680 12968 20686 12980
rect 22373 12971 22431 12977
rect 22373 12968 22385 12971
rect 20680 12940 22385 12968
rect 20680 12928 20686 12940
rect 22373 12937 22385 12940
rect 22419 12937 22431 12971
rect 22373 12931 22431 12937
rect 13998 12900 14004 12912
rect 13959 12872 14004 12900
rect 13998 12860 14004 12872
rect 14056 12860 14062 12912
rect 14093 12903 14151 12909
rect 14093 12869 14105 12903
rect 14139 12900 14151 12903
rect 14139 12872 14688 12900
rect 14139 12869 14151 12872
rect 14093 12863 14151 12869
rect 14660 12841 14688 12872
rect 16298 12860 16304 12912
rect 16356 12900 16362 12912
rect 16577 12903 16635 12909
rect 16577 12900 16589 12903
rect 16356 12872 16589 12900
rect 16356 12860 16362 12872
rect 16577 12869 16589 12872
rect 16623 12869 16635 12903
rect 17681 12903 17739 12909
rect 17681 12900 17693 12903
rect 16577 12863 16635 12869
rect 16684 12872 17693 12900
rect 14645 12835 14703 12841
rect 13639 12804 14228 12832
rect 10045 12795 10103 12801
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12733 1455 12767
rect 1397 12727 1455 12733
rect 1412 12628 1440 12727
rect 1578 12724 1584 12776
rect 1636 12764 1642 12776
rect 1949 12767 2007 12773
rect 1949 12764 1961 12767
rect 1636 12736 1961 12764
rect 1636 12724 1642 12736
rect 1949 12733 1961 12736
rect 1995 12764 2007 12767
rect 3605 12767 3663 12773
rect 3605 12764 3617 12767
rect 1995 12736 3617 12764
rect 1995 12733 2007 12736
rect 1949 12727 2007 12733
rect 3605 12733 3617 12736
rect 3651 12764 3663 12767
rect 4338 12764 4344 12776
rect 3651 12736 4344 12764
rect 3651 12733 3663 12736
rect 3605 12727 3663 12733
rect 4338 12724 4344 12736
rect 4396 12724 4402 12776
rect 5534 12724 5540 12776
rect 5592 12764 5598 12776
rect 5629 12767 5687 12773
rect 5629 12764 5641 12767
rect 5592 12736 5641 12764
rect 5592 12724 5598 12736
rect 5629 12733 5641 12736
rect 5675 12733 5687 12767
rect 6273 12767 6331 12773
rect 6273 12764 6285 12767
rect 5629 12727 5687 12733
rect 5828 12736 6285 12764
rect 2216 12699 2274 12705
rect 2216 12665 2228 12699
rect 2262 12696 2274 12699
rect 2958 12696 2964 12708
rect 2262 12668 2964 12696
rect 2262 12665 2274 12668
rect 2216 12659 2274 12665
rect 2958 12656 2964 12668
rect 3016 12656 3022 12708
rect 3850 12699 3908 12705
rect 3850 12696 3862 12699
rect 3344 12668 3862 12696
rect 2866 12628 2872 12640
rect 1412 12600 2872 12628
rect 2866 12588 2872 12600
rect 2924 12588 2930 12640
rect 3344 12637 3372 12668
rect 3850 12665 3862 12668
rect 3896 12696 3908 12699
rect 4430 12696 4436 12708
rect 3896 12668 4436 12696
rect 3896 12665 3908 12668
rect 3850 12659 3908 12665
rect 4430 12656 4436 12668
rect 4488 12656 4494 12708
rect 5828 12696 5856 12736
rect 6273 12733 6285 12736
rect 6319 12733 6331 12767
rect 6822 12764 6828 12776
rect 6783 12736 6828 12764
rect 6273 12727 6331 12733
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 9861 12767 9919 12773
rect 9861 12764 9873 12767
rect 7024 12736 9873 12764
rect 7024 12696 7052 12736
rect 9861 12733 9873 12736
rect 9907 12733 9919 12767
rect 9861 12727 9919 12733
rect 10321 12767 10379 12773
rect 10321 12733 10333 12767
rect 10367 12733 10379 12767
rect 10321 12727 10379 12733
rect 10588 12767 10646 12773
rect 10588 12733 10600 12767
rect 10634 12764 10646 12767
rect 11698 12764 11704 12776
rect 10634 12736 11704 12764
rect 10634 12733 10646 12736
rect 10588 12727 10646 12733
rect 4543 12668 5856 12696
rect 6196 12668 7052 12696
rect 7092 12699 7150 12705
rect 3329 12631 3387 12637
rect 3329 12597 3341 12631
rect 3375 12597 3387 12631
rect 3329 12591 3387 12597
rect 3418 12588 3424 12640
rect 3476 12628 3482 12640
rect 4543 12628 4571 12668
rect 3476 12600 4571 12628
rect 5261 12631 5319 12637
rect 3476 12588 3482 12600
rect 5261 12597 5273 12631
rect 5307 12628 5319 12631
rect 6196 12628 6224 12668
rect 7092 12665 7104 12699
rect 7138 12696 7150 12699
rect 7466 12696 7472 12708
rect 7138 12668 7472 12696
rect 7138 12665 7150 12668
rect 7092 12659 7150 12665
rect 7466 12656 7472 12668
rect 7524 12656 7530 12708
rect 10336 12640 10364 12727
rect 10502 12656 10508 12708
rect 10560 12696 10566 12708
rect 10603 12696 10631 12727
rect 11698 12724 11704 12736
rect 11756 12724 11762 12776
rect 11882 12764 11888 12776
rect 11843 12736 11888 12764
rect 11882 12724 11888 12736
rect 11940 12724 11946 12776
rect 11974 12724 11980 12776
rect 12032 12764 12038 12776
rect 12069 12767 12127 12773
rect 12069 12764 12081 12767
rect 12032 12736 12081 12764
rect 12032 12724 12038 12736
rect 12069 12733 12081 12736
rect 12115 12733 12127 12767
rect 12069 12727 12127 12733
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 12621 12767 12679 12773
rect 12621 12764 12633 12767
rect 12492 12736 12633 12764
rect 12492 12724 12498 12736
rect 12621 12733 12633 12736
rect 12667 12733 12679 12767
rect 12621 12727 12679 12733
rect 13354 12724 13360 12776
rect 13412 12764 13418 12776
rect 14093 12767 14151 12773
rect 14093 12764 14105 12767
rect 13412 12736 14105 12764
rect 13412 12724 13418 12736
rect 14093 12733 14105 12736
rect 14139 12733 14151 12767
rect 14093 12727 14151 12733
rect 10560 12668 10631 12696
rect 10560 12656 10566 12668
rect 11514 12656 11520 12708
rect 11572 12656 11578 12708
rect 12888 12699 12946 12705
rect 12888 12665 12900 12699
rect 12934 12665 12946 12699
rect 12888 12659 12946 12665
rect 5307 12600 6224 12628
rect 5307 12597 5319 12600
rect 5261 12591 5319 12597
rect 7374 12588 7380 12640
rect 7432 12628 7438 12640
rect 8205 12631 8263 12637
rect 8205 12628 8217 12631
rect 7432 12600 8217 12628
rect 7432 12588 7438 12600
rect 8205 12597 8217 12600
rect 8251 12597 8263 12631
rect 8846 12628 8852 12640
rect 8807 12600 8852 12628
rect 8205 12591 8263 12597
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 8938 12588 8944 12640
rect 8996 12628 9002 12640
rect 8996 12600 9041 12628
rect 8996 12588 9002 12600
rect 9122 12588 9128 12640
rect 9180 12628 9186 12640
rect 9493 12631 9551 12637
rect 9493 12628 9505 12631
rect 9180 12600 9505 12628
rect 9180 12588 9186 12600
rect 9493 12597 9505 12600
rect 9539 12597 9551 12631
rect 9950 12628 9956 12640
rect 9911 12600 9956 12628
rect 9493 12591 9551 12597
rect 9950 12588 9956 12600
rect 10008 12588 10014 12640
rect 10318 12628 10324 12640
rect 10231 12600 10324 12628
rect 10318 12588 10324 12600
rect 10376 12628 10382 12640
rect 10686 12628 10692 12640
rect 10376 12600 10692 12628
rect 10376 12588 10382 12600
rect 10686 12588 10692 12600
rect 10744 12588 10750 12640
rect 11532 12628 11560 12656
rect 11882 12628 11888 12640
rect 11532 12600 11888 12628
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 11974 12588 11980 12640
rect 12032 12628 12038 12640
rect 12253 12631 12311 12637
rect 12253 12628 12265 12631
rect 12032 12600 12265 12628
rect 12032 12588 12038 12600
rect 12253 12597 12265 12600
rect 12299 12597 12311 12631
rect 12903 12628 12931 12659
rect 13262 12656 13268 12708
rect 13320 12696 13326 12708
rect 13722 12696 13728 12708
rect 13320 12668 13728 12696
rect 13320 12656 13326 12668
rect 13722 12656 13728 12668
rect 13780 12656 13786 12708
rect 14200 12696 14228 12804
rect 14645 12801 14657 12835
rect 14691 12801 14703 12835
rect 14645 12795 14703 12801
rect 14737 12835 14795 12841
rect 14737 12801 14749 12835
rect 14783 12801 14795 12835
rect 14737 12795 14795 12801
rect 14366 12724 14372 12776
rect 14424 12764 14430 12776
rect 14752 12764 14780 12795
rect 14424 12736 14780 12764
rect 14424 12724 14430 12736
rect 14918 12724 14924 12776
rect 14976 12764 14982 12776
rect 15197 12767 15255 12773
rect 15197 12764 15209 12767
rect 14976 12736 15209 12764
rect 14976 12724 14982 12736
rect 15197 12733 15209 12736
rect 15243 12764 15255 12767
rect 16684 12764 16712 12872
rect 17681 12869 17693 12872
rect 17727 12869 17739 12903
rect 17681 12863 17739 12869
rect 17862 12860 17868 12912
rect 17920 12860 17926 12912
rect 18230 12900 18236 12912
rect 18191 12872 18236 12900
rect 18230 12860 18236 12872
rect 18288 12860 18294 12912
rect 21177 12903 21235 12909
rect 21177 12869 21189 12903
rect 21223 12900 21235 12903
rect 22186 12900 22192 12912
rect 21223 12872 22192 12900
rect 21223 12869 21235 12872
rect 21177 12863 21235 12869
rect 22186 12860 22192 12872
rect 22244 12860 22250 12912
rect 16850 12792 16856 12844
rect 16908 12832 16914 12844
rect 17126 12832 17132 12844
rect 16908 12804 17132 12832
rect 16908 12792 16914 12804
rect 17126 12792 17132 12804
rect 17184 12792 17190 12844
rect 17313 12835 17371 12841
rect 17313 12801 17325 12835
rect 17359 12832 17371 12835
rect 17497 12835 17555 12841
rect 17497 12832 17509 12835
rect 17359 12804 17509 12832
rect 17359 12801 17371 12804
rect 17313 12795 17371 12801
rect 17497 12801 17509 12804
rect 17543 12801 17555 12835
rect 17497 12795 17555 12801
rect 17589 12835 17647 12841
rect 17589 12801 17601 12835
rect 17635 12801 17647 12835
rect 17880 12832 17908 12860
rect 17880 12804 18092 12832
rect 17589 12795 17647 12801
rect 15243 12736 16712 12764
rect 15243 12733 15255 12736
rect 15197 12727 15255 12733
rect 14553 12699 14611 12705
rect 14553 12696 14565 12699
rect 14200 12668 14565 12696
rect 14553 12665 14565 12668
rect 14599 12665 14611 12699
rect 14553 12659 14611 12665
rect 15378 12656 15384 12708
rect 15436 12705 15442 12708
rect 15436 12699 15500 12705
rect 15436 12665 15454 12699
rect 15488 12665 15500 12699
rect 17037 12699 17095 12705
rect 17037 12696 17049 12699
rect 15436 12659 15500 12665
rect 15571 12668 17049 12696
rect 15436 12656 15442 12659
rect 13906 12628 13912 12640
rect 12903 12600 13912 12628
rect 12253 12591 12311 12597
rect 13906 12588 13912 12600
rect 13964 12588 13970 12640
rect 14918 12588 14924 12640
rect 14976 12628 14982 12640
rect 15571 12628 15599 12668
rect 17037 12665 17049 12668
rect 17083 12665 17095 12699
rect 17037 12659 17095 12665
rect 17129 12699 17187 12705
rect 17129 12665 17141 12699
rect 17175 12696 17187 12699
rect 17604 12696 17632 12795
rect 17862 12764 17868 12776
rect 17823 12736 17868 12764
rect 17862 12724 17868 12736
rect 17920 12724 17926 12776
rect 18064 12773 18092 12804
rect 20898 12792 20904 12844
rect 20956 12832 20962 12844
rect 21637 12835 21695 12841
rect 21637 12832 21649 12835
rect 20956 12804 21649 12832
rect 20956 12792 20962 12804
rect 21637 12801 21649 12804
rect 21683 12832 21695 12835
rect 21726 12832 21732 12844
rect 21683 12804 21732 12832
rect 21683 12801 21695 12804
rect 21637 12795 21695 12801
rect 21726 12792 21732 12804
rect 21784 12792 21790 12844
rect 21821 12835 21879 12841
rect 21821 12801 21833 12835
rect 21867 12832 21879 12835
rect 22002 12832 22008 12844
rect 21867 12804 22008 12832
rect 21867 12801 21879 12804
rect 21821 12795 21879 12801
rect 22002 12792 22008 12804
rect 22060 12792 22066 12844
rect 18049 12767 18107 12773
rect 18049 12733 18061 12767
rect 18095 12733 18107 12767
rect 18598 12764 18604 12776
rect 18511 12736 18604 12764
rect 18049 12727 18107 12733
rect 18598 12724 18604 12736
rect 18656 12724 18662 12776
rect 18868 12767 18926 12773
rect 18868 12733 18880 12767
rect 18914 12764 18926 12767
rect 19334 12764 19340 12776
rect 18914 12736 19340 12764
rect 18914 12733 18926 12736
rect 18868 12727 18926 12733
rect 19334 12724 19340 12736
rect 19392 12724 19398 12776
rect 20162 12724 20168 12776
rect 20220 12764 20226 12776
rect 20257 12767 20315 12773
rect 20257 12764 20269 12767
rect 20220 12736 20269 12764
rect 20220 12724 20226 12736
rect 20257 12733 20269 12736
rect 20303 12733 20315 12767
rect 20257 12727 20315 12733
rect 22189 12767 22247 12773
rect 22189 12733 22201 12767
rect 22235 12764 22247 12767
rect 22235 12736 22784 12764
rect 22235 12733 22247 12736
rect 22189 12727 22247 12733
rect 17175 12668 17632 12696
rect 17175 12665 17187 12668
rect 17129 12659 17187 12665
rect 14976 12600 15599 12628
rect 14976 12588 14982 12600
rect 16574 12588 16580 12640
rect 16632 12628 16638 12640
rect 16669 12631 16727 12637
rect 16669 12628 16681 12631
rect 16632 12600 16681 12628
rect 16632 12588 16638 12600
rect 16669 12597 16681 12600
rect 16715 12597 16727 12631
rect 16669 12591 16727 12597
rect 17218 12588 17224 12640
rect 17276 12628 17282 12640
rect 17497 12631 17555 12637
rect 17497 12628 17509 12631
rect 17276 12600 17509 12628
rect 17276 12588 17282 12600
rect 17497 12597 17509 12600
rect 17543 12597 17555 12631
rect 17497 12591 17555 12597
rect 17862 12588 17868 12640
rect 17920 12628 17926 12640
rect 18616 12628 18644 12724
rect 18690 12656 18696 12708
rect 18748 12696 18754 12708
rect 19702 12696 19708 12708
rect 18748 12668 19708 12696
rect 18748 12656 18754 12668
rect 19702 12656 19708 12668
rect 19760 12656 19766 12708
rect 20990 12696 20996 12708
rect 19812 12668 20996 12696
rect 19812 12628 19840 12668
rect 20990 12656 20996 12668
rect 21048 12656 21054 12708
rect 22756 12640 22784 12736
rect 19978 12628 19984 12640
rect 17920 12600 19840 12628
rect 19939 12600 19984 12628
rect 17920 12588 17926 12600
rect 19978 12588 19984 12600
rect 20036 12588 20042 12640
rect 20346 12588 20352 12640
rect 20404 12628 20410 12640
rect 21545 12631 21603 12637
rect 21545 12628 21557 12631
rect 20404 12600 21557 12628
rect 20404 12588 20410 12600
rect 21545 12597 21557 12600
rect 21591 12597 21603 12631
rect 21545 12591 21603 12597
rect 22738 12588 22744 12640
rect 22796 12588 22802 12640
rect 1104 12538 23276 12560
rect 1104 12486 8379 12538
rect 8431 12486 8443 12538
rect 8495 12486 8507 12538
rect 8559 12486 8571 12538
rect 8623 12486 15776 12538
rect 15828 12486 15840 12538
rect 15892 12486 15904 12538
rect 15956 12486 15968 12538
rect 16020 12486 23276 12538
rect 1104 12464 23276 12486
rect 2958 12424 2964 12436
rect 2919 12396 2964 12424
rect 2958 12384 2964 12396
rect 3016 12384 3022 12436
rect 3605 12427 3663 12433
rect 3605 12393 3617 12427
rect 3651 12393 3663 12427
rect 4430 12424 4436 12436
rect 4391 12396 4436 12424
rect 3605 12387 3663 12393
rect 3620 12356 3648 12387
rect 4430 12384 4436 12396
rect 4488 12384 4494 12436
rect 5721 12427 5779 12433
rect 5721 12393 5733 12427
rect 5767 12424 5779 12427
rect 6914 12424 6920 12436
rect 5767 12396 6920 12424
rect 5767 12393 5779 12396
rect 5721 12387 5779 12393
rect 6914 12384 6920 12396
rect 6972 12384 6978 12436
rect 8202 12424 8208 12436
rect 7031 12396 8208 12424
rect 5534 12356 5540 12368
rect 3620 12328 5540 12356
rect 5534 12316 5540 12328
rect 5592 12316 5598 12368
rect 5810 12316 5816 12368
rect 5868 12356 5874 12368
rect 6638 12356 6644 12368
rect 5868 12328 5913 12356
rect 6472 12328 6644 12356
rect 5868 12316 5874 12328
rect 1578 12288 1584 12300
rect 1539 12260 1584 12288
rect 1578 12248 1584 12260
rect 1636 12248 1642 12300
rect 1848 12291 1906 12297
rect 1848 12257 1860 12291
rect 1894 12288 1906 12291
rect 2774 12288 2780 12300
rect 1894 12260 2780 12288
rect 1894 12257 1906 12260
rect 1848 12251 1906 12257
rect 2774 12248 2780 12260
rect 2832 12248 2838 12300
rect 3421 12291 3479 12297
rect 3421 12257 3433 12291
rect 3467 12288 3479 12291
rect 5074 12288 5080 12300
rect 3467 12260 5080 12288
rect 3467 12257 3479 12260
rect 3421 12251 3479 12257
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 6472 12297 6500 12328
rect 6638 12316 6644 12328
rect 6696 12316 6702 12368
rect 6822 12316 6828 12368
rect 6880 12356 6886 12368
rect 7031 12356 7059 12396
rect 8202 12384 8208 12396
rect 8260 12424 8266 12436
rect 8665 12427 8723 12433
rect 8665 12424 8677 12427
rect 8260 12396 8677 12424
rect 8260 12384 8266 12396
rect 8665 12393 8677 12396
rect 8711 12393 8723 12427
rect 8665 12387 8723 12393
rect 9122 12384 9128 12436
rect 9180 12424 9186 12436
rect 9217 12427 9275 12433
rect 9217 12424 9229 12427
rect 9180 12396 9229 12424
rect 9180 12384 9186 12396
rect 9217 12393 9229 12396
rect 9263 12424 9275 12427
rect 9306 12424 9312 12436
rect 9263 12396 9312 12424
rect 9263 12393 9275 12396
rect 9217 12387 9275 12393
rect 9306 12384 9312 12396
rect 9364 12384 9370 12436
rect 9858 12384 9864 12436
rect 9916 12424 9922 12436
rect 9953 12427 10011 12433
rect 9953 12424 9965 12427
rect 9916 12396 9965 12424
rect 9916 12384 9922 12396
rect 9953 12393 9965 12396
rect 9999 12393 10011 12427
rect 9953 12387 10011 12393
rect 10505 12427 10563 12433
rect 10505 12393 10517 12427
rect 10551 12424 10563 12427
rect 10781 12427 10839 12433
rect 10781 12424 10793 12427
rect 10551 12396 10793 12424
rect 10551 12393 10563 12396
rect 10505 12387 10563 12393
rect 10781 12393 10793 12396
rect 10827 12393 10839 12427
rect 11422 12424 11428 12436
rect 10781 12387 10839 12393
rect 10980 12396 11428 12424
rect 6880 12328 7059 12356
rect 6880 12316 6886 12328
rect 7031 12297 7059 12328
rect 7276 12359 7334 12365
rect 7276 12325 7288 12359
rect 7322 12356 7334 12359
rect 7374 12356 7380 12368
rect 7322 12328 7380 12356
rect 7322 12325 7334 12328
rect 7276 12319 7334 12325
rect 7374 12316 7380 12328
rect 7432 12316 7438 12368
rect 7742 12316 7748 12368
rect 7800 12356 7806 12368
rect 8018 12356 8024 12368
rect 7800 12328 8024 12356
rect 7800 12316 7806 12328
rect 8018 12316 8024 12328
rect 8076 12316 8082 12368
rect 10980 12356 11008 12396
rect 11422 12384 11428 12396
rect 11480 12384 11486 12436
rect 13446 12384 13452 12436
rect 13504 12384 13510 12436
rect 14090 12384 14096 12436
rect 14148 12424 14154 12436
rect 14645 12427 14703 12433
rect 14645 12424 14657 12427
rect 14148 12396 14657 12424
rect 14148 12384 14154 12396
rect 14645 12393 14657 12396
rect 14691 12393 14703 12427
rect 14645 12387 14703 12393
rect 14734 12384 14740 12436
rect 14792 12424 14798 12436
rect 14921 12427 14979 12433
rect 14921 12424 14933 12427
rect 14792 12396 14933 12424
rect 14792 12384 14798 12396
rect 14921 12393 14933 12396
rect 14967 12424 14979 12427
rect 14967 12396 15608 12424
rect 14967 12393 14979 12396
rect 14921 12387 14979 12393
rect 9048 12328 11008 12356
rect 9048 12297 9076 12328
rect 5261 12291 5319 12297
rect 5261 12257 5273 12291
rect 5307 12288 5319 12291
rect 6457 12291 6515 12297
rect 5307 12260 6408 12288
rect 5307 12257 5319 12260
rect 5261 12251 5319 12257
rect 6380 12232 6408 12260
rect 6457 12257 6469 12291
rect 6503 12257 6515 12291
rect 6457 12251 6515 12257
rect 7009 12291 7067 12297
rect 7009 12257 7021 12291
rect 7055 12257 7067 12291
rect 8849 12291 8907 12297
rect 8849 12288 8861 12291
rect 7009 12251 7067 12257
rect 7107 12260 8861 12288
rect 2958 12180 2964 12232
rect 3016 12220 3022 12232
rect 4525 12223 4583 12229
rect 4525 12220 4537 12223
rect 3016 12192 4537 12220
rect 3016 12180 3022 12192
rect 4525 12189 4537 12192
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12220 4767 12223
rect 4893 12223 4951 12229
rect 4893 12220 4905 12223
rect 4755 12192 4905 12220
rect 4755 12189 4767 12192
rect 4709 12183 4767 12189
rect 4893 12189 4905 12192
rect 4939 12220 4951 12223
rect 5350 12220 5356 12232
rect 4939 12192 5356 12220
rect 4939 12189 4951 12192
rect 4893 12183 4951 12189
rect 5350 12180 5356 12192
rect 5408 12220 5414 12232
rect 5905 12223 5963 12229
rect 5905 12220 5917 12223
rect 5408 12192 5917 12220
rect 5408 12180 5414 12192
rect 5905 12189 5917 12192
rect 5951 12189 5963 12223
rect 5905 12183 5963 12189
rect 6362 12180 6368 12232
rect 6420 12180 6426 12232
rect 7107 12220 7135 12260
rect 8849 12257 8861 12260
rect 8895 12257 8907 12291
rect 8849 12251 8907 12257
rect 9033 12291 9091 12297
rect 9033 12257 9045 12291
rect 9079 12257 9091 12291
rect 9033 12251 9091 12257
rect 9214 12248 9220 12300
rect 9272 12248 9278 12300
rect 9766 12288 9772 12300
rect 9727 12260 9772 12288
rect 9766 12248 9772 12260
rect 9824 12248 9830 12300
rect 10689 12291 10747 12297
rect 10689 12257 10701 12291
rect 10735 12257 10747 12291
rect 10689 12251 10747 12257
rect 10781 12291 10839 12297
rect 10781 12257 10793 12291
rect 10827 12288 10839 12291
rect 10962 12288 10968 12300
rect 10827 12260 10968 12288
rect 10827 12257 10839 12260
rect 10781 12251 10839 12257
rect 6472 12192 7135 12220
rect 3510 12112 3516 12164
rect 3568 12152 3574 12164
rect 5077 12155 5135 12161
rect 5077 12152 5089 12155
rect 3568 12124 5089 12152
rect 3568 12112 3574 12124
rect 5077 12121 5089 12124
rect 5123 12152 5135 12155
rect 6472 12152 6500 12192
rect 9232 12152 9260 12248
rect 10704 12220 10732 12251
rect 10962 12248 10968 12260
rect 11020 12248 11026 12300
rect 11149 12291 11207 12297
rect 11149 12257 11161 12291
rect 11195 12288 11207 12291
rect 11241 12291 11299 12297
rect 11241 12288 11253 12291
rect 11195 12260 11253 12288
rect 11195 12257 11207 12260
rect 11149 12251 11207 12257
rect 11241 12257 11253 12260
rect 11287 12257 11299 12291
rect 11241 12251 11299 12257
rect 11333 12291 11391 12297
rect 11333 12257 11345 12291
rect 11379 12288 11391 12291
rect 11425 12291 11483 12297
rect 11425 12288 11437 12291
rect 11379 12260 11437 12288
rect 11379 12257 11391 12260
rect 11333 12251 11391 12257
rect 11425 12257 11437 12260
rect 11471 12257 11483 12291
rect 13464 12288 13492 12384
rect 15286 12316 15292 12368
rect 15344 12316 15350 12368
rect 13521 12291 13579 12297
rect 13521 12288 13533 12291
rect 13464 12260 13533 12288
rect 11425 12251 11483 12257
rect 13521 12257 13533 12260
rect 13567 12257 13579 12291
rect 13521 12251 13579 12257
rect 13998 12248 14004 12300
rect 14056 12288 14062 12300
rect 15105 12291 15163 12297
rect 15105 12288 15117 12291
rect 14056 12260 15117 12288
rect 14056 12248 14062 12260
rect 15105 12257 15117 12260
rect 15151 12257 15163 12291
rect 15105 12251 15163 12257
rect 13170 12220 13176 12232
rect 10704 12192 13176 12220
rect 13170 12180 13176 12192
rect 13228 12180 13234 12232
rect 13265 12223 13323 12229
rect 13265 12189 13277 12223
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 11333 12155 11391 12161
rect 11333 12152 11345 12155
rect 5123 12124 6500 12152
rect 7944 12124 9260 12152
rect 9324 12124 11345 12152
rect 5123 12121 5135 12124
rect 5077 12115 5135 12121
rect 4062 12084 4068 12096
rect 4023 12056 4068 12084
rect 4062 12044 4068 12056
rect 4120 12044 4126 12096
rect 4430 12044 4436 12096
rect 4488 12084 4494 12096
rect 4893 12087 4951 12093
rect 4893 12084 4905 12087
rect 4488 12056 4905 12084
rect 4488 12044 4494 12056
rect 4893 12053 4905 12056
rect 4939 12053 4951 12087
rect 5350 12084 5356 12096
rect 5311 12056 5356 12084
rect 4893 12047 4951 12053
rect 5350 12044 5356 12056
rect 5408 12044 5414 12096
rect 6641 12087 6699 12093
rect 6641 12053 6653 12087
rect 6687 12084 6699 12087
rect 7944 12084 7972 12124
rect 8386 12084 8392 12096
rect 6687 12056 7972 12084
rect 8347 12056 8392 12084
rect 6687 12053 6699 12056
rect 6641 12047 6699 12053
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 8570 12044 8576 12096
rect 8628 12084 8634 12096
rect 9324 12084 9352 12124
rect 11333 12121 11345 12124
rect 11379 12121 11391 12155
rect 11333 12115 11391 12121
rect 8628 12056 9352 12084
rect 8628 12044 8634 12056
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 10965 12087 11023 12093
rect 10965 12084 10977 12087
rect 9732 12056 10977 12084
rect 9732 12044 9738 12056
rect 10965 12053 10977 12056
rect 11011 12053 11023 12087
rect 10965 12047 11023 12053
rect 11241 12087 11299 12093
rect 11241 12053 11253 12087
rect 11287 12084 11299 12087
rect 12526 12084 12532 12096
rect 11287 12056 12532 12084
rect 11287 12053 11299 12056
rect 11241 12047 11299 12053
rect 12526 12044 12532 12056
rect 12584 12084 12590 12096
rect 12713 12087 12771 12093
rect 12713 12084 12725 12087
rect 12584 12056 12725 12084
rect 12584 12044 12590 12056
rect 12713 12053 12725 12056
rect 12759 12053 12771 12087
rect 13280 12084 13308 12183
rect 14274 12180 14280 12232
rect 14332 12220 14338 12232
rect 15304 12220 15332 12316
rect 15470 12288 15476 12300
rect 15431 12260 15476 12288
rect 15470 12248 15476 12260
rect 15528 12248 15534 12300
rect 14332 12192 15332 12220
rect 15580 12220 15608 12396
rect 15654 12384 15660 12436
rect 15712 12424 15718 12436
rect 16390 12424 16396 12436
rect 15712 12396 15757 12424
rect 16351 12396 16396 12424
rect 15712 12384 15718 12396
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 17037 12427 17095 12433
rect 17037 12393 17049 12427
rect 17083 12424 17095 12427
rect 17083 12396 20484 12424
rect 17083 12393 17095 12396
rect 17037 12387 17095 12393
rect 20456 12368 20484 12396
rect 16485 12359 16543 12365
rect 16485 12356 16497 12359
rect 16224 12328 16497 12356
rect 15746 12248 15752 12300
rect 15804 12288 15810 12300
rect 16224 12288 16252 12328
rect 16485 12325 16497 12328
rect 16531 12325 16543 12359
rect 17862 12356 17868 12368
rect 16485 12319 16543 12325
rect 17512 12328 17868 12356
rect 17218 12288 17224 12300
rect 15804 12260 16252 12288
rect 16316 12260 17224 12288
rect 15804 12248 15810 12260
rect 16316 12220 16344 12260
rect 17218 12248 17224 12260
rect 17276 12248 17282 12300
rect 17512 12297 17540 12328
rect 17862 12316 17868 12328
rect 17920 12316 17926 12368
rect 19886 12316 19892 12368
rect 19944 12356 19950 12368
rect 19944 12328 20208 12356
rect 19944 12316 19950 12328
rect 17497 12291 17555 12297
rect 17497 12257 17509 12291
rect 17543 12257 17555 12291
rect 17497 12251 17555 12257
rect 17764 12291 17822 12297
rect 17764 12257 17776 12291
rect 17810 12288 17822 12291
rect 18690 12288 18696 12300
rect 17810 12260 18696 12288
rect 17810 12257 17822 12260
rect 17764 12251 17822 12257
rect 18690 12248 18696 12260
rect 18748 12248 18754 12300
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 19794 12288 19800 12300
rect 19392 12260 19800 12288
rect 19392 12248 19398 12260
rect 19794 12248 19800 12260
rect 19852 12248 19858 12300
rect 20180 12232 20208 12328
rect 20438 12316 20444 12368
rect 20496 12316 20502 12368
rect 20901 12291 20959 12297
rect 20901 12257 20913 12291
rect 20947 12288 20959 12291
rect 20990 12288 20996 12300
rect 20947 12260 20996 12288
rect 20947 12257 20959 12260
rect 20901 12251 20959 12257
rect 20990 12248 20996 12260
rect 21048 12248 21054 12300
rect 21174 12297 21180 12300
rect 21168 12251 21180 12297
rect 21232 12288 21238 12300
rect 21232 12260 21268 12288
rect 21174 12248 21180 12251
rect 21232 12248 21238 12260
rect 16577 12223 16635 12229
rect 16577 12220 16589 12223
rect 15580 12192 16344 12220
rect 16408 12192 16589 12220
rect 14332 12180 14338 12192
rect 15470 12112 15476 12164
rect 15528 12152 15534 12164
rect 16408 12152 16436 12192
rect 16577 12189 16589 12192
rect 16623 12189 16635 12223
rect 19886 12220 19892 12232
rect 19847 12192 19892 12220
rect 16577 12183 16635 12189
rect 19886 12180 19892 12192
rect 19944 12180 19950 12232
rect 19978 12180 19984 12232
rect 20036 12220 20042 12232
rect 20036 12192 20081 12220
rect 20036 12180 20042 12192
rect 20162 12180 20168 12232
rect 20220 12180 20226 12232
rect 22554 12220 22560 12232
rect 22515 12192 22560 12220
rect 22554 12180 22560 12192
rect 22612 12180 22618 12232
rect 15528 12124 16436 12152
rect 15528 12112 15534 12124
rect 18782 12112 18788 12164
rect 18840 12152 18846 12164
rect 18877 12155 18935 12161
rect 18877 12152 18889 12155
rect 18840 12124 18889 12152
rect 18840 12112 18846 12124
rect 18877 12121 18889 12124
rect 18923 12121 18935 12155
rect 18877 12115 18935 12121
rect 14182 12084 14188 12096
rect 13280 12056 14188 12084
rect 12713 12047 12771 12053
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 15286 12044 15292 12096
rect 15344 12084 15350 12096
rect 16025 12087 16083 12093
rect 16025 12084 16037 12087
rect 15344 12056 16037 12084
rect 15344 12044 15350 12056
rect 16025 12053 16037 12056
rect 16071 12053 16083 12087
rect 16025 12047 16083 12053
rect 19429 12087 19487 12093
rect 19429 12053 19441 12087
rect 19475 12084 19487 12087
rect 21634 12084 21640 12096
rect 19475 12056 21640 12084
rect 19475 12053 19487 12056
rect 19429 12047 19487 12053
rect 21634 12044 21640 12056
rect 21692 12044 21698 12096
rect 21818 12044 21824 12096
rect 21876 12084 21882 12096
rect 22002 12084 22008 12096
rect 21876 12056 22008 12084
rect 21876 12044 21882 12056
rect 22002 12044 22008 12056
rect 22060 12084 22066 12096
rect 22281 12087 22339 12093
rect 22281 12084 22293 12087
rect 22060 12056 22293 12084
rect 22060 12044 22066 12056
rect 22281 12053 22293 12056
rect 22327 12053 22339 12087
rect 22281 12047 22339 12053
rect 1104 11994 23276 12016
rect 1104 11942 4680 11994
rect 4732 11942 4744 11994
rect 4796 11942 4808 11994
rect 4860 11942 4872 11994
rect 4924 11942 12078 11994
rect 12130 11942 12142 11994
rect 12194 11942 12206 11994
rect 12258 11942 12270 11994
rect 12322 11942 19475 11994
rect 19527 11942 19539 11994
rect 19591 11942 19603 11994
rect 19655 11942 19667 11994
rect 19719 11942 23276 11994
rect 1104 11920 23276 11942
rect 6457 11883 6515 11889
rect 6457 11880 6469 11883
rect 3528 11852 6469 11880
rect 3326 11704 3332 11756
rect 3384 11744 3390 11756
rect 3528 11753 3556 11852
rect 6457 11849 6469 11852
rect 6503 11849 6515 11883
rect 8849 11883 8907 11889
rect 8849 11880 8861 11883
rect 6457 11843 6515 11849
rect 7208 11852 8861 11880
rect 4338 11772 4344 11824
rect 4396 11812 4402 11824
rect 4396 11784 4936 11812
rect 4396 11772 4402 11784
rect 3513 11747 3571 11753
rect 3513 11744 3525 11747
rect 3384 11716 3525 11744
rect 3384 11704 3390 11716
rect 3513 11713 3525 11716
rect 3559 11713 3571 11747
rect 3513 11707 3571 11713
rect 3697 11747 3755 11753
rect 3697 11713 3709 11747
rect 3743 11744 3755 11747
rect 4430 11744 4436 11756
rect 3743 11716 4436 11744
rect 3743 11713 3755 11716
rect 3697 11707 3755 11713
rect 4430 11704 4436 11716
rect 4488 11744 4494 11756
rect 4706 11744 4712 11756
rect 4488 11716 4712 11744
rect 4488 11704 4494 11716
rect 4706 11704 4712 11716
rect 4764 11704 4770 11756
rect 4908 11688 4936 11784
rect 6362 11772 6368 11824
rect 6420 11812 6426 11824
rect 7208 11812 7236 11852
rect 8849 11849 8861 11852
rect 8895 11849 8907 11883
rect 8849 11843 8907 11849
rect 9309 11883 9367 11889
rect 9309 11849 9321 11883
rect 9355 11880 9367 11883
rect 10686 11880 10692 11892
rect 9355 11852 10692 11880
rect 9355 11849 9367 11852
rect 9309 11843 9367 11849
rect 6420 11784 7236 11812
rect 8864 11812 8892 11843
rect 10686 11840 10692 11852
rect 10744 11840 10750 11892
rect 11698 11880 11704 11892
rect 11659 11852 11704 11880
rect 11698 11840 11704 11852
rect 11756 11840 11762 11892
rect 12618 11840 12624 11892
rect 12676 11880 12682 11892
rect 12802 11880 12808 11892
rect 12676 11852 12808 11880
rect 12676 11840 12682 11852
rect 12802 11840 12808 11852
rect 12860 11840 12866 11892
rect 13170 11840 13176 11892
rect 13228 11880 13234 11892
rect 13909 11883 13967 11889
rect 13909 11880 13921 11883
rect 13228 11852 13921 11880
rect 13228 11840 13234 11852
rect 13909 11849 13921 11852
rect 13955 11880 13967 11883
rect 13998 11880 14004 11892
rect 13955 11852 14004 11880
rect 13955 11849 13967 11852
rect 13909 11843 13967 11849
rect 13998 11840 14004 11852
rect 14056 11840 14062 11892
rect 14182 11840 14188 11892
rect 14240 11880 14246 11892
rect 14826 11880 14832 11892
rect 14240 11852 14832 11880
rect 14240 11840 14246 11852
rect 14826 11840 14832 11852
rect 14884 11840 14890 11892
rect 14918 11840 14924 11892
rect 14976 11880 14982 11892
rect 15194 11880 15200 11892
rect 14976 11852 15200 11880
rect 14976 11840 14982 11852
rect 15194 11840 15200 11852
rect 15252 11840 15258 11892
rect 15473 11883 15531 11889
rect 15473 11849 15485 11883
rect 15519 11880 15531 11883
rect 16114 11880 16120 11892
rect 15519 11852 16120 11880
rect 15519 11849 15531 11852
rect 15473 11843 15531 11849
rect 16114 11840 16120 11852
rect 16172 11840 16178 11892
rect 16758 11840 16764 11892
rect 16816 11880 16822 11892
rect 17310 11880 17316 11892
rect 16816 11852 17316 11880
rect 16816 11840 16822 11852
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 20898 11880 20904 11892
rect 19076 11852 20484 11880
rect 20859 11852 20904 11880
rect 9766 11812 9772 11824
rect 8864 11784 9772 11812
rect 6420 11772 6426 11784
rect 9766 11772 9772 11784
rect 9824 11772 9830 11824
rect 11606 11772 11612 11824
rect 11664 11812 11670 11824
rect 12161 11815 12219 11821
rect 12161 11812 12173 11815
rect 11664 11784 12173 11812
rect 11664 11772 11670 11784
rect 12161 11781 12173 11784
rect 12207 11781 12219 11815
rect 12161 11775 12219 11781
rect 12526 11772 12532 11824
rect 12584 11812 12590 11824
rect 15933 11815 15991 11821
rect 15933 11812 15945 11815
rect 12584 11784 15945 11812
rect 12584 11772 12590 11784
rect 15933 11781 15945 11784
rect 15979 11781 15991 11815
rect 15933 11775 15991 11781
rect 16390 11772 16396 11824
rect 16448 11812 16454 11824
rect 16666 11812 16672 11824
rect 16448 11784 16672 11812
rect 16448 11772 16454 11784
rect 16666 11772 16672 11784
rect 16724 11772 16730 11824
rect 6822 11704 6828 11756
rect 6880 11744 6886 11756
rect 7193 11747 7251 11753
rect 7193 11744 7205 11747
rect 6880 11716 7205 11744
rect 6880 11704 6886 11716
rect 7193 11713 7205 11716
rect 7239 11713 7251 11747
rect 7193 11707 7251 11713
rect 8662 11704 8668 11756
rect 8720 11744 8726 11756
rect 8846 11744 8852 11756
rect 8720 11716 8852 11744
rect 8720 11704 8726 11716
rect 8846 11704 8852 11716
rect 8904 11704 8910 11756
rect 9858 11744 9864 11756
rect 9819 11716 9864 11744
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 10318 11744 10324 11756
rect 10279 11716 10324 11744
rect 10318 11704 10324 11716
rect 10376 11704 10382 11756
rect 15105 11747 15163 11753
rect 11440 11716 14964 11744
rect 1394 11676 1400 11688
rect 1355 11648 1400 11676
rect 1394 11636 1400 11648
rect 1452 11636 1458 11688
rect 1664 11679 1722 11685
rect 1664 11645 1676 11679
rect 1710 11676 1722 11679
rect 2958 11676 2964 11688
rect 1710 11648 2964 11676
rect 1710 11645 1722 11648
rect 1664 11639 1722 11645
rect 2958 11636 2964 11648
rect 3016 11676 3022 11688
rect 4525 11679 4583 11685
rect 4525 11676 4537 11679
rect 3016 11648 4537 11676
rect 3016 11636 3022 11648
rect 4525 11645 4537 11648
rect 4571 11645 4583 11679
rect 4525 11639 4583 11645
rect 4890 11636 4896 11688
rect 4948 11676 4954 11688
rect 5077 11679 5135 11685
rect 5077 11676 5089 11679
rect 4948 11648 5089 11676
rect 4948 11636 4954 11648
rect 5077 11645 5089 11648
rect 5123 11676 5135 11679
rect 6840 11676 6868 11704
rect 9030 11676 9036 11688
rect 5123 11648 6868 11676
rect 8991 11648 9036 11676
rect 5123 11645 5135 11648
rect 5077 11639 5135 11645
rect 9030 11636 9036 11648
rect 9088 11636 9094 11688
rect 10962 11636 10968 11688
rect 11020 11676 11026 11688
rect 11440 11676 11468 11716
rect 11974 11676 11980 11688
rect 11020 11648 11468 11676
rect 11935 11648 11980 11676
rect 11020 11636 11026 11648
rect 11974 11636 11980 11648
rect 12032 11636 12038 11688
rect 14826 11676 14832 11688
rect 14787 11648 14832 11676
rect 14826 11636 14832 11648
rect 14884 11636 14890 11688
rect 14936 11676 14964 11716
rect 15105 11713 15117 11747
rect 15151 11744 15163 11747
rect 15654 11744 15660 11756
rect 15151 11716 15660 11744
rect 15151 11713 15163 11716
rect 15105 11707 15163 11713
rect 15654 11704 15660 11716
rect 15712 11704 15718 11756
rect 16022 11704 16028 11756
rect 16080 11744 16086 11756
rect 16485 11747 16543 11753
rect 16485 11744 16497 11747
rect 16080 11716 16497 11744
rect 16080 11704 16086 11716
rect 16485 11713 16497 11716
rect 16531 11713 16543 11747
rect 17494 11744 17500 11756
rect 17455 11716 17500 11744
rect 16485 11707 16543 11713
rect 17494 11704 17500 11716
rect 17552 11704 17558 11756
rect 18690 11744 18696 11756
rect 18603 11716 18696 11744
rect 18690 11704 18696 11716
rect 18748 11744 18754 11756
rect 19076 11744 19104 11852
rect 20456 11812 20484 11852
rect 20898 11840 20904 11852
rect 20956 11840 20962 11892
rect 22741 11883 22799 11889
rect 22741 11880 22753 11883
rect 21008 11852 22753 11880
rect 21008 11812 21036 11852
rect 22741 11849 22753 11852
rect 22787 11849 22799 11883
rect 22741 11843 22799 11849
rect 20456 11784 21036 11812
rect 18748 11716 19104 11744
rect 18748 11704 18754 11716
rect 19242 11704 19248 11756
rect 19300 11704 19306 11756
rect 19524 11747 19582 11753
rect 19524 11713 19536 11747
rect 19570 11744 19582 11747
rect 19702 11744 19708 11756
rect 19570 11716 19708 11744
rect 19570 11713 19582 11716
rect 19524 11707 19582 11713
rect 19702 11704 19708 11716
rect 19760 11704 19766 11756
rect 15289 11679 15347 11685
rect 15289 11676 15301 11679
rect 14936 11648 15301 11676
rect 15289 11645 15301 11648
rect 15335 11645 15347 11679
rect 15289 11639 15347 11645
rect 16758 11636 16764 11688
rect 16816 11676 16822 11688
rect 17405 11679 17463 11685
rect 17405 11676 17417 11679
rect 16816 11648 17417 11676
rect 16816 11636 16822 11648
rect 17405 11645 17417 11648
rect 17451 11645 17463 11679
rect 17405 11639 17463 11645
rect 18417 11679 18475 11685
rect 18417 11645 18429 11679
rect 18463 11676 18475 11679
rect 18598 11676 18604 11688
rect 18463 11648 18604 11676
rect 18463 11645 18475 11648
rect 18417 11639 18475 11645
rect 18598 11636 18604 11648
rect 18656 11636 18662 11688
rect 19058 11676 19064 11688
rect 18971 11648 19064 11676
rect 19058 11636 19064 11648
rect 19116 11676 19122 11688
rect 19260 11676 19288 11704
rect 19116 11648 19288 11676
rect 19797 11679 19855 11685
rect 19116 11636 19122 11648
rect 19797 11645 19809 11679
rect 19843 11676 19855 11679
rect 19886 11676 19892 11688
rect 19843 11648 19892 11676
rect 19843 11645 19855 11648
rect 19797 11639 19855 11645
rect 19886 11636 19892 11648
rect 19944 11636 19950 11688
rect 21266 11636 21272 11688
rect 21324 11676 21330 11688
rect 21361 11679 21419 11685
rect 21361 11676 21373 11679
rect 21324 11648 21373 11676
rect 21324 11636 21330 11648
rect 21361 11645 21373 11648
rect 21407 11645 21419 11679
rect 21361 11639 21419 11645
rect 4433 11611 4491 11617
rect 4433 11608 4445 11611
rect 2976 11580 4445 11608
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 2976 11540 3004 11580
rect 4433 11577 4445 11580
rect 4479 11577 4491 11611
rect 4433 11571 4491 11577
rect 5344 11611 5402 11617
rect 5344 11577 5356 11611
rect 5390 11608 5402 11611
rect 6914 11608 6920 11620
rect 5390 11580 6920 11608
rect 5390 11577 5402 11580
rect 5344 11571 5402 11577
rect 6914 11568 6920 11580
rect 6972 11568 6978 11620
rect 7466 11617 7472 11620
rect 7460 11608 7472 11617
rect 7427 11580 7472 11608
rect 7460 11571 7472 11580
rect 7524 11608 7530 11620
rect 8386 11608 8392 11620
rect 7524 11580 8392 11608
rect 7466 11568 7472 11571
rect 7524 11568 7530 11580
rect 8386 11568 8392 11580
rect 8444 11568 8450 11620
rect 9677 11611 9735 11617
rect 9677 11577 9689 11611
rect 9723 11608 9735 11611
rect 10588 11611 10646 11617
rect 10588 11608 10600 11611
rect 9723 11580 10600 11608
rect 9723 11577 9735 11580
rect 9677 11571 9735 11577
rect 10588 11577 10600 11580
rect 10634 11608 10646 11611
rect 11790 11608 11796 11620
rect 10634 11580 11796 11608
rect 10634 11577 10646 11580
rect 10588 11571 10646 11577
rect 11790 11568 11796 11580
rect 11848 11568 11854 11620
rect 12621 11611 12679 11617
rect 12621 11577 12633 11611
rect 12667 11608 12679 11611
rect 13170 11608 13176 11620
rect 12667 11580 13176 11608
rect 12667 11577 12679 11580
rect 12621 11571 12679 11577
rect 13170 11568 13176 11580
rect 13228 11568 13234 11620
rect 14642 11568 14648 11620
rect 14700 11608 14706 11620
rect 14921 11611 14979 11617
rect 14921 11608 14933 11611
rect 14700 11580 14933 11608
rect 14700 11568 14706 11580
rect 14921 11577 14933 11580
rect 14967 11577 14979 11611
rect 14921 11571 14979 11577
rect 17313 11611 17371 11617
rect 17313 11577 17325 11611
rect 17359 11608 17371 11611
rect 18690 11608 18696 11620
rect 17359 11580 18696 11608
rect 17359 11577 17371 11580
rect 17313 11571 17371 11577
rect 18690 11568 18696 11580
rect 18748 11568 18754 11620
rect 21628 11611 21686 11617
rect 21628 11577 21640 11611
rect 21674 11608 21686 11611
rect 22646 11608 22652 11620
rect 21674 11580 22652 11608
rect 21674 11577 21686 11580
rect 21628 11571 21686 11577
rect 22646 11568 22652 11580
rect 22704 11568 22710 11620
rect 2832 11512 3004 11540
rect 2832 11500 2838 11512
rect 3050 11500 3056 11552
rect 3108 11540 3114 11552
rect 3418 11540 3424 11552
rect 3108 11512 3153 11540
rect 3379 11512 3424 11540
rect 3108 11500 3114 11512
rect 3418 11500 3424 11512
rect 3476 11500 3482 11552
rect 3694 11500 3700 11552
rect 3752 11540 3758 11552
rect 4065 11543 4123 11549
rect 4065 11540 4077 11543
rect 3752 11512 4077 11540
rect 3752 11500 3758 11512
rect 4065 11509 4077 11512
rect 4111 11509 4123 11543
rect 4065 11503 4123 11509
rect 7834 11500 7840 11552
rect 7892 11540 7898 11552
rect 8573 11543 8631 11549
rect 8573 11540 8585 11543
rect 7892 11512 8585 11540
rect 7892 11500 7898 11512
rect 8573 11509 8585 11512
rect 8619 11509 8631 11543
rect 8573 11503 8631 11509
rect 8754 11500 8760 11552
rect 8812 11540 8818 11552
rect 9030 11540 9036 11552
rect 8812 11512 9036 11540
rect 8812 11500 8818 11512
rect 9030 11500 9036 11512
rect 9088 11500 9094 11552
rect 9769 11543 9827 11549
rect 9769 11509 9781 11543
rect 9815 11540 9827 11543
rect 11422 11540 11428 11552
rect 9815 11512 11428 11540
rect 9815 11509 9827 11512
rect 9769 11503 9827 11509
rect 11422 11500 11428 11512
rect 11480 11500 11486 11552
rect 11606 11500 11612 11552
rect 11664 11540 11670 11552
rect 14461 11543 14519 11549
rect 14461 11540 14473 11543
rect 11664 11512 14473 11540
rect 11664 11500 11670 11512
rect 14461 11509 14473 11512
rect 14507 11509 14519 11543
rect 14461 11503 14519 11509
rect 16114 11500 16120 11552
rect 16172 11540 16178 11552
rect 16301 11543 16359 11549
rect 16301 11540 16313 11543
rect 16172 11512 16313 11540
rect 16172 11500 16178 11512
rect 16301 11509 16313 11512
rect 16347 11509 16359 11543
rect 16301 11503 16359 11509
rect 16390 11500 16396 11552
rect 16448 11540 16454 11552
rect 16942 11540 16948 11552
rect 16448 11512 16493 11540
rect 16903 11512 16948 11540
rect 16448 11500 16454 11512
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 18046 11540 18052 11552
rect 18007 11512 18052 11540
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 18509 11543 18567 11549
rect 18509 11509 18521 11543
rect 18555 11540 18567 11543
rect 19334 11540 19340 11552
rect 18555 11512 19340 11540
rect 18555 11509 18567 11512
rect 18509 11503 18567 11509
rect 19334 11500 19340 11512
rect 19392 11500 19398 11552
rect 19426 11500 19432 11552
rect 19484 11540 19490 11552
rect 19527 11543 19585 11549
rect 19527 11540 19539 11543
rect 19484 11512 19539 11540
rect 19484 11500 19490 11512
rect 19527 11509 19539 11512
rect 19573 11540 19585 11543
rect 20070 11540 20076 11552
rect 19573 11512 20076 11540
rect 19573 11509 19585 11512
rect 19527 11503 19585 11509
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 1104 11450 23276 11472
rect 1104 11398 8379 11450
rect 8431 11398 8443 11450
rect 8495 11398 8507 11450
rect 8559 11398 8571 11450
rect 8623 11398 15776 11450
rect 15828 11398 15840 11450
rect 15892 11398 15904 11450
rect 15956 11398 15968 11450
rect 16020 11398 23276 11450
rect 1104 11376 23276 11398
rect 2777 11339 2835 11345
rect 2777 11305 2789 11339
rect 2823 11336 2835 11339
rect 2958 11336 2964 11348
rect 2823 11308 2964 11336
rect 2823 11305 2835 11308
rect 2777 11299 2835 11305
rect 2958 11296 2964 11308
rect 3016 11296 3022 11348
rect 3142 11296 3148 11348
rect 3200 11336 3206 11348
rect 3418 11336 3424 11348
rect 3200 11308 3424 11336
rect 3200 11296 3206 11308
rect 3418 11296 3424 11308
rect 3476 11296 3482 11348
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 4120 11308 4476 11336
rect 4120 11296 4126 11308
rect 3510 11268 3516 11280
rect 3344 11240 3516 11268
rect 1664 11203 1722 11209
rect 1664 11169 1676 11203
rect 1710 11200 1722 11203
rect 3142 11200 3148 11212
rect 1710 11172 3148 11200
rect 1710 11169 1722 11172
rect 1664 11163 1722 11169
rect 3142 11160 3148 11172
rect 3200 11160 3206 11212
rect 3344 11209 3372 11240
rect 3510 11228 3516 11240
rect 3568 11228 3574 11280
rect 4448 11268 4476 11308
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 6549 11339 6607 11345
rect 6549 11336 6561 11339
rect 5868 11308 6561 11336
rect 5868 11296 5874 11308
rect 6549 11305 6561 11308
rect 6595 11305 6607 11339
rect 6549 11299 6607 11305
rect 7742 11296 7748 11348
rect 7800 11336 7806 11348
rect 8665 11339 8723 11345
rect 8665 11336 8677 11339
rect 7800 11308 8677 11336
rect 7800 11296 7806 11308
rect 8665 11305 8677 11308
rect 8711 11305 8723 11339
rect 8665 11299 8723 11305
rect 9217 11339 9275 11345
rect 9217 11305 9229 11339
rect 9263 11305 9275 11339
rect 9217 11299 9275 11305
rect 10045 11339 10103 11345
rect 10045 11305 10057 11339
rect 10091 11336 10103 11339
rect 10410 11336 10416 11348
rect 10091 11308 10416 11336
rect 10091 11305 10103 11308
rect 10045 11299 10103 11305
rect 9232 11268 9260 11299
rect 10410 11296 10416 11308
rect 10468 11296 10474 11348
rect 11790 11336 11796 11348
rect 11751 11308 11796 11336
rect 11790 11296 11796 11308
rect 11848 11296 11854 11348
rect 12621 11339 12679 11345
rect 12621 11305 12633 11339
rect 12667 11336 12679 11339
rect 14274 11336 14280 11348
rect 12667 11308 14280 11336
rect 12667 11305 12679 11308
rect 12621 11299 12679 11305
rect 14274 11296 14280 11308
rect 14332 11296 14338 11348
rect 14829 11339 14887 11345
rect 14829 11305 14841 11339
rect 14875 11336 14887 11339
rect 15194 11336 15200 11348
rect 14875 11308 15200 11336
rect 14875 11305 14887 11308
rect 14829 11299 14887 11305
rect 15194 11296 15200 11308
rect 15252 11296 15258 11348
rect 17129 11339 17187 11345
rect 17129 11305 17141 11339
rect 17175 11305 17187 11339
rect 17129 11299 17187 11305
rect 11054 11268 11060 11280
rect 4448 11240 9168 11268
rect 9232 11240 11060 11268
rect 3329 11203 3387 11209
rect 3329 11169 3341 11203
rect 3375 11169 3387 11203
rect 3329 11163 3387 11169
rect 3418 11160 3424 11212
rect 3476 11200 3482 11212
rect 4430 11200 4436 11212
rect 3476 11172 3521 11200
rect 4391 11172 4436 11200
rect 3476 11160 3482 11172
rect 4430 11160 4436 11172
rect 4488 11160 4494 11212
rect 4890 11160 4896 11212
rect 4948 11200 4954 11212
rect 5169 11203 5227 11209
rect 5169 11200 5181 11203
rect 4948 11172 5181 11200
rect 4948 11160 4954 11172
rect 5169 11169 5181 11172
rect 5215 11169 5227 11203
rect 5169 11163 5227 11169
rect 5436 11203 5494 11209
rect 5436 11169 5448 11203
rect 5482 11200 5494 11203
rect 6454 11200 6460 11212
rect 5482 11172 6460 11200
rect 5482 11169 5494 11172
rect 5436 11163 5494 11169
rect 6454 11160 6460 11172
rect 6512 11160 6518 11212
rect 6638 11160 6644 11212
rect 6696 11200 6702 11212
rect 7285 11203 7343 11209
rect 7285 11200 7297 11203
rect 6696 11172 7297 11200
rect 6696 11160 6702 11172
rect 7285 11169 7297 11172
rect 7331 11169 7343 11203
rect 7285 11163 7343 11169
rect 7552 11203 7610 11209
rect 7552 11169 7564 11203
rect 7598 11200 7610 11203
rect 7834 11200 7840 11212
rect 7598 11172 7840 11200
rect 7598 11169 7610 11172
rect 7552 11163 7610 11169
rect 7834 11160 7840 11172
rect 7892 11160 7898 11212
rect 7926 11160 7932 11212
rect 7984 11200 7990 11212
rect 9033 11203 9091 11209
rect 9033 11200 9045 11203
rect 7984 11172 9045 11200
rect 7984 11160 7990 11172
rect 9033 11169 9045 11172
rect 9079 11169 9091 11203
rect 9140 11200 9168 11240
rect 11054 11228 11060 11240
rect 11112 11228 11118 11280
rect 11698 11228 11704 11280
rect 11756 11268 11762 11280
rect 17144 11268 17172 11299
rect 17218 11296 17224 11348
rect 17276 11296 17282 11348
rect 18423 11339 18481 11345
rect 18423 11305 18435 11339
rect 18469 11336 18481 11339
rect 19426 11336 19432 11348
rect 18469 11308 19432 11336
rect 18469 11305 18481 11308
rect 18423 11299 18481 11305
rect 19426 11296 19432 11308
rect 19484 11296 19490 11348
rect 19797 11339 19855 11345
rect 19797 11305 19809 11339
rect 19843 11336 19855 11339
rect 19886 11336 19892 11348
rect 19843 11308 19892 11336
rect 19843 11305 19855 11308
rect 19797 11299 19855 11305
rect 19886 11296 19892 11308
rect 19944 11296 19950 11348
rect 20254 11296 20260 11348
rect 20312 11296 20318 11348
rect 22094 11296 22100 11348
rect 22152 11336 22158 11348
rect 22278 11336 22284 11348
rect 22152 11308 22284 11336
rect 22152 11296 22158 11308
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 22646 11336 22652 11348
rect 22607 11308 22652 11336
rect 22646 11296 22652 11308
rect 22704 11296 22710 11348
rect 11756 11240 17172 11268
rect 17236 11268 17264 11296
rect 20272 11268 20300 11296
rect 17236 11240 18000 11268
rect 11756 11228 11762 11240
rect 9674 11200 9680 11212
rect 9140 11172 9680 11200
rect 9033 11163 9091 11169
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 9861 11203 9919 11209
rect 9861 11169 9873 11203
rect 9907 11200 9919 11203
rect 10042 11200 10048 11212
rect 9907 11172 10048 11200
rect 9907 11169 9919 11172
rect 9861 11163 9919 11169
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 10318 11160 10324 11212
rect 10376 11200 10382 11212
rect 10413 11203 10471 11209
rect 10413 11200 10425 11203
rect 10376 11172 10425 11200
rect 10376 11160 10382 11172
rect 10413 11169 10425 11172
rect 10459 11169 10471 11203
rect 10413 11163 10471 11169
rect 10680 11203 10738 11209
rect 10680 11169 10692 11203
rect 10726 11200 10738 11203
rect 11422 11200 11428 11212
rect 10726 11172 11428 11200
rect 10726 11169 10738 11172
rect 10680 11163 10738 11169
rect 11422 11160 11428 11172
rect 11480 11160 11486 11212
rect 11514 11160 11520 11212
rect 11572 11200 11578 11212
rect 12253 11203 12311 11209
rect 12253 11200 12265 11203
rect 11572 11172 12265 11200
rect 11572 11160 11578 11172
rect 12253 11169 12265 11172
rect 12299 11169 12311 11203
rect 12253 11163 12311 11169
rect 12434 11160 12440 11212
rect 12492 11200 12498 11212
rect 12805 11203 12863 11209
rect 12805 11200 12817 11203
rect 12492 11172 12817 11200
rect 12492 11160 12498 11172
rect 12805 11169 12817 11172
rect 12851 11169 12863 11203
rect 12805 11163 12863 11169
rect 13072 11203 13130 11209
rect 13072 11169 13084 11203
rect 13118 11200 13130 11203
rect 13998 11200 14004 11212
rect 13118 11172 14004 11200
rect 13118 11169 13130 11172
rect 13072 11163 13130 11169
rect 13998 11160 14004 11172
rect 14056 11160 14062 11212
rect 14366 11160 14372 11212
rect 14424 11200 14430 11212
rect 15930 11209 15936 11212
rect 14645 11203 14703 11209
rect 14645 11200 14657 11203
rect 14424 11172 14657 11200
rect 14424 11160 14430 11172
rect 14645 11169 14657 11172
rect 14691 11169 14703 11203
rect 15913 11203 15936 11209
rect 15913 11200 15925 11203
rect 14645 11163 14703 11169
rect 14936 11172 15925 11200
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 4154 11092 4160 11144
rect 4212 11132 4218 11144
rect 4525 11135 4583 11141
rect 4525 11132 4537 11135
rect 4212 11104 4537 11132
rect 4212 11092 4218 11104
rect 4525 11101 4537 11104
rect 4571 11101 4583 11135
rect 4706 11132 4712 11144
rect 4667 11104 4712 11132
rect 4525 11095 4583 11101
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 6822 11132 6828 11144
rect 6783 11104 6828 11132
rect 6822 11092 6828 11104
rect 6880 11092 6886 11144
rect 8662 11092 8668 11144
rect 8720 11132 8726 11144
rect 8720 11104 10364 11132
rect 8720 11092 8726 11104
rect 4065 11067 4123 11073
rect 4065 11033 4077 11067
rect 4111 11064 4123 11067
rect 4338 11064 4344 11076
rect 4111 11036 4344 11064
rect 4111 11033 4123 11036
rect 4065 11027 4123 11033
rect 4338 11024 4344 11036
rect 4396 11024 4402 11076
rect 9950 11064 9956 11076
rect 9784 11036 9956 11064
rect 3145 10999 3203 11005
rect 3145 10965 3157 10999
rect 3191 10996 3203 10999
rect 3510 10996 3516 11008
rect 3191 10968 3516 10996
rect 3191 10965 3203 10968
rect 3145 10959 3203 10965
rect 3510 10956 3516 10968
rect 3568 10956 3574 11008
rect 3605 10999 3663 11005
rect 3605 10965 3617 10999
rect 3651 10996 3663 10999
rect 5534 10996 5540 11008
rect 3651 10968 5540 10996
rect 3651 10965 3663 10968
rect 3605 10959 3663 10965
rect 5534 10956 5540 10968
rect 5592 10956 5598 11008
rect 8570 10956 8576 11008
rect 8628 10996 8634 11008
rect 9784 10996 9812 11036
rect 9950 11024 9956 11036
rect 10008 11024 10014 11076
rect 8628 10968 9812 10996
rect 8628 10956 8634 10968
rect 10042 10956 10048 11008
rect 10100 10996 10106 11008
rect 10226 10996 10232 11008
rect 10100 10968 10232 10996
rect 10100 10956 10106 10968
rect 10226 10956 10232 10968
rect 10284 10956 10290 11008
rect 10336 10996 10364 11104
rect 12437 11067 12495 11073
rect 12437 11033 12449 11067
rect 12483 11064 12495 11067
rect 12621 11067 12679 11073
rect 12621 11064 12633 11067
rect 12483 11036 12633 11064
rect 12483 11033 12495 11036
rect 12437 11027 12495 11033
rect 12621 11033 12633 11036
rect 12667 11033 12679 11067
rect 14936 11064 14964 11172
rect 15913 11169 15925 11172
rect 15988 11200 15994 11212
rect 15988 11172 16061 11200
rect 15913 11163 15936 11169
rect 15930 11160 15936 11163
rect 15988 11160 15994 11172
rect 17218 11160 17224 11212
rect 17276 11200 17282 11212
rect 17497 11203 17555 11209
rect 17497 11200 17509 11203
rect 17276 11172 17509 11200
rect 17276 11160 17282 11172
rect 17497 11169 17509 11172
rect 17543 11169 17555 11203
rect 17497 11163 17555 11169
rect 17589 11203 17647 11209
rect 17589 11169 17601 11203
rect 17635 11200 17647 11203
rect 17862 11200 17868 11212
rect 17635 11172 17868 11200
rect 17635 11169 17647 11172
rect 17589 11163 17647 11169
rect 17862 11160 17868 11172
rect 17920 11160 17926 11212
rect 17972 11209 18000 11240
rect 19628 11240 20300 11268
rect 21536 11271 21594 11277
rect 17957 11203 18015 11209
rect 17957 11169 17969 11203
rect 18003 11200 18015 11203
rect 19058 11200 19064 11212
rect 18003 11172 19064 11200
rect 18003 11169 18015 11172
rect 17957 11163 18015 11169
rect 19058 11160 19064 11172
rect 19116 11200 19122 11212
rect 19334 11200 19340 11212
rect 19116 11172 19340 11200
rect 19116 11160 19122 11172
rect 19334 11160 19340 11172
rect 19392 11160 19398 11212
rect 15194 11092 15200 11144
rect 15252 11132 15258 11144
rect 15657 11135 15715 11141
rect 15657 11132 15669 11135
rect 15252 11104 15669 11132
rect 15252 11092 15258 11104
rect 15657 11101 15669 11104
rect 15703 11101 15715 11135
rect 17678 11132 17684 11144
rect 17639 11104 17684 11132
rect 15657 11095 15715 11101
rect 17678 11092 17684 11104
rect 17736 11092 17742 11144
rect 18414 11092 18420 11144
rect 18472 11132 18478 11144
rect 18472 11104 18517 11132
rect 18472 11092 18478 11104
rect 18598 11092 18604 11144
rect 18656 11132 18662 11144
rect 18693 11135 18751 11141
rect 18693 11132 18705 11135
rect 18656 11104 18705 11132
rect 18656 11092 18662 11104
rect 18693 11101 18705 11104
rect 18739 11101 18751 11135
rect 18693 11095 18751 11101
rect 12621 11027 12679 11033
rect 13740 11036 14964 11064
rect 13740 11008 13768 11036
rect 12986 10996 12992 11008
rect 10336 10968 12992 10996
rect 12986 10956 12992 10968
rect 13044 10956 13050 11008
rect 13722 10956 13728 11008
rect 13780 10956 13786 11008
rect 13906 10956 13912 11008
rect 13964 10996 13970 11008
rect 14185 10999 14243 11005
rect 14185 10996 14197 10999
rect 13964 10968 14197 10996
rect 13964 10956 13970 10968
rect 14185 10965 14197 10968
rect 14231 10965 14243 10999
rect 14185 10959 14243 10965
rect 14274 10956 14280 11008
rect 14332 10996 14338 11008
rect 17037 10999 17095 11005
rect 17037 10996 17049 10999
rect 14332 10968 17049 10996
rect 14332 10956 14338 10968
rect 17037 10965 17049 10968
rect 17083 10965 17095 10999
rect 17037 10959 17095 10965
rect 17218 10956 17224 11008
rect 17276 10996 17282 11008
rect 19628 10996 19656 11240
rect 21536 11237 21548 11271
rect 21582 11268 21594 11271
rect 21818 11268 21824 11280
rect 21582 11240 21824 11268
rect 21582 11237 21594 11240
rect 21536 11231 21594 11237
rect 21818 11228 21824 11240
rect 21876 11228 21882 11280
rect 20254 11200 20260 11212
rect 20215 11172 20260 11200
rect 20254 11160 20260 11172
rect 20312 11160 20318 11212
rect 20714 11092 20720 11144
rect 20772 11132 20778 11144
rect 21266 11132 21272 11144
rect 20772 11104 21272 11132
rect 20772 11092 20778 11104
rect 21266 11092 21272 11104
rect 21324 11092 21330 11144
rect 20346 11024 20352 11076
rect 20404 11064 20410 11076
rect 20441 11067 20499 11073
rect 20441 11064 20453 11067
rect 20404 11036 20453 11064
rect 20404 11024 20410 11036
rect 20441 11033 20453 11036
rect 20487 11033 20499 11067
rect 20441 11027 20499 11033
rect 17276 10968 19656 10996
rect 17276 10956 17282 10968
rect 1104 10906 23276 10928
rect 1104 10854 4680 10906
rect 4732 10854 4744 10906
rect 4796 10854 4808 10906
rect 4860 10854 4872 10906
rect 4924 10854 12078 10906
rect 12130 10854 12142 10906
rect 12194 10854 12206 10906
rect 12258 10854 12270 10906
rect 12322 10854 19475 10906
rect 19527 10854 19539 10906
rect 19591 10854 19603 10906
rect 19655 10854 19667 10906
rect 19719 10854 23276 10906
rect 1104 10832 23276 10854
rect 3142 10792 3148 10804
rect 3103 10764 3148 10792
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 4430 10752 4436 10804
rect 4488 10792 4494 10804
rect 4801 10795 4859 10801
rect 4801 10792 4813 10795
rect 4488 10764 4813 10792
rect 4488 10752 4494 10764
rect 4801 10761 4813 10764
rect 4847 10761 4859 10795
rect 6454 10792 6460 10804
rect 6415 10764 6460 10792
rect 4801 10755 4859 10761
rect 6454 10752 6460 10764
rect 6512 10752 6518 10804
rect 7009 10795 7067 10801
rect 7009 10761 7021 10795
rect 7055 10792 7067 10795
rect 7282 10792 7288 10804
rect 7055 10764 7288 10792
rect 7055 10761 7067 10764
rect 7009 10755 7067 10761
rect 7282 10752 7288 10764
rect 7340 10752 7346 10804
rect 8570 10792 8576 10804
rect 7392 10764 8576 10792
rect 1394 10548 1400 10600
rect 1452 10588 1458 10600
rect 1765 10591 1823 10597
rect 1765 10588 1777 10591
rect 1452 10560 1777 10588
rect 1452 10548 1458 10560
rect 1765 10557 1777 10560
rect 1811 10557 1823 10591
rect 1765 10551 1823 10557
rect 2032 10591 2090 10597
rect 2032 10557 2044 10591
rect 2078 10588 2090 10591
rect 3326 10588 3332 10600
rect 2078 10560 3332 10588
rect 2078 10557 2090 10560
rect 2032 10551 2090 10557
rect 1780 10520 1808 10551
rect 3326 10548 3332 10560
rect 3384 10548 3390 10600
rect 3421 10591 3479 10597
rect 3421 10557 3433 10591
rect 3467 10588 3479 10591
rect 3510 10588 3516 10600
rect 3467 10560 3516 10588
rect 3467 10557 3479 10560
rect 3421 10551 3479 10557
rect 3510 10548 3516 10560
rect 3568 10548 3574 10600
rect 3688 10591 3746 10597
rect 3688 10557 3700 10591
rect 3734 10588 3746 10591
rect 4154 10588 4160 10600
rect 3734 10560 4160 10588
rect 3734 10557 3746 10560
rect 3688 10551 3746 10557
rect 4154 10548 4160 10560
rect 4212 10548 4218 10600
rect 5077 10591 5135 10597
rect 5077 10557 5089 10591
rect 5123 10588 5135 10591
rect 5123 10560 5672 10588
rect 5123 10557 5135 10560
rect 5077 10551 5135 10557
rect 2130 10520 2136 10532
rect 1780 10492 2136 10520
rect 2130 10480 2136 10492
rect 2188 10480 2194 10532
rect 5344 10523 5402 10529
rect 5344 10489 5356 10523
rect 5390 10520 5402 10523
rect 5534 10520 5540 10532
rect 5390 10492 5540 10520
rect 5390 10489 5402 10492
rect 5344 10483 5402 10489
rect 5534 10480 5540 10492
rect 5592 10480 5598 10532
rect 5644 10520 5672 10560
rect 6270 10548 6276 10600
rect 6328 10588 6334 10600
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 6328 10560 6837 10588
rect 6328 10548 6334 10560
rect 6825 10557 6837 10560
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 6638 10520 6644 10532
rect 5644 10492 6644 10520
rect 6638 10480 6644 10492
rect 6696 10480 6702 10532
rect 3602 10412 3608 10464
rect 3660 10452 3666 10464
rect 7392 10452 7420 10764
rect 8570 10752 8576 10764
rect 8628 10752 8634 10804
rect 9309 10795 9367 10801
rect 9309 10761 9321 10795
rect 9355 10792 9367 10795
rect 9490 10792 9496 10804
rect 9355 10764 9496 10792
rect 9355 10761 9367 10764
rect 9309 10755 9367 10761
rect 9490 10752 9496 10764
rect 9548 10752 9554 10804
rect 10318 10792 10324 10804
rect 9968 10764 10324 10792
rect 9674 10724 9680 10736
rect 9635 10696 9680 10724
rect 9674 10684 9680 10696
rect 9732 10684 9738 10736
rect 9858 10684 9864 10736
rect 9916 10724 9922 10736
rect 9968 10724 9996 10764
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 10686 10752 10692 10804
rect 10744 10792 10750 10804
rect 10744 10764 10916 10792
rect 10744 10752 10750 10764
rect 9916 10696 9996 10724
rect 10888 10724 10916 10764
rect 11790 10752 11796 10804
rect 11848 10792 11854 10804
rect 17497 10795 17555 10801
rect 11848 10764 16804 10792
rect 11848 10752 11854 10764
rect 11977 10727 12035 10733
rect 11977 10724 11989 10727
rect 10888 10696 11989 10724
rect 9916 10684 9922 10696
rect 9968 10665 9996 10696
rect 11977 10693 11989 10696
rect 12023 10693 12035 10727
rect 11977 10687 12035 10693
rect 12434 10684 12440 10736
rect 12492 10724 12498 10736
rect 12492 10696 12572 10724
rect 12492 10684 12498 10696
rect 12544 10665 12572 10696
rect 15194 10684 15200 10736
rect 15252 10724 15258 10736
rect 16776 10724 16804 10764
rect 17497 10761 17509 10795
rect 17543 10792 17555 10795
rect 17678 10792 17684 10804
rect 17543 10764 17684 10792
rect 17543 10761 17555 10764
rect 17497 10755 17555 10761
rect 17678 10752 17684 10764
rect 17736 10752 17742 10804
rect 18233 10795 18291 10801
rect 18233 10761 18245 10795
rect 18279 10792 18291 10795
rect 18414 10792 18420 10804
rect 18279 10764 18420 10792
rect 18279 10761 18291 10764
rect 18233 10755 18291 10761
rect 18414 10752 18420 10764
rect 18472 10752 18478 10804
rect 21085 10795 21143 10801
rect 21085 10761 21097 10795
rect 21131 10792 21143 10795
rect 21174 10792 21180 10804
rect 21131 10764 21180 10792
rect 21131 10761 21143 10764
rect 21085 10755 21143 10761
rect 21174 10752 21180 10764
rect 21232 10752 21238 10804
rect 19058 10724 19064 10736
rect 15252 10696 15884 10724
rect 16776 10696 19064 10724
rect 15252 10684 15258 10696
rect 15856 10665 15884 10696
rect 19058 10684 19064 10696
rect 19116 10684 19122 10736
rect 9953 10659 10011 10665
rect 9953 10656 9965 10659
rect 8680 10628 9965 10656
rect 7469 10591 7527 10597
rect 7469 10557 7481 10591
rect 7515 10588 7527 10591
rect 8680 10588 8708 10628
rect 9953 10625 9965 10628
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 12529 10659 12587 10665
rect 12529 10625 12541 10659
rect 12575 10625 12587 10659
rect 15841 10659 15899 10665
rect 12529 10619 12587 10625
rect 13740 10628 14320 10656
rect 7515 10560 8708 10588
rect 7515 10557 7527 10560
rect 7469 10551 7527 10557
rect 8754 10548 8760 10600
rect 8812 10588 8818 10600
rect 9125 10591 9183 10597
rect 9125 10588 9137 10591
rect 8812 10560 9137 10588
rect 8812 10548 8818 10560
rect 9125 10557 9137 10560
rect 9171 10557 9183 10591
rect 9125 10551 9183 10557
rect 9766 10548 9772 10600
rect 9824 10588 9830 10600
rect 9861 10591 9919 10597
rect 9861 10588 9873 10591
rect 9824 10560 9873 10588
rect 9824 10548 9830 10560
rect 9861 10557 9873 10560
rect 9907 10557 9919 10591
rect 11146 10588 11152 10600
rect 9861 10551 9919 10557
rect 10060 10560 11152 10588
rect 7742 10529 7748 10532
rect 7736 10520 7748 10529
rect 7703 10492 7748 10520
rect 7736 10483 7748 10492
rect 7742 10480 7748 10483
rect 7800 10480 7806 10532
rect 9674 10480 9680 10532
rect 9732 10520 9738 10532
rect 10060 10520 10088 10560
rect 11146 10548 11152 10560
rect 11204 10548 11210 10600
rect 11793 10591 11851 10597
rect 11793 10557 11805 10591
rect 11839 10588 11851 10591
rect 12434 10588 12440 10600
rect 11839 10560 12440 10588
rect 11839 10557 11851 10560
rect 11793 10551 11851 10557
rect 12434 10548 12440 10560
rect 12492 10548 12498 10600
rect 10226 10529 10232 10532
rect 10220 10520 10232 10529
rect 9732 10492 10088 10520
rect 10187 10492 10232 10520
rect 9732 10480 9738 10492
rect 10220 10483 10232 10492
rect 10226 10480 10232 10483
rect 10284 10480 10290 10532
rect 12544 10520 12572 10619
rect 12618 10548 12624 10600
rect 12676 10588 12682 10600
rect 12785 10591 12843 10597
rect 12785 10588 12797 10591
rect 12676 10560 12797 10588
rect 12676 10548 12682 10560
rect 12785 10557 12797 10560
rect 12831 10588 12843 10591
rect 13740 10588 13768 10628
rect 14292 10600 14320 10628
rect 15841 10625 15853 10659
rect 15887 10625 15899 10659
rect 15841 10619 15899 10625
rect 14185 10591 14243 10597
rect 14185 10588 14197 10591
rect 12831 10560 13768 10588
rect 13823 10560 14197 10588
rect 12831 10557 12843 10560
rect 12785 10551 12843 10557
rect 13823 10520 13851 10560
rect 14185 10557 14197 10560
rect 14231 10557 14243 10591
rect 14185 10551 14243 10557
rect 14274 10548 14280 10600
rect 14332 10548 14338 10600
rect 15856 10588 15884 10619
rect 18046 10616 18052 10668
rect 18104 10656 18110 10668
rect 18693 10659 18751 10665
rect 18693 10656 18705 10659
rect 18104 10628 18705 10656
rect 18104 10616 18110 10628
rect 18693 10625 18705 10628
rect 18739 10625 18751 10659
rect 18874 10656 18880 10668
rect 18835 10628 18880 10656
rect 18693 10619 18751 10625
rect 18874 10616 18880 10628
rect 18932 10616 18938 10668
rect 21192 10656 21220 10752
rect 21913 10659 21971 10665
rect 21913 10656 21925 10659
rect 21192 10628 21925 10656
rect 21913 10625 21925 10628
rect 21959 10625 21971 10659
rect 21913 10619 21971 10625
rect 17313 10591 17371 10597
rect 15856 10560 16344 10588
rect 16316 10532 16344 10560
rect 17313 10557 17325 10591
rect 17359 10588 17371 10591
rect 19150 10588 19156 10600
rect 17359 10560 19156 10588
rect 17359 10557 17371 10560
rect 17313 10551 17371 10557
rect 19150 10548 19156 10560
rect 19208 10548 19214 10600
rect 19702 10588 19708 10600
rect 19663 10560 19708 10588
rect 19702 10548 19708 10560
rect 19760 10548 19766 10600
rect 19978 10597 19984 10600
rect 19972 10551 19984 10597
rect 20036 10588 20042 10600
rect 20036 10560 20072 10588
rect 19978 10548 19984 10551
rect 20036 10548 20042 10560
rect 21634 10548 21640 10600
rect 21692 10588 21698 10600
rect 21821 10591 21879 10597
rect 21821 10588 21833 10591
rect 21692 10560 21833 10588
rect 21692 10548 21698 10560
rect 21821 10557 21833 10560
rect 21867 10557 21879 10591
rect 22370 10588 22376 10600
rect 22331 10560 22376 10588
rect 21821 10551 21879 10557
rect 22370 10548 22376 10560
rect 22428 10548 22434 10600
rect 14430 10523 14488 10529
rect 14430 10520 14442 10523
rect 10428 10492 12480 10520
rect 12544 10492 13851 10520
rect 13924 10492 14442 10520
rect 3660 10424 7420 10452
rect 3660 10412 3666 10424
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 8849 10455 8907 10461
rect 8849 10452 8861 10455
rect 8260 10424 8861 10452
rect 8260 10412 8266 10424
rect 8849 10421 8861 10424
rect 8895 10421 8907 10455
rect 8849 10415 8907 10421
rect 9398 10412 9404 10464
rect 9456 10452 9462 10464
rect 10428 10452 10456 10492
rect 9456 10424 10456 10452
rect 9456 10412 9462 10424
rect 10502 10412 10508 10464
rect 10560 10452 10566 10464
rect 11333 10455 11391 10461
rect 11333 10452 11345 10455
rect 10560 10424 11345 10452
rect 10560 10412 10566 10424
rect 11333 10421 11345 10424
rect 11379 10421 11391 10455
rect 12452 10452 12480 10492
rect 13924 10461 13952 10492
rect 14430 10489 14442 10492
rect 14476 10489 14488 10523
rect 14430 10483 14488 10489
rect 15930 10480 15936 10532
rect 15988 10480 15994 10532
rect 16114 10529 16120 10532
rect 16108 10520 16120 10529
rect 16075 10492 16120 10520
rect 16108 10483 16120 10492
rect 16114 10480 16120 10483
rect 16172 10480 16178 10532
rect 16298 10480 16304 10532
rect 16356 10480 16362 10532
rect 16574 10480 16580 10532
rect 16632 10520 16638 10532
rect 17586 10520 17592 10532
rect 16632 10492 17592 10520
rect 16632 10480 16638 10492
rect 17586 10480 17592 10492
rect 17644 10480 17650 10532
rect 18601 10523 18659 10529
rect 18601 10489 18613 10523
rect 18647 10520 18659 10523
rect 19245 10523 19303 10529
rect 19245 10520 19257 10523
rect 18647 10492 19257 10520
rect 18647 10489 18659 10492
rect 18601 10483 18659 10489
rect 19245 10489 19257 10492
rect 19291 10489 19303 10523
rect 19245 10483 19303 10489
rect 19794 10480 19800 10532
rect 19852 10520 19858 10532
rect 21729 10523 21787 10529
rect 21729 10520 21741 10523
rect 19852 10492 21741 10520
rect 19852 10480 19858 10492
rect 21729 10489 21741 10492
rect 21775 10489 21787 10523
rect 21729 10483 21787 10489
rect 13909 10455 13967 10461
rect 13909 10452 13921 10455
rect 12452 10424 13921 10452
rect 11333 10415 11391 10421
rect 13909 10421 13921 10424
rect 13955 10421 13967 10455
rect 13909 10415 13967 10421
rect 14274 10412 14280 10464
rect 14332 10452 14338 10464
rect 15565 10455 15623 10461
rect 15565 10452 15577 10455
rect 14332 10424 15577 10452
rect 14332 10412 14338 10424
rect 15565 10421 15577 10424
rect 15611 10421 15623 10455
rect 15948 10452 15976 10480
rect 17221 10455 17279 10461
rect 17221 10452 17233 10455
rect 15948 10424 17233 10452
rect 15565 10415 15623 10421
rect 17221 10421 17233 10424
rect 17267 10421 17279 10455
rect 17678 10452 17684 10464
rect 17639 10424 17684 10452
rect 17221 10415 17279 10421
rect 17678 10412 17684 10424
rect 17736 10412 17742 10464
rect 20530 10412 20536 10464
rect 20588 10452 20594 10464
rect 21361 10455 21419 10461
rect 21361 10452 21373 10455
rect 20588 10424 21373 10452
rect 20588 10412 20594 10424
rect 21361 10421 21373 10424
rect 21407 10421 21419 10455
rect 21361 10415 21419 10421
rect 21450 10412 21456 10464
rect 21508 10452 21514 10464
rect 22557 10455 22615 10461
rect 22557 10452 22569 10455
rect 21508 10424 22569 10452
rect 21508 10412 21514 10424
rect 22557 10421 22569 10424
rect 22603 10421 22615 10455
rect 22557 10415 22615 10421
rect 1104 10362 23276 10384
rect 1104 10310 8379 10362
rect 8431 10310 8443 10362
rect 8495 10310 8507 10362
rect 8559 10310 8571 10362
rect 8623 10310 15776 10362
rect 15828 10310 15840 10362
rect 15892 10310 15904 10362
rect 15956 10310 15968 10362
rect 16020 10310 23276 10362
rect 1104 10288 23276 10310
rect 1673 10251 1731 10257
rect 1673 10217 1685 10251
rect 1719 10248 1731 10251
rect 1762 10248 1768 10260
rect 1719 10220 1768 10248
rect 1719 10217 1731 10220
rect 1673 10211 1731 10217
rect 1762 10208 1768 10220
rect 1820 10208 1826 10260
rect 1949 10251 2007 10257
rect 1949 10217 1961 10251
rect 1995 10248 2007 10251
rect 4798 10248 4804 10260
rect 1995 10220 4804 10248
rect 1995 10217 2007 10220
rect 1949 10211 2007 10217
rect 1489 10115 1547 10121
rect 1489 10081 1501 10115
rect 1535 10112 1547 10115
rect 1964 10112 1992 10211
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 5534 10248 5540 10260
rect 5495 10220 5540 10248
rect 5534 10208 5540 10220
rect 5592 10208 5598 10260
rect 6914 10208 6920 10260
rect 6972 10248 6978 10260
rect 7193 10251 7251 10257
rect 7193 10248 7205 10251
rect 6972 10220 7205 10248
rect 6972 10208 6978 10220
rect 7193 10217 7205 10220
rect 7239 10217 7251 10251
rect 7193 10211 7251 10217
rect 9306 10208 9312 10260
rect 9364 10248 9370 10260
rect 10226 10248 10232 10260
rect 9364 10220 10232 10248
rect 9364 10208 9370 10220
rect 10226 10208 10232 10220
rect 10284 10248 10290 10260
rect 11057 10251 11115 10257
rect 11057 10248 11069 10251
rect 10284 10220 11069 10248
rect 10284 10208 10290 10220
rect 11057 10217 11069 10220
rect 11103 10217 11115 10251
rect 11057 10211 11115 10217
rect 11624 10220 13001 10248
rect 2130 10180 2136 10192
rect 2043 10152 2136 10180
rect 2056 10121 2084 10152
rect 2130 10140 2136 10152
rect 2188 10180 2194 10192
rect 4430 10189 4436 10192
rect 4424 10180 4436 10189
rect 2188 10152 3556 10180
rect 4391 10152 4436 10180
rect 2188 10140 2194 10152
rect 3528 10124 3556 10152
rect 4424 10143 4436 10152
rect 4430 10140 4436 10143
rect 4488 10140 4494 10192
rect 5810 10140 5816 10192
rect 5868 10180 5874 10192
rect 6058 10183 6116 10189
rect 6058 10180 6070 10183
rect 5868 10152 6070 10180
rect 5868 10140 5874 10152
rect 6058 10149 6070 10152
rect 6104 10149 6116 10183
rect 6058 10143 6116 10149
rect 7558 10140 7564 10192
rect 7616 10180 7622 10192
rect 8294 10180 8300 10192
rect 7616 10152 8300 10180
rect 7616 10140 7622 10152
rect 8294 10140 8300 10152
rect 8352 10140 8358 10192
rect 8386 10140 8392 10192
rect 8444 10180 8450 10192
rect 8938 10180 8944 10192
rect 8444 10152 8944 10180
rect 8444 10140 8450 10152
rect 8938 10140 8944 10152
rect 8996 10140 9002 10192
rect 9858 10140 9864 10192
rect 9916 10180 9922 10192
rect 11624 10180 11652 10220
rect 9916 10152 11652 10180
rect 9916 10140 9922 10152
rect 11698 10140 11704 10192
rect 11756 10180 11762 10192
rect 12161 10183 12219 10189
rect 12161 10180 12173 10183
rect 11756 10152 12173 10180
rect 11756 10140 11762 10152
rect 12161 10149 12173 10152
rect 12207 10149 12219 10183
rect 12161 10143 12219 10149
rect 12342 10140 12348 10192
rect 12400 10180 12406 10192
rect 12973 10189 13001 10220
rect 13170 10208 13176 10260
rect 13228 10248 13234 10260
rect 13998 10248 14004 10260
rect 13228 10220 14004 10248
rect 13228 10208 13234 10220
rect 13998 10208 14004 10220
rect 14056 10248 14062 10260
rect 14093 10251 14151 10257
rect 14093 10248 14105 10251
rect 14056 10220 14105 10248
rect 14056 10208 14062 10220
rect 14093 10217 14105 10220
rect 14139 10217 14151 10251
rect 14550 10248 14556 10260
rect 14511 10220 14556 10248
rect 14093 10211 14151 10217
rect 14550 10208 14556 10220
rect 14608 10208 14614 10260
rect 14642 10208 14648 10260
rect 14700 10248 14706 10260
rect 14737 10251 14795 10257
rect 14737 10248 14749 10251
rect 14700 10220 14749 10248
rect 14700 10208 14706 10220
rect 14737 10217 14749 10220
rect 14783 10217 14795 10251
rect 14737 10211 14795 10217
rect 16114 10208 16120 10260
rect 16172 10248 16178 10260
rect 16853 10251 16911 10257
rect 16853 10248 16865 10251
rect 16172 10220 16865 10248
rect 16172 10208 16178 10220
rect 16853 10217 16865 10220
rect 16899 10217 16911 10251
rect 16853 10211 16911 10217
rect 17310 10208 17316 10260
rect 17368 10248 17374 10260
rect 18414 10248 18420 10260
rect 17368 10220 18420 10248
rect 17368 10208 17374 10220
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 18690 10208 18696 10260
rect 18748 10248 18754 10260
rect 20073 10251 20131 10257
rect 20073 10248 20085 10251
rect 18748 10220 20085 10248
rect 18748 10208 18754 10220
rect 20073 10217 20085 10220
rect 20119 10217 20131 10251
rect 20073 10211 20131 10217
rect 20349 10251 20407 10257
rect 20349 10217 20361 10251
rect 20395 10248 20407 10251
rect 21726 10248 21732 10260
rect 20395 10220 21732 10248
rect 20395 10217 20407 10220
rect 20349 10211 20407 10217
rect 21726 10208 21732 10220
rect 21784 10208 21790 10260
rect 22278 10248 22284 10260
rect 22239 10220 22284 10248
rect 22278 10208 22284 10220
rect 22336 10208 22342 10260
rect 12621 10183 12679 10189
rect 12621 10180 12633 10183
rect 12400 10152 12633 10180
rect 12400 10140 12406 10152
rect 12621 10149 12633 10152
rect 12667 10180 12679 10183
rect 12958 10183 13016 10189
rect 12667 10152 12756 10180
rect 12667 10149 12679 10152
rect 12621 10143 12679 10149
rect 1535 10084 1992 10112
rect 2041 10115 2099 10121
rect 1535 10081 1547 10084
rect 1489 10075 1547 10081
rect 2041 10081 2053 10115
rect 2087 10081 2099 10115
rect 2041 10075 2099 10081
rect 2308 10115 2366 10121
rect 2308 10081 2320 10115
rect 2354 10112 2366 10115
rect 2774 10112 2780 10124
rect 2354 10084 2780 10112
rect 2354 10081 2366 10084
rect 2308 10075 2366 10081
rect 2774 10072 2780 10084
rect 2832 10072 2838 10124
rect 3510 10072 3516 10124
rect 3568 10112 3574 10124
rect 4157 10115 4215 10121
rect 4157 10112 4169 10115
rect 3568 10084 4169 10112
rect 3568 10072 3574 10084
rect 4157 10081 4169 10084
rect 4203 10112 4215 10115
rect 6638 10112 6644 10124
rect 4203 10084 6644 10112
rect 4203 10081 4215 10084
rect 4157 10075 4215 10081
rect 5828 10053 5856 10084
rect 6638 10072 6644 10084
rect 6696 10072 6702 10124
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 8202 10121 8208 10124
rect 8185 10115 8208 10121
rect 8185 10112 8197 10115
rect 6972 10084 8197 10112
rect 6972 10072 6978 10084
rect 8185 10081 8197 10084
rect 8260 10112 8266 10124
rect 9944 10115 10002 10121
rect 8260 10084 8333 10112
rect 8185 10075 8208 10081
rect 8202 10072 8208 10075
rect 8260 10072 8266 10084
rect 9944 10081 9956 10115
rect 9990 10112 10002 10115
rect 10226 10112 10232 10124
rect 9990 10084 10232 10112
rect 9990 10081 10002 10084
rect 9944 10075 10002 10081
rect 10226 10072 10232 10084
rect 10284 10072 10290 10124
rect 11790 10072 11796 10124
rect 11848 10112 11854 10124
rect 12728 10121 12756 10152
rect 12958 10149 12970 10183
rect 13004 10180 13016 10183
rect 14274 10180 14280 10192
rect 13004 10152 14280 10180
rect 13004 10149 13016 10152
rect 12958 10143 13016 10149
rect 14274 10140 14280 10152
rect 14332 10140 14338 10192
rect 15740 10183 15798 10189
rect 14384 10152 15700 10180
rect 14384 10121 14412 10152
rect 12069 10115 12127 10121
rect 12069 10112 12081 10115
rect 11848 10084 12081 10112
rect 11848 10072 11854 10084
rect 12069 10081 12081 10084
rect 12115 10081 12127 10115
rect 12069 10075 12127 10081
rect 12713 10115 12771 10121
rect 12713 10081 12725 10115
rect 12759 10081 12771 10115
rect 14369 10115 14427 10121
rect 12713 10075 12771 10081
rect 12820 10084 13768 10112
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10013 5871 10047
rect 5813 10007 5871 10013
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10013 7987 10047
rect 9674 10044 9680 10056
rect 9635 10016 9680 10044
rect 7929 10007 7987 10013
rect 3326 9868 3332 9920
rect 3384 9908 3390 9920
rect 3421 9911 3479 9917
rect 3421 9908 3433 9911
rect 3384 9880 3433 9908
rect 3384 9868 3390 9880
rect 3421 9877 3433 9880
rect 3467 9877 3479 9911
rect 3421 9871 3479 9877
rect 4062 9868 4068 9920
rect 4120 9908 4126 9920
rect 4430 9908 4436 9920
rect 4120 9880 4436 9908
rect 4120 9868 4126 9880
rect 4430 9868 4436 9880
rect 4488 9868 4494 9920
rect 7944 9908 7972 10007
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 12345 10047 12403 10053
rect 12345 10013 12357 10047
rect 12391 10044 12403 10047
rect 12434 10044 12440 10056
rect 12391 10016 12440 10044
rect 12391 10013 12403 10016
rect 12345 10007 12403 10013
rect 12434 10004 12440 10016
rect 12492 10044 12498 10056
rect 12820 10044 12848 10084
rect 12492 10016 12848 10044
rect 13740 10044 13768 10084
rect 14369 10081 14381 10115
rect 14415 10081 14427 10115
rect 14918 10112 14924 10124
rect 14369 10075 14427 10081
rect 14660 10084 14924 10112
rect 14660 10056 14688 10084
rect 14918 10072 14924 10084
rect 14976 10072 14982 10124
rect 15102 10112 15108 10124
rect 15063 10084 15108 10112
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 15672 10112 15700 10152
rect 15740 10149 15752 10183
rect 15786 10180 15798 10183
rect 16390 10180 16396 10192
rect 15786 10152 16396 10180
rect 15786 10149 15798 10152
rect 15740 10143 15798 10149
rect 16390 10140 16396 10152
rect 16448 10140 16454 10192
rect 19794 10180 19800 10192
rect 18340 10152 19800 10180
rect 17034 10112 17040 10124
rect 15672 10084 17040 10112
rect 17034 10072 17040 10084
rect 17092 10072 17098 10124
rect 17586 10112 17592 10124
rect 17547 10084 17592 10112
rect 17586 10072 17592 10084
rect 17644 10072 17650 10124
rect 17681 10115 17739 10121
rect 17681 10081 17693 10115
rect 17727 10112 17739 10115
rect 17862 10112 17868 10124
rect 17727 10084 17868 10112
rect 17727 10081 17739 10084
rect 17681 10075 17739 10081
rect 17862 10072 17868 10084
rect 17920 10072 17926 10124
rect 18230 10112 18236 10124
rect 18191 10084 18236 10112
rect 18230 10072 18236 10084
rect 18288 10072 18294 10124
rect 14642 10044 14648 10056
rect 13740 10016 14648 10044
rect 12492 10004 12498 10016
rect 14642 10004 14648 10016
rect 14700 10004 14706 10056
rect 14734 10004 14740 10056
rect 14792 10044 14798 10056
rect 15473 10047 15531 10053
rect 15473 10044 15485 10047
rect 14792 10016 15485 10044
rect 14792 10004 14798 10016
rect 15473 10013 15485 10016
rect 15519 10013 15531 10047
rect 15473 10007 15531 10013
rect 17773 10047 17831 10053
rect 17773 10013 17785 10047
rect 17819 10044 17831 10047
rect 18340 10044 18368 10152
rect 19794 10140 19800 10152
rect 19852 10140 19858 10192
rect 20438 10140 20444 10192
rect 20496 10180 20502 10192
rect 22189 10183 22247 10189
rect 22189 10180 22201 10183
rect 20496 10152 22201 10180
rect 20496 10140 20502 10152
rect 22189 10149 22201 10152
rect 22235 10149 22247 10183
rect 22189 10143 22247 10149
rect 18500 10115 18558 10121
rect 18500 10081 18512 10115
rect 18546 10112 18558 10115
rect 18782 10112 18788 10124
rect 18546 10084 18788 10112
rect 18546 10081 18558 10084
rect 18500 10075 18558 10081
rect 18782 10072 18788 10084
rect 18840 10072 18846 10124
rect 18874 10072 18880 10124
rect 18932 10112 18938 10124
rect 19889 10115 19947 10121
rect 19889 10112 19901 10115
rect 18932 10084 19901 10112
rect 18932 10072 18938 10084
rect 19889 10081 19901 10084
rect 19935 10081 19947 10115
rect 19889 10075 19947 10081
rect 19978 10072 19984 10124
rect 20036 10112 20042 10124
rect 20625 10115 20683 10121
rect 20625 10112 20637 10115
rect 20036 10084 20637 10112
rect 20036 10072 20042 10084
rect 20625 10081 20637 10084
rect 20671 10081 20683 10115
rect 21266 10112 21272 10124
rect 21227 10084 21272 10112
rect 20625 10075 20683 10081
rect 21266 10072 21272 10084
rect 21324 10072 21330 10124
rect 17819 10016 18368 10044
rect 17819 10013 17831 10016
rect 17773 10007 17831 10013
rect 19702 10004 19708 10056
rect 19760 10044 19766 10056
rect 20714 10044 20720 10056
rect 19760 10016 20720 10044
rect 19760 10004 19766 10016
rect 9692 9976 9720 10004
rect 20456 9985 20484 10016
rect 20714 10004 20720 10016
rect 20772 10004 20778 10056
rect 22465 10047 22523 10053
rect 22465 10013 22477 10047
rect 22511 10044 22523 10047
rect 22646 10044 22652 10056
rect 22511 10016 22652 10044
rect 22511 10013 22523 10016
rect 22465 10007 22523 10013
rect 22646 10004 22652 10016
rect 22704 10004 22710 10056
rect 20349 9979 20407 9985
rect 20349 9976 20361 9979
rect 8864 9948 9720 9976
rect 16408 9948 18283 9976
rect 8864 9908 8892 9948
rect 7944 9880 8892 9908
rect 8938 9868 8944 9920
rect 8996 9908 9002 9920
rect 9309 9911 9367 9917
rect 9309 9908 9321 9911
rect 8996 9880 9321 9908
rect 8996 9868 9002 9880
rect 9309 9877 9321 9880
rect 9355 9877 9367 9911
rect 9309 9871 9367 9877
rect 9490 9868 9496 9920
rect 9548 9908 9554 9920
rect 11701 9911 11759 9917
rect 11701 9908 11713 9911
rect 9548 9880 11713 9908
rect 9548 9868 9554 9880
rect 11701 9877 11713 9880
rect 11747 9877 11759 9911
rect 11701 9871 11759 9877
rect 12621 9911 12679 9917
rect 12621 9877 12633 9911
rect 12667 9908 12679 9911
rect 12986 9908 12992 9920
rect 12667 9880 12992 9908
rect 12667 9877 12679 9880
rect 12621 9871 12679 9877
rect 12986 9868 12992 9880
rect 13044 9868 13050 9920
rect 14090 9868 14096 9920
rect 14148 9908 14154 9920
rect 14737 9911 14795 9917
rect 14737 9908 14749 9911
rect 14148 9880 14749 9908
rect 14148 9868 14154 9880
rect 14737 9877 14749 9880
rect 14783 9877 14795 9911
rect 14918 9908 14924 9920
rect 14879 9880 14924 9908
rect 14737 9871 14795 9877
rect 14918 9868 14924 9880
rect 14976 9868 14982 9920
rect 15194 9868 15200 9920
rect 15252 9908 15258 9920
rect 16408 9908 16436 9948
rect 17218 9908 17224 9920
rect 15252 9880 16436 9908
rect 17179 9880 17224 9908
rect 15252 9868 15258 9880
rect 17218 9868 17224 9880
rect 17276 9868 17282 9920
rect 18255 9908 18283 9948
rect 19168 9948 20361 9976
rect 19168 9908 19196 9948
rect 20349 9945 20361 9948
rect 20395 9945 20407 9979
rect 20349 9939 20407 9945
rect 20441 9979 20499 9985
rect 20441 9945 20453 9979
rect 20487 9945 20499 9979
rect 20441 9939 20499 9945
rect 20622 9936 20628 9988
rect 20680 9976 20686 9988
rect 20680 9948 21772 9976
rect 20680 9936 20686 9948
rect 21744 9920 21772 9948
rect 18255 9880 19196 9908
rect 19334 9868 19340 9920
rect 19392 9908 19398 9920
rect 19613 9911 19671 9917
rect 19613 9908 19625 9911
rect 19392 9880 19625 9908
rect 19392 9868 19398 9880
rect 19613 9877 19625 9880
rect 19659 9877 19671 9911
rect 19613 9871 19671 9877
rect 20898 9868 20904 9920
rect 20956 9908 20962 9920
rect 21453 9911 21511 9917
rect 21453 9908 21465 9911
rect 20956 9880 21465 9908
rect 20956 9868 20962 9880
rect 21453 9877 21465 9880
rect 21499 9877 21511 9911
rect 21453 9871 21511 9877
rect 21726 9868 21732 9920
rect 21784 9908 21790 9920
rect 21821 9911 21879 9917
rect 21821 9908 21833 9911
rect 21784 9880 21833 9908
rect 21784 9868 21790 9880
rect 21821 9877 21833 9880
rect 21867 9877 21879 9911
rect 21821 9871 21879 9877
rect 1104 9818 23276 9840
rect 1104 9766 4680 9818
rect 4732 9766 4744 9818
rect 4796 9766 4808 9818
rect 4860 9766 4872 9818
rect 4924 9766 12078 9818
rect 12130 9766 12142 9818
rect 12194 9766 12206 9818
rect 12258 9766 12270 9818
rect 12322 9766 19475 9818
rect 19527 9766 19539 9818
rect 19591 9766 19603 9818
rect 19655 9766 19667 9818
rect 19719 9766 23276 9818
rect 1104 9744 23276 9766
rect 2130 9704 2136 9716
rect 1412 9676 2136 9704
rect 1412 9577 1440 9676
rect 2130 9664 2136 9676
rect 2188 9664 2194 9716
rect 7006 9704 7012 9716
rect 6932 9676 7012 9704
rect 2774 9596 2780 9648
rect 2832 9636 2838 9648
rect 2832 9608 2877 9636
rect 2832 9596 2838 9608
rect 4154 9596 4160 9648
rect 4212 9636 4218 9648
rect 4433 9639 4491 9645
rect 4433 9636 4445 9639
rect 4212 9608 4445 9636
rect 4212 9596 4218 9608
rect 4433 9605 4445 9608
rect 4479 9605 4491 9639
rect 4433 9599 4491 9605
rect 5810 9596 5816 9648
rect 5868 9636 5874 9648
rect 6932 9636 6960 9676
rect 7006 9664 7012 9676
rect 7064 9664 7070 9716
rect 7653 9707 7711 9713
rect 7653 9673 7665 9707
rect 7699 9704 7711 9707
rect 7926 9704 7932 9716
rect 7699 9676 7932 9704
rect 7699 9673 7711 9676
rect 7653 9667 7711 9673
rect 7926 9664 7932 9676
rect 7984 9664 7990 9716
rect 8386 9664 8392 9716
rect 8444 9704 8450 9716
rect 8444 9676 9904 9704
rect 8444 9664 8450 9676
rect 5868 9608 6960 9636
rect 7285 9639 7343 9645
rect 5868 9596 5874 9608
rect 7285 9605 7297 9639
rect 7331 9636 7343 9639
rect 7469 9639 7527 9645
rect 7469 9636 7481 9639
rect 7331 9608 7481 9636
rect 7331 9605 7343 9608
rect 7285 9599 7343 9605
rect 7469 9605 7481 9608
rect 7515 9605 7527 9639
rect 8662 9636 8668 9648
rect 7469 9599 7527 9605
rect 8220 9608 8668 9636
rect 1397 9571 1455 9577
rect 1397 9537 1409 9571
rect 1443 9537 1455 9571
rect 1397 9531 1455 9537
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9568 4767 9571
rect 5258 9568 5264 9580
rect 4755 9540 5264 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 5258 9528 5264 9540
rect 5316 9528 5322 9580
rect 5534 9528 5540 9580
rect 5592 9568 5598 9580
rect 5629 9571 5687 9577
rect 5629 9568 5641 9571
rect 5592 9540 5641 9568
rect 5592 9528 5598 9540
rect 5629 9537 5641 9540
rect 5675 9537 5687 9571
rect 5629 9531 5687 9537
rect 5721 9571 5779 9577
rect 5721 9537 5733 9571
rect 5767 9537 5779 9571
rect 8220 9568 8248 9608
rect 8662 9596 8668 9608
rect 8720 9596 8726 9648
rect 5721 9531 5779 9537
rect 6196 9540 8248 9568
rect 8297 9571 8355 9577
rect 3326 9509 3332 9512
rect 3053 9503 3111 9509
rect 3053 9469 3065 9503
rect 3099 9469 3111 9503
rect 3320 9500 3332 9509
rect 3287 9472 3332 9500
rect 3053 9463 3111 9469
rect 3320 9463 3332 9472
rect 1486 9392 1492 9444
rect 1544 9432 1550 9444
rect 1642 9435 1700 9441
rect 1642 9432 1654 9435
rect 1544 9404 1654 9432
rect 1544 9392 1550 9404
rect 1642 9401 1654 9404
rect 1688 9401 1700 9435
rect 3068 9432 3096 9463
rect 3326 9460 3332 9463
rect 3384 9460 3390 9512
rect 4890 9460 4896 9512
rect 4948 9500 4954 9512
rect 5736 9500 5764 9531
rect 6196 9509 6224 9540
rect 8297 9537 8309 9571
rect 8343 9568 8355 9571
rect 9876 9568 9904 9676
rect 9950 9664 9956 9716
rect 10008 9704 10014 9716
rect 10318 9704 10324 9716
rect 10008 9676 10324 9704
rect 10008 9664 10014 9676
rect 10318 9664 10324 9676
rect 10376 9664 10382 9716
rect 11790 9664 11796 9716
rect 11848 9704 11854 9716
rect 12526 9704 12532 9716
rect 11848 9676 12532 9704
rect 11848 9664 11854 9676
rect 12526 9664 12532 9676
rect 12584 9664 12590 9716
rect 12986 9704 12992 9716
rect 12719 9676 12992 9704
rect 10045 9639 10103 9645
rect 10045 9605 10057 9639
rect 10091 9636 10103 9639
rect 10226 9636 10232 9648
rect 10091 9608 10232 9636
rect 10091 9605 10103 9608
rect 10045 9599 10103 9605
rect 10226 9596 10232 9608
rect 10284 9596 10290 9648
rect 11422 9596 11428 9648
rect 11480 9636 11486 9648
rect 11701 9639 11759 9645
rect 11701 9636 11713 9639
rect 11480 9608 11713 9636
rect 11480 9596 11486 9608
rect 11701 9605 11713 9608
rect 11747 9605 11759 9639
rect 11701 9599 11759 9605
rect 12069 9639 12127 9645
rect 12069 9605 12081 9639
rect 12115 9636 12127 9639
rect 12719 9636 12747 9676
rect 12986 9664 12992 9676
rect 13044 9704 13050 9716
rect 14369 9707 14427 9713
rect 13044 9676 13768 9704
rect 13044 9664 13050 9676
rect 12115 9608 12747 9636
rect 12115 9605 12127 9608
rect 12069 9599 12127 9605
rect 12618 9568 12624 9580
rect 8343 9540 8800 9568
rect 9876 9540 10456 9568
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 4948 9472 5764 9500
rect 6181 9503 6239 9509
rect 4948 9460 4954 9472
rect 6181 9469 6193 9503
rect 6227 9469 6239 9503
rect 6181 9463 6239 9469
rect 7006 9460 7012 9512
rect 7064 9500 7070 9512
rect 7101 9503 7159 9509
rect 7101 9500 7113 9503
rect 7064 9472 7113 9500
rect 7064 9460 7070 9472
rect 7101 9469 7113 9472
rect 7147 9469 7159 9503
rect 8113 9503 8171 9509
rect 8113 9500 8125 9503
rect 7101 9463 7159 9469
rect 7484 9472 8125 9500
rect 3510 9432 3516 9444
rect 3068 9404 3516 9432
rect 1642 9395 1700 9401
rect 3510 9392 3516 9404
rect 3568 9392 3574 9444
rect 5537 9435 5595 9441
rect 5537 9401 5549 9435
rect 5583 9432 5595 9435
rect 6454 9432 6460 9444
rect 5583 9404 6460 9432
rect 5583 9401 5595 9404
rect 5537 9395 5595 9401
rect 6454 9392 6460 9404
rect 6512 9392 6518 9444
rect 6638 9392 6644 9444
rect 6696 9432 6702 9444
rect 7484 9432 7512 9472
rect 8113 9469 8125 9472
rect 8159 9469 8171 9503
rect 8478 9500 8484 9512
rect 8113 9463 8171 9469
rect 8220 9472 8484 9500
rect 8220 9432 8248 9472
rect 8478 9460 8484 9472
rect 8536 9460 8542 9512
rect 8665 9503 8723 9509
rect 8665 9469 8677 9503
rect 8711 9469 8723 9503
rect 8665 9463 8723 9469
rect 6696 9404 7512 9432
rect 7944 9404 8248 9432
rect 6696 9392 6702 9404
rect 2314 9324 2320 9376
rect 2372 9364 2378 9376
rect 4798 9364 4804 9376
rect 2372 9336 4804 9364
rect 2372 9324 2378 9336
rect 4798 9324 4804 9336
rect 4856 9324 4862 9376
rect 5169 9367 5227 9373
rect 5169 9333 5181 9367
rect 5215 9364 5227 9367
rect 5258 9364 5264 9376
rect 5215 9336 5264 9364
rect 5215 9333 5227 9336
rect 5169 9327 5227 9333
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 6362 9364 6368 9376
rect 6323 9336 6368 9364
rect 6362 9324 6368 9336
rect 6420 9324 6426 9376
rect 7006 9324 7012 9376
rect 7064 9364 7070 9376
rect 7282 9364 7288 9376
rect 7064 9336 7288 9364
rect 7064 9324 7070 9336
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 7469 9367 7527 9373
rect 7469 9333 7481 9367
rect 7515 9364 7527 9367
rect 7944 9364 7972 9404
rect 8570 9392 8576 9444
rect 8628 9392 8634 9444
rect 7515 9336 7972 9364
rect 8021 9367 8079 9373
rect 7515 9333 7527 9336
rect 7469 9327 7527 9333
rect 8021 9333 8033 9367
rect 8067 9364 8079 9367
rect 8588 9364 8616 9392
rect 8067 9336 8616 9364
rect 8680 9364 8708 9463
rect 8772 9444 8800 9540
rect 8938 9509 8944 9512
rect 8932 9500 8944 9509
rect 8899 9472 8944 9500
rect 8932 9463 8944 9472
rect 8938 9460 8944 9463
rect 8996 9460 9002 9512
rect 10321 9503 10379 9509
rect 10321 9500 10333 9503
rect 9959 9472 10333 9500
rect 8754 9392 8760 9444
rect 8812 9432 8818 9444
rect 9122 9432 9128 9444
rect 8812 9404 9128 9432
rect 8812 9392 8818 9404
rect 9122 9392 9128 9404
rect 9180 9392 9186 9444
rect 9766 9364 9772 9376
rect 8680 9336 9772 9364
rect 8067 9333 8079 9336
rect 8021 9327 8079 9333
rect 9766 9324 9772 9336
rect 9824 9364 9830 9376
rect 9959 9364 9987 9472
rect 10321 9469 10333 9472
rect 10367 9469 10379 9503
rect 10428 9500 10456 9540
rect 12176 9540 12624 9568
rect 12176 9500 12204 9540
rect 12618 9528 12624 9540
rect 12676 9528 12682 9580
rect 12719 9577 12747 9608
rect 12713 9571 12771 9577
rect 12713 9537 12725 9571
rect 12759 9537 12771 9571
rect 13740 9568 13768 9676
rect 14369 9673 14381 9707
rect 14415 9704 14427 9707
rect 15102 9704 15108 9716
rect 14415 9676 15108 9704
rect 14415 9673 14427 9676
rect 14369 9667 14427 9673
rect 15102 9664 15108 9676
rect 15160 9664 15166 9716
rect 18598 9704 18604 9716
rect 17512 9676 18604 9704
rect 14090 9636 14096 9648
rect 14051 9608 14096 9636
rect 14090 9596 14096 9608
rect 14148 9596 14154 9648
rect 16390 9596 16396 9648
rect 16448 9636 16454 9648
rect 16669 9639 16727 9645
rect 16669 9636 16681 9639
rect 16448 9608 16681 9636
rect 16448 9596 16454 9608
rect 16669 9605 16681 9608
rect 16715 9605 16727 9639
rect 16669 9599 16727 9605
rect 14734 9568 14740 9580
rect 13740 9540 14740 9568
rect 12713 9531 12771 9537
rect 14734 9528 14740 9540
rect 14792 9568 14798 9580
rect 15289 9571 15347 9577
rect 15289 9568 15301 9571
rect 14792 9540 15301 9568
rect 14792 9528 14798 9540
rect 15289 9537 15301 9540
rect 15335 9537 15347 9571
rect 15289 9531 15347 9537
rect 17405 9571 17463 9577
rect 17405 9537 17417 9571
rect 17451 9568 17463 9571
rect 17512 9568 17540 9676
rect 18598 9664 18604 9676
rect 18656 9704 18662 9716
rect 18656 9676 20576 9704
rect 18656 9664 18662 9676
rect 17862 9596 17868 9648
rect 17920 9636 17926 9648
rect 20548 9636 20576 9676
rect 20993 9639 21051 9645
rect 20993 9636 21005 9639
rect 17920 9608 18911 9636
rect 20548 9608 21005 9636
rect 17920 9596 17926 9608
rect 17451 9540 17540 9568
rect 17589 9571 17647 9577
rect 17451 9537 17463 9540
rect 17405 9531 17463 9537
rect 17589 9537 17601 9571
rect 17635 9568 17647 9571
rect 17770 9568 17776 9580
rect 17635 9540 17776 9568
rect 17635 9537 17647 9540
rect 17589 9531 17647 9537
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 18785 9571 18843 9577
rect 18785 9537 18797 9571
rect 18831 9537 18843 9571
rect 18785 9531 18843 9537
rect 10428 9472 12204 9500
rect 12253 9503 12311 9509
rect 10321 9463 10379 9469
rect 12253 9469 12265 9503
rect 12299 9500 12311 9503
rect 12434 9500 12440 9512
rect 12299 9472 12440 9500
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 12434 9460 12440 9472
rect 12492 9460 12498 9512
rect 12526 9460 12532 9512
rect 12584 9500 12590 9512
rect 12584 9472 13023 9500
rect 12584 9460 12590 9472
rect 10502 9392 10508 9444
rect 10560 9441 10566 9444
rect 12995 9441 13023 9472
rect 13262 9460 13268 9512
rect 13320 9500 13326 9512
rect 14553 9503 14611 9509
rect 14553 9500 14565 9503
rect 13320 9472 14565 9500
rect 13320 9460 13326 9472
rect 14553 9469 14565 9472
rect 14599 9469 14611 9503
rect 14553 9463 14611 9469
rect 14645 9503 14703 9509
rect 14645 9469 14657 9503
rect 14691 9500 14703 9503
rect 15010 9500 15016 9512
rect 14691 9472 15016 9500
rect 14691 9469 14703 9472
rect 14645 9463 14703 9469
rect 15010 9460 15016 9472
rect 15068 9460 15074 9512
rect 15556 9503 15614 9509
rect 15556 9469 15568 9503
rect 15602 9500 15614 9503
rect 18690 9500 18696 9512
rect 15602 9472 18696 9500
rect 15602 9469 15614 9472
rect 15556 9463 15614 9469
rect 18690 9460 18696 9472
rect 18748 9500 18754 9512
rect 18800 9500 18828 9531
rect 18748 9472 18828 9500
rect 18748 9460 18754 9472
rect 10560 9435 10624 9441
rect 10560 9401 10578 9435
rect 10612 9401 10624 9435
rect 10560 9395 10624 9401
rect 12980 9435 13038 9441
rect 12980 9401 12992 9435
rect 13026 9432 13038 9435
rect 14458 9432 14464 9444
rect 13026 9404 14464 9432
rect 13026 9401 13038 9404
rect 12980 9395 13038 9401
rect 10560 9392 10566 9395
rect 14458 9392 14464 9404
rect 14516 9392 14522 9444
rect 14734 9392 14740 9444
rect 14792 9432 14798 9444
rect 14829 9435 14887 9441
rect 14829 9432 14841 9435
rect 14792 9404 14841 9432
rect 14792 9392 14798 9404
rect 14829 9401 14841 9404
rect 14875 9401 14887 9435
rect 18883 9432 18911 9608
rect 20993 9605 21005 9608
rect 21039 9605 21051 9639
rect 20993 9599 21051 9605
rect 19150 9568 19156 9580
rect 19111 9540 19156 9568
rect 19150 9528 19156 9540
rect 19208 9528 19214 9580
rect 19702 9577 19708 9580
rect 19659 9571 19708 9577
rect 19659 9537 19671 9571
rect 19705 9537 19708 9571
rect 19659 9531 19708 9537
rect 19702 9528 19708 9531
rect 19760 9528 19766 9580
rect 19886 9568 19892 9580
rect 19847 9540 19892 9568
rect 19886 9528 19892 9540
rect 19944 9528 19950 9580
rect 20714 9528 20720 9580
rect 20772 9568 20778 9580
rect 21361 9571 21419 9577
rect 21361 9568 21373 9571
rect 20772 9540 21373 9568
rect 20772 9528 20778 9540
rect 21361 9537 21373 9540
rect 21407 9537 21419 9571
rect 21361 9531 21419 9537
rect 18966 9460 18972 9512
rect 19024 9500 19030 9512
rect 19476 9503 19534 9509
rect 19476 9500 19488 9503
rect 19024 9472 19488 9500
rect 19024 9460 19030 9472
rect 19476 9469 19488 9472
rect 19522 9469 19534 9503
rect 19476 9463 19534 9469
rect 19058 9432 19064 9444
rect 14829 9395 14887 9401
rect 16960 9404 17816 9432
rect 18883 9404 19064 9432
rect 9824 9336 9987 9364
rect 9824 9324 9830 9336
rect 10410 9324 10416 9376
rect 10468 9364 10474 9376
rect 11330 9364 11336 9376
rect 10468 9336 11336 9364
rect 10468 9324 10474 9336
rect 11330 9324 11336 9336
rect 11388 9324 11394 9376
rect 15010 9364 15016 9376
rect 14971 9336 15016 9364
rect 15010 9324 15016 9336
rect 15068 9324 15074 9376
rect 16960 9373 16988 9404
rect 17788 9376 17816 9404
rect 19058 9392 19064 9404
rect 19116 9392 19122 9444
rect 21628 9435 21686 9441
rect 20548 9404 21128 9432
rect 16945 9367 17003 9373
rect 16945 9333 16957 9367
rect 16991 9333 17003 9367
rect 17310 9364 17316 9376
rect 17271 9336 17316 9364
rect 16945 9327 17003 9333
rect 17310 9324 17316 9336
rect 17368 9324 17374 9376
rect 17770 9324 17776 9376
rect 17828 9324 17834 9376
rect 18138 9364 18144 9376
rect 18099 9336 18144 9364
rect 18138 9324 18144 9336
rect 18196 9324 18202 9376
rect 18230 9324 18236 9376
rect 18288 9364 18294 9376
rect 18509 9367 18567 9373
rect 18509 9364 18521 9367
rect 18288 9336 18521 9364
rect 18288 9324 18294 9336
rect 18509 9333 18521 9336
rect 18555 9333 18567 9367
rect 18509 9327 18567 9333
rect 18598 9324 18604 9376
rect 18656 9364 18662 9376
rect 18656 9336 18701 9364
rect 18656 9324 18662 9336
rect 18782 9324 18788 9376
rect 18840 9364 18846 9376
rect 20548 9364 20576 9404
rect 18840 9336 20576 9364
rect 21100 9364 21128 9404
rect 21628 9401 21640 9435
rect 21674 9432 21686 9435
rect 22646 9432 22652 9444
rect 21674 9404 22652 9432
rect 21674 9401 21686 9404
rect 21628 9395 21686 9401
rect 22646 9392 22652 9404
rect 22704 9392 22710 9444
rect 22741 9367 22799 9373
rect 22741 9364 22753 9367
rect 21100 9336 22753 9364
rect 18840 9324 18846 9336
rect 22741 9333 22753 9336
rect 22787 9333 22799 9367
rect 22741 9327 22799 9333
rect 1104 9274 23276 9296
rect 1104 9222 8379 9274
rect 8431 9222 8443 9274
rect 8495 9222 8507 9274
rect 8559 9222 8571 9274
rect 8623 9222 15776 9274
rect 15828 9222 15840 9274
rect 15892 9222 15904 9274
rect 15956 9222 15968 9274
rect 16020 9222 23276 9274
rect 1104 9200 23276 9222
rect 2314 9160 2320 9172
rect 2275 9132 2320 9160
rect 2314 9120 2320 9132
rect 2372 9120 2378 9172
rect 3237 9163 3295 9169
rect 3237 9129 3249 9163
rect 3283 9160 3295 9163
rect 3326 9160 3332 9172
rect 3283 9132 3332 9160
rect 3283 9129 3295 9132
rect 3237 9123 3295 9129
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 3418 9120 3424 9172
rect 3476 9160 3482 9172
rect 4065 9163 4123 9169
rect 4065 9160 4077 9163
rect 3476 9132 4077 9160
rect 3476 9120 3482 9132
rect 4065 9129 4077 9132
rect 4111 9129 4123 9163
rect 4065 9123 4123 9129
rect 4338 9120 4344 9172
rect 4396 9160 4402 9172
rect 4433 9163 4491 9169
rect 4433 9160 4445 9163
rect 4396 9132 4445 9160
rect 4396 9120 4402 9132
rect 4433 9129 4445 9132
rect 4479 9129 4491 9163
rect 5074 9160 5080 9172
rect 5035 9132 5080 9160
rect 4433 9123 4491 9129
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 5350 9120 5356 9172
rect 5408 9160 5414 9172
rect 5445 9163 5503 9169
rect 5445 9160 5457 9163
rect 5408 9132 5457 9160
rect 5408 9120 5414 9132
rect 5445 9129 5457 9132
rect 5491 9129 5503 9163
rect 7006 9160 7012 9172
rect 5445 9123 5503 9129
rect 5828 9132 7012 9160
rect 2225 9095 2283 9101
rect 2225 9061 2237 9095
rect 2271 9092 2283 9095
rect 2498 9092 2504 9104
rect 2271 9064 2504 9092
rect 2271 9061 2283 9064
rect 2225 9055 2283 9061
rect 2498 9052 2504 9064
rect 2556 9052 2562 9104
rect 3970 9092 3976 9104
rect 3436 9064 3976 9092
rect 2774 8984 2780 9036
rect 2832 9024 2838 9036
rect 3329 9027 3387 9033
rect 3329 9024 3341 9027
rect 2832 8996 3341 9024
rect 2832 8984 2838 8996
rect 3329 8993 3341 8996
rect 3375 8993 3387 9027
rect 3329 8987 3387 8993
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8956 2559 8959
rect 3436 8956 3464 9064
rect 3970 9052 3976 9064
rect 4028 9052 4034 9104
rect 5258 9052 5264 9104
rect 5316 9092 5322 9104
rect 5537 9095 5595 9101
rect 5537 9092 5549 9095
rect 5316 9064 5549 9092
rect 5316 9052 5322 9064
rect 5537 9061 5549 9064
rect 5583 9061 5595 9095
rect 5537 9055 5595 9061
rect 4890 9024 4896 9036
rect 3528 8996 4896 9024
rect 3528 8965 3556 8996
rect 4890 8984 4896 8996
rect 4948 9024 4954 9036
rect 5074 9024 5080 9036
rect 4948 8996 5080 9024
rect 4948 8984 4954 8996
rect 5074 8984 5080 8996
rect 5132 8984 5138 9036
rect 2547 8928 3464 8956
rect 3513 8959 3571 8965
rect 2547 8925 2559 8928
rect 2501 8919 2559 8925
rect 3513 8925 3525 8959
rect 3559 8925 3571 8959
rect 3513 8919 3571 8925
rect 4525 8959 4583 8965
rect 4525 8925 4537 8959
rect 4571 8925 4583 8959
rect 4525 8919 4583 8925
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8956 4767 8959
rect 5350 8956 5356 8968
rect 4755 8928 5356 8956
rect 4755 8925 4767 8928
rect 4709 8919 4767 8925
rect 2869 8891 2927 8897
rect 2869 8857 2881 8891
rect 2915 8888 2927 8891
rect 4540 8888 4568 8919
rect 5350 8916 5356 8928
rect 5408 8956 5414 8968
rect 5721 8959 5779 8965
rect 5721 8956 5733 8959
rect 5408 8928 5733 8956
rect 5408 8916 5414 8928
rect 5721 8925 5733 8928
rect 5767 8956 5779 8959
rect 5828 8956 5856 9132
rect 7006 9120 7012 9132
rect 7064 9120 7070 9172
rect 7282 9120 7288 9172
rect 7340 9160 7346 9172
rect 7929 9163 7987 9169
rect 7929 9160 7941 9163
rect 7340 9132 7941 9160
rect 7340 9120 7346 9132
rect 7929 9129 7941 9132
rect 7975 9129 7987 9163
rect 7929 9123 7987 9129
rect 8021 9163 8079 9169
rect 8021 9129 8033 9163
rect 8067 9160 8079 9163
rect 8573 9163 8631 9169
rect 8067 9132 8524 9160
rect 8067 9129 8079 9132
rect 8021 9123 8079 9129
rect 8496 9104 8524 9132
rect 8573 9129 8585 9163
rect 8619 9129 8631 9163
rect 8938 9160 8944 9172
rect 8899 9132 8944 9160
rect 8573 9123 8631 9129
rect 8389 9095 8447 9101
rect 8389 9092 8401 9095
rect 7392 9064 8401 9092
rect 6917 9027 6975 9033
rect 6917 8993 6929 9027
rect 6963 9024 6975 9027
rect 6963 8996 7144 9024
rect 6963 8993 6975 8996
rect 6917 8987 6975 8993
rect 5767 8928 5856 8956
rect 5767 8925 5779 8928
rect 5721 8919 5779 8925
rect 6362 8916 6368 8968
rect 6420 8956 6426 8968
rect 6546 8956 6552 8968
rect 6420 8928 6552 8956
rect 6420 8916 6426 8928
rect 6546 8916 6552 8928
rect 6604 8916 6610 8968
rect 7006 8956 7012 8968
rect 6967 8928 7012 8956
rect 7006 8916 7012 8928
rect 7064 8916 7070 8968
rect 2915 8860 4568 8888
rect 7116 8888 7144 8996
rect 7193 8959 7251 8965
rect 7193 8925 7205 8959
rect 7239 8956 7251 8959
rect 7392 8956 7420 9064
rect 8389 9061 8401 9064
rect 8435 9061 8447 9095
rect 8389 9055 8447 9061
rect 8478 9052 8484 9104
rect 8536 9052 8542 9104
rect 8588 9092 8616 9123
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 9490 9160 9496 9172
rect 9048 9132 9496 9160
rect 9048 9101 9076 9132
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 10229 9163 10287 9169
rect 10229 9129 10241 9163
rect 10275 9160 10287 9163
rect 10410 9160 10416 9172
rect 10275 9132 10416 9160
rect 10275 9129 10287 9132
rect 10229 9123 10287 9129
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 11609 9163 11667 9169
rect 11609 9129 11621 9163
rect 11655 9129 11667 9163
rect 12986 9160 12992 9172
rect 11609 9123 11667 9129
rect 12820 9132 12992 9160
rect 9033 9095 9091 9101
rect 8588 9064 8984 9092
rect 8018 8984 8024 9036
rect 8076 9024 8082 9036
rect 8662 9024 8668 9036
rect 8076 8996 8668 9024
rect 8076 8984 8082 8996
rect 8662 8984 8668 8996
rect 8720 8984 8726 9036
rect 8956 9024 8984 9064
rect 9033 9061 9045 9095
rect 9079 9061 9091 9095
rect 9033 9055 9091 9061
rect 9122 9052 9128 9104
rect 9180 9092 9186 9104
rect 11624 9092 11652 9123
rect 11977 9095 12035 9101
rect 11977 9092 11989 9095
rect 9180 9064 11652 9092
rect 11900 9064 11989 9092
rect 9180 9052 9186 9064
rect 10045 9027 10103 9033
rect 10045 9024 10057 9027
rect 8956 8996 10057 9024
rect 10045 8993 10057 8996
rect 10091 8993 10103 9027
rect 10045 8987 10103 8993
rect 10870 8984 10876 9036
rect 10928 9024 10934 9036
rect 10965 9027 11023 9033
rect 10965 9024 10977 9027
rect 10928 8996 10977 9024
rect 10928 8984 10934 8996
rect 10965 8993 10977 8996
rect 11011 8993 11023 9027
rect 10965 8987 11023 8993
rect 11330 8984 11336 9036
rect 11388 9024 11394 9036
rect 11900 9024 11928 9064
rect 11977 9061 11989 9064
rect 12023 9061 12035 9095
rect 11977 9055 12035 9061
rect 12069 9027 12127 9033
rect 12069 9024 12081 9027
rect 11388 8996 11928 9024
rect 11992 8996 12081 9024
rect 11388 8984 11394 8996
rect 8113 8959 8171 8965
rect 7239 8928 7420 8956
rect 7484 8928 8064 8956
rect 7239 8925 7251 8928
rect 7193 8919 7251 8925
rect 7484 8888 7512 8928
rect 7116 8860 7512 8888
rect 7561 8891 7619 8897
rect 2915 8857 2927 8860
rect 2869 8851 2927 8857
rect 7561 8857 7573 8891
rect 7607 8888 7619 8891
rect 7650 8888 7656 8900
rect 7607 8860 7656 8888
rect 7607 8857 7619 8860
rect 7561 8851 7619 8857
rect 7650 8848 7656 8860
rect 7708 8848 7714 8900
rect 8036 8888 8064 8928
rect 8113 8925 8125 8959
rect 8159 8956 8171 8959
rect 8754 8956 8760 8968
rect 8159 8928 8760 8956
rect 8159 8925 8171 8928
rect 8113 8919 8171 8925
rect 8754 8916 8760 8928
rect 8812 8916 8818 8968
rect 9214 8956 9220 8968
rect 9175 8928 9220 8956
rect 9214 8916 9220 8928
rect 9272 8916 9278 8968
rect 10134 8916 10140 8968
rect 10192 8956 10198 8968
rect 11057 8959 11115 8965
rect 11057 8956 11069 8959
rect 10192 8928 11069 8956
rect 10192 8916 10198 8928
rect 11057 8925 11069 8928
rect 11103 8925 11115 8959
rect 11057 8919 11115 8925
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 8202 8888 8208 8900
rect 8036 8860 8208 8888
rect 8202 8848 8208 8860
rect 8260 8848 8266 8900
rect 8386 8848 8392 8900
rect 8444 8888 8450 8900
rect 8444 8860 8489 8888
rect 8444 8848 8450 8860
rect 8662 8848 8668 8900
rect 8720 8888 8726 8900
rect 9858 8888 9864 8900
rect 8720 8860 9864 8888
rect 8720 8848 8726 8860
rect 9858 8848 9864 8860
rect 9916 8848 9922 8900
rect 11146 8848 11152 8900
rect 11204 8848 11210 8900
rect 11256 8888 11284 8919
rect 11422 8916 11428 8968
rect 11480 8956 11486 8968
rect 11992 8956 12020 8996
rect 12069 8993 12081 8996
rect 12115 8993 12127 9027
rect 12069 8987 12127 8993
rect 11480 8928 12020 8956
rect 12253 8959 12311 8965
rect 11480 8916 11486 8928
rect 12253 8925 12265 8959
rect 12299 8956 12311 8959
rect 12342 8956 12348 8968
rect 12299 8928 12348 8956
rect 12299 8925 12311 8928
rect 12253 8919 12311 8925
rect 12268 8888 12296 8919
rect 12342 8916 12348 8928
rect 12400 8916 12406 8968
rect 12820 8956 12848 9132
rect 12986 9120 12992 9132
rect 13044 9120 13050 9172
rect 13173 9163 13231 9169
rect 13173 9129 13185 9163
rect 13219 9160 13231 9163
rect 13354 9160 13360 9172
rect 13219 9132 13360 9160
rect 13219 9129 13231 9132
rect 13173 9123 13231 9129
rect 13354 9120 13360 9132
rect 13412 9120 13418 9172
rect 13630 9120 13636 9172
rect 13688 9160 13694 9172
rect 15841 9163 15899 9169
rect 13688 9132 15240 9160
rect 13688 9120 13694 9132
rect 15212 9104 15240 9132
rect 15841 9129 15853 9163
rect 15887 9160 15899 9163
rect 22278 9160 22284 9172
rect 15887 9132 22284 9160
rect 15887 9129 15899 9132
rect 15841 9123 15899 9129
rect 22278 9120 22284 9132
rect 22336 9120 22342 9172
rect 22646 9160 22652 9172
rect 22607 9132 22652 9160
rect 22646 9120 22652 9132
rect 22704 9120 22710 9172
rect 13262 9092 13268 9104
rect 12912 9064 13268 9092
rect 12912 9033 12940 9064
rect 13262 9052 13268 9064
rect 13320 9092 13326 9104
rect 14918 9092 14924 9104
rect 13320 9064 14924 9092
rect 13320 9052 13326 9064
rect 14918 9052 14924 9064
rect 14976 9052 14982 9104
rect 15194 9052 15200 9104
rect 15252 9052 15258 9104
rect 15933 9095 15991 9101
rect 15933 9061 15945 9095
rect 15979 9092 15991 9095
rect 17218 9092 17224 9104
rect 15979 9064 17224 9092
rect 15979 9061 15991 9064
rect 15933 9055 15991 9061
rect 17218 9052 17224 9064
rect 17276 9052 17282 9104
rect 17586 9052 17592 9104
rect 17644 9092 17650 9104
rect 17862 9092 17868 9104
rect 17644 9064 17868 9092
rect 17644 9052 17650 9064
rect 17862 9052 17868 9064
rect 17920 9052 17926 9104
rect 12897 9027 12955 9033
rect 12897 8993 12909 9027
rect 12943 8993 12955 9027
rect 12897 8987 12955 8993
rect 12986 8984 12992 9036
rect 13044 9024 13050 9036
rect 13808 9027 13866 9033
rect 13044 8996 13089 9024
rect 13044 8984 13050 8996
rect 13808 8993 13820 9027
rect 13854 9024 13866 9027
rect 14826 9024 14832 9036
rect 13854 8996 14832 9024
rect 13854 8993 13866 8996
rect 13808 8987 13866 8993
rect 14826 8984 14832 8996
rect 14884 8984 14890 9036
rect 16390 8984 16396 9036
rect 16448 9024 16454 9036
rect 16485 9027 16543 9033
rect 16485 9024 16497 9027
rect 16448 8996 16497 9024
rect 16448 8984 16454 8996
rect 16485 8993 16497 8996
rect 16531 8993 16543 9027
rect 16485 8987 16543 8993
rect 16752 9027 16810 9033
rect 16752 8993 16764 9027
rect 16798 9024 16810 9027
rect 17494 9024 17500 9036
rect 16798 8996 17500 9024
rect 16798 8993 16810 8996
rect 16752 8987 16810 8993
rect 17494 8984 17500 8996
rect 17552 8984 17558 9036
rect 18046 8984 18052 9036
rect 18104 9024 18110 9036
rect 18690 9033 18696 9036
rect 18648 9027 18696 9033
rect 18648 9024 18660 9027
rect 18104 8996 18368 9024
rect 18603 8996 18660 9024
rect 18104 8984 18110 8996
rect 13354 8956 13360 8968
rect 12820 8928 13360 8956
rect 13354 8916 13360 8928
rect 13412 8956 13418 8968
rect 13541 8959 13599 8965
rect 13541 8956 13553 8959
rect 13412 8928 13553 8956
rect 13412 8916 13418 8928
rect 13541 8925 13553 8928
rect 13587 8925 13599 8959
rect 13541 8919 13599 8925
rect 16117 8959 16175 8965
rect 16117 8925 16129 8959
rect 16163 8956 16175 8959
rect 16298 8956 16304 8968
rect 16163 8928 16304 8956
rect 16163 8925 16175 8928
rect 16117 8919 16175 8925
rect 16298 8916 16304 8928
rect 16356 8916 16362 8968
rect 18230 8956 18236 8968
rect 17512 8928 18236 8956
rect 11256 8860 12296 8888
rect 14734 8848 14740 8900
rect 14792 8888 14798 8900
rect 14792 8860 15599 8888
rect 14792 8848 14798 8860
rect 1857 8823 1915 8829
rect 1857 8789 1869 8823
rect 1903 8820 1915 8823
rect 6362 8820 6368 8832
rect 1903 8792 6368 8820
rect 1903 8789 1915 8792
rect 1857 8783 1915 8789
rect 6362 8780 6368 8792
rect 6420 8780 6426 8832
rect 6549 8823 6607 8829
rect 6549 8789 6561 8823
rect 6595 8820 6607 8823
rect 8754 8820 8760 8832
rect 6595 8792 8760 8820
rect 6595 8789 6607 8792
rect 6549 8783 6607 8789
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 10597 8823 10655 8829
rect 10597 8820 10609 8823
rect 9732 8792 10609 8820
rect 9732 8780 9738 8792
rect 10597 8789 10609 8792
rect 10643 8789 10655 8823
rect 11164 8820 11192 8848
rect 11606 8820 11612 8832
rect 11164 8792 11612 8820
rect 10597 8783 10655 8789
rect 11606 8780 11612 8792
rect 11664 8780 11670 8832
rect 12710 8820 12716 8832
rect 12671 8792 12716 8820
rect 12710 8780 12716 8792
rect 12768 8780 12774 8832
rect 14918 8820 14924 8832
rect 14879 8792 14924 8820
rect 14918 8780 14924 8792
rect 14976 8780 14982 8832
rect 15194 8780 15200 8832
rect 15252 8820 15258 8832
rect 15473 8823 15531 8829
rect 15473 8820 15485 8823
rect 15252 8792 15485 8820
rect 15252 8780 15258 8792
rect 15473 8789 15485 8792
rect 15519 8789 15531 8823
rect 15571 8820 15599 8860
rect 17512 8820 17540 8928
rect 18230 8916 18236 8928
rect 18288 8916 18294 8968
rect 18340 8965 18368 8996
rect 18648 8993 18660 8996
rect 18694 8993 18696 9027
rect 18648 8987 18696 8993
rect 18690 8984 18696 8987
rect 18748 9024 18754 9036
rect 18966 9024 18972 9036
rect 18748 8996 18972 9024
rect 18748 8984 18754 8996
rect 18966 8984 18972 8996
rect 19024 8984 19030 9036
rect 19150 8984 19156 9036
rect 19208 9024 19214 9036
rect 21525 9027 21583 9033
rect 21525 9024 21537 9027
rect 19208 8996 21537 9024
rect 19208 8984 19214 8996
rect 21525 8993 21537 8996
rect 21571 9024 21583 9027
rect 22094 9024 22100 9036
rect 21571 8996 22100 9024
rect 21571 8993 21583 8996
rect 21525 8987 21583 8993
rect 22094 8984 22100 8996
rect 22152 8984 22158 9036
rect 18325 8959 18383 8965
rect 18325 8925 18337 8959
rect 18371 8956 18383 8959
rect 18506 8956 18512 8968
rect 18371 8928 18512 8956
rect 18371 8925 18383 8928
rect 18325 8919 18383 8925
rect 18506 8916 18512 8928
rect 18564 8916 18570 8968
rect 18874 8965 18880 8968
rect 18831 8959 18880 8965
rect 18831 8925 18843 8959
rect 18877 8925 18880 8959
rect 18831 8919 18880 8925
rect 18874 8916 18880 8919
rect 18932 8916 18938 8968
rect 19058 8956 19064 8968
rect 19019 8928 19064 8956
rect 19058 8916 19064 8928
rect 19116 8916 19122 8968
rect 20714 8916 20720 8968
rect 20772 8956 20778 8968
rect 21269 8959 21327 8965
rect 21269 8956 21281 8959
rect 20772 8928 21281 8956
rect 20772 8916 20778 8928
rect 21269 8925 21281 8928
rect 21315 8925 21327 8959
rect 21269 8919 21327 8925
rect 17770 8848 17776 8900
rect 17828 8888 17834 8900
rect 20162 8888 20168 8900
rect 17828 8860 18184 8888
rect 20123 8860 20168 8888
rect 17828 8848 17834 8860
rect 15571 8792 17540 8820
rect 15473 8783 15531 8789
rect 17586 8780 17592 8832
rect 17644 8820 17650 8832
rect 17865 8823 17923 8829
rect 17865 8820 17877 8823
rect 17644 8792 17877 8820
rect 17644 8780 17650 8792
rect 17865 8789 17877 8792
rect 17911 8789 17923 8823
rect 18156 8820 18184 8860
rect 20162 8848 20168 8860
rect 20220 8848 20226 8900
rect 22186 8820 22192 8832
rect 18156 8792 22192 8820
rect 17865 8783 17923 8789
rect 22186 8780 22192 8792
rect 22244 8780 22250 8832
rect 1104 8730 23276 8752
rect 1104 8678 4680 8730
rect 4732 8678 4744 8730
rect 4796 8678 4808 8730
rect 4860 8678 4872 8730
rect 4924 8678 12078 8730
rect 12130 8678 12142 8730
rect 12194 8678 12206 8730
rect 12258 8678 12270 8730
rect 12322 8678 19475 8730
rect 19527 8678 19539 8730
rect 19591 8678 19603 8730
rect 19655 8678 19667 8730
rect 19719 8678 23276 8730
rect 1104 8656 23276 8678
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 2961 8619 3019 8625
rect 2961 8616 2973 8619
rect 2924 8588 2973 8616
rect 2924 8576 2930 8588
rect 2961 8585 2973 8588
rect 3007 8585 3019 8619
rect 2961 8579 3019 8585
rect 3602 8576 3608 8628
rect 3660 8616 3666 8628
rect 3789 8619 3847 8625
rect 3789 8616 3801 8619
rect 3660 8588 3801 8616
rect 3660 8576 3666 8588
rect 3789 8585 3801 8588
rect 3835 8585 3847 8619
rect 3789 8579 3847 8585
rect 3878 8576 3884 8628
rect 3936 8616 3942 8628
rect 4157 8619 4215 8625
rect 4157 8616 4169 8619
rect 3936 8588 4169 8616
rect 3936 8576 3942 8588
rect 4157 8585 4169 8588
rect 4203 8585 4215 8619
rect 4157 8579 4215 8585
rect 4709 8619 4767 8625
rect 4709 8585 4721 8619
rect 4755 8616 4767 8619
rect 6730 8616 6736 8628
rect 4755 8588 6736 8616
rect 4755 8585 4767 8588
rect 4709 8579 4767 8585
rect 6730 8576 6736 8588
rect 6788 8576 6794 8628
rect 7009 8619 7067 8625
rect 7009 8585 7021 8619
rect 7055 8616 7067 8619
rect 7558 8616 7564 8628
rect 7055 8588 7564 8616
rect 7055 8585 7067 8588
rect 7009 8579 7067 8585
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 7745 8619 7803 8625
rect 7745 8585 7757 8619
rect 7791 8616 7803 8619
rect 8662 8616 8668 8628
rect 7791 8588 8668 8616
rect 7791 8585 7803 8588
rect 7745 8579 7803 8585
rect 8662 8576 8668 8588
rect 8720 8576 8726 8628
rect 9398 8616 9404 8628
rect 8864 8588 9404 8616
rect 1949 8551 2007 8557
rect 1949 8517 1961 8551
rect 1995 8548 2007 8551
rect 4062 8548 4068 8560
rect 1995 8520 4068 8548
rect 1995 8517 2007 8520
rect 1949 8511 2007 8517
rect 4062 8508 4068 8520
rect 4120 8508 4126 8560
rect 5350 8548 5356 8560
rect 5000 8520 5356 8548
rect 2590 8480 2596 8492
rect 2551 8452 2596 8480
rect 2590 8440 2596 8452
rect 2648 8440 2654 8492
rect 3050 8440 3056 8492
rect 3108 8480 3114 8492
rect 3421 8483 3479 8489
rect 3421 8480 3433 8483
rect 3108 8452 3433 8480
rect 3108 8440 3114 8452
rect 3421 8449 3433 8452
rect 3467 8449 3479 8483
rect 3421 8443 3479 8449
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8480 3663 8483
rect 5000 8480 5028 8520
rect 5350 8508 5356 8520
rect 5408 8508 5414 8560
rect 5721 8551 5779 8557
rect 5721 8517 5733 8551
rect 5767 8548 5779 8551
rect 8202 8548 8208 8560
rect 5767 8520 8208 8548
rect 5767 8517 5779 8520
rect 5721 8511 5779 8517
rect 8202 8508 8208 8520
rect 8260 8508 8266 8560
rect 5166 8480 5172 8492
rect 3651 8452 5028 8480
rect 5127 8452 5172 8480
rect 3651 8449 3663 8452
rect 3605 8443 3663 8449
rect 5166 8440 5172 8452
rect 5224 8440 5230 8492
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 5534 8480 5540 8492
rect 5307 8452 5540 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8480 6423 8483
rect 8294 8480 8300 8492
rect 6411 8452 8300 8480
rect 6411 8449 6423 8452
rect 6365 8443 6423 8449
rect 8294 8440 8300 8452
rect 8352 8440 8358 8492
rect 8386 8440 8392 8492
rect 8444 8480 8450 8492
rect 8864 8480 8892 8588
rect 9398 8576 9404 8588
rect 9456 8576 9462 8628
rect 9585 8619 9643 8625
rect 9585 8585 9597 8619
rect 9631 8616 9643 8619
rect 9674 8616 9680 8628
rect 9631 8588 9680 8616
rect 9631 8585 9643 8588
rect 9585 8579 9643 8585
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 9766 8576 9772 8628
rect 9824 8616 9830 8628
rect 11977 8619 12035 8625
rect 11977 8616 11989 8619
rect 9824 8588 11989 8616
rect 9824 8576 9830 8588
rect 11977 8585 11989 8588
rect 12023 8585 12035 8619
rect 11977 8579 12035 8585
rect 12526 8576 12532 8628
rect 12584 8616 12590 8628
rect 13081 8619 13139 8625
rect 13081 8616 13093 8619
rect 12584 8588 13093 8616
rect 12584 8576 12590 8588
rect 13081 8585 13093 8588
rect 13127 8616 13139 8619
rect 13998 8616 14004 8628
rect 13127 8588 14004 8616
rect 13127 8585 13139 8588
rect 13081 8579 13139 8585
rect 13998 8576 14004 8588
rect 14056 8576 14062 8628
rect 14737 8619 14795 8625
rect 14737 8585 14749 8619
rect 14783 8616 14795 8619
rect 14826 8616 14832 8628
rect 14783 8588 14832 8616
rect 14783 8585 14795 8588
rect 14737 8579 14795 8585
rect 14826 8576 14832 8588
rect 14884 8576 14890 8628
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8616 15255 8619
rect 15470 8616 15476 8628
rect 15243 8588 15476 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 16298 8576 16304 8628
rect 16356 8616 16362 8628
rect 16945 8619 17003 8625
rect 16356 8588 16896 8616
rect 16356 8576 16362 8588
rect 9214 8508 9220 8560
rect 9272 8548 9278 8560
rect 11149 8551 11207 8557
rect 9272 8520 9352 8548
rect 9272 8508 9278 8520
rect 9324 8489 9352 8520
rect 11149 8517 11161 8551
rect 11195 8548 11207 8551
rect 11238 8548 11244 8560
rect 11195 8520 11244 8548
rect 11195 8517 11207 8520
rect 11149 8511 11207 8517
rect 11238 8508 11244 8520
rect 11296 8508 11302 8560
rect 11422 8508 11428 8560
rect 11480 8548 11486 8560
rect 12621 8551 12679 8557
rect 12621 8548 12633 8551
rect 11480 8520 12633 8548
rect 11480 8508 11486 8520
rect 12621 8517 12633 8520
rect 12667 8517 12679 8551
rect 12621 8511 12679 8517
rect 14918 8508 14924 8560
rect 14976 8548 14982 8560
rect 15381 8551 15439 8557
rect 15381 8548 15393 8551
rect 14976 8520 15393 8548
rect 14976 8508 14982 8520
rect 15381 8517 15393 8520
rect 15427 8517 15439 8551
rect 16868 8548 16896 8588
rect 16945 8585 16957 8619
rect 16991 8616 17003 8619
rect 17494 8616 17500 8628
rect 16991 8588 17500 8616
rect 16991 8585 17003 8588
rect 16945 8579 17003 8585
rect 17494 8576 17500 8588
rect 17552 8576 17558 8628
rect 18141 8619 18199 8625
rect 18141 8585 18153 8619
rect 18187 8616 18199 8619
rect 18598 8616 18604 8628
rect 18187 8588 18604 8616
rect 18187 8585 18199 8588
rect 18141 8579 18199 8585
rect 18598 8576 18604 8588
rect 18656 8576 18662 8628
rect 20533 8619 20591 8625
rect 20533 8616 20545 8619
rect 19168 8588 20545 8616
rect 19168 8548 19196 8588
rect 20533 8585 20545 8588
rect 20579 8585 20591 8619
rect 20533 8579 20591 8585
rect 16868 8520 19196 8548
rect 15381 8511 15439 8517
rect 8444 8452 8489 8480
rect 8680 8452 8892 8480
rect 9309 8483 9367 8489
rect 8444 8440 8450 8452
rect 2317 8415 2375 8421
rect 2317 8381 2329 8415
rect 2363 8412 2375 8415
rect 3234 8412 3240 8424
rect 2363 8384 3240 8412
rect 2363 8381 2375 8384
rect 2317 8375 2375 8381
rect 3234 8372 3240 8384
rect 3292 8372 3298 8424
rect 3329 8415 3387 8421
rect 3329 8381 3341 8415
rect 3375 8412 3387 8415
rect 3694 8412 3700 8424
rect 3375 8384 3700 8412
rect 3375 8381 3387 8384
rect 3329 8375 3387 8381
rect 3694 8372 3700 8384
rect 3752 8372 3758 8424
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8412 3847 8415
rect 3973 8415 4031 8421
rect 3973 8412 3985 8415
rect 3835 8384 3985 8412
rect 3835 8381 3847 8384
rect 3789 8375 3847 8381
rect 3973 8381 3985 8384
rect 4019 8381 4031 8415
rect 3973 8375 4031 8381
rect 5077 8415 5135 8421
rect 5077 8381 5089 8415
rect 5123 8412 5135 8415
rect 5626 8412 5632 8424
rect 5123 8384 5632 8412
rect 5123 8381 5135 8384
rect 5077 8375 5135 8381
rect 5626 8372 5632 8384
rect 5684 8372 5690 8424
rect 6730 8372 6736 8424
rect 6788 8412 6794 8424
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 6788 8384 6837 8412
rect 6788 8372 6794 8384
rect 6825 8381 6837 8384
rect 6871 8381 6883 8415
rect 6825 8375 6883 8381
rect 7650 8372 7656 8424
rect 7708 8412 7714 8424
rect 8478 8412 8484 8424
rect 7708 8384 8484 8412
rect 7708 8372 7714 8384
rect 8478 8372 8484 8384
rect 8536 8372 8542 8424
rect 2409 8347 2467 8353
rect 2409 8313 2421 8347
rect 2455 8344 2467 8347
rect 4154 8344 4160 8356
rect 2455 8316 4160 8344
rect 2455 8313 2467 8316
rect 2409 8307 2467 8313
rect 4154 8304 4160 8316
rect 4212 8304 4218 8356
rect 6089 8347 6147 8353
rect 6089 8313 6101 8347
rect 6135 8344 6147 8347
rect 7926 8344 7932 8356
rect 6135 8316 7932 8344
rect 6135 8313 6147 8316
rect 6089 8307 6147 8313
rect 7926 8304 7932 8316
rect 7984 8304 7990 8356
rect 8113 8347 8171 8353
rect 8113 8313 8125 8347
rect 8159 8344 8171 8347
rect 8570 8344 8576 8356
rect 8159 8316 8576 8344
rect 8159 8313 8171 8316
rect 8113 8307 8171 8313
rect 8570 8304 8576 8316
rect 8628 8304 8634 8356
rect 6181 8279 6239 8285
rect 6181 8245 6193 8279
rect 6227 8276 6239 8279
rect 6730 8276 6736 8288
rect 6227 8248 6736 8276
rect 6227 8245 6239 8248
rect 6181 8239 6239 8245
rect 6730 8236 6736 8248
rect 6788 8236 6794 8288
rect 8205 8279 8263 8285
rect 8205 8245 8217 8279
rect 8251 8276 8263 8279
rect 8680 8276 8708 8452
rect 9309 8449 9321 8483
rect 9355 8449 9367 8483
rect 9766 8480 9772 8492
rect 9727 8452 9772 8480
rect 9309 8443 9367 8449
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 10870 8440 10876 8492
rect 10928 8480 10934 8492
rect 12066 8480 12072 8492
rect 10928 8452 12072 8480
rect 10928 8440 10934 8452
rect 12066 8440 12072 8452
rect 12124 8440 12130 8492
rect 13354 8480 13360 8492
rect 13315 8452 13360 8480
rect 13354 8440 13360 8452
rect 13412 8440 13418 8492
rect 15102 8440 15108 8492
rect 15160 8480 15166 8492
rect 15160 8452 15700 8480
rect 15160 8440 15166 8452
rect 11425 8415 11483 8421
rect 11425 8412 11437 8415
rect 9048 8384 11437 8412
rect 9048 8344 9076 8384
rect 11425 8381 11437 8384
rect 11471 8381 11483 8415
rect 11425 8375 11483 8381
rect 11606 8372 11612 8424
rect 11664 8412 11670 8424
rect 12161 8415 12219 8421
rect 12161 8412 12173 8415
rect 11664 8384 12173 8412
rect 11664 8372 11670 8384
rect 12161 8381 12173 8384
rect 12207 8381 12219 8415
rect 12161 8375 12219 8381
rect 12434 8372 12440 8424
rect 12492 8412 12498 8424
rect 13262 8412 13268 8424
rect 12492 8384 12537 8412
rect 13223 8384 13268 8412
rect 12492 8372 12498 8384
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 13624 8415 13682 8421
rect 13624 8381 13636 8415
rect 13670 8412 13682 8415
rect 14090 8412 14096 8424
rect 13670 8384 14096 8412
rect 13670 8381 13682 8384
rect 13624 8375 13682 8381
rect 14090 8372 14096 8384
rect 14148 8372 14154 8424
rect 15010 8412 15016 8424
rect 14971 8384 15016 8412
rect 15010 8372 15016 8384
rect 15068 8372 15074 8424
rect 15470 8372 15476 8424
rect 15528 8412 15534 8424
rect 15565 8415 15623 8421
rect 15565 8412 15577 8415
rect 15528 8384 15577 8412
rect 15528 8372 15534 8384
rect 15565 8381 15577 8384
rect 15611 8381 15623 8415
rect 15672 8412 15700 8452
rect 16850 8440 16856 8492
rect 16908 8480 16914 8492
rect 17405 8483 17463 8489
rect 17405 8480 17417 8483
rect 16908 8452 17417 8480
rect 16908 8440 16914 8452
rect 17405 8449 17417 8452
rect 17451 8449 17463 8483
rect 18782 8480 18788 8492
rect 18743 8452 18788 8480
rect 17405 8443 17463 8449
rect 18782 8440 18788 8452
rect 18840 8440 18846 8492
rect 20548 8480 20576 8579
rect 22094 8576 22100 8628
rect 22152 8616 22158 8628
rect 22189 8619 22247 8625
rect 22189 8616 22201 8619
rect 22152 8588 22201 8616
rect 22152 8576 22158 8588
rect 22189 8585 22201 8588
rect 22235 8585 22247 8619
rect 22189 8579 22247 8585
rect 22649 8551 22707 8557
rect 22649 8517 22661 8551
rect 22695 8517 22707 8551
rect 22649 8511 22707 8517
rect 22664 8480 22692 8511
rect 20548 8452 20944 8480
rect 17218 8412 17224 8424
rect 15672 8384 17224 8412
rect 15565 8375 15623 8381
rect 17218 8372 17224 8384
rect 17276 8372 17282 8424
rect 18509 8415 18567 8421
rect 18509 8381 18521 8415
rect 18555 8412 18567 8415
rect 19150 8412 19156 8424
rect 18555 8384 19012 8412
rect 19111 8384 19156 8412
rect 18555 8381 18567 8384
rect 18509 8375 18567 8381
rect 8772 8316 9076 8344
rect 8772 8285 8800 8316
rect 9122 8304 9128 8356
rect 9180 8344 9186 8356
rect 9585 8347 9643 8353
rect 9585 8344 9597 8347
rect 9180 8316 9225 8344
rect 9324 8316 9597 8344
rect 9180 8304 9186 8316
rect 8251 8248 8708 8276
rect 8757 8279 8815 8285
rect 8251 8245 8263 8248
rect 8205 8239 8263 8245
rect 8757 8245 8769 8279
rect 8803 8245 8815 8279
rect 8757 8239 8815 8245
rect 9217 8279 9275 8285
rect 9217 8245 9229 8279
rect 9263 8276 9275 8279
rect 9324 8276 9352 8316
rect 9585 8313 9597 8316
rect 9631 8313 9643 8347
rect 9585 8307 9643 8313
rect 10036 8347 10094 8353
rect 10036 8313 10048 8347
rect 10082 8344 10094 8347
rect 10870 8344 10876 8356
rect 10082 8316 10876 8344
rect 10082 8313 10094 8316
rect 10036 8307 10094 8313
rect 10870 8304 10876 8316
rect 10928 8304 10934 8356
rect 12710 8304 12716 8356
rect 12768 8344 12774 8356
rect 15381 8347 15439 8353
rect 12768 8316 15332 8344
rect 12768 8304 12774 8316
rect 11606 8276 11612 8288
rect 9263 8248 9352 8276
rect 11567 8248 11612 8276
rect 9263 8245 9275 8248
rect 9217 8239 9275 8245
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 15304 8276 15332 8316
rect 15381 8313 15393 8347
rect 15427 8344 15439 8347
rect 15810 8347 15868 8353
rect 15810 8344 15822 8347
rect 15427 8316 15822 8344
rect 15427 8313 15439 8316
rect 15381 8307 15439 8313
rect 15810 8313 15822 8316
rect 15856 8313 15868 8347
rect 15810 8307 15868 8313
rect 15948 8316 17816 8344
rect 15948 8276 15976 8316
rect 15304 8248 15976 8276
rect 17788 8276 17816 8316
rect 17862 8304 17868 8356
rect 17920 8344 17926 8356
rect 18601 8347 18659 8353
rect 18601 8344 18613 8347
rect 17920 8316 18613 8344
rect 17920 8304 17926 8316
rect 18601 8313 18613 8316
rect 18647 8313 18659 8347
rect 18984 8344 19012 8384
rect 19150 8372 19156 8384
rect 19208 8372 19214 8424
rect 19426 8421 19432 8424
rect 19420 8412 19432 8421
rect 19339 8384 19432 8412
rect 19420 8375 19432 8384
rect 19484 8412 19490 8424
rect 19794 8412 19800 8424
rect 19484 8384 19800 8412
rect 19426 8372 19432 8375
rect 19484 8372 19490 8384
rect 19794 8372 19800 8384
rect 19852 8372 19858 8424
rect 20714 8372 20720 8424
rect 20772 8412 20778 8424
rect 20809 8415 20867 8421
rect 20809 8412 20821 8415
rect 20772 8384 20821 8412
rect 20772 8372 20778 8384
rect 20809 8381 20821 8384
rect 20855 8381 20867 8415
rect 20916 8412 20944 8452
rect 22112 8452 22692 8480
rect 21065 8415 21123 8421
rect 21065 8412 21077 8415
rect 20916 8384 21077 8412
rect 20809 8375 20867 8381
rect 21065 8381 21077 8384
rect 21111 8381 21123 8415
rect 21065 8375 21123 8381
rect 21358 8372 21364 8424
rect 21416 8412 21422 8424
rect 22112 8412 22140 8452
rect 22462 8412 22468 8424
rect 21416 8384 22140 8412
rect 22423 8384 22468 8412
rect 21416 8372 21422 8384
rect 22462 8372 22468 8384
rect 22520 8372 22526 8424
rect 19058 8344 19064 8356
rect 18971 8316 19064 8344
rect 18601 8307 18659 8313
rect 19058 8304 19064 8316
rect 19116 8344 19122 8356
rect 19886 8344 19892 8356
rect 19116 8316 19892 8344
rect 19116 8304 19122 8316
rect 19886 8304 19892 8316
rect 19944 8304 19950 8356
rect 20438 8344 20444 8356
rect 19996 8316 20444 8344
rect 19996 8288 20024 8316
rect 20438 8304 20444 8316
rect 20496 8304 20502 8356
rect 19978 8276 19984 8288
rect 17788 8248 19984 8276
rect 19978 8236 19984 8248
rect 20036 8236 20042 8288
rect 1104 8186 23276 8208
rect 1104 8134 8379 8186
rect 8431 8134 8443 8186
rect 8495 8134 8507 8186
rect 8559 8134 8571 8186
rect 8623 8134 15776 8186
rect 15828 8134 15840 8186
rect 15892 8134 15904 8186
rect 15956 8134 15968 8186
rect 16020 8134 23276 8186
rect 1104 8112 23276 8134
rect 5074 8032 5080 8084
rect 5132 8072 5138 8084
rect 5905 8075 5963 8081
rect 5905 8072 5917 8075
rect 5132 8044 5917 8072
rect 5132 8032 5138 8044
rect 5905 8041 5917 8044
rect 5951 8041 5963 8075
rect 5905 8035 5963 8041
rect 6917 8075 6975 8081
rect 6917 8041 6929 8075
rect 6963 8072 6975 8075
rect 7006 8072 7012 8084
rect 6963 8044 7012 8072
rect 6963 8041 6975 8044
rect 6917 8035 6975 8041
rect 7006 8032 7012 8044
rect 7064 8032 7070 8084
rect 8938 8072 8944 8084
rect 8899 8044 8944 8072
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 9033 8075 9091 8081
rect 9033 8041 9045 8075
rect 9079 8072 9091 8075
rect 11606 8072 11612 8084
rect 9079 8044 11612 8072
rect 9079 8041 9091 8044
rect 9033 8035 9091 8041
rect 11606 8032 11612 8044
rect 11664 8032 11670 8084
rect 11698 8032 11704 8084
rect 11756 8032 11762 8084
rect 12066 8032 12072 8084
rect 12124 8072 12130 8084
rect 12805 8075 12863 8081
rect 12805 8072 12817 8075
rect 12124 8044 12817 8072
rect 12124 8032 12130 8044
rect 12805 8041 12817 8044
rect 12851 8041 12863 8075
rect 12805 8035 12863 8041
rect 12989 8075 13047 8081
rect 12989 8041 13001 8075
rect 13035 8072 13047 8075
rect 13906 8072 13912 8084
rect 13035 8044 13912 8072
rect 13035 8041 13047 8044
rect 12989 8035 13047 8041
rect 13906 8032 13912 8044
rect 13964 8032 13970 8084
rect 14458 8072 14464 8084
rect 14419 8044 14464 8072
rect 14458 8032 14464 8044
rect 14516 8032 14522 8084
rect 14734 8072 14740 8084
rect 14695 8044 14740 8072
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 17310 8032 17316 8084
rect 17368 8072 17374 8084
rect 17497 8075 17555 8081
rect 17497 8072 17509 8075
rect 17368 8044 17509 8072
rect 17368 8032 17374 8044
rect 17497 8041 17509 8044
rect 17543 8041 17555 8075
rect 17497 8035 17555 8041
rect 18322 8032 18328 8084
rect 18380 8072 18386 8084
rect 19150 8072 19156 8084
rect 18380 8044 19156 8072
rect 18380 8032 18386 8044
rect 19150 8032 19156 8044
rect 19208 8032 19214 8084
rect 19337 8075 19395 8081
rect 19337 8041 19349 8075
rect 19383 8072 19395 8075
rect 19426 8072 19432 8084
rect 19383 8044 19432 8072
rect 19383 8041 19395 8044
rect 19337 8035 19395 8041
rect 19426 8032 19432 8044
rect 19484 8032 19490 8084
rect 19613 8075 19671 8081
rect 19613 8041 19625 8075
rect 19659 8072 19671 8075
rect 19794 8072 19800 8084
rect 19659 8044 19800 8072
rect 19659 8041 19671 8044
rect 19613 8035 19671 8041
rect 19794 8032 19800 8044
rect 19852 8032 19858 8084
rect 22186 8072 22192 8084
rect 22147 8044 22192 8072
rect 22186 8032 22192 8044
rect 22244 8032 22250 8084
rect 7926 8004 7932 8016
rect 2516 7976 5856 8004
rect 7887 7976 7932 8004
rect 1762 7896 1768 7948
rect 1820 7936 1826 7948
rect 2516 7945 2544 7976
rect 2501 7939 2559 7945
rect 2501 7936 2513 7939
rect 1820 7908 2513 7936
rect 1820 7896 1826 7908
rect 2501 7905 2513 7908
rect 2547 7905 2559 7939
rect 3142 7936 3148 7948
rect 3103 7908 3148 7936
rect 2501 7899 2559 7905
rect 3142 7896 3148 7908
rect 3200 7896 3206 7948
rect 4338 7896 4344 7948
rect 4396 7936 4402 7948
rect 4433 7939 4491 7945
rect 4433 7936 4445 7939
rect 4396 7908 4445 7936
rect 4396 7896 4402 7908
rect 4433 7905 4445 7908
rect 4479 7905 4491 7939
rect 5721 7939 5779 7945
rect 5721 7936 5733 7939
rect 4433 7899 4491 7905
rect 4540 7908 5733 7936
rect 3786 7828 3792 7880
rect 3844 7868 3850 7880
rect 4540 7868 4568 7908
rect 5721 7905 5733 7908
rect 5767 7905 5779 7939
rect 5828 7936 5856 7976
rect 7926 7964 7932 7976
rect 7984 7964 7990 8016
rect 8021 8007 8079 8013
rect 8021 7973 8033 8007
rect 8067 8004 8079 8007
rect 8067 7976 8616 8004
rect 8067 7973 8079 7976
rect 8021 7967 8079 7973
rect 8588 7936 8616 7976
rect 8754 7964 8760 8016
rect 8812 8004 8818 8016
rect 9214 8004 9220 8016
rect 8812 7976 9220 8004
rect 8812 7964 8818 7976
rect 9214 7964 9220 7976
rect 9272 7964 9278 8016
rect 10036 8007 10094 8013
rect 10036 7973 10048 8007
rect 10082 8004 10094 8007
rect 11238 8004 11244 8016
rect 10082 7976 11244 8004
rect 10082 7973 10094 7976
rect 10036 7967 10094 7973
rect 11238 7964 11244 7976
rect 11296 7964 11302 8016
rect 11716 8004 11744 8032
rect 11716 7976 12296 8004
rect 5828 7908 8340 7936
rect 8588 7908 9628 7936
rect 5721 7899 5779 7905
rect 4982 7868 4988 7880
rect 3844 7840 4568 7868
rect 4943 7840 4988 7868
rect 3844 7828 3850 7840
rect 4982 7828 4988 7840
rect 5040 7828 5046 7880
rect 7006 7868 7012 7880
rect 6967 7840 7012 7868
rect 7006 7828 7012 7840
rect 7064 7828 7070 7880
rect 7190 7868 7196 7880
rect 7151 7840 7196 7868
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 7926 7828 7932 7880
rect 7984 7868 7990 7880
rect 8113 7871 8171 7877
rect 8113 7868 8125 7871
rect 7984 7840 8125 7868
rect 7984 7828 7990 7840
rect 8113 7837 8125 7840
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 5074 7760 5080 7812
rect 5132 7800 5138 7812
rect 7558 7800 7564 7812
rect 5132 7772 6684 7800
rect 7519 7772 7564 7800
rect 5132 7760 5138 7772
rect 5626 7692 5632 7744
rect 5684 7732 5690 7744
rect 6549 7735 6607 7741
rect 6549 7732 6561 7735
rect 5684 7704 6561 7732
rect 5684 7692 5690 7704
rect 6549 7701 6561 7704
rect 6595 7701 6607 7735
rect 6656 7732 6684 7772
rect 7558 7760 7564 7772
rect 7616 7760 7622 7812
rect 8312 7800 8340 7908
rect 9600 7880 9628 7908
rect 9674 7896 9680 7948
rect 9732 7936 9738 7948
rect 9769 7939 9827 7945
rect 9769 7936 9781 7939
rect 9732 7908 9781 7936
rect 9732 7896 9738 7908
rect 9769 7905 9781 7908
rect 9815 7905 9827 7939
rect 9769 7899 9827 7905
rect 9858 7896 9864 7948
rect 9916 7936 9922 7948
rect 11681 7939 11739 7945
rect 11681 7936 11693 7939
rect 9916 7908 11693 7936
rect 9916 7896 9922 7908
rect 11681 7905 11693 7908
rect 11727 7905 11739 7939
rect 12268 7936 12296 7976
rect 12342 7964 12348 8016
rect 12400 8004 12406 8016
rect 20622 8004 20628 8016
rect 12400 7976 20628 8004
rect 12400 7964 12406 7976
rect 20622 7964 20628 7976
rect 20680 7964 20686 8016
rect 21266 8004 21272 8016
rect 21227 7976 21272 8004
rect 21266 7964 21272 7976
rect 21324 7964 21330 8016
rect 22097 8007 22155 8013
rect 22097 7973 22109 8007
rect 22143 8004 22155 8007
rect 22554 8004 22560 8016
rect 22143 7976 22560 8004
rect 22143 7973 22155 7976
rect 22097 7967 22155 7973
rect 22554 7964 22560 7976
rect 22612 7964 22618 8016
rect 13348 7939 13406 7945
rect 13348 7936 13360 7939
rect 12268 7908 13360 7936
rect 11681 7899 11739 7905
rect 13348 7905 13360 7908
rect 13394 7936 13406 7939
rect 14918 7936 14924 7948
rect 13394 7908 14924 7936
rect 13394 7905 13406 7908
rect 13348 7899 13406 7905
rect 14918 7896 14924 7908
rect 14976 7896 14982 7948
rect 15924 7939 15982 7945
rect 15924 7905 15936 7939
rect 15970 7936 15982 7939
rect 16390 7936 16396 7948
rect 15970 7908 16396 7936
rect 15970 7905 15982 7908
rect 15924 7899 15982 7905
rect 16390 7896 16396 7908
rect 16448 7896 16454 7948
rect 16666 7896 16672 7948
rect 16724 7936 16730 7948
rect 17313 7939 17371 7945
rect 17313 7936 17325 7939
rect 16724 7908 17325 7936
rect 16724 7896 16730 7908
rect 17313 7905 17325 7908
rect 17359 7905 17371 7939
rect 17313 7899 17371 7905
rect 17586 7896 17592 7948
rect 17644 7936 17650 7948
rect 18213 7939 18271 7945
rect 18213 7936 18225 7939
rect 17644 7908 18225 7936
rect 17644 7896 17650 7908
rect 18213 7905 18225 7908
rect 18259 7905 18271 7939
rect 18213 7899 18271 7905
rect 18506 7896 18512 7948
rect 18564 7936 18570 7948
rect 19978 7936 19984 7948
rect 18564 7908 19104 7936
rect 19939 7908 19984 7936
rect 18564 7896 18570 7908
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7868 9275 7871
rect 9401 7871 9459 7877
rect 9401 7868 9413 7871
rect 9263 7840 9413 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 9401 7837 9413 7840
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 9582 7828 9588 7880
rect 9640 7828 9646 7880
rect 11422 7868 11428 7880
rect 11383 7840 11428 7868
rect 11422 7828 11428 7840
rect 11480 7828 11486 7880
rect 12618 7828 12624 7880
rect 12676 7868 12682 7880
rect 12989 7871 13047 7877
rect 12989 7868 13001 7871
rect 12676 7840 13001 7868
rect 12676 7828 12682 7840
rect 12989 7837 13001 7840
rect 13035 7837 13047 7871
rect 12989 7831 13047 7837
rect 13081 7871 13139 7877
rect 13081 7837 13093 7871
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 9122 7800 9128 7812
rect 8312 7772 9128 7800
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 9674 7800 9680 7812
rect 9223 7772 9680 7800
rect 7190 7732 7196 7744
rect 6656 7704 7196 7732
rect 6549 7695 6607 7701
rect 7190 7692 7196 7704
rect 7248 7692 7254 7744
rect 8570 7732 8576 7744
rect 8531 7704 8576 7732
rect 8570 7692 8576 7704
rect 8628 7692 8634 7744
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 9223 7732 9251 7772
rect 9674 7760 9680 7772
rect 9732 7760 9738 7812
rect 10870 7760 10876 7812
rect 10928 7800 10934 7812
rect 11149 7803 11207 7809
rect 11149 7800 11161 7803
rect 10928 7772 11161 7800
rect 10928 7760 10934 7772
rect 11149 7769 11161 7772
rect 11195 7800 11207 7803
rect 11330 7800 11336 7812
rect 11195 7772 11336 7800
rect 11195 7769 11207 7772
rect 11149 7763 11207 7769
rect 11330 7760 11336 7772
rect 11388 7760 11394 7812
rect 12526 7760 12532 7812
rect 12584 7800 12590 7812
rect 13096 7800 13124 7831
rect 14734 7828 14740 7880
rect 14792 7868 14798 7880
rect 15470 7868 15476 7880
rect 14792 7840 15476 7868
rect 14792 7828 14798 7840
rect 15470 7828 15476 7840
rect 15528 7868 15534 7880
rect 15657 7871 15715 7877
rect 15657 7868 15669 7871
rect 15528 7840 15669 7868
rect 15528 7828 15534 7840
rect 15657 7837 15669 7840
rect 15703 7837 15715 7871
rect 15657 7831 15715 7837
rect 17957 7871 18015 7877
rect 17957 7837 17969 7871
rect 18003 7837 18015 7871
rect 17957 7831 18015 7837
rect 12584 7772 13124 7800
rect 12584 7760 12590 7772
rect 8720 7704 9251 7732
rect 9401 7735 9459 7741
rect 8720 7692 8726 7704
rect 9401 7701 9413 7735
rect 9447 7732 9459 7735
rect 11790 7732 11796 7744
rect 9447 7704 11796 7732
rect 9447 7701 9459 7704
rect 9401 7695 9459 7701
rect 11790 7692 11796 7704
rect 11848 7692 11854 7744
rect 12710 7692 12716 7744
rect 12768 7732 12774 7744
rect 13722 7732 13728 7744
rect 12768 7704 13728 7732
rect 12768 7692 12774 7704
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 15654 7692 15660 7744
rect 15712 7732 15718 7744
rect 16022 7732 16028 7744
rect 15712 7704 16028 7732
rect 15712 7692 15718 7704
rect 16022 7692 16028 7704
rect 16080 7692 16086 7744
rect 16298 7692 16304 7744
rect 16356 7732 16362 7744
rect 17037 7735 17095 7741
rect 17037 7732 17049 7735
rect 16356 7704 17049 7732
rect 16356 7692 16362 7704
rect 17037 7701 17049 7704
rect 17083 7701 17095 7735
rect 17972 7732 18000 7831
rect 19076 7800 19104 7908
rect 19978 7896 19984 7908
rect 20036 7896 20042 7948
rect 20990 7936 20996 7948
rect 20951 7908 20996 7936
rect 20990 7896 20996 7908
rect 21048 7896 21054 7948
rect 22186 7936 22192 7948
rect 21744 7908 22192 7936
rect 19150 7828 19156 7880
rect 19208 7868 19214 7880
rect 20073 7871 20131 7877
rect 20073 7868 20085 7871
rect 19208 7840 20085 7868
rect 19208 7828 19214 7840
rect 20073 7837 20085 7840
rect 20119 7837 20131 7871
rect 20073 7831 20131 7837
rect 20162 7828 20168 7880
rect 20220 7868 20226 7880
rect 20220 7840 20265 7868
rect 20220 7828 20226 7840
rect 21744 7809 21772 7908
rect 22186 7896 22192 7908
rect 22244 7896 22250 7948
rect 22373 7871 22431 7877
rect 22373 7837 22385 7871
rect 22419 7868 22431 7871
rect 22646 7868 22652 7880
rect 22419 7840 22652 7868
rect 22419 7837 22431 7840
rect 22373 7831 22431 7837
rect 22646 7828 22652 7840
rect 22704 7828 22710 7880
rect 21729 7803 21787 7809
rect 21729 7800 21741 7803
rect 19076 7772 21741 7800
rect 21729 7769 21741 7772
rect 21775 7769 21787 7803
rect 21729 7763 21787 7769
rect 18322 7732 18328 7744
rect 17972 7704 18328 7732
rect 17037 7695 17095 7701
rect 18322 7692 18328 7704
rect 18380 7692 18386 7744
rect 18598 7692 18604 7744
rect 18656 7732 18662 7744
rect 23014 7732 23020 7744
rect 18656 7704 23020 7732
rect 18656 7692 18662 7704
rect 23014 7692 23020 7704
rect 23072 7692 23078 7744
rect 1104 7642 23276 7664
rect 1104 7590 4680 7642
rect 4732 7590 4744 7642
rect 4796 7590 4808 7642
rect 4860 7590 4872 7642
rect 4924 7590 12078 7642
rect 12130 7590 12142 7642
rect 12194 7590 12206 7642
rect 12258 7590 12270 7642
rect 12322 7590 19475 7642
rect 19527 7590 19539 7642
rect 19591 7590 19603 7642
rect 19655 7590 19667 7642
rect 19719 7590 23276 7642
rect 1104 7568 23276 7590
rect 4709 7531 4767 7537
rect 4709 7497 4721 7531
rect 4755 7528 4767 7531
rect 5074 7528 5080 7540
rect 4755 7500 5080 7528
rect 4755 7497 4767 7500
rect 4709 7491 4767 7497
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 5721 7531 5779 7537
rect 5721 7497 5733 7531
rect 5767 7528 5779 7531
rect 6638 7528 6644 7540
rect 5767 7500 6644 7528
rect 5767 7497 5779 7500
rect 5721 7491 5779 7497
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 7561 7531 7619 7537
rect 7561 7497 7573 7531
rect 7607 7528 7619 7531
rect 7926 7528 7932 7540
rect 7607 7500 7932 7528
rect 7607 7497 7619 7500
rect 7561 7491 7619 7497
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 8570 7488 8576 7540
rect 8628 7528 8634 7540
rect 12618 7528 12624 7540
rect 8628 7500 12624 7528
rect 8628 7488 8634 7500
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 16298 7528 16304 7540
rect 13556 7500 16304 7528
rect 3697 7463 3755 7469
rect 3697 7429 3709 7463
rect 3743 7460 3755 7463
rect 4982 7460 4988 7472
rect 3743 7432 4988 7460
rect 3743 7429 3755 7432
rect 3697 7423 3755 7429
rect 4982 7420 4988 7432
rect 5040 7420 5046 7472
rect 5626 7460 5632 7472
rect 5092 7432 5632 7460
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 5092 7392 5120 7432
rect 5626 7420 5632 7432
rect 5684 7420 5690 7472
rect 9858 7420 9864 7472
rect 9916 7460 9922 7472
rect 9953 7463 10011 7469
rect 9953 7460 9965 7463
rect 9916 7432 9965 7460
rect 9916 7420 9922 7432
rect 9953 7429 9965 7432
rect 9999 7460 10011 7463
rect 10134 7460 10140 7472
rect 9999 7432 10140 7460
rect 9999 7429 10011 7432
rect 9953 7423 10011 7429
rect 10134 7420 10140 7432
rect 10192 7420 10198 7472
rect 11422 7420 11428 7472
rect 11480 7460 11486 7472
rect 12526 7460 12532 7472
rect 11480 7432 12532 7460
rect 11480 7420 11486 7432
rect 12526 7420 12532 7432
rect 12584 7420 12590 7472
rect 4387 7364 5120 7392
rect 5353 7395 5411 7401
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 5353 7361 5365 7395
rect 5399 7392 5411 7395
rect 6273 7395 6331 7401
rect 6273 7392 6285 7395
rect 5399 7364 6285 7392
rect 5399 7361 5411 7364
rect 5353 7355 5411 7361
rect 6273 7361 6285 7364
rect 6319 7392 6331 7395
rect 6638 7392 6644 7404
rect 6319 7364 6644 7392
rect 6319 7361 6331 7364
rect 6273 7355 6331 7361
rect 6638 7352 6644 7364
rect 6696 7352 6702 7404
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7392 8263 7395
rect 8386 7392 8392 7404
rect 8251 7364 8392 7392
rect 8251 7361 8263 7364
rect 8205 7355 8263 7361
rect 8386 7352 8392 7364
rect 8444 7352 8450 7404
rect 8570 7392 8576 7404
rect 8531 7364 8576 7392
rect 8570 7352 8576 7364
rect 8628 7352 8634 7404
rect 9674 7352 9680 7404
rect 9732 7392 9738 7404
rect 10226 7392 10232 7404
rect 9732 7364 10232 7392
rect 9732 7352 9738 7364
rect 10226 7352 10232 7364
rect 10284 7352 10290 7404
rect 4157 7327 4215 7333
rect 4157 7293 4169 7327
rect 4203 7324 4215 7327
rect 6086 7324 6092 7336
rect 4203 7296 6092 7324
rect 4203 7293 4215 7296
rect 4157 7287 4215 7293
rect 6086 7284 6092 7296
rect 6144 7284 6150 7336
rect 8021 7327 8079 7333
rect 8021 7293 8033 7327
rect 8067 7324 8079 7327
rect 9858 7324 9864 7336
rect 8067 7296 9864 7324
rect 8067 7293 8079 7296
rect 8021 7287 8079 7293
rect 9858 7284 9864 7296
rect 9916 7284 9922 7336
rect 10496 7327 10554 7333
rect 10496 7293 10508 7327
rect 10542 7324 10554 7327
rect 10870 7324 10876 7336
rect 10542 7296 10876 7324
rect 10542 7293 10554 7296
rect 10496 7287 10554 7293
rect 10870 7284 10876 7296
rect 10928 7284 10934 7336
rect 12544 7324 12572 7420
rect 13173 7395 13231 7401
rect 13173 7361 13185 7395
rect 13219 7392 13231 7395
rect 13556 7392 13584 7500
rect 16298 7488 16304 7500
rect 16356 7488 16362 7540
rect 17681 7531 17739 7537
rect 17681 7497 17693 7531
rect 17727 7528 17739 7531
rect 19150 7528 19156 7540
rect 17727 7500 19156 7528
rect 17727 7497 17739 7500
rect 17681 7491 17739 7497
rect 19150 7488 19156 7500
rect 19208 7488 19214 7540
rect 19886 7488 19892 7540
rect 19944 7528 19950 7540
rect 20257 7531 20315 7537
rect 20257 7528 20269 7531
rect 19944 7500 20269 7528
rect 19944 7488 19950 7500
rect 20257 7497 20269 7500
rect 20303 7528 20315 7531
rect 20714 7528 20720 7540
rect 20303 7500 20720 7528
rect 20303 7497 20315 7500
rect 20257 7491 20315 7497
rect 20714 7488 20720 7500
rect 20772 7488 20778 7540
rect 14918 7460 14924 7472
rect 14879 7432 14924 7460
rect 14918 7420 14924 7432
rect 14976 7420 14982 7472
rect 15838 7392 15844 7404
rect 13219 7364 13584 7392
rect 15799 7364 15844 7392
rect 13219 7361 13231 7364
rect 13173 7355 13231 7361
rect 15838 7352 15844 7364
rect 15896 7352 15902 7404
rect 16114 7352 16120 7404
rect 16172 7392 16178 7404
rect 16304 7395 16362 7401
rect 16304 7392 16316 7395
rect 16172 7364 16316 7392
rect 16172 7352 16178 7364
rect 16304 7361 16316 7364
rect 16350 7361 16362 7395
rect 16758 7392 16764 7404
rect 16304 7355 16362 7361
rect 16408 7364 16764 7392
rect 13262 7324 13268 7336
rect 12544 7296 13268 7324
rect 13262 7284 13268 7296
rect 13320 7324 13326 7336
rect 13541 7327 13599 7333
rect 13541 7324 13553 7327
rect 13320 7296 13553 7324
rect 13320 7284 13326 7296
rect 13541 7293 13553 7296
rect 13587 7293 13599 7327
rect 15102 7324 15108 7336
rect 13541 7287 13599 7293
rect 13740 7296 15108 7324
rect 4246 7216 4252 7268
rect 4304 7256 4310 7268
rect 5169 7259 5227 7265
rect 5169 7256 5181 7259
rect 4304 7228 5181 7256
rect 4304 7216 4310 7228
rect 5169 7225 5181 7228
rect 5215 7225 5227 7259
rect 5169 7219 5227 7225
rect 6181 7259 6239 7265
rect 6181 7225 6193 7259
rect 6227 7256 6239 7259
rect 7558 7256 7564 7268
rect 6227 7228 7564 7256
rect 6227 7225 6239 7228
rect 6181 7219 6239 7225
rect 7558 7216 7564 7228
rect 7616 7216 7622 7268
rect 7929 7259 7987 7265
rect 7929 7225 7941 7259
rect 7975 7256 7987 7259
rect 8840 7259 8898 7265
rect 7975 7228 8708 7256
rect 7975 7225 7987 7228
rect 7929 7219 7987 7225
rect 1946 7148 1952 7200
rect 2004 7188 2010 7200
rect 2958 7188 2964 7200
rect 2004 7160 2964 7188
rect 2004 7148 2010 7160
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 4062 7188 4068 7200
rect 4023 7160 4068 7188
rect 4062 7148 4068 7160
rect 4120 7148 4126 7200
rect 5077 7191 5135 7197
rect 5077 7157 5089 7191
rect 5123 7188 5135 7191
rect 5810 7188 5816 7200
rect 5123 7160 5816 7188
rect 5123 7157 5135 7160
rect 5077 7151 5135 7157
rect 5810 7148 5816 7160
rect 5868 7148 5874 7200
rect 6089 7191 6147 7197
rect 6089 7157 6101 7191
rect 6135 7188 6147 7191
rect 7190 7188 7196 7200
rect 6135 7160 7196 7188
rect 6135 7157 6147 7160
rect 6089 7151 6147 7157
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 8680 7188 8708 7228
rect 8840 7225 8852 7259
rect 8886 7256 8898 7259
rect 12342 7256 12348 7268
rect 8886 7228 10364 7256
rect 8886 7225 8898 7228
rect 8840 7219 8898 7225
rect 9122 7188 9128 7200
rect 8680 7160 9128 7188
rect 9122 7148 9128 7160
rect 9180 7148 9186 7200
rect 10336 7188 10364 7228
rect 11440 7228 12348 7256
rect 11440 7188 11468 7228
rect 12342 7216 12348 7228
rect 12400 7216 12406 7268
rect 13740 7256 13768 7296
rect 15102 7284 15108 7296
rect 15160 7284 15166 7336
rect 15286 7324 15292 7336
rect 15247 7296 15292 7324
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 16408 7324 16436 7364
rect 16758 7352 16764 7364
rect 16816 7352 16822 7404
rect 18414 7392 18420 7404
rect 18375 7364 18420 7392
rect 18414 7352 18420 7364
rect 18472 7352 18478 7404
rect 18880 7395 18938 7401
rect 18880 7361 18892 7395
rect 18926 7361 18938 7395
rect 19150 7392 19156 7404
rect 19111 7364 19156 7392
rect 18880 7355 18938 7361
rect 15948 7296 16436 7324
rect 16577 7327 16635 7333
rect 12544 7228 13768 7256
rect 13808 7259 13866 7265
rect 11606 7188 11612 7200
rect 10336 7160 11468 7188
rect 11567 7160 11612 7188
rect 11606 7148 11612 7160
rect 11664 7148 11670 7200
rect 12544 7197 12572 7228
rect 13808 7225 13820 7259
rect 13854 7256 13866 7259
rect 14826 7256 14832 7268
rect 13854 7228 14832 7256
rect 13854 7225 13866 7228
rect 13808 7219 13866 7225
rect 14826 7216 14832 7228
rect 14884 7216 14890 7268
rect 12529 7191 12587 7197
rect 12529 7157 12541 7191
rect 12575 7157 12587 7191
rect 12529 7151 12587 7157
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 12897 7191 12955 7197
rect 12897 7188 12909 7191
rect 12676 7160 12909 7188
rect 12676 7148 12682 7160
rect 12897 7157 12909 7160
rect 12943 7157 12955 7191
rect 12897 7151 12955 7157
rect 12989 7191 13047 7197
rect 12989 7157 13001 7191
rect 13035 7188 13047 7191
rect 15286 7188 15292 7200
rect 13035 7160 15292 7188
rect 13035 7157 13047 7160
rect 12989 7151 13047 7157
rect 15286 7148 15292 7160
rect 15344 7148 15350 7200
rect 15473 7191 15531 7197
rect 15473 7157 15485 7191
rect 15519 7188 15531 7191
rect 15948 7188 15976 7296
rect 16577 7293 16589 7327
rect 16623 7324 16635 7327
rect 16850 7324 16856 7336
rect 16623 7296 16856 7324
rect 16623 7293 16635 7296
rect 16577 7287 16635 7293
rect 16850 7284 16856 7296
rect 16908 7324 16914 7336
rect 17034 7324 17040 7336
rect 16908 7296 17040 7324
rect 16908 7284 16914 7296
rect 17034 7284 17040 7296
rect 17092 7284 17098 7336
rect 18892 7324 18920 7355
rect 19150 7352 19156 7364
rect 19208 7352 19214 7404
rect 20254 7324 20260 7336
rect 18892 7296 20260 7324
rect 20254 7284 20260 7296
rect 20312 7284 20318 7336
rect 20533 7327 20591 7333
rect 20533 7293 20545 7327
rect 20579 7293 20591 7327
rect 20533 7287 20591 7293
rect 20548 7256 20576 7287
rect 20622 7284 20628 7336
rect 20680 7324 20686 7336
rect 22189 7327 22247 7333
rect 22189 7324 22201 7327
rect 20680 7296 22201 7324
rect 20680 7284 20686 7296
rect 22189 7293 22201 7296
rect 22235 7324 22247 7327
rect 22738 7324 22744 7336
rect 22235 7296 22744 7324
rect 22235 7293 22247 7296
rect 22189 7287 22247 7293
rect 22738 7284 22744 7296
rect 22796 7284 22802 7336
rect 20548 7228 20668 7256
rect 15519 7160 15976 7188
rect 16307 7191 16365 7197
rect 15519 7157 15531 7160
rect 15473 7151 15531 7157
rect 16307 7157 16319 7191
rect 16353 7188 16365 7191
rect 18690 7188 18696 7200
rect 16353 7160 18696 7188
rect 16353 7157 16365 7160
rect 16307 7151 16365 7157
rect 18690 7148 18696 7160
rect 18748 7188 18754 7200
rect 18883 7191 18941 7197
rect 18883 7188 18895 7191
rect 18748 7160 18895 7188
rect 18748 7148 18754 7160
rect 18883 7157 18895 7160
rect 18929 7157 18941 7191
rect 20640 7188 20668 7228
rect 20714 7216 20720 7268
rect 20772 7265 20778 7268
rect 20772 7259 20836 7265
rect 20772 7225 20790 7259
rect 20824 7225 20836 7259
rect 22462 7256 22468 7268
rect 22423 7228 22468 7256
rect 20772 7219 20836 7225
rect 20772 7216 20778 7219
rect 22462 7216 22468 7228
rect 22520 7216 22526 7268
rect 20990 7188 20996 7200
rect 20640 7160 20996 7188
rect 18883 7151 18941 7157
rect 20990 7148 20996 7160
rect 21048 7148 21054 7200
rect 21082 7148 21088 7200
rect 21140 7188 21146 7200
rect 21913 7191 21971 7197
rect 21913 7188 21925 7191
rect 21140 7160 21925 7188
rect 21140 7148 21146 7160
rect 21913 7157 21925 7160
rect 21959 7157 21971 7191
rect 21913 7151 21971 7157
rect 1104 7098 23276 7120
rect 1104 7046 8379 7098
rect 8431 7046 8443 7098
rect 8495 7046 8507 7098
rect 8559 7046 8571 7098
rect 8623 7046 15776 7098
rect 15828 7046 15840 7098
rect 15892 7046 15904 7098
rect 15956 7046 15968 7098
rect 16020 7046 23276 7098
rect 1104 7024 23276 7046
rect 5905 6987 5963 6993
rect 5905 6953 5917 6987
rect 5951 6984 5963 6987
rect 6178 6984 6184 6996
rect 5951 6956 6184 6984
rect 5951 6953 5963 6956
rect 5905 6947 5963 6953
rect 6178 6944 6184 6956
rect 6236 6944 6242 6996
rect 6546 6984 6552 6996
rect 6507 6956 6552 6984
rect 6546 6944 6552 6956
rect 6604 6944 6610 6996
rect 6914 6984 6920 6996
rect 6875 6956 6920 6984
rect 6914 6944 6920 6956
rect 6972 6944 6978 6996
rect 7006 6944 7012 6996
rect 7064 6984 7070 6996
rect 7558 6984 7564 6996
rect 7064 6956 7564 6984
rect 7064 6944 7070 6956
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 7926 6984 7932 6996
rect 7887 6956 7932 6984
rect 7926 6944 7932 6956
rect 7984 6944 7990 6996
rect 8021 6987 8079 6993
rect 8021 6953 8033 6987
rect 8067 6984 8079 6987
rect 8662 6984 8668 6996
rect 8067 6956 8668 6984
rect 8067 6953 8079 6956
rect 8021 6947 8079 6953
rect 8662 6944 8668 6956
rect 8720 6944 8726 6996
rect 8938 6984 8944 6996
rect 8899 6956 8944 6984
rect 8938 6944 8944 6956
rect 8996 6944 9002 6996
rect 9582 6944 9588 6996
rect 9640 6984 9646 6996
rect 11790 6984 11796 6996
rect 9640 6956 11796 6984
rect 9640 6944 9646 6956
rect 11790 6944 11796 6956
rect 11848 6944 11854 6996
rect 13262 6944 13268 6996
rect 13320 6984 13326 6996
rect 13449 6987 13507 6993
rect 13449 6984 13461 6987
rect 13320 6956 13461 6984
rect 13320 6944 13326 6956
rect 13449 6953 13461 6956
rect 13495 6953 13507 6987
rect 13449 6947 13507 6953
rect 14090 6944 14096 6996
rect 14148 6984 14154 6996
rect 14366 6984 14372 6996
rect 14148 6956 14372 6984
rect 14148 6944 14154 6956
rect 14366 6944 14372 6956
rect 14424 6944 14430 6996
rect 14826 6944 14832 6996
rect 14884 6984 14890 6996
rect 14921 6987 14979 6993
rect 14921 6984 14933 6987
rect 14884 6956 14933 6984
rect 14884 6944 14890 6956
rect 14921 6953 14933 6956
rect 14967 6953 14979 6987
rect 14921 6947 14979 6953
rect 15286 6944 15292 6996
rect 15344 6984 15350 6996
rect 19429 6987 19487 6993
rect 19429 6984 19441 6987
rect 15344 6956 19441 6984
rect 15344 6944 15350 6956
rect 19429 6953 19441 6956
rect 19475 6984 19487 6987
rect 19978 6984 19984 6996
rect 19475 6956 19984 6984
rect 19475 6953 19487 6956
rect 19429 6947 19487 6953
rect 19978 6944 19984 6956
rect 20036 6944 20042 6996
rect 20990 6984 20996 6996
rect 20916 6956 20996 6984
rect 4893 6919 4951 6925
rect 4893 6885 4905 6919
rect 4939 6916 4951 6919
rect 6822 6916 6828 6928
rect 4939 6888 6828 6916
rect 4939 6885 4951 6888
rect 4893 6879 4951 6885
rect 6822 6876 6828 6888
rect 6880 6876 6886 6928
rect 7190 6876 7196 6928
rect 7248 6916 7254 6928
rect 10410 6916 10416 6928
rect 7248 6888 10416 6916
rect 7248 6876 7254 6888
rect 10410 6876 10416 6888
rect 10468 6876 10474 6928
rect 12897 6919 12955 6925
rect 10520 6888 10824 6916
rect 4982 6848 4988 6860
rect 4943 6820 4988 6848
rect 4982 6808 4988 6820
rect 5040 6808 5046 6860
rect 7009 6851 7067 6857
rect 7009 6817 7021 6851
rect 7055 6848 7067 6851
rect 7742 6848 7748 6860
rect 7055 6820 7748 6848
rect 7055 6817 7067 6820
rect 7009 6811 7067 6817
rect 7742 6808 7748 6820
rect 7800 6808 7806 6860
rect 9861 6851 9919 6857
rect 8220 6820 9168 6848
rect 8220 6792 8248 6820
rect 5166 6780 5172 6792
rect 5127 6752 5172 6780
rect 5166 6740 5172 6752
rect 5224 6740 5230 6792
rect 5626 6740 5632 6792
rect 5684 6780 5690 6792
rect 5997 6783 6055 6789
rect 5997 6780 6009 6783
rect 5684 6752 6009 6780
rect 5684 6740 5690 6752
rect 5997 6749 6009 6752
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 6181 6783 6239 6789
rect 6181 6749 6193 6783
rect 6227 6780 6239 6783
rect 6914 6780 6920 6792
rect 6227 6752 6920 6780
rect 6227 6749 6239 6752
rect 6181 6743 6239 6749
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 7101 6783 7159 6789
rect 7101 6749 7113 6783
rect 7147 6749 7159 6783
rect 8202 6780 8208 6792
rect 8163 6752 8208 6780
rect 7101 6743 7159 6749
rect 4522 6712 4528 6724
rect 4483 6684 4528 6712
rect 4522 6672 4528 6684
rect 4580 6672 4586 6724
rect 5442 6672 5448 6724
rect 5500 6712 5506 6724
rect 5537 6715 5595 6721
rect 5537 6712 5549 6715
rect 5500 6684 5549 6712
rect 5500 6672 5506 6684
rect 5537 6681 5549 6684
rect 5583 6681 5595 6715
rect 5537 6675 5595 6681
rect 6638 6672 6644 6724
rect 6696 6712 6702 6724
rect 7116 6712 7144 6743
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 9140 6789 9168 6820
rect 9861 6817 9873 6851
rect 9907 6848 9919 6851
rect 10520 6848 10548 6888
rect 10686 6857 10692 6860
rect 10680 6848 10692 6857
rect 9907 6820 10548 6848
rect 10647 6820 10692 6848
rect 9907 6817 9919 6820
rect 9861 6811 9919 6817
rect 10680 6811 10692 6820
rect 10686 6808 10692 6811
rect 10744 6808 10750 6860
rect 10796 6848 10824 6888
rect 12897 6885 12909 6919
rect 12943 6916 12955 6919
rect 13630 6916 13636 6928
rect 12943 6888 13636 6916
rect 12943 6885 12955 6888
rect 12897 6879 12955 6885
rect 13630 6876 13636 6888
rect 13688 6876 13694 6928
rect 18874 6916 18880 6928
rect 13740 6888 14504 6916
rect 13078 6848 13084 6860
rect 10796 6820 13084 6848
rect 13078 6808 13084 6820
rect 13136 6808 13142 6860
rect 13740 6848 13768 6888
rect 13188 6820 13768 6848
rect 13808 6851 13866 6857
rect 9033 6783 9091 6789
rect 9033 6749 9045 6783
rect 9079 6749 9091 6783
rect 9033 6743 9091 6749
rect 9125 6783 9183 6789
rect 9125 6749 9137 6783
rect 9171 6749 9183 6783
rect 10134 6780 10140 6792
rect 9125 6743 9183 6749
rect 9416 6752 10140 6780
rect 7926 6712 7932 6724
rect 6696 6684 7932 6712
rect 6696 6672 6702 6684
rect 7926 6672 7932 6684
rect 7984 6672 7990 6724
rect 8570 6712 8576 6724
rect 8531 6684 8576 6712
rect 8570 6672 8576 6684
rect 8628 6672 8634 6724
rect 9048 6712 9076 6743
rect 9416 6712 9444 6752
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10226 6740 10232 6792
rect 10284 6780 10290 6792
rect 10410 6780 10416 6792
rect 10284 6752 10416 6780
rect 10284 6740 10290 6752
rect 10410 6740 10416 6752
rect 10468 6740 10474 6792
rect 13188 6789 13216 6820
rect 13808 6817 13820 6851
rect 13854 6848 13866 6851
rect 14366 6848 14372 6860
rect 13854 6820 14372 6848
rect 13854 6817 13866 6820
rect 13808 6811 13866 6817
rect 14366 6808 14372 6820
rect 14424 6808 14430 6860
rect 14476 6848 14504 6888
rect 15212 6888 16436 6916
rect 15212 6848 15240 6888
rect 16408 6860 16436 6888
rect 17972 6888 18880 6916
rect 14476 6820 15240 6848
rect 15657 6851 15715 6857
rect 15657 6817 15669 6851
rect 15703 6848 15715 6851
rect 15746 6848 15752 6860
rect 15703 6820 15752 6848
rect 15703 6817 15715 6820
rect 15657 6811 15715 6817
rect 15746 6808 15752 6820
rect 15804 6808 15810 6860
rect 15924 6851 15982 6857
rect 15924 6817 15936 6851
rect 15970 6848 15982 6851
rect 16298 6848 16304 6860
rect 15970 6820 16304 6848
rect 15970 6817 15982 6820
rect 15924 6811 15982 6817
rect 16298 6808 16304 6820
rect 16356 6808 16362 6860
rect 16390 6808 16396 6860
rect 16448 6848 16454 6860
rect 17972 6848 18000 6888
rect 18874 6876 18880 6888
rect 18932 6876 18938 6928
rect 19058 6876 19064 6928
rect 19116 6916 19122 6928
rect 19797 6919 19855 6925
rect 19797 6916 19809 6919
rect 19116 6888 19809 6916
rect 19116 6876 19122 6888
rect 19797 6885 19809 6888
rect 19843 6885 19855 6919
rect 19797 6879 19855 6885
rect 16448 6820 18000 6848
rect 18040 6851 18098 6857
rect 16448 6808 16454 6820
rect 18040 6817 18052 6851
rect 18086 6848 18098 6851
rect 18506 6848 18512 6860
rect 18086 6820 18512 6848
rect 18086 6817 18098 6820
rect 18040 6811 18098 6817
rect 18506 6808 18512 6820
rect 18564 6848 18570 6860
rect 18564 6820 20024 6848
rect 18564 6808 18570 6820
rect 12989 6783 13047 6789
rect 12989 6749 13001 6783
rect 13035 6749 13047 6783
rect 12989 6743 13047 6749
rect 13173 6783 13231 6789
rect 13173 6749 13185 6783
rect 13219 6749 13231 6783
rect 13173 6743 13231 6749
rect 13449 6783 13507 6789
rect 13449 6749 13461 6783
rect 13495 6780 13507 6783
rect 13541 6783 13599 6789
rect 13541 6780 13553 6783
rect 13495 6752 13553 6780
rect 13495 6749 13507 6752
rect 13449 6743 13507 6749
rect 13541 6749 13553 6752
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 10042 6712 10048 6724
rect 9048 6684 9444 6712
rect 10003 6684 10048 6712
rect 10042 6672 10048 6684
rect 10100 6672 10106 6724
rect 13004 6712 13032 6743
rect 16666 6740 16672 6792
rect 16724 6780 16730 6792
rect 17129 6783 17187 6789
rect 17129 6780 17141 6783
rect 16724 6752 17141 6780
rect 16724 6740 16730 6752
rect 17129 6749 17141 6752
rect 17175 6749 17187 6783
rect 17310 6780 17316 6792
rect 17271 6752 17316 6780
rect 17129 6743 17187 6749
rect 17310 6740 17316 6752
rect 17368 6740 17374 6792
rect 17681 6783 17739 6789
rect 17681 6749 17693 6783
rect 17727 6780 17739 6783
rect 17773 6783 17831 6789
rect 17773 6780 17785 6783
rect 17727 6752 17785 6780
rect 17727 6749 17739 6752
rect 17681 6743 17739 6749
rect 17773 6749 17785 6752
rect 17819 6749 17831 6783
rect 17773 6743 17831 6749
rect 18782 6740 18788 6792
rect 18840 6780 18846 6792
rect 19996 6789 20024 6820
rect 20438 6808 20444 6860
rect 20496 6848 20502 6860
rect 20625 6851 20683 6857
rect 20625 6848 20637 6851
rect 20496 6820 20637 6848
rect 20496 6808 20502 6820
rect 20625 6817 20637 6820
rect 20671 6817 20683 6851
rect 20625 6811 20683 6817
rect 20916 6789 20944 6956
rect 20990 6944 20996 6956
rect 21048 6944 21054 6996
rect 21082 6876 21088 6928
rect 21140 6925 21146 6928
rect 21140 6919 21204 6925
rect 21140 6885 21158 6919
rect 21192 6885 21204 6919
rect 21140 6879 21204 6885
rect 21140 6876 21146 6879
rect 20990 6808 20996 6860
rect 21048 6848 21054 6860
rect 21048 6820 22232 6848
rect 21048 6808 21054 6820
rect 19889 6783 19947 6789
rect 19889 6780 19901 6783
rect 18840 6752 19901 6780
rect 18840 6740 18846 6752
rect 19889 6749 19901 6752
rect 19935 6749 19947 6783
rect 19889 6743 19947 6749
rect 19981 6783 20039 6789
rect 19981 6749 19993 6783
rect 20027 6749 20039 6783
rect 19981 6743 20039 6749
rect 20349 6783 20407 6789
rect 20349 6749 20361 6783
rect 20395 6780 20407 6783
rect 20901 6783 20959 6789
rect 20901 6780 20913 6783
rect 20395 6752 20913 6780
rect 20395 6749 20407 6752
rect 20349 6743 20407 6749
rect 20901 6749 20913 6752
rect 20947 6749 20959 6783
rect 20901 6743 20959 6749
rect 13262 6712 13268 6724
rect 13004 6684 13268 6712
rect 13262 6672 13268 6684
rect 13320 6672 13326 6724
rect 14642 6672 14648 6724
rect 14700 6712 14706 6724
rect 14918 6712 14924 6724
rect 14700 6684 14924 6712
rect 14700 6672 14706 6684
rect 14918 6672 14924 6684
rect 14976 6672 14982 6724
rect 16960 6684 17816 6712
rect 6362 6604 6368 6656
rect 6420 6644 6426 6656
rect 7006 6644 7012 6656
rect 6420 6616 7012 6644
rect 6420 6604 6426 6616
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 7561 6647 7619 6653
rect 7561 6613 7573 6647
rect 7607 6644 7619 6647
rect 9950 6644 9956 6656
rect 7607 6616 9956 6644
rect 7607 6613 7619 6616
rect 7561 6607 7619 6613
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 10686 6604 10692 6656
rect 10744 6644 10750 6656
rect 11606 6644 11612 6656
rect 10744 6616 11612 6644
rect 10744 6604 10750 6616
rect 11606 6604 11612 6616
rect 11664 6604 11670 6656
rect 11790 6644 11796 6656
rect 11751 6616 11796 6644
rect 11790 6604 11796 6616
rect 11848 6604 11854 6656
rect 12529 6647 12587 6653
rect 12529 6613 12541 6647
rect 12575 6644 12587 6647
rect 16960 6644 16988 6684
rect 12575 6616 16988 6644
rect 12575 6613 12587 6616
rect 12529 6607 12587 6613
rect 17034 6604 17040 6656
rect 17092 6644 17098 6656
rect 17092 6616 17137 6644
rect 17092 6604 17098 6616
rect 17218 6604 17224 6656
rect 17276 6644 17282 6656
rect 17681 6647 17739 6653
rect 17681 6644 17693 6647
rect 17276 6616 17693 6644
rect 17276 6604 17282 6616
rect 17681 6613 17693 6616
rect 17727 6613 17739 6647
rect 17788 6644 17816 6684
rect 18874 6672 18880 6724
rect 18932 6712 18938 6724
rect 18932 6684 19104 6712
rect 18932 6672 18938 6684
rect 18690 6644 18696 6656
rect 17788 6616 18696 6644
rect 17681 6607 17739 6613
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 19076 6644 19104 6684
rect 19150 6672 19156 6724
rect 19208 6712 19214 6724
rect 20162 6712 20168 6724
rect 19208 6684 20168 6712
rect 19208 6672 19214 6684
rect 20162 6672 20168 6684
rect 20220 6672 20226 6724
rect 22204 6712 22232 6820
rect 22278 6808 22284 6860
rect 22336 6848 22342 6860
rect 22557 6851 22615 6857
rect 22557 6848 22569 6851
rect 22336 6820 22569 6848
rect 22336 6808 22342 6820
rect 22557 6817 22569 6820
rect 22603 6817 22615 6851
rect 22557 6811 22615 6817
rect 22922 6712 22928 6724
rect 20272 6684 20576 6712
rect 22204 6684 22928 6712
rect 20272 6644 20300 6684
rect 19076 6616 20300 6644
rect 20349 6647 20407 6653
rect 20349 6613 20361 6647
rect 20395 6644 20407 6647
rect 20438 6644 20444 6656
rect 20395 6616 20444 6644
rect 20395 6613 20407 6616
rect 20349 6607 20407 6613
rect 20438 6604 20444 6616
rect 20496 6604 20502 6656
rect 20548 6644 20576 6684
rect 22922 6672 22928 6684
rect 22980 6672 22986 6724
rect 22281 6647 22339 6653
rect 22281 6644 22293 6647
rect 20548 6616 22293 6644
rect 22281 6613 22293 6616
rect 22327 6613 22339 6647
rect 22281 6607 22339 6613
rect 1104 6554 23276 6576
rect 1104 6502 4680 6554
rect 4732 6502 4744 6554
rect 4796 6502 4808 6554
rect 4860 6502 4872 6554
rect 4924 6502 12078 6554
rect 12130 6502 12142 6554
rect 12194 6502 12206 6554
rect 12258 6502 12270 6554
rect 12322 6502 19475 6554
rect 19527 6502 19539 6554
rect 19591 6502 19603 6554
rect 19655 6502 19667 6554
rect 19719 6502 23276 6554
rect 1104 6480 23276 6502
rect 5626 6440 5632 6452
rect 5587 6412 5632 6440
rect 5626 6400 5632 6412
rect 5684 6400 5690 6452
rect 7653 6443 7711 6449
rect 7653 6409 7665 6443
rect 7699 6440 7711 6443
rect 8018 6440 8024 6452
rect 7699 6412 8024 6440
rect 7699 6409 7711 6412
rect 7653 6403 7711 6409
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 9677 6443 9735 6449
rect 8128 6412 9352 6440
rect 7926 6332 7932 6384
rect 7984 6372 7990 6384
rect 8128 6372 8156 6412
rect 8662 6372 8668 6384
rect 7984 6344 8156 6372
rect 8623 6344 8668 6372
rect 7984 6332 7990 6344
rect 8662 6332 8668 6344
rect 8720 6332 8726 6384
rect 9324 6372 9352 6412
rect 9677 6409 9689 6443
rect 9723 6440 9735 6443
rect 12434 6440 12440 6452
rect 9723 6412 12440 6440
rect 9723 6409 9735 6412
rect 9677 6403 9735 6409
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 21085 6443 21143 6449
rect 21085 6440 21097 6443
rect 12544 6412 21097 6440
rect 10134 6372 10140 6384
rect 9324 6344 10140 6372
rect 10134 6332 10140 6344
rect 10192 6332 10198 6384
rect 4062 6264 4068 6316
rect 4120 6304 4126 6316
rect 6089 6307 6147 6313
rect 6089 6304 6101 6307
rect 4120 6276 6101 6304
rect 4120 6264 4126 6276
rect 6089 6273 6101 6276
rect 6135 6273 6147 6307
rect 6089 6267 6147 6273
rect 6273 6307 6331 6313
rect 6273 6273 6285 6307
rect 6319 6304 6331 6307
rect 7282 6304 7288 6316
rect 6319 6276 7288 6304
rect 6319 6273 6331 6276
rect 6273 6267 6331 6273
rect 7282 6264 7288 6276
rect 7340 6264 7346 6316
rect 7742 6264 7748 6316
rect 7800 6304 7806 6316
rect 7944 6304 7972 6332
rect 8205 6307 8263 6313
rect 8205 6304 8217 6307
rect 7800 6276 8217 6304
rect 7800 6264 7806 6276
rect 8205 6273 8217 6276
rect 8251 6273 8263 6307
rect 8205 6267 8263 6273
rect 8294 6264 8300 6316
rect 8352 6304 8358 6316
rect 9125 6307 9183 6313
rect 9125 6304 9137 6307
rect 8352 6276 9137 6304
rect 8352 6264 8358 6276
rect 9125 6273 9137 6276
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 9309 6307 9367 6313
rect 9309 6273 9321 6307
rect 9355 6304 9367 6307
rect 9674 6304 9680 6316
rect 9355 6276 9680 6304
rect 9355 6273 9367 6276
rect 9309 6267 9367 6273
rect 9674 6264 9680 6276
rect 9732 6264 9738 6316
rect 10318 6304 10324 6316
rect 10279 6276 10324 6304
rect 10318 6264 10324 6276
rect 10376 6264 10382 6316
rect 5994 6236 6000 6248
rect 5955 6208 6000 6236
rect 5994 6196 6000 6208
rect 6052 6196 6058 6248
rect 8021 6239 8079 6245
rect 8021 6205 8033 6239
rect 8067 6236 8079 6239
rect 8386 6236 8392 6248
rect 8067 6208 8392 6236
rect 8067 6205 8079 6208
rect 8021 6199 8079 6205
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 9033 6239 9091 6245
rect 9033 6205 9045 6239
rect 9079 6236 9091 6239
rect 9398 6236 9404 6248
rect 9079 6208 9404 6236
rect 9079 6205 9091 6208
rect 9033 6199 9091 6205
rect 9398 6196 9404 6208
rect 9456 6196 9462 6248
rect 10410 6196 10416 6248
rect 10468 6236 10474 6248
rect 10686 6236 10692 6248
rect 10468 6208 10692 6236
rect 10468 6196 10474 6208
rect 10686 6196 10692 6208
rect 10744 6196 10750 6248
rect 11330 6236 11336 6248
rect 10888 6208 11336 6236
rect 8113 6171 8171 6177
rect 8113 6137 8125 6171
rect 8159 6168 8171 6171
rect 9306 6168 9312 6180
rect 8159 6140 9312 6168
rect 8159 6137 8171 6140
rect 8113 6131 8171 6137
rect 9306 6128 9312 6140
rect 9364 6128 9370 6180
rect 10045 6171 10103 6177
rect 10045 6137 10057 6171
rect 10091 6168 10103 6171
rect 10888 6168 10916 6208
rect 11330 6196 11336 6208
rect 11388 6196 11394 6248
rect 12544 6245 12572 6412
rect 21085 6409 21097 6412
rect 21131 6409 21143 6443
rect 21085 6403 21143 6409
rect 14645 6375 14703 6381
rect 14645 6372 14657 6375
rect 14108 6344 14657 6372
rect 12618 6264 12624 6316
rect 12676 6304 12682 6316
rect 13078 6304 13084 6316
rect 12676 6276 13084 6304
rect 12676 6264 12682 6276
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 12529 6239 12587 6245
rect 12529 6205 12541 6239
rect 12575 6205 12587 6239
rect 13096 6236 13124 6264
rect 14108 6236 14136 6344
rect 14645 6341 14657 6344
rect 14691 6341 14703 6375
rect 14645 6335 14703 6341
rect 15746 6332 15752 6384
rect 15804 6372 15810 6384
rect 16574 6372 16580 6384
rect 15804 6344 16580 6372
rect 15804 6332 15810 6344
rect 16574 6332 16580 6344
rect 16632 6332 16638 6384
rect 16758 6332 16764 6384
rect 16816 6372 16822 6384
rect 20165 6375 20223 6381
rect 20165 6372 20177 6375
rect 16816 6344 18828 6372
rect 16816 6332 16822 6344
rect 16666 6304 16672 6316
rect 13096 6208 14136 6236
rect 14200 6276 14872 6304
rect 12529 6199 12587 6205
rect 10091 6140 10916 6168
rect 10956 6171 11014 6177
rect 10091 6137 10103 6140
rect 10045 6131 10103 6137
rect 10956 6137 10968 6171
rect 11002 6168 11014 6171
rect 11514 6168 11520 6180
rect 11002 6140 11520 6168
rect 11002 6137 11014 6140
rect 10956 6131 11014 6137
rect 11514 6128 11520 6140
rect 11572 6168 11578 6180
rect 11790 6168 11796 6180
rect 11572 6140 11796 6168
rect 11572 6128 11578 6140
rect 11790 6128 11796 6140
rect 11848 6128 11854 6180
rect 13348 6171 13406 6177
rect 13348 6137 13360 6171
rect 13394 6168 13406 6171
rect 13630 6168 13636 6180
rect 13394 6140 13636 6168
rect 13394 6137 13406 6140
rect 13348 6131 13406 6137
rect 13630 6128 13636 6140
rect 13688 6128 13694 6180
rect 10137 6103 10195 6109
rect 10137 6069 10149 6103
rect 10183 6100 10195 6103
rect 11146 6100 11152 6112
rect 10183 6072 11152 6100
rect 10183 6069 10195 6072
rect 10137 6063 10195 6069
rect 11146 6060 11152 6072
rect 11204 6060 11210 6112
rect 12069 6103 12127 6109
rect 12069 6069 12081 6103
rect 12115 6100 12127 6103
rect 12434 6100 12440 6112
rect 12115 6072 12440 6100
rect 12115 6069 12127 6072
rect 12069 6063 12127 6069
rect 12434 6060 12440 6072
rect 12492 6060 12498 6112
rect 12713 6103 12771 6109
rect 12713 6069 12725 6103
rect 12759 6100 12771 6103
rect 14200 6100 14228 6276
rect 14645 6239 14703 6245
rect 14645 6205 14657 6239
rect 14691 6236 14703 6239
rect 14734 6236 14740 6248
rect 14691 6208 14740 6236
rect 14691 6205 14703 6208
rect 14645 6199 14703 6205
rect 14734 6196 14740 6208
rect 14792 6196 14798 6248
rect 14844 6236 14872 6276
rect 16316 6276 16672 6304
rect 16316 6236 16344 6276
rect 16666 6264 16672 6276
rect 16724 6264 16730 6316
rect 16942 6264 16948 6316
rect 17000 6304 17006 6316
rect 17405 6307 17463 6313
rect 17405 6304 17417 6307
rect 17000 6276 17417 6304
rect 17000 6264 17006 6276
rect 17405 6273 17417 6276
rect 17451 6273 17463 6307
rect 17586 6304 17592 6316
rect 17547 6276 17592 6304
rect 17405 6267 17463 6273
rect 17586 6264 17592 6276
rect 17644 6264 17650 6316
rect 18800 6304 18828 6344
rect 19812 6344 20177 6372
rect 18800 6276 18920 6304
rect 14844 6208 16344 6236
rect 16393 6239 16451 6245
rect 16393 6205 16405 6239
rect 16439 6236 16451 6239
rect 16850 6236 16856 6248
rect 16439 6208 16856 6236
rect 16439 6205 16451 6208
rect 16393 6199 16451 6205
rect 16850 6196 16856 6208
rect 16908 6196 16914 6248
rect 17313 6239 17371 6245
rect 17313 6205 17325 6239
rect 17359 6236 17371 6239
rect 17678 6236 17684 6248
rect 17359 6208 17684 6236
rect 17359 6205 17371 6208
rect 17313 6199 17371 6205
rect 17678 6196 17684 6208
rect 17736 6196 17742 6248
rect 18230 6236 18236 6248
rect 18191 6208 18236 6236
rect 18230 6196 18236 6208
rect 18288 6196 18294 6248
rect 18322 6196 18328 6248
rect 18380 6236 18386 6248
rect 18785 6239 18843 6245
rect 18785 6236 18797 6239
rect 18380 6208 18797 6236
rect 18380 6196 18386 6208
rect 18785 6205 18797 6208
rect 18831 6205 18843 6239
rect 18892 6236 18920 6276
rect 19812 6236 19840 6344
rect 20165 6341 20177 6344
rect 20211 6372 20223 6375
rect 20714 6372 20720 6384
rect 20211 6344 20720 6372
rect 20211 6341 20223 6344
rect 20165 6335 20223 6341
rect 20714 6332 20720 6344
rect 20772 6332 20778 6384
rect 20438 6264 20444 6316
rect 20496 6304 20502 6316
rect 20496 6276 21220 6304
rect 20496 6264 20502 6276
rect 21192 6248 21220 6276
rect 18892 6208 19840 6236
rect 20717 6239 20775 6245
rect 18785 6199 18843 6205
rect 20717 6205 20729 6239
rect 20763 6236 20775 6239
rect 20806 6236 20812 6248
rect 20763 6208 20812 6236
rect 20763 6205 20775 6208
rect 20717 6199 20775 6205
rect 20806 6196 20812 6208
rect 20864 6196 20870 6248
rect 21174 6196 21180 6248
rect 21232 6236 21238 6248
rect 21361 6239 21419 6245
rect 21361 6236 21373 6239
rect 21232 6208 21373 6236
rect 21232 6196 21238 6208
rect 21361 6205 21373 6208
rect 21407 6205 21419 6239
rect 21361 6199 21419 6205
rect 14982 6171 15040 6177
rect 14982 6168 14994 6171
rect 14476 6140 14994 6168
rect 12759 6072 14228 6100
rect 12759 6069 12771 6072
rect 12713 6063 12771 6069
rect 14274 6060 14280 6112
rect 14332 6100 14338 6112
rect 14476 6109 14504 6140
rect 14982 6137 14994 6140
rect 15028 6137 15040 6171
rect 14982 6131 15040 6137
rect 15286 6128 15292 6180
rect 15344 6168 15350 6180
rect 15746 6168 15752 6180
rect 15344 6140 15752 6168
rect 15344 6128 15350 6140
rect 15746 6128 15752 6140
rect 15804 6128 15810 6180
rect 18138 6168 18144 6180
rect 16592 6140 18144 6168
rect 14461 6103 14519 6109
rect 14461 6100 14473 6103
rect 14332 6072 14473 6100
rect 14332 6060 14338 6072
rect 14461 6069 14473 6072
rect 14507 6069 14519 6103
rect 14461 6063 14519 6069
rect 14550 6060 14556 6112
rect 14608 6100 14614 6112
rect 16592 6109 16620 6140
rect 18138 6128 18144 6140
rect 18196 6128 18202 6180
rect 19052 6171 19110 6177
rect 19052 6137 19064 6171
rect 19098 6168 19110 6171
rect 19150 6168 19156 6180
rect 19098 6140 19156 6168
rect 19098 6137 19110 6140
rect 19052 6131 19110 6137
rect 19150 6128 19156 6140
rect 19208 6128 19214 6180
rect 20901 6171 20959 6177
rect 19260 6140 19932 6168
rect 16117 6103 16175 6109
rect 16117 6100 16129 6103
rect 14608 6072 16129 6100
rect 14608 6060 14614 6072
rect 16117 6069 16129 6072
rect 16163 6069 16175 6103
rect 16117 6063 16175 6069
rect 16577 6103 16635 6109
rect 16577 6069 16589 6103
rect 16623 6069 16635 6103
rect 16577 6063 16635 6069
rect 16945 6103 17003 6109
rect 16945 6069 16957 6103
rect 16991 6100 17003 6103
rect 17862 6100 17868 6112
rect 16991 6072 17868 6100
rect 16991 6069 17003 6072
rect 16945 6063 17003 6069
rect 17862 6060 17868 6072
rect 17920 6060 17926 6112
rect 18417 6103 18475 6109
rect 18417 6069 18429 6103
rect 18463 6100 18475 6103
rect 18598 6100 18604 6112
rect 18463 6072 18604 6100
rect 18463 6069 18475 6072
rect 18417 6063 18475 6069
rect 18598 6060 18604 6072
rect 18656 6060 18662 6112
rect 18690 6060 18696 6112
rect 18748 6100 18754 6112
rect 19260 6100 19288 6140
rect 18748 6072 19288 6100
rect 18748 6060 18754 6072
rect 19334 6060 19340 6112
rect 19392 6100 19398 6112
rect 19794 6100 19800 6112
rect 19392 6072 19800 6100
rect 19392 6060 19398 6072
rect 19794 6060 19800 6072
rect 19852 6060 19858 6112
rect 19904 6100 19932 6140
rect 20901 6137 20913 6171
rect 20947 6168 20959 6171
rect 21628 6171 21686 6177
rect 21628 6168 21640 6171
rect 20947 6140 21640 6168
rect 20947 6137 20959 6140
rect 20901 6131 20959 6137
rect 21628 6137 21640 6140
rect 21674 6168 21686 6171
rect 21818 6168 21824 6180
rect 21674 6140 21824 6168
rect 21674 6137 21686 6140
rect 21628 6131 21686 6137
rect 21818 6128 21824 6140
rect 21876 6128 21882 6180
rect 22646 6100 22652 6112
rect 19904 6072 22652 6100
rect 22646 6060 22652 6072
rect 22704 6060 22710 6112
rect 22738 6060 22744 6112
rect 22796 6100 22802 6112
rect 22796 6072 22841 6100
rect 22796 6060 22802 6072
rect 1104 6010 23276 6032
rect 1104 5958 8379 6010
rect 8431 5958 8443 6010
rect 8495 5958 8507 6010
rect 8559 5958 8571 6010
rect 8623 5958 15776 6010
rect 15828 5958 15840 6010
rect 15892 5958 15904 6010
rect 15956 5958 15968 6010
rect 16020 5958 23276 6010
rect 1104 5936 23276 5958
rect 4154 5856 4160 5908
rect 4212 5896 4218 5908
rect 5537 5899 5595 5905
rect 5537 5896 5549 5899
rect 4212 5868 5549 5896
rect 4212 5856 4218 5868
rect 5537 5865 5549 5868
rect 5583 5865 5595 5899
rect 6546 5896 6552 5908
rect 6507 5868 6552 5896
rect 5537 5859 5595 5865
rect 6546 5856 6552 5868
rect 6604 5856 6610 5908
rect 7006 5896 7012 5908
rect 6967 5868 7012 5896
rect 7006 5856 7012 5868
rect 7064 5856 7070 5908
rect 7561 5899 7619 5905
rect 7561 5865 7573 5899
rect 7607 5896 7619 5899
rect 7650 5896 7656 5908
rect 7607 5868 7656 5896
rect 7607 5865 7619 5868
rect 7561 5859 7619 5865
rect 7650 5856 7656 5868
rect 7708 5856 7714 5908
rect 7834 5856 7840 5908
rect 7892 5896 7898 5908
rect 7929 5899 7987 5905
rect 7929 5896 7941 5899
rect 7892 5868 7941 5896
rect 7892 5856 7898 5868
rect 7929 5865 7941 5868
rect 7975 5865 7987 5899
rect 7929 5859 7987 5865
rect 9033 5899 9091 5905
rect 9033 5865 9045 5899
rect 9079 5896 9091 5899
rect 9398 5896 9404 5908
rect 9079 5868 9404 5896
rect 9079 5865 9091 5868
rect 9033 5859 9091 5865
rect 9398 5856 9404 5868
rect 9456 5856 9462 5908
rect 11977 5899 12035 5905
rect 11977 5865 11989 5899
rect 12023 5865 12035 5899
rect 13630 5896 13636 5908
rect 13591 5868 13636 5896
rect 11977 5859 12035 5865
rect 4430 5788 4436 5840
rect 4488 5828 4494 5840
rect 5905 5831 5963 5837
rect 5905 5828 5917 5831
rect 4488 5800 5917 5828
rect 4488 5788 4494 5800
rect 5905 5797 5917 5800
rect 5951 5797 5963 5831
rect 5905 5791 5963 5797
rect 5997 5831 6055 5837
rect 5997 5797 6009 5831
rect 6043 5828 6055 5831
rect 6454 5828 6460 5840
rect 6043 5800 6460 5828
rect 6043 5797 6055 5800
rect 5997 5791 6055 5797
rect 6454 5788 6460 5800
rect 6512 5788 6518 5840
rect 7466 5788 7472 5840
rect 7524 5828 7530 5840
rect 8021 5831 8079 5837
rect 8021 5828 8033 5831
rect 7524 5800 8033 5828
rect 7524 5788 7530 5800
rect 8021 5797 8033 5800
rect 8067 5797 8079 5831
rect 8021 5791 8079 5797
rect 8941 5831 8999 5837
rect 8941 5797 8953 5831
rect 8987 5828 8999 5831
rect 9306 5828 9312 5840
rect 8987 5800 9312 5828
rect 8987 5797 8999 5800
rect 8941 5791 8999 5797
rect 9306 5788 9312 5800
rect 9364 5788 9370 5840
rect 11992 5828 12020 5859
rect 13630 5856 13636 5868
rect 13688 5856 13694 5908
rect 14274 5896 14280 5908
rect 14235 5868 14280 5896
rect 14274 5856 14280 5868
rect 14332 5856 14338 5908
rect 14734 5856 14740 5908
rect 14792 5896 14798 5908
rect 14921 5899 14979 5905
rect 14921 5896 14933 5899
rect 14792 5868 14933 5896
rect 14792 5856 14798 5868
rect 14921 5865 14933 5868
rect 14967 5865 14979 5899
rect 14921 5859 14979 5865
rect 15749 5899 15807 5905
rect 15749 5865 15761 5899
rect 15795 5896 15807 5899
rect 18506 5896 18512 5908
rect 15795 5868 18000 5896
rect 18467 5868 18512 5896
rect 15795 5865 15807 5868
rect 15749 5859 15807 5865
rect 12520 5831 12578 5837
rect 12520 5828 12532 5831
rect 11992 5800 12532 5828
rect 12520 5797 12532 5800
rect 12566 5828 12578 5831
rect 12802 5828 12808 5840
rect 12566 5800 12808 5828
rect 12566 5797 12578 5800
rect 12520 5791 12578 5797
rect 12802 5788 12808 5800
rect 12860 5788 12866 5840
rect 13648 5828 13676 5856
rect 14369 5831 14427 5837
rect 14369 5828 14381 5831
rect 13648 5800 14381 5828
rect 14369 5797 14381 5800
rect 14415 5797 14427 5831
rect 14369 5791 14427 5797
rect 16485 5831 16543 5837
rect 16485 5797 16497 5831
rect 16531 5828 16543 5831
rect 17862 5828 17868 5840
rect 16531 5800 17868 5828
rect 16531 5797 16543 5800
rect 16485 5791 16543 5797
rect 17862 5788 17868 5800
rect 17920 5788 17926 5840
rect 17972 5828 18000 5868
rect 18506 5856 18512 5868
rect 18564 5856 18570 5908
rect 18598 5856 18604 5908
rect 18656 5896 18662 5908
rect 19153 5899 19211 5905
rect 19153 5896 19165 5899
rect 18656 5868 19165 5896
rect 18656 5856 18662 5868
rect 19153 5865 19165 5868
rect 19199 5865 19211 5899
rect 19153 5859 19211 5865
rect 20257 5899 20315 5905
rect 20257 5865 20269 5899
rect 20303 5896 20315 5899
rect 22649 5899 22707 5905
rect 22649 5896 22661 5899
rect 20303 5868 22661 5896
rect 20303 5865 20315 5868
rect 20257 5859 20315 5865
rect 22649 5865 22661 5868
rect 22695 5865 22707 5899
rect 22649 5859 22707 5865
rect 20165 5831 20223 5837
rect 20165 5828 20177 5831
rect 17972 5800 20177 5828
rect 20165 5797 20177 5800
rect 20211 5797 20223 5831
rect 20165 5791 20223 5797
rect 20714 5788 20720 5840
rect 20772 5828 20778 5840
rect 20772 5800 22508 5828
rect 20772 5788 20778 5800
rect 6917 5763 6975 5769
rect 6917 5729 6929 5763
rect 6963 5760 6975 5763
rect 9030 5760 9036 5772
rect 6963 5732 9036 5760
rect 6963 5729 6975 5732
rect 6917 5723 6975 5729
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 10597 5763 10655 5769
rect 10597 5729 10609 5763
rect 10643 5760 10655 5763
rect 10686 5760 10692 5772
rect 10643 5732 10692 5760
rect 10643 5729 10655 5732
rect 10597 5723 10655 5729
rect 10686 5720 10692 5732
rect 10744 5720 10750 5772
rect 10864 5763 10922 5769
rect 10864 5729 10876 5763
rect 10910 5760 10922 5763
rect 12342 5760 12348 5772
rect 10910 5732 12348 5760
rect 10910 5729 10922 5732
rect 10864 5723 10922 5729
rect 12342 5720 12348 5732
rect 12400 5720 12406 5772
rect 12894 5720 12900 5772
rect 12952 5760 12958 5772
rect 12952 5732 13952 5760
rect 12952 5720 12958 5732
rect 5902 5652 5908 5704
rect 5960 5692 5966 5704
rect 6089 5695 6147 5701
rect 6089 5692 6101 5695
rect 5960 5664 6101 5692
rect 5960 5652 5966 5664
rect 6089 5661 6101 5664
rect 6135 5661 6147 5695
rect 6089 5655 6147 5661
rect 6270 5652 6276 5704
rect 6328 5692 6334 5704
rect 7101 5695 7159 5701
rect 7101 5692 7113 5695
rect 6328 5664 7113 5692
rect 6328 5652 6334 5664
rect 7101 5661 7113 5664
rect 7147 5661 7159 5695
rect 7101 5655 7159 5661
rect 7742 5652 7748 5704
rect 7800 5692 7806 5704
rect 8205 5695 8263 5701
rect 8205 5692 8217 5695
rect 7800 5664 8217 5692
rect 7800 5652 7806 5664
rect 8205 5661 8217 5664
rect 8251 5661 8263 5695
rect 8205 5655 8263 5661
rect 8846 5652 8852 5704
rect 8904 5692 8910 5704
rect 9217 5695 9275 5701
rect 9217 5692 9229 5695
rect 8904 5664 9229 5692
rect 8904 5652 8910 5664
rect 9217 5661 9229 5664
rect 9263 5692 9275 5695
rect 9398 5692 9404 5704
rect 9263 5664 9404 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 9398 5652 9404 5664
rect 9456 5652 9462 5704
rect 12250 5692 12256 5704
rect 12211 5664 12256 5692
rect 12250 5652 12256 5664
rect 12308 5652 12314 5704
rect 13924 5692 13952 5732
rect 13998 5720 14004 5772
rect 14056 5760 14062 5772
rect 15105 5763 15163 5769
rect 15105 5760 15117 5763
rect 14056 5732 15117 5760
rect 14056 5720 14062 5732
rect 15105 5729 15117 5732
rect 15151 5729 15163 5763
rect 15105 5723 15163 5729
rect 15565 5763 15623 5769
rect 15565 5729 15577 5763
rect 15611 5760 15623 5763
rect 17034 5760 17040 5772
rect 15611 5732 17040 5760
rect 15611 5729 15623 5732
rect 15565 5723 15623 5729
rect 17034 5720 17040 5732
rect 17092 5720 17098 5772
rect 17129 5763 17187 5769
rect 17129 5729 17141 5763
rect 17175 5760 17187 5763
rect 17218 5760 17224 5772
rect 17175 5732 17224 5760
rect 17175 5729 17187 5732
rect 17129 5723 17187 5729
rect 17218 5720 17224 5732
rect 17276 5720 17282 5772
rect 17396 5763 17454 5769
rect 17396 5729 17408 5763
rect 17442 5760 17454 5763
rect 19245 5763 19303 5769
rect 17442 5732 19196 5760
rect 17442 5729 17454 5732
rect 17396 5723 17454 5729
rect 14366 5692 14372 5704
rect 13924 5664 14372 5692
rect 14366 5652 14372 5664
rect 14424 5652 14430 5704
rect 14458 5652 14464 5704
rect 14516 5692 14522 5704
rect 14553 5695 14611 5701
rect 14553 5692 14565 5695
rect 14516 5664 14565 5692
rect 14516 5652 14522 5664
rect 14553 5661 14565 5664
rect 14599 5692 14611 5695
rect 14918 5692 14924 5704
rect 14599 5664 14924 5692
rect 14599 5661 14611 5664
rect 14553 5655 14611 5661
rect 14918 5652 14924 5664
rect 14976 5652 14982 5704
rect 16577 5695 16635 5701
rect 16577 5661 16589 5695
rect 16623 5661 16635 5695
rect 16758 5692 16764 5704
rect 16719 5664 16764 5692
rect 16577 5655 16635 5661
rect 8573 5627 8631 5633
rect 8573 5593 8585 5627
rect 8619 5624 8631 5627
rect 9582 5624 9588 5636
rect 8619 5596 9588 5624
rect 8619 5593 8631 5596
rect 8573 5587 8631 5593
rect 9582 5584 9588 5596
rect 9640 5584 9646 5636
rect 13262 5584 13268 5636
rect 13320 5624 13326 5636
rect 16022 5624 16028 5636
rect 13320 5596 16028 5624
rect 13320 5584 13326 5596
rect 16022 5584 16028 5596
rect 16080 5584 16086 5636
rect 16592 5624 16620 5655
rect 16758 5652 16764 5664
rect 16816 5652 16822 5704
rect 19168 5692 19196 5732
rect 19245 5729 19257 5763
rect 19291 5760 19303 5763
rect 20070 5760 20076 5772
rect 19291 5732 20076 5760
rect 19291 5729 19303 5732
rect 19245 5723 19303 5729
rect 20070 5720 20076 5732
rect 20128 5720 20134 5772
rect 20901 5763 20959 5769
rect 20901 5760 20913 5763
rect 20180 5732 20913 5760
rect 19429 5695 19487 5701
rect 19429 5692 19441 5695
rect 19168 5664 19441 5692
rect 19429 5661 19441 5664
rect 19475 5661 19487 5695
rect 19429 5655 19487 5661
rect 18782 5624 18788 5636
rect 16592 5596 16712 5624
rect 18743 5596 18788 5624
rect 10318 5516 10324 5568
rect 10376 5556 10382 5568
rect 12894 5556 12900 5568
rect 10376 5528 12900 5556
rect 10376 5516 10382 5528
rect 12894 5516 12900 5528
rect 12952 5516 12958 5568
rect 13909 5559 13967 5565
rect 13909 5525 13921 5559
rect 13955 5556 13967 5559
rect 13998 5556 14004 5568
rect 13955 5528 14004 5556
rect 13955 5525 13967 5528
rect 13909 5519 13967 5525
rect 13998 5516 14004 5528
rect 14056 5516 14062 5568
rect 14366 5516 14372 5568
rect 14424 5556 14430 5568
rect 16117 5559 16175 5565
rect 16117 5556 16129 5559
rect 14424 5528 16129 5556
rect 14424 5516 14430 5528
rect 16117 5525 16129 5528
rect 16163 5556 16175 5559
rect 16390 5556 16396 5568
rect 16163 5528 16396 5556
rect 16163 5525 16175 5528
rect 16117 5519 16175 5525
rect 16390 5516 16396 5528
rect 16448 5516 16454 5568
rect 16684 5556 16712 5596
rect 18782 5584 18788 5596
rect 18840 5584 18846 5636
rect 19444 5624 19472 5655
rect 19794 5652 19800 5704
rect 19852 5692 19858 5704
rect 20180 5692 20208 5732
rect 20901 5729 20913 5732
rect 20947 5729 20959 5763
rect 20901 5723 20959 5729
rect 21634 5720 21640 5772
rect 21692 5760 21698 5772
rect 21821 5763 21879 5769
rect 21821 5760 21833 5763
rect 21692 5732 21833 5760
rect 21692 5720 21698 5732
rect 21821 5729 21833 5732
rect 21867 5729 21879 5763
rect 21821 5723 21879 5729
rect 21913 5763 21971 5769
rect 21913 5729 21925 5763
rect 21959 5760 21971 5763
rect 22278 5760 22284 5772
rect 21959 5732 22284 5760
rect 21959 5729 21971 5732
rect 21913 5723 21971 5729
rect 22278 5720 22284 5732
rect 22336 5720 22342 5772
rect 22480 5769 22508 5800
rect 22465 5763 22523 5769
rect 22465 5729 22477 5763
rect 22511 5729 22523 5763
rect 22465 5723 22523 5729
rect 20346 5692 20352 5704
rect 19852 5664 20208 5692
rect 20307 5664 20352 5692
rect 19852 5652 19858 5664
rect 20346 5652 20352 5664
rect 20404 5652 20410 5704
rect 20438 5652 20444 5704
rect 20496 5692 20502 5704
rect 21269 5695 21327 5701
rect 21269 5692 21281 5695
rect 20496 5664 21281 5692
rect 20496 5652 20502 5664
rect 21269 5661 21281 5664
rect 21315 5661 21327 5695
rect 22094 5692 22100 5704
rect 22055 5664 22100 5692
rect 21269 5655 21327 5661
rect 22094 5652 22100 5664
rect 22152 5652 22158 5704
rect 19444 5596 21588 5624
rect 19334 5556 19340 5568
rect 16684 5528 19340 5556
rect 19334 5516 19340 5528
rect 19392 5516 19398 5568
rect 19794 5556 19800 5568
rect 19755 5528 19800 5556
rect 19794 5516 19800 5528
rect 19852 5516 19858 5568
rect 19978 5516 19984 5568
rect 20036 5556 20042 5568
rect 20254 5556 20260 5568
rect 20036 5528 20260 5556
rect 20036 5516 20042 5528
rect 20254 5516 20260 5528
rect 20312 5556 20318 5568
rect 21085 5559 21143 5565
rect 21085 5556 21097 5559
rect 20312 5528 21097 5556
rect 20312 5516 20318 5528
rect 21085 5525 21097 5528
rect 21131 5525 21143 5559
rect 21085 5519 21143 5525
rect 21269 5559 21327 5565
rect 21269 5525 21281 5559
rect 21315 5556 21327 5559
rect 21453 5559 21511 5565
rect 21453 5556 21465 5559
rect 21315 5528 21465 5556
rect 21315 5525 21327 5528
rect 21269 5519 21327 5525
rect 21453 5525 21465 5528
rect 21499 5525 21511 5559
rect 21560 5556 21588 5596
rect 22738 5556 22744 5568
rect 21560 5528 22744 5556
rect 21453 5519 21511 5525
rect 22738 5516 22744 5528
rect 22796 5516 22802 5568
rect 1104 5466 23276 5488
rect 1104 5414 4680 5466
rect 4732 5414 4744 5466
rect 4796 5414 4808 5466
rect 4860 5414 4872 5466
rect 4924 5414 12078 5466
rect 12130 5414 12142 5466
rect 12194 5414 12206 5466
rect 12258 5414 12270 5466
rect 12322 5414 19475 5466
rect 19527 5414 19539 5466
rect 19591 5414 19603 5466
rect 19655 5414 19667 5466
rect 19719 5414 23276 5466
rect 1104 5392 23276 5414
rect 7653 5355 7711 5361
rect 7653 5321 7665 5355
rect 7699 5352 7711 5355
rect 8938 5352 8944 5364
rect 7699 5324 8944 5352
rect 7699 5321 7711 5324
rect 7653 5315 7711 5321
rect 8938 5312 8944 5324
rect 8996 5312 9002 5364
rect 9122 5352 9128 5364
rect 9083 5324 9128 5352
rect 9122 5312 9128 5324
rect 9180 5312 9186 5364
rect 9858 5312 9864 5364
rect 9916 5352 9922 5364
rect 10137 5355 10195 5361
rect 10137 5352 10149 5355
rect 9916 5324 10149 5352
rect 9916 5312 9922 5324
rect 10137 5321 10149 5324
rect 10183 5321 10195 5355
rect 10686 5352 10692 5364
rect 10137 5315 10195 5321
rect 10336 5324 10692 5352
rect 10336 5284 10364 5324
rect 10686 5312 10692 5324
rect 10744 5312 10750 5364
rect 11146 5352 11152 5364
rect 11107 5324 11152 5352
rect 11146 5312 11152 5324
rect 11204 5312 11210 5364
rect 11330 5312 11336 5364
rect 11388 5352 11394 5364
rect 12437 5355 12495 5361
rect 12437 5352 12449 5355
rect 11388 5324 12449 5352
rect 11388 5312 11394 5324
rect 12437 5321 12449 5324
rect 12483 5321 12495 5355
rect 12437 5315 12495 5321
rect 13078 5312 13084 5364
rect 13136 5352 13142 5364
rect 13354 5352 13360 5364
rect 13136 5324 13360 5352
rect 13136 5312 13142 5324
rect 13354 5312 13360 5324
rect 13412 5312 13418 5364
rect 14458 5352 14464 5364
rect 13556 5324 14464 5352
rect 13446 5284 13452 5296
rect 9784 5256 10364 5284
rect 10520 5256 13452 5284
rect 9784 5228 9812 5256
rect 7742 5176 7748 5228
rect 7800 5216 7806 5228
rect 8205 5219 8263 5225
rect 8205 5216 8217 5219
rect 7800 5188 8217 5216
rect 7800 5176 7806 5188
rect 8205 5185 8217 5188
rect 8251 5185 8263 5219
rect 9766 5216 9772 5228
rect 9727 5188 9772 5216
rect 8205 5179 8263 5185
rect 9766 5176 9772 5188
rect 9824 5176 9830 5228
rect 7374 5108 7380 5160
rect 7432 5148 7438 5160
rect 10520 5157 10548 5256
rect 13446 5244 13452 5256
rect 13504 5244 13510 5296
rect 10686 5216 10692 5228
rect 10647 5188 10692 5216
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 11606 5216 11612 5228
rect 11567 5188 11612 5216
rect 11606 5176 11612 5188
rect 11664 5176 11670 5228
rect 11793 5219 11851 5225
rect 11793 5185 11805 5219
rect 11839 5185 11851 5219
rect 11793 5179 11851 5185
rect 8021 5151 8079 5157
rect 8021 5148 8033 5151
rect 7432 5120 8033 5148
rect 7432 5108 7438 5120
rect 8021 5117 8033 5120
rect 8067 5117 8079 5151
rect 8021 5111 8079 5117
rect 10505 5151 10563 5157
rect 10505 5117 10517 5151
rect 10551 5117 10563 5151
rect 10505 5111 10563 5117
rect 10597 5151 10655 5157
rect 10597 5117 10609 5151
rect 10643 5148 10655 5151
rect 11514 5148 11520 5160
rect 10643 5120 11376 5148
rect 11475 5120 11520 5148
rect 10643 5117 10655 5120
rect 10597 5111 10655 5117
rect 7926 5040 7932 5092
rect 7984 5080 7990 5092
rect 8113 5083 8171 5089
rect 8113 5080 8125 5083
rect 7984 5052 8125 5080
rect 7984 5040 7990 5052
rect 8113 5049 8125 5052
rect 8159 5049 8171 5083
rect 8113 5043 8171 5049
rect 9493 5083 9551 5089
rect 9493 5049 9505 5083
rect 9539 5080 9551 5083
rect 11348 5080 11376 5120
rect 11514 5108 11520 5120
rect 11572 5108 11578 5160
rect 11808 5148 11836 5179
rect 12434 5176 12440 5228
rect 12492 5216 12498 5228
rect 12897 5219 12955 5225
rect 12897 5216 12909 5219
rect 12492 5188 12909 5216
rect 12492 5176 12498 5188
rect 12897 5185 12909 5188
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5216 13139 5219
rect 13556 5216 13584 5324
rect 14458 5312 14464 5324
rect 14516 5312 14522 5364
rect 14918 5312 14924 5364
rect 14976 5352 14982 5364
rect 16577 5355 16635 5361
rect 16577 5352 16589 5355
rect 14976 5324 16589 5352
rect 14976 5312 14982 5324
rect 16577 5321 16589 5324
rect 16623 5321 16635 5355
rect 16850 5352 16856 5364
rect 16811 5324 16856 5352
rect 16577 5315 16635 5321
rect 16850 5312 16856 5324
rect 16908 5312 16914 5364
rect 18230 5312 18236 5364
rect 18288 5352 18294 5364
rect 18509 5355 18567 5361
rect 18509 5352 18521 5355
rect 18288 5324 18521 5352
rect 18288 5312 18294 5324
rect 18509 5321 18521 5324
rect 18555 5321 18567 5355
rect 18509 5315 18567 5321
rect 20070 5312 20076 5364
rect 20128 5352 20134 5364
rect 20809 5355 20867 5361
rect 20809 5352 20821 5355
rect 20128 5324 20821 5352
rect 20128 5312 20134 5324
rect 20809 5321 20821 5324
rect 20855 5321 20867 5355
rect 20809 5315 20867 5321
rect 21818 5312 21824 5364
rect 21876 5352 21882 5364
rect 22557 5355 22615 5361
rect 22557 5352 22569 5355
rect 21876 5324 22569 5352
rect 21876 5312 21882 5324
rect 22557 5321 22569 5324
rect 22603 5321 22615 5355
rect 22557 5315 22615 5321
rect 19613 5287 19671 5293
rect 19613 5253 19625 5287
rect 19659 5284 19671 5287
rect 20714 5284 20720 5296
rect 19659 5256 20720 5284
rect 19659 5253 19671 5256
rect 19613 5247 19671 5253
rect 20714 5244 20720 5256
rect 20772 5244 20778 5296
rect 13127 5188 13584 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 13096 5148 13124 5179
rect 14734 5176 14740 5228
rect 14792 5216 14798 5228
rect 15197 5219 15255 5225
rect 15197 5216 15209 5219
rect 14792 5188 15209 5216
rect 14792 5176 14798 5188
rect 15197 5185 15209 5188
rect 15243 5185 15255 5219
rect 15197 5179 15255 5185
rect 17497 5219 17555 5225
rect 17497 5185 17509 5219
rect 17543 5216 17555 5219
rect 17586 5216 17592 5228
rect 17543 5188 17592 5216
rect 17543 5185 17555 5188
rect 17497 5179 17555 5185
rect 17586 5176 17592 5188
rect 17644 5176 17650 5228
rect 17862 5176 17868 5228
rect 17920 5216 17926 5228
rect 18049 5219 18107 5225
rect 18049 5216 18061 5219
rect 17920 5188 18061 5216
rect 17920 5176 17926 5188
rect 18049 5185 18061 5188
rect 18095 5185 18107 5219
rect 18049 5179 18107 5185
rect 18138 5176 18144 5228
rect 18196 5216 18202 5228
rect 18969 5219 19027 5225
rect 18969 5216 18981 5219
rect 18196 5188 18981 5216
rect 18196 5176 18202 5188
rect 18969 5185 18981 5188
rect 19015 5185 19027 5219
rect 19150 5216 19156 5228
rect 19111 5188 19156 5216
rect 18969 5179 19027 5185
rect 19150 5176 19156 5188
rect 19208 5176 19214 5228
rect 20254 5216 20260 5228
rect 20167 5188 20260 5216
rect 20254 5176 20260 5188
rect 20312 5216 20318 5228
rect 20898 5216 20904 5228
rect 20312 5188 20904 5216
rect 20312 5176 20318 5188
rect 20898 5176 20904 5188
rect 20956 5176 20962 5228
rect 11808 5120 13124 5148
rect 13354 5108 13360 5160
rect 13412 5148 13418 5160
rect 13541 5151 13599 5157
rect 13541 5148 13553 5151
rect 13412 5120 13553 5148
rect 13412 5108 13418 5120
rect 13541 5117 13553 5120
rect 13587 5117 13599 5151
rect 13541 5111 13599 5117
rect 13808 5151 13866 5157
rect 13808 5117 13820 5151
rect 13854 5148 13866 5151
rect 14182 5148 14188 5160
rect 13854 5120 14188 5148
rect 13854 5117 13866 5120
rect 13808 5111 13866 5117
rect 14182 5108 14188 5120
rect 14240 5108 14246 5160
rect 16022 5108 16028 5160
rect 16080 5148 16086 5160
rect 16080 5120 17724 5148
rect 16080 5108 16086 5120
rect 12618 5080 12624 5092
rect 9539 5052 10631 5080
rect 11348 5052 12624 5080
rect 9539 5049 9551 5052
rect 9493 5043 9551 5049
rect 9582 5012 9588 5024
rect 9543 4984 9588 5012
rect 9582 4972 9588 4984
rect 9640 4972 9646 5024
rect 10603 5012 10631 5052
rect 12618 5040 12624 5052
rect 12676 5040 12682 5092
rect 15442 5083 15500 5089
rect 12728 5052 13768 5080
rect 12250 5012 12256 5024
rect 10603 4984 12256 5012
rect 12250 4972 12256 4984
rect 12308 4972 12314 5024
rect 12342 4972 12348 5024
rect 12400 5012 12406 5024
rect 12728 5012 12756 5052
rect 12400 4984 12756 5012
rect 12400 4972 12406 4984
rect 12802 4972 12808 5024
rect 12860 5012 12866 5024
rect 13740 5012 13768 5052
rect 15442 5049 15454 5083
rect 15488 5049 15500 5083
rect 15442 5043 15500 5049
rect 14921 5015 14979 5021
rect 14921 5012 14933 5015
rect 12860 4984 12905 5012
rect 13740 4984 14933 5012
rect 12860 4972 12866 4984
rect 14921 4981 14933 4984
rect 14967 5012 14979 5015
rect 15457 5012 15485 5043
rect 15562 5040 15568 5092
rect 15620 5080 15626 5092
rect 17313 5083 17371 5089
rect 17313 5080 17325 5083
rect 15620 5052 17325 5080
rect 15620 5040 15626 5052
rect 17313 5049 17325 5052
rect 17359 5049 17371 5083
rect 17696 5080 17724 5120
rect 17770 5108 17776 5160
rect 17828 5148 17834 5160
rect 19426 5148 19432 5160
rect 17828 5120 19432 5148
rect 17828 5108 17834 5120
rect 19426 5108 19432 5120
rect 19484 5108 19490 5160
rect 20625 5151 20683 5157
rect 20625 5117 20637 5151
rect 20671 5148 20683 5151
rect 20714 5148 20720 5160
rect 20671 5120 20720 5148
rect 20671 5117 20683 5120
rect 20625 5111 20683 5117
rect 20714 5108 20720 5120
rect 20772 5108 20778 5160
rect 21174 5148 21180 5160
rect 21135 5120 21180 5148
rect 21174 5108 21180 5120
rect 21232 5108 21238 5160
rect 17862 5080 17868 5092
rect 17696 5052 17868 5080
rect 17313 5043 17371 5049
rect 17862 5040 17868 5052
rect 17920 5040 17926 5092
rect 18322 5040 18328 5092
rect 18380 5080 18386 5092
rect 18380 5052 19012 5080
rect 18380 5040 18386 5052
rect 17218 5012 17224 5024
rect 14967 4984 15485 5012
rect 17179 4984 17224 5012
rect 14967 4981 14979 4984
rect 14921 4975 14979 4981
rect 17218 4972 17224 4984
rect 17276 4972 17282 5024
rect 17494 4972 17500 5024
rect 17552 5012 17558 5024
rect 18877 5015 18935 5021
rect 18877 5012 18889 5015
rect 17552 4984 18889 5012
rect 17552 4972 17558 4984
rect 18877 4981 18889 4984
rect 18923 4981 18935 5015
rect 18984 5012 19012 5052
rect 19334 5040 19340 5092
rect 19392 5080 19398 5092
rect 19981 5083 20039 5089
rect 19981 5080 19993 5083
rect 19392 5052 19993 5080
rect 19392 5040 19398 5052
rect 19981 5049 19993 5052
rect 20027 5049 20039 5083
rect 19981 5043 20039 5049
rect 21444 5083 21502 5089
rect 21444 5049 21456 5083
rect 21490 5080 21502 5083
rect 22094 5080 22100 5092
rect 21490 5052 22100 5080
rect 21490 5049 21502 5052
rect 21444 5043 21502 5049
rect 22094 5040 22100 5052
rect 22152 5040 22158 5092
rect 20073 5015 20131 5021
rect 20073 5012 20085 5015
rect 18984 4984 20085 5012
rect 18877 4975 18935 4981
rect 20073 4981 20085 4984
rect 20119 4981 20131 5015
rect 20073 4975 20131 4981
rect 1104 4922 23276 4944
rect 1104 4870 8379 4922
rect 8431 4870 8443 4922
rect 8495 4870 8507 4922
rect 8559 4870 8571 4922
rect 8623 4870 15776 4922
rect 15828 4870 15840 4922
rect 15892 4870 15904 4922
rect 15956 4870 15968 4922
rect 16020 4870 23276 4922
rect 1104 4848 23276 4870
rect 9858 4808 9864 4820
rect 9819 4780 9864 4808
rect 9858 4768 9864 4780
rect 9916 4768 9922 4820
rect 10229 4811 10287 4817
rect 10229 4777 10241 4811
rect 10275 4808 10287 4811
rect 10778 4808 10784 4820
rect 10275 4780 10784 4808
rect 10275 4777 10287 4780
rect 10229 4771 10287 4777
rect 10778 4768 10784 4780
rect 10836 4768 10842 4820
rect 11333 4811 11391 4817
rect 11333 4777 11345 4811
rect 11379 4808 11391 4811
rect 11698 4808 11704 4820
rect 11379 4780 11704 4808
rect 11379 4777 11391 4780
rect 11333 4771 11391 4777
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 11882 4808 11888 4820
rect 11843 4780 11888 4808
rect 11882 4768 11888 4780
rect 11940 4768 11946 4820
rect 11974 4768 11980 4820
rect 12032 4808 12038 4820
rect 12345 4811 12403 4817
rect 12345 4808 12357 4811
rect 12032 4780 12357 4808
rect 12032 4768 12038 4780
rect 12345 4777 12357 4780
rect 12391 4777 12403 4811
rect 12345 4771 12403 4777
rect 12897 4811 12955 4817
rect 12897 4777 12909 4811
rect 12943 4808 12955 4811
rect 12986 4808 12992 4820
rect 12943 4780 12992 4808
rect 12943 4777 12955 4780
rect 12897 4771 12955 4777
rect 12986 4768 12992 4780
rect 13044 4768 13050 4820
rect 13265 4811 13323 4817
rect 13265 4777 13277 4811
rect 13311 4808 13323 4811
rect 13909 4811 13967 4817
rect 13909 4808 13921 4811
rect 13311 4780 13921 4808
rect 13311 4777 13323 4780
rect 13265 4771 13323 4777
rect 13909 4777 13921 4780
rect 13955 4777 13967 4811
rect 13909 4771 13967 4777
rect 14277 4811 14335 4817
rect 14277 4777 14289 4811
rect 14323 4808 14335 4811
rect 14826 4808 14832 4820
rect 14323 4780 14832 4808
rect 14323 4777 14335 4780
rect 14277 4771 14335 4777
rect 14826 4768 14832 4780
rect 14884 4768 14890 4820
rect 15473 4811 15531 4817
rect 15473 4777 15485 4811
rect 15519 4808 15531 4811
rect 17494 4808 17500 4820
rect 15519 4780 17500 4808
rect 15519 4777 15531 4780
rect 15473 4771 15531 4777
rect 17494 4768 17500 4780
rect 17552 4768 17558 4820
rect 17770 4808 17776 4820
rect 17731 4780 17776 4808
rect 17770 4768 17776 4780
rect 17828 4768 17834 4820
rect 18230 4808 18236 4820
rect 18191 4780 18236 4808
rect 18230 4768 18236 4780
rect 18288 4768 18294 4820
rect 19153 4811 19211 4817
rect 19153 4777 19165 4811
rect 19199 4808 19211 4811
rect 19797 4811 19855 4817
rect 19797 4808 19809 4811
rect 19199 4780 19809 4808
rect 19199 4777 19211 4780
rect 19153 4771 19211 4777
rect 19797 4777 19809 4780
rect 19843 4777 19855 4811
rect 19797 4771 19855 4777
rect 20165 4811 20223 4817
rect 20165 4777 20177 4811
rect 20211 4808 20223 4811
rect 22094 4808 22100 4820
rect 20211 4780 22100 4808
rect 20211 4777 20223 4780
rect 20165 4771 20223 4777
rect 22094 4768 22100 4780
rect 22152 4808 22158 4820
rect 22465 4811 22523 4817
rect 22465 4808 22477 4811
rect 22152 4780 22477 4808
rect 22152 4768 22158 4780
rect 22465 4777 22477 4780
rect 22511 4777 22523 4811
rect 22465 4771 22523 4777
rect 10318 4740 10324 4752
rect 10279 4712 10324 4740
rect 10318 4700 10324 4712
rect 10376 4700 10382 4752
rect 13354 4740 13360 4752
rect 13315 4712 13360 4740
rect 13354 4700 13360 4712
rect 13412 4700 13418 4752
rect 14369 4743 14427 4749
rect 14369 4709 14381 4743
rect 14415 4740 14427 4743
rect 14550 4740 14556 4752
rect 14415 4712 14556 4740
rect 14415 4709 14427 4712
rect 14369 4703 14427 4709
rect 14550 4700 14556 4712
rect 14608 4700 14614 4752
rect 18046 4740 18052 4752
rect 15304 4712 18052 4740
rect 11241 4675 11299 4681
rect 11241 4641 11253 4675
rect 11287 4672 11299 4675
rect 11882 4672 11888 4684
rect 11287 4644 11888 4672
rect 11287 4641 11299 4644
rect 11241 4635 11299 4641
rect 11882 4632 11888 4644
rect 11940 4632 11946 4684
rect 12253 4675 12311 4681
rect 12253 4672 12265 4675
rect 11992 4644 12265 4672
rect 10505 4607 10563 4613
rect 10505 4573 10517 4607
rect 10551 4604 10563 4607
rect 10686 4604 10692 4616
rect 10551 4576 10692 4604
rect 10551 4573 10563 4576
rect 10505 4567 10563 4573
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 11517 4607 11575 4613
rect 11517 4573 11529 4607
rect 11563 4604 11575 4607
rect 11606 4604 11612 4616
rect 11563 4576 11612 4604
rect 11563 4573 11575 4576
rect 11517 4567 11575 4573
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 11793 4607 11851 4613
rect 11793 4573 11805 4607
rect 11839 4604 11851 4607
rect 11992 4604 12020 4644
rect 12253 4641 12265 4644
rect 12299 4672 12311 4675
rect 14182 4672 14188 4684
rect 12299 4644 14188 4672
rect 12299 4641 12311 4644
rect 12253 4635 12311 4641
rect 14182 4632 14188 4644
rect 14240 4632 14246 4684
rect 15304 4681 15332 4712
rect 18046 4700 18052 4712
rect 18104 4700 18110 4752
rect 19245 4743 19303 4749
rect 19245 4709 19257 4743
rect 19291 4740 19303 4743
rect 20438 4740 20444 4752
rect 19291 4712 20444 4740
rect 19291 4709 19303 4712
rect 19245 4703 19303 4709
rect 20438 4700 20444 4712
rect 20496 4700 20502 4752
rect 21008 4712 21312 4740
rect 15289 4675 15347 4681
rect 15289 4641 15301 4675
rect 15335 4641 15347 4675
rect 15289 4635 15347 4641
rect 15654 4632 15660 4684
rect 15712 4672 15718 4684
rect 16097 4675 16155 4681
rect 16097 4672 16109 4675
rect 15712 4644 16109 4672
rect 15712 4632 15718 4644
rect 16097 4641 16109 4644
rect 16143 4641 16155 4675
rect 16097 4635 16155 4641
rect 16666 4632 16672 4684
rect 16724 4672 16730 4684
rect 16724 4644 16896 4672
rect 16724 4632 16730 4644
rect 11839 4576 12020 4604
rect 11839 4573 11851 4576
rect 11793 4567 11851 4573
rect 12434 4564 12440 4616
rect 12492 4604 12498 4616
rect 12492 4576 12537 4604
rect 12492 4564 12498 4576
rect 12894 4564 12900 4616
rect 12952 4604 12958 4616
rect 13449 4607 13507 4613
rect 13449 4604 13461 4607
rect 12952 4576 13461 4604
rect 12952 4564 12958 4576
rect 13449 4573 13461 4576
rect 13495 4573 13507 4607
rect 14458 4604 14464 4616
rect 14419 4576 14464 4604
rect 13449 4567 13507 4573
rect 14458 4564 14464 4576
rect 14516 4564 14522 4616
rect 15841 4607 15899 4613
rect 15841 4573 15853 4607
rect 15887 4573 15899 4607
rect 16868 4604 16896 4644
rect 16942 4632 16948 4684
rect 17000 4672 17006 4684
rect 17310 4672 17316 4684
rect 17000 4644 17316 4672
rect 17000 4632 17006 4644
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 18141 4675 18199 4681
rect 18141 4641 18153 4675
rect 18187 4672 18199 4675
rect 19794 4672 19800 4684
rect 18187 4644 19800 4672
rect 18187 4641 18199 4644
rect 18141 4635 18199 4641
rect 19794 4632 19800 4644
rect 19852 4632 19858 4684
rect 20257 4675 20315 4681
rect 20257 4641 20269 4675
rect 20303 4672 20315 4675
rect 21008 4672 21036 4712
rect 20303 4644 21036 4672
rect 21085 4675 21143 4681
rect 20303 4641 20315 4644
rect 20257 4635 20315 4641
rect 21085 4641 21097 4675
rect 21131 4672 21143 4675
rect 21174 4672 21180 4684
rect 21131 4644 21180 4672
rect 21131 4641 21143 4644
rect 21085 4635 21143 4641
rect 21174 4632 21180 4644
rect 21232 4632 21238 4684
rect 21284 4672 21312 4712
rect 21358 4681 21364 4684
rect 21352 4672 21364 4681
rect 21284 4644 21364 4672
rect 21352 4635 21364 4644
rect 21358 4632 21364 4635
rect 21416 4632 21422 4684
rect 18325 4607 18383 4613
rect 18325 4604 18337 4607
rect 16868 4576 18337 4604
rect 15841 4567 15899 4573
rect 18325 4573 18337 4576
rect 18371 4573 18383 4607
rect 18325 4567 18383 4573
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 10873 4539 10931 4545
rect 10873 4505 10885 4539
rect 10919 4536 10931 4539
rect 15562 4536 15568 4548
rect 10919 4508 15568 4536
rect 10919 4505 10931 4508
rect 10873 4499 10931 4505
rect 15562 4496 15568 4508
rect 15620 4496 15626 4548
rect 15856 4480 15884 4567
rect 17034 4496 17040 4548
rect 17092 4536 17098 4548
rect 18785 4539 18843 4545
rect 18785 4536 18797 4539
rect 17092 4508 18797 4536
rect 17092 4496 17098 4508
rect 18785 4505 18797 4508
rect 18831 4505 18843 4539
rect 18785 4499 18843 4505
rect 18874 4496 18880 4548
rect 18932 4536 18938 4548
rect 19444 4536 19472 4567
rect 20070 4564 20076 4616
rect 20128 4604 20134 4616
rect 20349 4607 20407 4613
rect 20349 4604 20361 4607
rect 20128 4576 20361 4604
rect 20128 4564 20134 4576
rect 20349 4573 20361 4576
rect 20395 4573 20407 4607
rect 20349 4567 20407 4573
rect 20254 4536 20260 4548
rect 18932 4508 20260 4536
rect 18932 4496 18938 4508
rect 20254 4496 20260 4508
rect 20312 4496 20318 4548
rect 6914 4428 6920 4480
rect 6972 4468 6978 4480
rect 11793 4471 11851 4477
rect 11793 4468 11805 4471
rect 6972 4440 11805 4468
rect 6972 4428 6978 4440
rect 11793 4437 11805 4440
rect 11839 4437 11851 4471
rect 11793 4431 11851 4437
rect 11974 4428 11980 4480
rect 12032 4468 12038 4480
rect 14918 4468 14924 4480
rect 12032 4440 14924 4468
rect 12032 4428 12038 4440
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 15286 4428 15292 4480
rect 15344 4468 15350 4480
rect 15838 4468 15844 4480
rect 15344 4440 15844 4468
rect 15344 4428 15350 4440
rect 15838 4428 15844 4440
rect 15896 4428 15902 4480
rect 16574 4428 16580 4480
rect 16632 4468 16638 4480
rect 17221 4471 17279 4477
rect 17221 4468 17233 4471
rect 16632 4440 17233 4468
rect 16632 4428 16638 4440
rect 17221 4437 17233 4440
rect 17267 4437 17279 4471
rect 17221 4431 17279 4437
rect 17678 4428 17684 4480
rect 17736 4468 17742 4480
rect 20806 4468 20812 4480
rect 17736 4440 20812 4468
rect 17736 4428 17742 4440
rect 20806 4428 20812 4440
rect 20864 4428 20870 4480
rect 1104 4378 23276 4400
rect 1104 4326 4680 4378
rect 4732 4326 4744 4378
rect 4796 4326 4808 4378
rect 4860 4326 4872 4378
rect 4924 4326 12078 4378
rect 12130 4326 12142 4378
rect 12194 4326 12206 4378
rect 12258 4326 12270 4378
rect 12322 4326 19475 4378
rect 19527 4326 19539 4378
rect 19591 4326 19603 4378
rect 19655 4326 19667 4378
rect 19719 4326 23276 4378
rect 1104 4304 23276 4326
rect 9582 4224 9588 4276
rect 9640 4264 9646 4276
rect 13262 4264 13268 4276
rect 9640 4236 13268 4264
rect 9640 4224 9646 4236
rect 13262 4224 13268 4236
rect 13320 4224 13326 4276
rect 13630 4264 13636 4276
rect 13591 4236 13636 4264
rect 13630 4224 13636 4236
rect 13688 4224 13694 4276
rect 14826 4264 14832 4276
rect 14660 4236 14832 4264
rect 8202 4156 8208 4208
rect 8260 4196 8266 4208
rect 14461 4199 14519 4205
rect 14461 4196 14473 4199
rect 8260 4168 14473 4196
rect 8260 4156 8266 4168
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 11793 4131 11851 4137
rect 11793 4128 11805 4131
rect 9272 4100 11805 4128
rect 9272 4088 9278 4100
rect 11793 4097 11805 4100
rect 11839 4097 11851 4131
rect 11793 4091 11851 4097
rect 11882 4088 11888 4140
rect 11940 4128 11946 4140
rect 13188 4137 13216 4168
rect 14461 4165 14473 4168
rect 14507 4165 14519 4199
rect 14461 4159 14519 4165
rect 13173 4131 13231 4137
rect 11940 4100 11985 4128
rect 11940 4088 11946 4100
rect 13173 4097 13185 4131
rect 13219 4097 13231 4131
rect 14090 4128 14096 4140
rect 13173 4091 13231 4097
rect 13280 4100 14096 4128
rect 13280 4060 13308 4100
rect 14090 4088 14096 4100
rect 14148 4088 14154 4140
rect 14277 4131 14335 4137
rect 14277 4097 14289 4131
rect 14323 4128 14335 4131
rect 14660 4128 14688 4236
rect 14826 4224 14832 4236
rect 14884 4264 14890 4276
rect 18046 4264 18052 4276
rect 14884 4236 17264 4264
rect 18007 4236 18052 4264
rect 14884 4224 14890 4236
rect 15654 4156 15660 4208
rect 15712 4196 15718 4208
rect 16025 4199 16083 4205
rect 16025 4196 16037 4199
rect 15712 4168 16037 4196
rect 15712 4156 15718 4168
rect 16025 4165 16037 4168
rect 16071 4165 16083 4199
rect 17236 4196 17264 4236
rect 18046 4224 18052 4236
rect 18104 4224 18110 4276
rect 22002 4264 22008 4276
rect 18156 4236 22008 4264
rect 18156 4196 18184 4236
rect 22002 4224 22008 4236
rect 22060 4224 22066 4276
rect 17236 4168 18184 4196
rect 16025 4159 16083 4165
rect 14323 4100 14688 4128
rect 14323 4097 14335 4100
rect 14277 4091 14335 4097
rect 15838 4088 15844 4140
rect 15896 4128 15902 4140
rect 16209 4131 16267 4137
rect 16209 4128 16221 4131
rect 15896 4100 16221 4128
rect 15896 4088 15902 4100
rect 16209 4097 16221 4100
rect 16255 4128 16267 4131
rect 16301 4131 16359 4137
rect 16301 4128 16313 4131
rect 16255 4100 16313 4128
rect 16255 4097 16267 4100
rect 16209 4091 16267 4097
rect 16301 4097 16313 4100
rect 16347 4097 16359 4131
rect 16301 4091 16359 4097
rect 17586 4088 17592 4140
rect 17644 4128 17650 4140
rect 18693 4131 18751 4137
rect 18693 4128 18705 4131
rect 17644 4100 18705 4128
rect 17644 4088 17650 4100
rect 18693 4097 18705 4100
rect 18739 4128 18751 4131
rect 18874 4128 18880 4140
rect 18739 4100 18880 4128
rect 18739 4097 18751 4100
rect 18693 4091 18751 4097
rect 18874 4088 18880 4100
rect 18932 4088 18938 4140
rect 19058 4128 19064 4140
rect 19019 4100 19064 4128
rect 19058 4088 19064 4100
rect 19116 4088 19122 4140
rect 20990 4088 20996 4140
rect 21048 4128 21054 4140
rect 21266 4128 21272 4140
rect 21048 4100 21272 4128
rect 21048 4088 21054 4100
rect 21266 4088 21272 4100
rect 21324 4088 21330 4140
rect 13998 4060 14004 4072
rect 12452 4032 13308 4060
rect 13959 4032 14004 4060
rect 12452 3992 12480 4032
rect 13998 4020 14004 4032
rect 14056 4020 14062 4072
rect 14645 4063 14703 4069
rect 14645 4029 14657 4063
rect 14691 4060 14703 4063
rect 14734 4060 14740 4072
rect 14691 4032 14740 4060
rect 14691 4029 14703 4032
rect 14645 4023 14703 4029
rect 14734 4020 14740 4032
rect 14792 4020 14798 4072
rect 14918 4069 14924 4072
rect 14912 4060 14924 4069
rect 14879 4032 14924 4060
rect 14912 4023 14924 4032
rect 14918 4020 14924 4023
rect 14976 4020 14982 4072
rect 18417 4063 18475 4069
rect 18417 4060 18429 4063
rect 15028 4032 18429 4060
rect 15028 3992 15056 4032
rect 18417 4029 18429 4032
rect 18463 4029 18475 4063
rect 18417 4023 18475 4029
rect 18966 4020 18972 4072
rect 19024 4060 19030 4072
rect 19521 4063 19579 4069
rect 19521 4060 19533 4063
rect 19024 4032 19533 4060
rect 19024 4020 19030 4032
rect 19521 4029 19533 4032
rect 19567 4060 19579 4063
rect 20346 4060 20352 4072
rect 19567 4032 20352 4060
rect 19567 4029 19579 4032
rect 19521 4023 19579 4029
rect 20346 4020 20352 4032
rect 20404 4060 20410 4072
rect 21174 4060 21180 4072
rect 20404 4032 21180 4060
rect 20404 4020 20410 4032
rect 21174 4020 21180 4032
rect 21232 4060 21238 4072
rect 21634 4069 21640 4072
rect 21361 4063 21419 4069
rect 21361 4060 21373 4063
rect 21232 4032 21373 4060
rect 21232 4020 21238 4032
rect 21361 4029 21373 4032
rect 21407 4029 21419 4063
rect 21628 4060 21640 4069
rect 21595 4032 21640 4060
rect 21361 4023 21419 4029
rect 21628 4023 21640 4032
rect 21634 4020 21640 4023
rect 21692 4020 21698 4072
rect 16574 4001 16580 4004
rect 11348 3964 12480 3992
rect 12544 3964 15056 3992
rect 11348 3933 11376 3964
rect 11333 3927 11391 3933
rect 11333 3893 11345 3927
rect 11379 3893 11391 3927
rect 11333 3887 11391 3893
rect 11422 3884 11428 3936
rect 11480 3924 11486 3936
rect 11701 3927 11759 3933
rect 11701 3924 11713 3927
rect 11480 3896 11713 3924
rect 11480 3884 11486 3896
rect 11701 3893 11713 3896
rect 11747 3893 11759 3927
rect 11701 3887 11759 3893
rect 12158 3884 12164 3936
rect 12216 3924 12222 3936
rect 12544 3924 12572 3964
rect 16568 3955 16580 4001
rect 16632 3992 16638 4004
rect 16632 3964 16668 3992
rect 16574 3952 16580 3955
rect 16632 3952 16638 3964
rect 19150 3952 19156 4004
rect 19208 3992 19214 4004
rect 19766 3995 19824 4001
rect 19766 3992 19778 3995
rect 19208 3964 19778 3992
rect 19208 3952 19214 3964
rect 19766 3961 19778 3964
rect 19812 3961 19824 3995
rect 19766 3955 19824 3961
rect 12216 3896 12572 3924
rect 12216 3884 12222 3896
rect 12618 3884 12624 3936
rect 12676 3924 12682 3936
rect 12986 3924 12992 3936
rect 12676 3896 12721 3924
rect 12947 3896 12992 3924
rect 12676 3884 12682 3896
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 13078 3884 13084 3936
rect 13136 3924 13142 3936
rect 14093 3927 14151 3933
rect 13136 3896 13181 3924
rect 13136 3884 13142 3896
rect 14093 3893 14105 3927
rect 14139 3924 14151 3927
rect 14366 3924 14372 3936
rect 14139 3896 14372 3924
rect 14139 3893 14151 3896
rect 14093 3887 14151 3893
rect 14366 3884 14372 3896
rect 14424 3884 14430 3936
rect 14461 3927 14519 3933
rect 14461 3893 14473 3927
rect 14507 3924 14519 3927
rect 15010 3924 15016 3936
rect 14507 3896 15016 3924
rect 14507 3893 14519 3896
rect 14461 3887 14519 3893
rect 15010 3884 15016 3896
rect 15068 3884 15074 3936
rect 16209 3927 16267 3933
rect 16209 3893 16221 3927
rect 16255 3924 16267 3927
rect 17034 3924 17040 3936
rect 16255 3896 17040 3924
rect 16255 3893 16267 3896
rect 16209 3887 16267 3893
rect 17034 3884 17040 3896
rect 17092 3884 17098 3936
rect 17678 3924 17684 3936
rect 17639 3896 17684 3924
rect 17678 3884 17684 3896
rect 17736 3884 17742 3936
rect 18506 3924 18512 3936
rect 18467 3896 18512 3924
rect 18506 3884 18512 3896
rect 18564 3884 18570 3936
rect 20901 3927 20959 3933
rect 20901 3893 20913 3927
rect 20947 3924 20959 3927
rect 21266 3924 21272 3936
rect 20947 3896 21272 3924
rect 20947 3893 20959 3896
rect 20901 3887 20959 3893
rect 21266 3884 21272 3896
rect 21324 3884 21330 3936
rect 21358 3884 21364 3936
rect 21416 3924 21422 3936
rect 22741 3927 22799 3933
rect 22741 3924 22753 3927
rect 21416 3896 22753 3924
rect 21416 3884 21422 3896
rect 22741 3893 22753 3896
rect 22787 3893 22799 3927
rect 22741 3887 22799 3893
rect 1104 3834 23276 3856
rect 1104 3782 8379 3834
rect 8431 3782 8443 3834
rect 8495 3782 8507 3834
rect 8559 3782 8571 3834
rect 8623 3782 15776 3834
rect 15828 3782 15840 3834
rect 15892 3782 15904 3834
rect 15956 3782 15968 3834
rect 16020 3782 23276 3834
rect 1104 3760 23276 3782
rect 11149 3723 11207 3729
rect 11149 3689 11161 3723
rect 11195 3720 11207 3723
rect 11422 3720 11428 3732
rect 11195 3692 11428 3720
rect 11195 3689 11207 3692
rect 11149 3683 11207 3689
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 11609 3723 11667 3729
rect 11609 3689 11621 3723
rect 11655 3720 11667 3723
rect 13170 3720 13176 3732
rect 11655 3692 13176 3720
rect 11655 3689 11667 3692
rect 11609 3683 11667 3689
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 13538 3720 13544 3732
rect 13499 3692 13544 3720
rect 13538 3680 13544 3692
rect 13596 3680 13602 3732
rect 13633 3723 13691 3729
rect 13633 3689 13645 3723
rect 13679 3720 13691 3723
rect 13722 3720 13728 3732
rect 13679 3692 13728 3720
rect 13679 3689 13691 3692
rect 13633 3683 13691 3689
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 14185 3723 14243 3729
rect 14185 3689 14197 3723
rect 14231 3720 14243 3723
rect 14274 3720 14280 3732
rect 14231 3692 14280 3720
rect 14231 3689 14243 3692
rect 14185 3683 14243 3689
rect 14274 3680 14280 3692
rect 14332 3680 14338 3732
rect 14553 3723 14611 3729
rect 14553 3689 14565 3723
rect 14599 3720 14611 3723
rect 15933 3723 15991 3729
rect 15933 3720 15945 3723
rect 14599 3692 15945 3720
rect 14599 3689 14611 3692
rect 14553 3683 14611 3689
rect 15933 3689 15945 3692
rect 15979 3689 15991 3723
rect 16114 3720 16120 3732
rect 16075 3692 16120 3720
rect 15933 3683 15991 3689
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 16485 3723 16543 3729
rect 16485 3689 16497 3723
rect 16531 3720 16543 3723
rect 16942 3720 16948 3732
rect 16531 3692 16948 3720
rect 16531 3689 16543 3692
rect 16485 3683 16543 3689
rect 16942 3680 16948 3692
rect 17000 3680 17006 3732
rect 18509 3723 18567 3729
rect 18509 3720 18521 3723
rect 17052 3692 18521 3720
rect 11517 3655 11575 3661
rect 11517 3621 11529 3655
rect 11563 3652 11575 3655
rect 12434 3652 12440 3664
rect 11563 3624 12440 3652
rect 11563 3621 11575 3624
rect 11517 3615 11575 3621
rect 12434 3612 12440 3624
rect 12492 3612 12498 3664
rect 12621 3655 12679 3661
rect 12621 3621 12633 3655
rect 12667 3652 12679 3655
rect 17052 3652 17080 3692
rect 18509 3689 18521 3692
rect 18555 3720 18567 3723
rect 18598 3720 18604 3732
rect 18555 3692 18604 3720
rect 18555 3689 18567 3692
rect 18509 3683 18567 3689
rect 18598 3680 18604 3692
rect 18656 3680 18662 3732
rect 20806 3680 20812 3732
rect 20864 3720 20870 3732
rect 20901 3723 20959 3729
rect 20901 3720 20913 3723
rect 20864 3692 20913 3720
rect 20864 3680 20870 3692
rect 20901 3689 20913 3692
rect 20947 3689 20959 3723
rect 20901 3683 20959 3689
rect 21634 3680 21640 3732
rect 21692 3720 21698 3732
rect 22741 3723 22799 3729
rect 22741 3720 22753 3723
rect 21692 3692 22753 3720
rect 21692 3680 21698 3692
rect 22741 3689 22753 3692
rect 22787 3689 22799 3723
rect 22741 3683 22799 3689
rect 12667 3624 17080 3652
rect 17396 3655 17454 3661
rect 12667 3621 12679 3624
rect 12621 3615 12679 3621
rect 17396 3621 17408 3655
rect 17442 3652 17454 3655
rect 17494 3652 17500 3664
rect 17442 3624 17500 3652
rect 17442 3621 17454 3624
rect 17396 3615 17454 3621
rect 17494 3612 17500 3624
rect 17552 3612 17558 3664
rect 17770 3612 17776 3664
rect 17828 3652 17834 3664
rect 20990 3652 20996 3664
rect 17828 3624 20996 3652
rect 17828 3612 17834 3624
rect 20990 3612 20996 3624
rect 21048 3612 21054 3664
rect 22278 3652 22284 3664
rect 21643 3624 22284 3652
rect 11606 3544 11612 3596
rect 11664 3584 11670 3596
rect 12526 3584 12532 3596
rect 11664 3556 11836 3584
rect 12487 3556 12532 3584
rect 11664 3544 11670 3556
rect 10686 3476 10692 3528
rect 10744 3516 10750 3528
rect 11698 3516 11704 3528
rect 10744 3488 11704 3516
rect 10744 3476 10750 3488
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 11808 3516 11836 3556
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 13998 3584 14004 3596
rect 12820 3556 14004 3584
rect 12820 3525 12848 3556
rect 13998 3544 14004 3556
rect 14056 3544 14062 3596
rect 14642 3584 14648 3596
rect 14603 3556 14648 3584
rect 14642 3544 14648 3556
rect 14700 3544 14706 3596
rect 15562 3584 15568 3596
rect 15523 3556 15568 3584
rect 15562 3544 15568 3556
rect 15620 3544 15626 3596
rect 16025 3587 16083 3593
rect 16025 3553 16037 3587
rect 16071 3584 16083 3587
rect 18506 3584 18512 3596
rect 16071 3556 18512 3584
rect 16071 3553 16083 3556
rect 16025 3547 16083 3553
rect 18506 3544 18512 3556
rect 18564 3544 18570 3596
rect 19242 3593 19248 3596
rect 19236 3547 19248 3593
rect 19300 3584 19306 3596
rect 19300 3556 19336 3584
rect 19242 3544 19248 3547
rect 19300 3544 19306 3556
rect 20346 3544 20352 3596
rect 20404 3584 20410 3596
rect 21643 3593 21671 3624
rect 22278 3612 22284 3624
rect 22336 3612 22342 3664
rect 21361 3587 21419 3593
rect 21361 3584 21373 3587
rect 20404 3556 21373 3584
rect 20404 3544 20410 3556
rect 21361 3553 21373 3556
rect 21407 3553 21419 3587
rect 21361 3547 21419 3553
rect 21628 3587 21686 3593
rect 21628 3553 21640 3587
rect 21674 3553 21686 3587
rect 21628 3547 21686 3553
rect 12805 3519 12863 3525
rect 12805 3516 12817 3519
rect 11808 3488 12817 3516
rect 12805 3485 12817 3488
rect 12851 3485 12863 3519
rect 13814 3516 13820 3528
rect 13775 3488 13820 3516
rect 12805 3479 12863 3485
rect 13814 3476 13820 3488
rect 13872 3476 13878 3528
rect 14826 3516 14832 3528
rect 14787 3488 14832 3516
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 15102 3476 15108 3528
rect 15160 3516 15166 3528
rect 16577 3519 16635 3525
rect 16577 3516 16589 3519
rect 15160 3488 16589 3516
rect 15160 3476 15166 3488
rect 16577 3485 16589 3488
rect 16623 3485 16635 3519
rect 16577 3479 16635 3485
rect 16669 3519 16727 3525
rect 16669 3485 16681 3519
rect 16715 3485 16727 3519
rect 16669 3479 16727 3485
rect 12158 3448 12164 3460
rect 12119 3420 12164 3448
rect 12158 3408 12164 3420
rect 12216 3408 12222 3460
rect 16025 3451 16083 3457
rect 16025 3448 16037 3451
rect 14016 3420 16037 3448
rect 7558 3340 7564 3392
rect 7616 3380 7622 3392
rect 13173 3383 13231 3389
rect 13173 3380 13185 3383
rect 7616 3352 13185 3380
rect 7616 3340 7622 3352
rect 13173 3349 13185 3352
rect 13219 3349 13231 3383
rect 13173 3343 13231 3349
rect 13262 3340 13268 3392
rect 13320 3380 13326 3392
rect 14016 3380 14044 3420
rect 16025 3417 16037 3420
rect 16071 3417 16083 3451
rect 16025 3411 16083 3417
rect 16298 3408 16304 3460
rect 16356 3448 16362 3460
rect 16684 3448 16712 3479
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17129 3519 17187 3525
rect 17129 3516 17141 3519
rect 17092 3488 17141 3516
rect 17092 3476 17098 3488
rect 17129 3485 17141 3488
rect 17175 3485 17187 3519
rect 17129 3479 17187 3485
rect 18138 3476 18144 3528
rect 18196 3516 18202 3528
rect 18966 3516 18972 3528
rect 18196 3488 18972 3516
rect 18196 3476 18202 3488
rect 18966 3476 18972 3488
rect 19024 3476 19030 3528
rect 16356 3420 16712 3448
rect 16356 3408 16362 3420
rect 18414 3408 18420 3460
rect 18472 3448 18478 3460
rect 18472 3420 19012 3448
rect 18472 3408 18478 3420
rect 13320 3352 14044 3380
rect 13320 3340 13326 3352
rect 15562 3340 15568 3392
rect 15620 3380 15626 3392
rect 15749 3383 15807 3389
rect 15749 3380 15761 3383
rect 15620 3352 15761 3380
rect 15620 3340 15626 3352
rect 15749 3349 15761 3352
rect 15795 3349 15807 3383
rect 15749 3343 15807 3349
rect 15933 3383 15991 3389
rect 15933 3349 15945 3383
rect 15979 3380 15991 3383
rect 17770 3380 17776 3392
rect 15979 3352 17776 3380
rect 15979 3349 15991 3352
rect 15933 3343 15991 3349
rect 17770 3340 17776 3352
rect 17828 3340 17834 3392
rect 18984 3380 19012 3420
rect 19150 3380 19156 3392
rect 18984 3352 19156 3380
rect 19150 3340 19156 3352
rect 19208 3380 19214 3392
rect 20349 3383 20407 3389
rect 20349 3380 20361 3383
rect 19208 3352 20361 3380
rect 19208 3340 19214 3352
rect 20349 3349 20361 3352
rect 20395 3349 20407 3383
rect 20349 3343 20407 3349
rect 20438 3340 20444 3392
rect 20496 3380 20502 3392
rect 21542 3380 21548 3392
rect 20496 3352 21548 3380
rect 20496 3340 20502 3352
rect 21542 3340 21548 3352
rect 21600 3340 21606 3392
rect 1104 3290 23276 3312
rect 1104 3238 4680 3290
rect 4732 3238 4744 3290
rect 4796 3238 4808 3290
rect 4860 3238 4872 3290
rect 4924 3238 12078 3290
rect 12130 3238 12142 3290
rect 12194 3238 12206 3290
rect 12258 3238 12270 3290
rect 12322 3238 19475 3290
rect 19527 3238 19539 3290
rect 19591 3238 19603 3290
rect 19655 3238 19667 3290
rect 19719 3238 23276 3290
rect 1104 3216 23276 3238
rect 13262 3176 13268 3188
rect 13223 3148 13268 3176
rect 13262 3136 13268 3148
rect 13320 3136 13326 3188
rect 14090 3176 14096 3188
rect 14051 3148 14096 3176
rect 14090 3136 14096 3148
rect 14148 3136 14154 3188
rect 14182 3136 14188 3188
rect 14240 3176 14246 3188
rect 15289 3179 15347 3185
rect 15289 3176 15301 3179
rect 14240 3148 15301 3176
rect 14240 3136 14246 3148
rect 15289 3145 15301 3148
rect 15335 3145 15347 3179
rect 15289 3139 15347 3145
rect 15378 3136 15384 3188
rect 15436 3176 15442 3188
rect 16117 3179 16175 3185
rect 15436 3148 15884 3176
rect 15436 3136 15442 3148
rect 2958 3068 2964 3120
rect 3016 3108 3022 3120
rect 3016 3080 15792 3108
rect 3016 3068 3022 3080
rect 1946 3040 1952 3052
rect 1907 3012 1952 3040
rect 1946 3000 1952 3012
rect 2004 3000 2010 3052
rect 11054 3040 11060 3052
rect 2516 3012 11060 3040
rect 1762 2972 1768 2984
rect 1723 2944 1768 2972
rect 1762 2932 1768 2944
rect 1820 2932 1826 2984
rect 2516 2981 2544 3012
rect 11054 3000 11060 3012
rect 11112 3040 11118 3052
rect 11974 3040 11980 3052
rect 11112 3012 11980 3040
rect 11112 3000 11118 3012
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 13909 3043 13967 3049
rect 13909 3009 13921 3043
rect 13955 3040 13967 3043
rect 13998 3040 14004 3052
rect 13955 3012 14004 3040
rect 13955 3009 13967 3012
rect 13909 3003 13967 3009
rect 13998 3000 14004 3012
rect 14056 3000 14062 3052
rect 14737 3043 14795 3049
rect 14737 3009 14749 3043
rect 14783 3040 14795 3043
rect 15010 3040 15016 3052
rect 14783 3012 15016 3040
rect 14783 3009 14795 3012
rect 14737 3003 14795 3009
rect 15010 3000 15016 3012
rect 15068 3000 15074 3052
rect 15764 3049 15792 3080
rect 15856 3049 15884 3148
rect 16117 3145 16129 3179
rect 16163 3176 16175 3179
rect 16482 3176 16488 3188
rect 16163 3148 16488 3176
rect 16163 3145 16175 3148
rect 16117 3139 16175 3145
rect 16482 3136 16488 3148
rect 16540 3136 16546 3188
rect 19150 3136 19156 3188
rect 19208 3136 19214 3188
rect 19242 3136 19248 3188
rect 19300 3176 19306 3188
rect 19613 3179 19671 3185
rect 19613 3176 19625 3179
rect 19300 3148 19625 3176
rect 19300 3136 19306 3148
rect 19613 3145 19625 3148
rect 19659 3145 19671 3179
rect 22097 3179 22155 3185
rect 19613 3139 19671 3145
rect 19720 3148 21680 3176
rect 19168 3108 19196 3136
rect 19720 3108 19748 3148
rect 19168 3080 19748 3108
rect 20346 3068 20352 3120
rect 20404 3108 20410 3120
rect 21652 3108 21680 3148
rect 22097 3145 22109 3179
rect 22143 3176 22155 3179
rect 22278 3176 22284 3188
rect 22143 3148 22284 3176
rect 22143 3145 22155 3148
rect 22097 3139 22155 3145
rect 22278 3136 22284 3148
rect 22336 3136 22342 3188
rect 22557 3111 22615 3117
rect 22557 3108 22569 3111
rect 20404 3080 20760 3108
rect 21652 3080 22569 3108
rect 20404 3068 20410 3080
rect 15749 3043 15807 3049
rect 15749 3009 15761 3043
rect 15795 3009 15807 3043
rect 15749 3003 15807 3009
rect 15841 3043 15899 3049
rect 15841 3009 15853 3043
rect 15887 3009 15899 3043
rect 15841 3003 15899 3009
rect 16040 3012 16436 3040
rect 2501 2975 2559 2981
rect 2501 2941 2513 2975
rect 2547 2941 2559 2975
rect 5074 2972 5080 2984
rect 5035 2944 5080 2972
rect 2501 2935 2559 2941
rect 5074 2932 5080 2944
rect 5132 2932 5138 2984
rect 13725 2975 13783 2981
rect 13725 2941 13737 2975
rect 13771 2972 13783 2975
rect 16040 2972 16068 3012
rect 13771 2944 16068 2972
rect 16301 2975 16359 2981
rect 13771 2941 13783 2944
rect 13725 2935 13783 2941
rect 16301 2941 16313 2975
rect 16347 2941 16359 2975
rect 16408 2972 16436 3012
rect 17310 3000 17316 3052
rect 17368 3040 17374 3052
rect 20438 3040 20444 3052
rect 17368 3012 18368 3040
rect 17368 3000 17374 3012
rect 16568 2975 16626 2981
rect 16568 2972 16580 2975
rect 16408 2944 16580 2972
rect 16301 2935 16359 2941
rect 16568 2941 16580 2944
rect 16614 2972 16626 2975
rect 17678 2972 17684 2984
rect 16614 2944 17684 2972
rect 16614 2941 16626 2944
rect 16568 2935 16626 2941
rect 13633 2907 13691 2913
rect 13633 2873 13645 2907
rect 13679 2904 13691 2907
rect 16316 2904 16344 2935
rect 17678 2932 17684 2944
rect 17736 2932 17742 2984
rect 18233 2975 18291 2981
rect 18233 2941 18245 2975
rect 18279 2941 18291 2975
rect 18340 2972 18368 3012
rect 19260 3012 20444 3040
rect 19260 2972 19288 3012
rect 20438 3000 20444 3012
rect 20496 3000 20502 3052
rect 20732 3049 20760 3080
rect 22557 3077 22569 3080
rect 22603 3077 22615 3111
rect 22557 3071 22615 3077
rect 20717 3043 20775 3049
rect 20717 3009 20729 3043
rect 20763 3009 20775 3043
rect 20717 3003 20775 3009
rect 18340 2944 19288 2972
rect 19981 2975 20039 2981
rect 18233 2935 18291 2941
rect 19981 2941 19993 2975
rect 20027 2972 20039 2975
rect 21450 2972 21456 2984
rect 20027 2944 21456 2972
rect 20027 2941 20039 2944
rect 19981 2935 20039 2941
rect 17034 2904 17040 2916
rect 13679 2876 16252 2904
rect 16316 2876 17040 2904
rect 13679 2873 13691 2876
rect 13633 2867 13691 2873
rect 1670 2796 1676 2848
rect 1728 2836 1734 2848
rect 2685 2839 2743 2845
rect 2685 2836 2697 2839
rect 1728 2808 2697 2836
rect 1728 2796 1734 2808
rect 2685 2805 2697 2808
rect 2731 2805 2743 2839
rect 2685 2799 2743 2805
rect 14366 2796 14372 2848
rect 14424 2836 14430 2848
rect 14461 2839 14519 2845
rect 14461 2836 14473 2839
rect 14424 2808 14473 2836
rect 14424 2796 14430 2808
rect 14461 2805 14473 2808
rect 14507 2805 14519 2839
rect 14461 2799 14519 2805
rect 14553 2839 14611 2845
rect 14553 2805 14565 2839
rect 14599 2836 14611 2839
rect 15102 2836 15108 2848
rect 14599 2808 15108 2836
rect 14599 2805 14611 2808
rect 14553 2799 14611 2805
rect 15102 2796 15108 2808
rect 15160 2796 15166 2848
rect 15197 2839 15255 2845
rect 15197 2805 15209 2839
rect 15243 2836 15255 2839
rect 15657 2839 15715 2845
rect 15657 2836 15669 2839
rect 15243 2808 15669 2836
rect 15243 2805 15255 2808
rect 15197 2799 15255 2805
rect 15657 2805 15669 2808
rect 15703 2836 15715 2839
rect 16117 2839 16175 2845
rect 16117 2836 16129 2839
rect 15703 2808 16129 2836
rect 15703 2805 15715 2808
rect 15657 2799 15715 2805
rect 16117 2805 16129 2808
rect 16163 2805 16175 2839
rect 16224 2836 16252 2876
rect 17034 2864 17040 2876
rect 17092 2904 17098 2916
rect 18138 2904 18144 2916
rect 17092 2876 18144 2904
rect 17092 2864 17098 2876
rect 18138 2864 18144 2876
rect 18196 2904 18202 2916
rect 18248 2904 18276 2935
rect 21450 2932 21456 2944
rect 21508 2972 21514 2984
rect 22373 2975 22431 2981
rect 22373 2972 22385 2975
rect 21508 2944 22385 2972
rect 21508 2932 21514 2944
rect 22373 2941 22385 2944
rect 22419 2941 22431 2975
rect 22373 2935 22431 2941
rect 18196 2876 18276 2904
rect 18196 2864 18202 2876
rect 18322 2864 18328 2916
rect 18380 2904 18386 2916
rect 18478 2907 18536 2913
rect 18478 2904 18490 2907
rect 18380 2876 18490 2904
rect 18380 2864 18386 2876
rect 18478 2873 18490 2876
rect 18524 2873 18536 2907
rect 18478 2867 18536 2873
rect 20257 2907 20315 2913
rect 20257 2873 20269 2907
rect 20303 2873 20315 2907
rect 20257 2867 20315 2873
rect 17494 2836 17500 2848
rect 16224 2808 17500 2836
rect 16117 2799 16175 2805
rect 17494 2796 17500 2808
rect 17552 2836 17558 2848
rect 17681 2839 17739 2845
rect 17681 2836 17693 2839
rect 17552 2808 17693 2836
rect 17552 2796 17558 2808
rect 17681 2805 17693 2808
rect 17727 2805 17739 2839
rect 17681 2799 17739 2805
rect 18046 2796 18052 2848
rect 18104 2836 18110 2848
rect 20070 2836 20076 2848
rect 18104 2808 20076 2836
rect 18104 2796 18110 2808
rect 20070 2796 20076 2808
rect 20128 2796 20134 2848
rect 20272 2836 20300 2867
rect 20898 2864 20904 2916
rect 20956 2913 20962 2916
rect 20956 2907 21020 2913
rect 20956 2873 20974 2907
rect 21008 2873 21020 2907
rect 20956 2867 21020 2873
rect 20956 2864 20962 2867
rect 22554 2836 22560 2848
rect 20272 2808 22560 2836
rect 22554 2796 22560 2808
rect 22612 2796 22618 2848
rect 1104 2746 23276 2768
rect 1104 2694 8379 2746
rect 8431 2694 8443 2746
rect 8495 2694 8507 2746
rect 8559 2694 8571 2746
rect 8623 2694 15776 2746
rect 15828 2694 15840 2746
rect 15892 2694 15904 2746
rect 15956 2694 15968 2746
rect 16020 2694 23276 2746
rect 1104 2672 23276 2694
rect 13725 2635 13783 2641
rect 13725 2601 13737 2635
rect 13771 2632 13783 2635
rect 13906 2632 13912 2644
rect 13771 2604 13912 2632
rect 13771 2601 13783 2604
rect 13725 2595 13783 2601
rect 13906 2592 13912 2604
rect 13964 2592 13970 2644
rect 14829 2635 14887 2641
rect 14829 2601 14841 2635
rect 14875 2632 14887 2635
rect 15654 2632 15660 2644
rect 14875 2604 15660 2632
rect 14875 2601 14887 2604
rect 14829 2595 14887 2601
rect 15654 2592 15660 2604
rect 15712 2592 15718 2644
rect 16577 2635 16635 2641
rect 16577 2601 16589 2635
rect 16623 2632 16635 2635
rect 17494 2632 17500 2644
rect 16623 2604 17500 2632
rect 16623 2601 16635 2604
rect 16577 2595 16635 2601
rect 17494 2592 17500 2604
rect 17552 2592 17558 2644
rect 18322 2592 18328 2644
rect 18380 2632 18386 2644
rect 19705 2635 19763 2641
rect 19705 2632 19717 2635
rect 18380 2604 19717 2632
rect 18380 2592 18386 2604
rect 19705 2601 19717 2604
rect 19751 2601 19763 2635
rect 19705 2595 19763 2601
rect 19978 2592 19984 2644
rect 20036 2632 20042 2644
rect 20441 2635 20499 2641
rect 20441 2632 20453 2635
rect 20036 2604 20453 2632
rect 20036 2592 20042 2604
rect 20441 2601 20453 2604
rect 20487 2601 20499 2635
rect 20441 2595 20499 2601
rect 20533 2635 20591 2641
rect 20533 2601 20545 2635
rect 20579 2632 20591 2635
rect 20622 2632 20628 2644
rect 20579 2604 20628 2632
rect 20579 2601 20591 2604
rect 20533 2595 20591 2601
rect 20622 2592 20628 2604
rect 20680 2592 20686 2644
rect 22557 2635 22615 2641
rect 22557 2601 22569 2635
rect 22603 2601 22615 2635
rect 22557 2595 22615 2601
rect 11698 2524 11704 2576
rect 11756 2564 11762 2576
rect 14737 2567 14795 2573
rect 11756 2536 13952 2564
rect 11756 2524 11762 2536
rect 13924 2437 13952 2536
rect 14737 2533 14749 2567
rect 14783 2564 14795 2567
rect 16482 2564 16488 2576
rect 14783 2536 16488 2564
rect 14783 2533 14795 2536
rect 14737 2527 14795 2533
rect 16482 2524 16488 2536
rect 16540 2524 16546 2576
rect 16669 2567 16727 2573
rect 16669 2533 16681 2567
rect 16715 2564 16727 2567
rect 16758 2564 16764 2576
rect 16715 2536 16764 2564
rect 16715 2533 16727 2536
rect 16669 2527 16727 2533
rect 16758 2524 16764 2536
rect 16816 2524 16822 2576
rect 17589 2567 17647 2573
rect 17589 2564 17601 2567
rect 17512 2536 17601 2564
rect 13998 2456 14004 2508
rect 14056 2496 14062 2508
rect 14056 2468 15056 2496
rect 14056 2456 14062 2468
rect 15028 2437 15056 2468
rect 17402 2456 17408 2508
rect 17460 2496 17466 2508
rect 17512 2496 17540 2536
rect 17589 2533 17601 2536
rect 17635 2533 17647 2567
rect 17589 2527 17647 2533
rect 17678 2524 17684 2576
rect 17736 2564 17742 2576
rect 18414 2564 18420 2576
rect 17736 2536 18420 2564
rect 17736 2524 17742 2536
rect 18414 2524 18420 2536
rect 18472 2524 18478 2576
rect 18598 2573 18604 2576
rect 18592 2564 18604 2573
rect 18559 2536 18604 2564
rect 18592 2527 18604 2536
rect 18598 2524 18604 2527
rect 18656 2524 18662 2576
rect 20898 2524 20904 2576
rect 20956 2564 20962 2576
rect 22572 2564 22600 2595
rect 20956 2536 22600 2564
rect 20956 2524 20962 2536
rect 17460 2468 17540 2496
rect 17604 2468 17908 2496
rect 17460 2456 17466 2468
rect 13817 2431 13875 2437
rect 13817 2397 13829 2431
rect 13863 2397 13875 2431
rect 13817 2391 13875 2397
rect 13909 2431 13967 2437
rect 13909 2397 13921 2431
rect 13955 2397 13967 2431
rect 15013 2431 15071 2437
rect 13909 2391 13967 2397
rect 14016 2400 14780 2428
rect 13832 2360 13860 2391
rect 14016 2360 14044 2400
rect 14366 2360 14372 2372
rect 13832 2332 14044 2360
rect 14327 2332 14372 2360
rect 14366 2320 14372 2332
rect 14424 2320 14430 2372
rect 14752 2360 14780 2400
rect 15013 2397 15025 2431
rect 15059 2428 15071 2431
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 15059 2400 16865 2428
rect 15059 2397 15071 2400
rect 15013 2391 15071 2397
rect 16853 2397 16865 2400
rect 16899 2428 16911 2431
rect 17604 2428 17632 2468
rect 17880 2437 17908 2468
rect 18138 2456 18144 2508
rect 18196 2496 18202 2508
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 18196 2468 18337 2496
rect 18196 2456 18202 2468
rect 18325 2465 18337 2468
rect 18371 2465 18383 2499
rect 19334 2496 19340 2508
rect 18325 2459 18383 2465
rect 18432 2468 19340 2496
rect 16899 2400 17632 2428
rect 17681 2431 17739 2437
rect 16899 2397 16911 2400
rect 16853 2391 16911 2397
rect 17681 2397 17693 2431
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 17865 2431 17923 2437
rect 17865 2397 17877 2431
rect 17911 2428 17923 2431
rect 18046 2428 18052 2440
rect 17911 2400 18052 2428
rect 17911 2397 17923 2400
rect 17865 2391 17923 2397
rect 16114 2360 16120 2372
rect 14752 2332 16120 2360
rect 16114 2320 16120 2332
rect 16172 2320 16178 2372
rect 17494 2320 17500 2372
rect 17552 2360 17558 2372
rect 17696 2360 17724 2391
rect 18046 2388 18052 2400
rect 18104 2388 18110 2440
rect 18432 2428 18460 2468
rect 19334 2456 19340 2468
rect 19392 2456 19398 2508
rect 20346 2456 20352 2508
rect 20404 2496 20410 2508
rect 21177 2499 21235 2505
rect 21177 2496 21189 2499
rect 20404 2468 21189 2496
rect 20404 2456 20410 2468
rect 21177 2465 21189 2468
rect 21223 2465 21235 2499
rect 21177 2459 21235 2465
rect 21266 2456 21272 2508
rect 21324 2496 21330 2508
rect 21433 2499 21491 2505
rect 21433 2496 21445 2499
rect 21324 2468 21445 2496
rect 21324 2456 21330 2468
rect 21433 2465 21445 2468
rect 21479 2465 21491 2499
rect 21433 2459 21491 2465
rect 18248 2400 18460 2428
rect 20625 2431 20683 2437
rect 18248 2360 18276 2400
rect 20625 2397 20637 2431
rect 20671 2428 20683 2431
rect 21082 2428 21088 2440
rect 20671 2400 21088 2428
rect 20671 2397 20683 2400
rect 20625 2391 20683 2397
rect 21082 2388 21088 2400
rect 21140 2388 21146 2440
rect 17552 2332 17724 2360
rect 17788 2332 18276 2360
rect 17552 2320 17558 2332
rect 13357 2295 13415 2301
rect 13357 2261 13369 2295
rect 13403 2292 13415 2295
rect 15470 2292 15476 2304
rect 13403 2264 15476 2292
rect 13403 2261 13415 2264
rect 13357 2255 13415 2261
rect 15470 2252 15476 2264
rect 15528 2252 15534 2304
rect 16209 2295 16267 2301
rect 16209 2261 16221 2295
rect 16255 2292 16267 2295
rect 16298 2292 16304 2304
rect 16255 2264 16304 2292
rect 16255 2261 16267 2264
rect 16209 2255 16267 2261
rect 16298 2252 16304 2264
rect 16356 2252 16362 2304
rect 17221 2295 17279 2301
rect 17221 2261 17233 2295
rect 17267 2292 17279 2295
rect 17788 2292 17816 2332
rect 17267 2264 17816 2292
rect 17267 2261 17279 2264
rect 17221 2255 17279 2261
rect 17862 2252 17868 2304
rect 17920 2292 17926 2304
rect 20073 2295 20131 2301
rect 20073 2292 20085 2295
rect 17920 2264 20085 2292
rect 17920 2252 17926 2264
rect 20073 2261 20085 2264
rect 20119 2261 20131 2295
rect 20073 2255 20131 2261
rect 1104 2202 23276 2224
rect 1104 2150 4680 2202
rect 4732 2150 4744 2202
rect 4796 2150 4808 2202
rect 4860 2150 4872 2202
rect 4924 2150 12078 2202
rect 12130 2150 12142 2202
rect 12194 2150 12206 2202
rect 12258 2150 12270 2202
rect 12322 2150 19475 2202
rect 19527 2150 19539 2202
rect 19591 2150 19603 2202
rect 19655 2150 19667 2202
rect 19719 2150 23276 2202
rect 1104 2128 23276 2150
rect 16758 2048 16764 2100
rect 16816 2088 16822 2100
rect 19242 2088 19248 2100
rect 16816 2060 19248 2088
rect 16816 2048 16822 2060
rect 19242 2048 19248 2060
rect 19300 2048 19306 2100
rect 14366 1980 14372 2032
rect 14424 2020 14430 2032
rect 17218 2020 17224 2032
rect 14424 1992 17224 2020
rect 14424 1980 14430 1992
rect 17218 1980 17224 1992
rect 17276 1980 17282 2032
rect 17402 1980 17408 2032
rect 17460 2020 17466 2032
rect 20898 2020 20904 2032
rect 17460 1992 20904 2020
rect 17460 1980 17466 1992
rect 20898 1980 20904 1992
rect 20956 1980 20962 2032
rect 17494 1912 17500 1964
rect 17552 1952 17558 1964
rect 21266 1952 21272 1964
rect 17552 1924 21272 1952
rect 17552 1912 17558 1924
rect 21266 1912 21272 1924
rect 21324 1912 21330 1964
rect 16298 1844 16304 1896
rect 16356 1884 16362 1896
rect 18230 1884 18236 1896
rect 16356 1856 18236 1884
rect 16356 1844 16362 1856
rect 18230 1844 18236 1856
rect 18288 1844 18294 1896
rect 15194 1776 15200 1828
rect 15252 1816 15258 1828
rect 19886 1816 19892 1828
rect 15252 1788 19892 1816
rect 15252 1776 15258 1788
rect 19886 1776 19892 1788
rect 19944 1776 19950 1828
rect 16390 1300 16396 1352
rect 16448 1340 16454 1352
rect 19334 1340 19340 1352
rect 16448 1312 19340 1340
rect 16448 1300 16454 1312
rect 19334 1300 19340 1312
rect 19392 1300 19398 1352
<< via1 >>
rect 7564 21972 7616 22024
rect 16672 21972 16724 22024
rect 9956 21904 10008 21956
rect 16948 21904 17000 21956
rect 18696 21904 18748 21956
rect 19524 21904 19576 21956
rect 18328 21836 18380 21888
rect 20076 21836 20128 21888
rect 4680 21734 4732 21786
rect 4744 21734 4796 21786
rect 4808 21734 4860 21786
rect 4872 21734 4924 21786
rect 12078 21734 12130 21786
rect 12142 21734 12194 21786
rect 12206 21734 12258 21786
rect 12270 21734 12322 21786
rect 19475 21734 19527 21786
rect 19539 21734 19591 21786
rect 19603 21734 19655 21786
rect 19667 21734 19719 21786
rect 1492 21632 1544 21684
rect 8116 21632 8168 21684
rect 8576 21632 8628 21684
rect 9956 21675 10008 21684
rect 9956 21641 9965 21675
rect 9965 21641 9999 21675
rect 9999 21641 10008 21675
rect 9956 21632 10008 21641
rect 14740 21632 14792 21684
rect 19800 21632 19852 21684
rect 7564 21564 7616 21616
rect 16764 21564 16816 21616
rect 5540 21496 5592 21548
rect 14188 21539 14240 21548
rect 14188 21505 14197 21539
rect 14197 21505 14231 21539
rect 14231 21505 14240 21539
rect 14188 21496 14240 21505
rect 2688 21360 2740 21412
rect 4160 21428 4212 21480
rect 9128 21428 9180 21480
rect 10416 21428 10468 21480
rect 12164 21428 12216 21480
rect 15568 21428 15620 21480
rect 16120 21539 16172 21548
rect 16120 21505 16129 21539
rect 16129 21505 16163 21539
rect 16163 21505 16172 21539
rect 16120 21496 16172 21505
rect 16488 21496 16540 21548
rect 17684 21564 17736 21616
rect 21916 21564 21968 21616
rect 18604 21496 18656 21548
rect 21824 21539 21876 21548
rect 21824 21505 21833 21539
rect 21833 21505 21867 21539
rect 21867 21505 21876 21539
rect 21824 21496 21876 21505
rect 18328 21471 18380 21480
rect 18328 21437 18337 21471
rect 18337 21437 18371 21471
rect 18371 21437 18380 21471
rect 18328 21428 18380 21437
rect 18880 21471 18932 21480
rect 18880 21437 18889 21471
rect 18889 21437 18923 21471
rect 18923 21437 18932 21471
rect 18880 21428 18932 21437
rect 6092 21360 6144 21412
rect 6460 21360 6512 21412
rect 7012 21360 7064 21412
rect 8852 21403 8904 21412
rect 8852 21369 8861 21403
rect 8861 21369 8895 21403
rect 8895 21369 8904 21403
rect 8852 21360 8904 21369
rect 11796 21360 11848 21412
rect 14464 21360 14516 21412
rect 19892 21428 19944 21480
rect 20536 21471 20588 21480
rect 20536 21437 20545 21471
rect 20545 21437 20579 21471
rect 20579 21437 20588 21471
rect 20536 21428 20588 21437
rect 22192 21471 22244 21480
rect 22192 21437 22201 21471
rect 22201 21437 22235 21471
rect 22235 21437 22244 21471
rect 22192 21428 22244 21437
rect 1952 21335 2004 21344
rect 1952 21301 1961 21335
rect 1961 21301 1995 21335
rect 1995 21301 2004 21335
rect 1952 21292 2004 21301
rect 2412 21335 2464 21344
rect 2412 21301 2421 21335
rect 2421 21301 2455 21335
rect 2455 21301 2464 21335
rect 2964 21335 3016 21344
rect 2412 21292 2464 21301
rect 2964 21301 2973 21335
rect 2973 21301 3007 21335
rect 3007 21301 3016 21335
rect 2964 21292 3016 21301
rect 3332 21335 3384 21344
rect 3332 21301 3341 21335
rect 3341 21301 3375 21335
rect 3375 21301 3384 21335
rect 3332 21292 3384 21301
rect 3424 21335 3476 21344
rect 3424 21301 3433 21335
rect 3433 21301 3467 21335
rect 3467 21301 3476 21335
rect 4068 21335 4120 21344
rect 3424 21292 3476 21301
rect 4068 21301 4077 21335
rect 4077 21301 4111 21335
rect 4111 21301 4120 21335
rect 4068 21292 4120 21301
rect 4436 21335 4488 21344
rect 4436 21301 4445 21335
rect 4445 21301 4479 21335
rect 4479 21301 4488 21335
rect 4436 21292 4488 21301
rect 4528 21335 4580 21344
rect 4528 21301 4537 21335
rect 4537 21301 4571 21335
rect 4571 21301 4580 21335
rect 5264 21335 5316 21344
rect 4528 21292 4580 21301
rect 5264 21301 5273 21335
rect 5273 21301 5307 21335
rect 5307 21301 5316 21335
rect 5264 21292 5316 21301
rect 5816 21335 5868 21344
rect 5816 21301 5825 21335
rect 5825 21301 5859 21335
rect 5859 21301 5868 21335
rect 5816 21292 5868 21301
rect 6276 21335 6328 21344
rect 6276 21301 6285 21335
rect 6285 21301 6319 21335
rect 6319 21301 6328 21335
rect 6276 21292 6328 21301
rect 6920 21335 6972 21344
rect 6920 21301 6929 21335
rect 6929 21301 6963 21335
rect 6963 21301 6972 21335
rect 6920 21292 6972 21301
rect 7288 21335 7340 21344
rect 7288 21301 7297 21335
rect 7297 21301 7331 21335
rect 7331 21301 7340 21335
rect 7288 21292 7340 21301
rect 7380 21335 7432 21344
rect 7380 21301 7389 21335
rect 7389 21301 7423 21335
rect 7423 21301 7432 21335
rect 7380 21292 7432 21301
rect 8668 21292 8720 21344
rect 8760 21335 8812 21344
rect 8760 21301 8769 21335
rect 8769 21301 8803 21335
rect 8803 21301 8812 21335
rect 12072 21335 12124 21344
rect 8760 21292 8812 21301
rect 12072 21301 12081 21335
rect 12081 21301 12115 21335
rect 12115 21301 12124 21335
rect 12072 21292 12124 21301
rect 12900 21292 12952 21344
rect 13728 21292 13780 21344
rect 19340 21360 19392 21412
rect 15108 21292 15160 21344
rect 16304 21292 16356 21344
rect 16856 21335 16908 21344
rect 16856 21301 16865 21335
rect 16865 21301 16899 21335
rect 16899 21301 16908 21335
rect 16856 21292 16908 21301
rect 16948 21335 17000 21344
rect 16948 21301 16957 21335
rect 16957 21301 16991 21335
rect 16991 21301 17000 21335
rect 16948 21292 17000 21301
rect 19248 21292 19300 21344
rect 20260 21335 20312 21344
rect 20260 21301 20269 21335
rect 20269 21301 20303 21335
rect 20303 21301 20312 21335
rect 20260 21292 20312 21301
rect 21088 21292 21140 21344
rect 21548 21335 21600 21344
rect 21548 21301 21557 21335
rect 21557 21301 21591 21335
rect 21591 21301 21600 21335
rect 21548 21292 21600 21301
rect 21640 21335 21692 21344
rect 21640 21301 21649 21335
rect 21649 21301 21683 21335
rect 21683 21301 21692 21335
rect 21640 21292 21692 21301
rect 22284 21292 22336 21344
rect 8379 21190 8431 21242
rect 8443 21190 8495 21242
rect 8507 21190 8559 21242
rect 8571 21190 8623 21242
rect 15776 21190 15828 21242
rect 15840 21190 15892 21242
rect 15904 21190 15956 21242
rect 15968 21190 16020 21242
rect 296 21088 348 21140
rect 4068 21088 4120 21140
rect 7380 21088 7432 21140
rect 8852 21088 8904 21140
rect 11520 21088 11572 21140
rect 16948 21088 17000 21140
rect 19156 21088 19208 21140
rect 2964 21020 3016 21072
rect 3424 20952 3476 21004
rect 1768 20884 1820 20936
rect 4344 20884 4396 20936
rect 5448 21020 5500 21072
rect 5172 20952 5224 21004
rect 7288 21020 7340 21072
rect 8208 21020 8260 21072
rect 8668 21020 8720 21072
rect 12072 21020 12124 21072
rect 6460 20952 6512 21004
rect 6828 20952 6880 21004
rect 10048 20995 10100 21004
rect 7564 20927 7616 20936
rect 3884 20816 3936 20868
rect 3332 20791 3384 20800
rect 3332 20757 3341 20791
rect 3341 20757 3375 20791
rect 3375 20757 3384 20791
rect 3332 20748 3384 20757
rect 3976 20748 4028 20800
rect 5080 20748 5132 20800
rect 7564 20893 7573 20927
rect 7573 20893 7607 20927
rect 7607 20893 7616 20927
rect 7564 20884 7616 20893
rect 10048 20961 10057 20995
rect 10057 20961 10091 20995
rect 10091 20961 10100 20995
rect 10048 20952 10100 20961
rect 13176 20952 13228 21004
rect 13728 21020 13780 21072
rect 13820 20952 13872 21004
rect 14648 20952 14700 21004
rect 18052 21020 18104 21072
rect 18880 21020 18932 21072
rect 20260 21020 20312 21072
rect 10416 20884 10468 20936
rect 15292 20927 15344 20936
rect 15292 20893 15301 20927
rect 15301 20893 15335 20927
rect 15335 20893 15344 20927
rect 15292 20884 15344 20893
rect 6552 20748 6604 20800
rect 9772 20748 9824 20800
rect 12440 20791 12492 20800
rect 12440 20757 12449 20791
rect 12449 20757 12483 20791
rect 12483 20757 12492 20791
rect 14464 20791 14516 20800
rect 12440 20748 12492 20757
rect 14464 20757 14473 20791
rect 14473 20757 14507 20791
rect 14507 20757 14516 20791
rect 14464 20748 14516 20757
rect 14556 20748 14608 20800
rect 15108 20748 15160 20800
rect 15200 20748 15252 20800
rect 19800 20952 19852 21004
rect 21640 21020 21692 21072
rect 20904 20927 20956 20936
rect 20904 20893 20913 20927
rect 20913 20893 20947 20927
rect 20947 20893 20956 20927
rect 20904 20884 20956 20893
rect 17776 20748 17828 20800
rect 19340 20748 19392 20800
rect 20168 20748 20220 20800
rect 21548 20748 21600 20800
rect 4680 20646 4732 20698
rect 4744 20646 4796 20698
rect 4808 20646 4860 20698
rect 4872 20646 4924 20698
rect 12078 20646 12130 20698
rect 12142 20646 12194 20698
rect 12206 20646 12258 20698
rect 12270 20646 12322 20698
rect 19475 20646 19527 20698
rect 19539 20646 19591 20698
rect 19603 20646 19655 20698
rect 19667 20646 19719 20698
rect 3424 20544 3476 20596
rect 4436 20544 4488 20596
rect 6460 20587 6512 20596
rect 6460 20553 6469 20587
rect 6469 20553 6503 20587
rect 6503 20553 6512 20587
rect 6460 20544 6512 20553
rect 6552 20544 6604 20596
rect 5080 20451 5132 20460
rect 5080 20417 5089 20451
rect 5089 20417 5123 20451
rect 5123 20417 5132 20451
rect 5080 20408 5132 20417
rect 7564 20544 7616 20596
rect 8208 20587 8260 20596
rect 8208 20553 8217 20587
rect 8217 20553 8251 20587
rect 8251 20553 8260 20587
rect 8208 20544 8260 20553
rect 8760 20544 8812 20596
rect 11796 20587 11848 20596
rect 9496 20476 9548 20528
rect 11796 20553 11805 20587
rect 11805 20553 11839 20587
rect 11839 20553 11848 20587
rect 11796 20544 11848 20553
rect 14648 20587 14700 20596
rect 13084 20476 13136 20528
rect 14648 20553 14657 20587
rect 14657 20553 14691 20587
rect 14691 20553 14700 20587
rect 14648 20544 14700 20553
rect 19064 20544 19116 20596
rect 19800 20544 19852 20596
rect 16212 20476 16264 20528
rect 11428 20408 11480 20460
rect 1768 20340 1820 20392
rect 3424 20383 3476 20392
rect 3424 20349 3433 20383
rect 3433 20349 3467 20383
rect 3467 20349 3476 20383
rect 3424 20340 3476 20349
rect 4528 20340 4580 20392
rect 6276 20340 6328 20392
rect 7380 20340 7432 20392
rect 8024 20340 8076 20392
rect 10416 20383 10468 20392
rect 10416 20349 10425 20383
rect 10425 20349 10459 20383
rect 10459 20349 10468 20383
rect 10416 20340 10468 20349
rect 11980 20340 12032 20392
rect 2044 20272 2096 20324
rect 4252 20272 4304 20324
rect 6644 20272 6696 20324
rect 8852 20272 8904 20324
rect 9036 20272 9088 20324
rect 11336 20272 11388 20324
rect 11428 20272 11480 20324
rect 12532 20272 12584 20324
rect 13176 20340 13228 20392
rect 16120 20408 16172 20460
rect 16580 20408 16632 20460
rect 16764 20408 16816 20460
rect 21824 20544 21876 20596
rect 20168 20451 20220 20460
rect 20168 20417 20177 20451
rect 20177 20417 20211 20451
rect 20211 20417 20220 20451
rect 20168 20408 20220 20417
rect 20352 20451 20404 20460
rect 20352 20417 20361 20451
rect 20361 20417 20395 20451
rect 20395 20417 20404 20451
rect 20352 20408 20404 20417
rect 13360 20272 13412 20324
rect 14464 20340 14516 20392
rect 15200 20383 15252 20392
rect 15200 20349 15234 20383
rect 15234 20349 15252 20383
rect 15200 20340 15252 20349
rect 18052 20383 18104 20392
rect 15476 20272 15528 20324
rect 18052 20349 18061 20383
rect 18061 20349 18095 20383
rect 18095 20349 18104 20383
rect 18052 20340 18104 20349
rect 19156 20272 19208 20324
rect 848 20204 900 20256
rect 5264 20204 5316 20256
rect 5448 20204 5500 20256
rect 12164 20204 12216 20256
rect 12256 20204 12308 20256
rect 12716 20204 12768 20256
rect 12808 20204 12860 20256
rect 13176 20204 13228 20256
rect 15292 20204 15344 20256
rect 16304 20247 16356 20256
rect 16304 20213 16313 20247
rect 16313 20213 16347 20247
rect 16347 20213 16356 20247
rect 16304 20204 16356 20213
rect 17040 20204 17092 20256
rect 17224 20204 17276 20256
rect 19984 20272 20036 20324
rect 20260 20272 20312 20324
rect 20904 20340 20956 20392
rect 21548 20340 21600 20392
rect 22560 20340 22612 20392
rect 21456 20272 21508 20324
rect 20168 20204 20220 20256
rect 20444 20204 20496 20256
rect 24032 20272 24084 20324
rect 21732 20204 21784 20256
rect 22928 20204 22980 20256
rect 8379 20102 8431 20154
rect 8443 20102 8495 20154
rect 8507 20102 8559 20154
rect 8571 20102 8623 20154
rect 15776 20102 15828 20154
rect 15840 20102 15892 20154
rect 15904 20102 15956 20154
rect 15968 20102 16020 20154
rect 2136 20000 2188 20052
rect 4160 20000 4212 20052
rect 1768 19932 1820 19984
rect 3792 19932 3844 19984
rect 4436 19932 4488 19984
rect 4988 20000 5040 20052
rect 5448 20000 5500 20052
rect 6920 20000 6972 20052
rect 9220 20000 9272 20052
rect 9864 20000 9916 20052
rect 11980 20000 12032 20052
rect 13728 20000 13780 20052
rect 13820 20000 13872 20052
rect 2780 19864 2832 19916
rect 1400 19839 1452 19848
rect 1400 19805 1409 19839
rect 1409 19805 1443 19839
rect 1443 19805 1452 19839
rect 1400 19796 1452 19805
rect 3424 19864 3476 19916
rect 4068 19796 4120 19848
rect 5080 19864 5132 19916
rect 5816 19932 5868 19984
rect 8024 19864 8076 19916
rect 8208 19907 8260 19916
rect 8208 19873 8242 19907
rect 8242 19873 8260 19907
rect 8208 19864 8260 19873
rect 5448 19796 5500 19848
rect 6828 19839 6880 19848
rect 6276 19728 6328 19780
rect 6828 19805 6837 19839
rect 6837 19805 6871 19839
rect 6871 19805 6880 19839
rect 6828 19796 6880 19805
rect 7656 19728 7708 19780
rect 9864 19907 9916 19916
rect 9864 19873 9873 19907
rect 9873 19873 9907 19907
rect 9907 19873 9916 19907
rect 9864 19864 9916 19873
rect 10416 19839 10468 19848
rect 10416 19805 10425 19839
rect 10425 19805 10459 19839
rect 10459 19805 10468 19839
rect 12164 19932 12216 19984
rect 16304 19932 16356 19984
rect 17408 20000 17460 20052
rect 18788 20000 18840 20052
rect 19156 20043 19208 20052
rect 19156 20009 19165 20043
rect 19165 20009 19199 20043
rect 19199 20009 19208 20043
rect 19156 20000 19208 20009
rect 18696 19932 18748 19984
rect 19800 19975 19852 19984
rect 19800 19941 19809 19975
rect 19809 19941 19843 19975
rect 19843 19941 19852 19975
rect 19800 19932 19852 19941
rect 10692 19907 10744 19916
rect 10692 19873 10726 19907
rect 10726 19873 10744 19907
rect 10692 19864 10744 19873
rect 11980 19864 12032 19916
rect 12348 19907 12400 19916
rect 12348 19873 12382 19907
rect 12382 19873 12400 19907
rect 12348 19864 12400 19873
rect 15016 19864 15068 19916
rect 17868 19864 17920 19916
rect 18880 19864 18932 19916
rect 14188 19839 14240 19848
rect 10416 19796 10468 19805
rect 14188 19805 14197 19839
rect 14197 19805 14231 19839
rect 14231 19805 14240 19839
rect 14188 19796 14240 19805
rect 14832 19796 14884 19848
rect 15292 19796 15344 19848
rect 18788 19796 18840 19848
rect 20812 19864 20864 19916
rect 21640 19907 21692 19916
rect 21640 19873 21649 19907
rect 21649 19873 21683 19907
rect 21683 19873 21692 19907
rect 21640 19864 21692 19873
rect 22008 19864 22060 19916
rect 22468 19907 22520 19916
rect 22468 19873 22477 19907
rect 22477 19873 22511 19907
rect 22511 19873 22520 19907
rect 22468 19864 22520 19873
rect 19800 19796 19852 19848
rect 20352 19796 20404 19848
rect 21732 19839 21784 19848
rect 21732 19805 21741 19839
rect 21741 19805 21775 19839
rect 21775 19805 21784 19839
rect 21732 19796 21784 19805
rect 21824 19839 21876 19848
rect 21824 19805 21833 19839
rect 21833 19805 21867 19839
rect 21867 19805 21876 19839
rect 21824 19796 21876 19805
rect 2044 19660 2096 19712
rect 5080 19660 5132 19712
rect 6000 19660 6052 19712
rect 7564 19703 7616 19712
rect 7564 19669 7573 19703
rect 7573 19669 7607 19703
rect 7607 19669 7616 19703
rect 7564 19660 7616 19669
rect 8300 19660 8352 19712
rect 9680 19660 9732 19712
rect 12072 19728 12124 19780
rect 11888 19660 11940 19712
rect 12440 19660 12492 19712
rect 12716 19660 12768 19712
rect 13544 19703 13596 19712
rect 13544 19669 13553 19703
rect 13553 19669 13587 19703
rect 13587 19669 13596 19703
rect 14924 19728 14976 19780
rect 17224 19728 17276 19780
rect 13544 19660 13596 19669
rect 16396 19660 16448 19712
rect 16672 19660 16724 19712
rect 17132 19660 17184 19712
rect 17960 19660 18012 19712
rect 19892 19728 19944 19780
rect 19248 19660 19300 19712
rect 21364 19660 21416 19712
rect 22652 19703 22704 19712
rect 22652 19669 22661 19703
rect 22661 19669 22695 19703
rect 22695 19669 22704 19703
rect 22652 19660 22704 19669
rect 4680 19558 4732 19610
rect 4744 19558 4796 19610
rect 4808 19558 4860 19610
rect 4872 19558 4924 19610
rect 12078 19558 12130 19610
rect 12142 19558 12194 19610
rect 12206 19558 12258 19610
rect 12270 19558 12322 19610
rect 19475 19558 19527 19610
rect 19539 19558 19591 19610
rect 19603 19558 19655 19610
rect 19667 19558 19719 19610
rect 3424 19456 3476 19508
rect 3792 19456 3844 19508
rect 4528 19456 4580 19508
rect 5356 19456 5408 19508
rect 5448 19456 5500 19508
rect 7840 19388 7892 19440
rect 1400 19295 1452 19304
rect 1400 19261 1409 19295
rect 1409 19261 1443 19295
rect 1443 19261 1452 19295
rect 1400 19252 1452 19261
rect 3332 19295 3384 19304
rect 3332 19261 3366 19295
rect 3366 19261 3384 19295
rect 3332 19252 3384 19261
rect 3700 19252 3752 19304
rect 5080 19295 5132 19304
rect 5080 19261 5089 19295
rect 5089 19261 5123 19295
rect 5123 19261 5132 19295
rect 5080 19252 5132 19261
rect 5540 19320 5592 19372
rect 6460 19320 6512 19372
rect 10140 19456 10192 19508
rect 12532 19456 12584 19508
rect 1676 19227 1728 19236
rect 1676 19193 1710 19227
rect 1710 19193 1728 19227
rect 1676 19184 1728 19193
rect 2320 19184 2372 19236
rect 2964 19184 3016 19236
rect 5264 19184 5316 19236
rect 8300 19252 8352 19304
rect 14188 19456 14240 19508
rect 15476 19456 15528 19508
rect 8484 19184 8536 19236
rect 10048 19252 10100 19304
rect 13084 19363 13136 19372
rect 13084 19329 13093 19363
rect 13093 19329 13127 19363
rect 13127 19329 13136 19363
rect 13084 19320 13136 19329
rect 8668 19184 8720 19236
rect 8760 19184 8812 19236
rect 9772 19184 9824 19236
rect 10232 19184 10284 19236
rect 2780 19159 2832 19168
rect 2780 19125 2789 19159
rect 2789 19125 2823 19159
rect 2823 19125 2832 19159
rect 2780 19116 2832 19125
rect 3240 19116 3292 19168
rect 4160 19116 4212 19168
rect 4712 19159 4764 19168
rect 4712 19125 4721 19159
rect 4721 19125 4755 19159
rect 4755 19125 4764 19159
rect 4712 19116 4764 19125
rect 5724 19159 5776 19168
rect 5724 19125 5733 19159
rect 5733 19125 5767 19159
rect 5767 19125 5776 19159
rect 5724 19116 5776 19125
rect 6828 19116 6880 19168
rect 7840 19116 7892 19168
rect 8116 19116 8168 19168
rect 13544 19252 13596 19304
rect 13636 19252 13688 19304
rect 19340 19456 19392 19508
rect 19432 19431 19484 19440
rect 19432 19397 19441 19431
rect 19441 19397 19475 19431
rect 19475 19397 19484 19431
rect 19432 19388 19484 19397
rect 14648 19320 14700 19372
rect 14924 19363 14976 19372
rect 14924 19329 14933 19363
rect 14933 19329 14967 19363
rect 14967 19329 14976 19363
rect 14924 19320 14976 19329
rect 15936 19320 15988 19372
rect 16580 19320 16632 19372
rect 19892 19320 19944 19372
rect 16120 19252 16172 19304
rect 16672 19295 16724 19304
rect 16672 19261 16681 19295
rect 16681 19261 16715 19295
rect 16715 19261 16724 19295
rect 16672 19252 16724 19261
rect 17408 19295 17460 19304
rect 17408 19261 17417 19295
rect 17417 19261 17451 19295
rect 17451 19261 17460 19295
rect 17408 19252 17460 19261
rect 18052 19295 18104 19304
rect 18052 19261 18061 19295
rect 18061 19261 18095 19295
rect 18095 19261 18104 19295
rect 18052 19252 18104 19261
rect 18696 19252 18748 19304
rect 20904 19252 20956 19304
rect 12900 19227 12952 19236
rect 10692 19159 10744 19168
rect 10692 19125 10701 19159
rect 10701 19125 10735 19159
rect 10735 19125 10744 19159
rect 10692 19116 10744 19125
rect 10784 19159 10836 19168
rect 10784 19125 10793 19159
rect 10793 19125 10827 19159
rect 10827 19125 10836 19159
rect 10784 19116 10836 19125
rect 11704 19159 11756 19168
rect 11704 19125 11713 19159
rect 11713 19125 11747 19159
rect 11747 19125 11756 19159
rect 11704 19116 11756 19125
rect 11796 19159 11848 19168
rect 11796 19125 11805 19159
rect 11805 19125 11839 19159
rect 11839 19125 11848 19159
rect 11796 19116 11848 19125
rect 12348 19116 12400 19168
rect 12900 19193 12909 19227
rect 12909 19193 12943 19227
rect 12943 19193 12952 19227
rect 12900 19184 12952 19193
rect 19248 19184 19300 19236
rect 15200 19116 15252 19168
rect 15292 19159 15344 19168
rect 15292 19125 15301 19159
rect 15301 19125 15335 19159
rect 15335 19125 15344 19159
rect 16304 19159 16356 19168
rect 15292 19116 15344 19125
rect 16304 19125 16313 19159
rect 16313 19125 16347 19159
rect 16347 19125 16356 19159
rect 16304 19116 16356 19125
rect 16764 19159 16816 19168
rect 16764 19125 16773 19159
rect 16773 19125 16807 19159
rect 16807 19125 16816 19159
rect 16764 19116 16816 19125
rect 17316 19116 17368 19168
rect 17960 19116 18012 19168
rect 20260 19116 20312 19168
rect 21732 19252 21784 19304
rect 21272 19116 21324 19168
rect 21640 19116 21692 19168
rect 8379 19014 8431 19066
rect 8443 19014 8495 19066
rect 8507 19014 8559 19066
rect 8571 19014 8623 19066
rect 15776 19014 15828 19066
rect 15840 19014 15892 19066
rect 15904 19014 15956 19066
rect 15968 19014 16020 19066
rect 1676 18912 1728 18964
rect 4712 18912 4764 18964
rect 4804 18912 4856 18964
rect 6828 18912 6880 18964
rect 9864 18912 9916 18964
rect 10692 18912 10744 18964
rect 5724 18844 5776 18896
rect 3700 18776 3752 18828
rect 4160 18776 4212 18828
rect 7932 18844 7984 18896
rect 8208 18887 8260 18896
rect 8208 18853 8242 18887
rect 8242 18853 8260 18887
rect 8208 18844 8260 18853
rect 8300 18844 8352 18896
rect 12532 18912 12584 18964
rect 16120 18912 16172 18964
rect 16856 18912 16908 18964
rect 18880 18955 18932 18964
rect 18880 18921 18889 18955
rect 18889 18921 18923 18955
rect 18923 18921 18932 18955
rect 18880 18912 18932 18921
rect 22468 18912 22520 18964
rect 16212 18844 16264 18896
rect 19432 18844 19484 18896
rect 21640 18844 21692 18896
rect 9496 18776 9548 18828
rect 9680 18819 9732 18828
rect 9680 18785 9689 18819
rect 9689 18785 9723 18819
rect 9723 18785 9732 18819
rect 9680 18776 9732 18785
rect 10784 18776 10836 18828
rect 11612 18776 11664 18828
rect 11980 18776 12032 18828
rect 12164 18819 12216 18828
rect 12164 18785 12198 18819
rect 12198 18785 12216 18819
rect 12164 18776 12216 18785
rect 12624 18776 12676 18828
rect 2320 18751 2372 18760
rect 2320 18717 2329 18751
rect 2329 18717 2363 18751
rect 2363 18717 2372 18751
rect 2320 18708 2372 18717
rect 4620 18751 4672 18760
rect 4620 18717 4629 18751
rect 4629 18717 4663 18751
rect 4663 18717 4672 18751
rect 4620 18708 4672 18717
rect 7288 18751 7340 18760
rect 5264 18640 5316 18692
rect 7288 18717 7297 18751
rect 7297 18717 7331 18751
rect 7331 18717 7340 18751
rect 7288 18708 7340 18717
rect 7564 18708 7616 18760
rect 7932 18751 7984 18760
rect 7932 18717 7941 18751
rect 7941 18717 7975 18751
rect 7975 18717 7984 18751
rect 7932 18708 7984 18717
rect 9772 18708 9824 18760
rect 13268 18776 13320 18828
rect 15108 18776 15160 18828
rect 15200 18776 15252 18828
rect 15384 18819 15436 18828
rect 15384 18785 15393 18819
rect 15393 18785 15427 18819
rect 15427 18785 15436 18819
rect 15384 18776 15436 18785
rect 15476 18776 15528 18828
rect 14924 18708 14976 18760
rect 17500 18751 17552 18760
rect 17500 18717 17509 18751
rect 17509 18717 17543 18751
rect 17543 18717 17552 18751
rect 17500 18708 17552 18717
rect 19800 18751 19852 18760
rect 19800 18717 19809 18751
rect 19809 18717 19843 18751
rect 19843 18717 19852 18751
rect 19800 18708 19852 18717
rect 5080 18615 5132 18624
rect 5080 18581 5089 18615
rect 5089 18581 5123 18615
rect 5123 18581 5132 18615
rect 5080 18572 5132 18581
rect 6460 18615 6512 18624
rect 6460 18581 6469 18615
rect 6469 18581 6503 18615
rect 6503 18581 6512 18615
rect 6460 18572 6512 18581
rect 6828 18615 6880 18624
rect 6828 18581 6837 18615
rect 6837 18581 6871 18615
rect 6871 18581 6880 18615
rect 6828 18572 6880 18581
rect 7564 18572 7616 18624
rect 10048 18572 10100 18624
rect 13084 18572 13136 18624
rect 13268 18615 13320 18624
rect 13268 18581 13277 18615
rect 13277 18581 13311 18615
rect 13311 18581 13320 18615
rect 13268 18572 13320 18581
rect 13544 18615 13596 18624
rect 13544 18581 13553 18615
rect 13553 18581 13587 18615
rect 13587 18581 13596 18615
rect 13544 18572 13596 18581
rect 15016 18640 15068 18692
rect 22100 18776 22152 18828
rect 21272 18751 21324 18760
rect 21272 18717 21281 18751
rect 21281 18717 21315 18751
rect 21315 18717 21324 18751
rect 21272 18708 21324 18717
rect 18512 18572 18564 18624
rect 20352 18615 20404 18624
rect 20352 18581 20361 18615
rect 20361 18581 20395 18615
rect 20395 18581 20404 18615
rect 20352 18572 20404 18581
rect 4680 18470 4732 18522
rect 4744 18470 4796 18522
rect 4808 18470 4860 18522
rect 4872 18470 4924 18522
rect 12078 18470 12130 18522
rect 12142 18470 12194 18522
rect 12206 18470 12258 18522
rect 12270 18470 12322 18522
rect 19475 18470 19527 18522
rect 19539 18470 19591 18522
rect 19603 18470 19655 18522
rect 19667 18470 19719 18522
rect 4160 18411 4212 18420
rect 3700 18343 3752 18352
rect 3700 18309 3709 18343
rect 3709 18309 3743 18343
rect 3743 18309 3752 18343
rect 3700 18300 3752 18309
rect 4160 18377 4169 18411
rect 4169 18377 4203 18411
rect 4203 18377 4212 18411
rect 4160 18368 4212 18377
rect 9588 18368 9640 18420
rect 9772 18368 9824 18420
rect 11612 18411 11664 18420
rect 11612 18377 11621 18411
rect 11621 18377 11655 18411
rect 11655 18377 11664 18411
rect 11612 18368 11664 18377
rect 7196 18300 7248 18352
rect 3424 18232 3476 18284
rect 3976 18207 4028 18216
rect 3608 18096 3660 18148
rect 3976 18173 3985 18207
rect 3985 18173 4019 18207
rect 4019 18173 4028 18207
rect 3976 18164 4028 18173
rect 7564 18232 7616 18284
rect 8300 18300 8352 18352
rect 10140 18300 10192 18352
rect 7932 18275 7984 18284
rect 7932 18241 7941 18275
rect 7941 18241 7975 18275
rect 7975 18241 7984 18275
rect 7932 18232 7984 18241
rect 2320 18028 2372 18080
rect 3424 18028 3476 18080
rect 5632 18096 5684 18148
rect 6828 18164 6880 18216
rect 8208 18164 8260 18216
rect 8392 18164 8444 18216
rect 9864 18164 9916 18216
rect 12072 18232 12124 18284
rect 14832 18368 14884 18420
rect 16396 18368 16448 18420
rect 18696 18368 18748 18420
rect 19340 18368 19392 18420
rect 14096 18300 14148 18352
rect 14924 18232 14976 18284
rect 16212 18275 16264 18284
rect 16212 18241 16221 18275
rect 16221 18241 16255 18275
rect 16255 18241 16264 18275
rect 16212 18232 16264 18241
rect 17500 18300 17552 18352
rect 20076 18300 20128 18352
rect 18052 18275 18104 18284
rect 18052 18241 18061 18275
rect 18061 18241 18095 18275
rect 18095 18241 18104 18275
rect 18052 18232 18104 18241
rect 10324 18164 10376 18216
rect 10784 18164 10836 18216
rect 12440 18207 12492 18216
rect 12440 18173 12449 18207
rect 12449 18173 12483 18207
rect 12483 18173 12492 18207
rect 12440 18164 12492 18173
rect 12808 18164 12860 18216
rect 5724 18028 5776 18080
rect 5908 18071 5960 18080
rect 5908 18037 5917 18071
rect 5917 18037 5951 18071
rect 5951 18037 5960 18071
rect 5908 18028 5960 18037
rect 6276 18028 6328 18080
rect 8944 18028 8996 18080
rect 11704 18096 11756 18148
rect 12348 18096 12400 18148
rect 14740 18164 14792 18216
rect 16856 18164 16908 18216
rect 17868 18207 17920 18216
rect 17868 18173 17877 18207
rect 17877 18173 17911 18207
rect 17911 18173 17920 18207
rect 17868 18164 17920 18173
rect 20076 18164 20128 18216
rect 14280 18096 14332 18148
rect 15384 18096 15436 18148
rect 16304 18096 16356 18148
rect 18788 18096 18840 18148
rect 20720 18232 20772 18284
rect 20812 18164 20864 18216
rect 21272 18164 21324 18216
rect 22468 18164 22520 18216
rect 22376 18096 22428 18148
rect 12532 18028 12584 18080
rect 13912 18028 13964 18080
rect 14924 18028 14976 18080
rect 16948 18028 17000 18080
rect 17500 18028 17552 18080
rect 19984 18071 20036 18080
rect 19984 18037 19993 18071
rect 19993 18037 20027 18071
rect 20027 18037 20036 18071
rect 19984 18028 20036 18037
rect 20352 18071 20404 18080
rect 20352 18037 20361 18071
rect 20361 18037 20395 18071
rect 20395 18037 20404 18071
rect 20352 18028 20404 18037
rect 20444 18028 20496 18080
rect 21180 18028 21232 18080
rect 8379 17926 8431 17978
rect 8443 17926 8495 17978
rect 8507 17926 8559 17978
rect 8571 17926 8623 17978
rect 15776 17926 15828 17978
rect 15840 17926 15892 17978
rect 15904 17926 15956 17978
rect 15968 17926 16020 17978
rect 2780 17824 2832 17876
rect 2596 17756 2648 17808
rect 2320 17688 2372 17740
rect 3516 17688 3568 17740
rect 3608 17595 3660 17604
rect 3608 17561 3617 17595
rect 3617 17561 3651 17595
rect 3651 17561 3660 17595
rect 3608 17552 3660 17561
rect 4068 17688 4120 17740
rect 4436 17688 4488 17740
rect 4160 17620 4212 17672
rect 5908 17688 5960 17740
rect 4804 17663 4856 17672
rect 4804 17629 4813 17663
rect 4813 17629 4847 17663
rect 4847 17629 4856 17663
rect 4804 17620 4856 17629
rect 4160 17484 4212 17536
rect 5448 17484 5500 17536
rect 6092 17484 6144 17536
rect 8760 17688 8812 17740
rect 11796 17756 11848 17808
rect 12072 17756 12124 17808
rect 12440 17756 12492 17808
rect 12716 17824 12768 17876
rect 13728 17824 13780 17876
rect 14280 17867 14332 17876
rect 14280 17833 14289 17867
rect 14289 17833 14323 17867
rect 14323 17833 14332 17867
rect 14280 17824 14332 17833
rect 16212 17824 16264 17876
rect 18788 17867 18840 17876
rect 18788 17833 18797 17867
rect 18797 17833 18831 17867
rect 18831 17833 18840 17867
rect 18788 17824 18840 17833
rect 15292 17756 15344 17808
rect 15476 17756 15528 17808
rect 16120 17756 16172 17808
rect 16304 17756 16356 17808
rect 12348 17731 12400 17740
rect 6460 17663 6512 17672
rect 6460 17629 6469 17663
rect 6469 17629 6503 17663
rect 6503 17629 6512 17663
rect 6460 17620 6512 17629
rect 8576 17663 8628 17672
rect 8576 17629 8585 17663
rect 8585 17629 8619 17663
rect 8619 17629 8628 17663
rect 8576 17620 8628 17629
rect 9036 17620 9088 17672
rect 9404 17620 9456 17672
rect 12348 17697 12357 17731
rect 12357 17697 12391 17731
rect 12391 17697 12400 17731
rect 12348 17688 12400 17697
rect 12808 17688 12860 17740
rect 10324 17663 10376 17672
rect 9496 17552 9548 17604
rect 10324 17629 10333 17663
rect 10333 17629 10367 17663
rect 10367 17629 10376 17663
rect 10324 17620 10376 17629
rect 17132 17688 17184 17740
rect 18052 17756 18104 17808
rect 19340 17756 19392 17808
rect 22652 17824 22704 17876
rect 21180 17799 21232 17808
rect 18972 17688 19024 17740
rect 19248 17688 19300 17740
rect 21180 17765 21214 17799
rect 21214 17765 21232 17799
rect 21180 17756 21232 17765
rect 14004 17620 14056 17672
rect 10232 17552 10284 17604
rect 11704 17595 11756 17604
rect 11704 17561 11713 17595
rect 11713 17561 11747 17595
rect 11747 17561 11756 17595
rect 11704 17552 11756 17561
rect 12900 17552 12952 17604
rect 14832 17552 14884 17604
rect 15108 17552 15160 17604
rect 18420 17620 18472 17672
rect 19892 17688 19944 17740
rect 20536 17688 20588 17740
rect 19800 17620 19852 17672
rect 20352 17620 20404 17672
rect 20812 17620 20864 17672
rect 7840 17527 7892 17536
rect 7840 17493 7849 17527
rect 7849 17493 7883 17527
rect 7883 17493 7892 17527
rect 7840 17484 7892 17493
rect 8024 17484 8076 17536
rect 9220 17484 9272 17536
rect 11520 17484 11572 17536
rect 16672 17527 16724 17536
rect 16672 17493 16681 17527
rect 16681 17493 16715 17527
rect 16715 17493 16724 17527
rect 16672 17484 16724 17493
rect 17408 17484 17460 17536
rect 19064 17527 19116 17536
rect 19064 17493 19073 17527
rect 19073 17493 19107 17527
rect 19107 17493 19116 17527
rect 19064 17484 19116 17493
rect 20168 17484 20220 17536
rect 21548 17484 21600 17536
rect 22008 17484 22060 17536
rect 4680 17382 4732 17434
rect 4744 17382 4796 17434
rect 4808 17382 4860 17434
rect 4872 17382 4924 17434
rect 12078 17382 12130 17434
rect 12142 17382 12194 17434
rect 12206 17382 12258 17434
rect 12270 17382 12322 17434
rect 19475 17382 19527 17434
rect 19539 17382 19591 17434
rect 19603 17382 19655 17434
rect 19667 17382 19719 17434
rect 1400 17280 1452 17332
rect 3516 17323 3568 17332
rect 3516 17289 3525 17323
rect 3525 17289 3559 17323
rect 3559 17289 3568 17323
rect 3516 17280 3568 17289
rect 4344 17280 4396 17332
rect 4436 17280 4488 17332
rect 5080 17280 5132 17332
rect 5172 17280 5224 17332
rect 5356 17280 5408 17332
rect 5540 17280 5592 17332
rect 3700 17212 3752 17264
rect 4068 17212 4120 17264
rect 4620 17212 4672 17264
rect 3608 17144 3660 17196
rect 4712 17144 4764 17196
rect 2228 17076 2280 17128
rect 4068 17076 4120 17128
rect 3332 17008 3384 17060
rect 4068 16940 4120 16992
rect 4252 16983 4304 16992
rect 4252 16949 4261 16983
rect 4261 16949 4295 16983
rect 4295 16949 4304 16983
rect 6828 17212 6880 17264
rect 6000 17144 6052 17196
rect 6000 17008 6052 17060
rect 6552 17076 6604 17128
rect 7840 17076 7892 17128
rect 8300 17076 8352 17128
rect 11980 17280 12032 17332
rect 14004 17323 14056 17332
rect 14004 17289 14013 17323
rect 14013 17289 14047 17323
rect 14047 17289 14056 17323
rect 14004 17280 14056 17289
rect 14924 17280 14976 17332
rect 16488 17323 16540 17332
rect 16488 17289 16497 17323
rect 16497 17289 16531 17323
rect 16531 17289 16540 17323
rect 16488 17280 16540 17289
rect 20444 17280 20496 17332
rect 12256 17212 12308 17264
rect 14832 17255 14884 17264
rect 14832 17221 14841 17255
rect 14841 17221 14875 17255
rect 14875 17221 14884 17255
rect 14832 17212 14884 17221
rect 17132 17212 17184 17264
rect 12624 17187 12676 17196
rect 12624 17153 12633 17187
rect 12633 17153 12667 17187
rect 12667 17153 12676 17187
rect 12624 17144 12676 17153
rect 10324 17119 10376 17128
rect 10324 17085 10333 17119
rect 10333 17085 10367 17119
rect 10367 17085 10376 17119
rect 10324 17076 10376 17085
rect 13268 17076 13320 17128
rect 14372 17076 14424 17128
rect 14464 17076 14516 17128
rect 15200 17076 15252 17128
rect 17408 17076 17460 17128
rect 4252 16940 4304 16949
rect 4804 16940 4856 16992
rect 5264 16983 5316 16992
rect 5264 16949 5273 16983
rect 5273 16949 5307 16983
rect 5307 16949 5316 16983
rect 5264 16940 5316 16949
rect 7288 16940 7340 16992
rect 7840 16940 7892 16992
rect 8944 17008 8996 17060
rect 11060 17008 11112 17060
rect 8852 16940 8904 16992
rect 13820 17008 13872 17060
rect 19800 17212 19852 17264
rect 19984 17144 20036 17196
rect 21180 17280 21232 17332
rect 18972 17119 19024 17128
rect 18972 17085 18981 17119
rect 18981 17085 19015 17119
rect 19015 17085 19024 17119
rect 18972 17076 19024 17085
rect 19800 17076 19852 17128
rect 20168 17119 20220 17128
rect 20168 17085 20177 17119
rect 20177 17085 20211 17119
rect 20211 17085 20220 17119
rect 20168 17076 20220 17085
rect 20812 17119 20864 17128
rect 20812 17085 20821 17119
rect 20821 17085 20855 17119
rect 20855 17085 20864 17119
rect 20812 17076 20864 17085
rect 22008 17076 22060 17128
rect 11520 16940 11572 16992
rect 13084 16940 13136 16992
rect 14924 16940 14976 16992
rect 15016 16940 15068 16992
rect 21640 17008 21692 17060
rect 22468 17119 22520 17128
rect 22468 17085 22477 17119
rect 22477 17085 22511 17119
rect 22511 17085 22520 17119
rect 22468 17076 22520 17085
rect 16672 16940 16724 16992
rect 18052 16940 18104 16992
rect 18328 16940 18380 16992
rect 18880 16940 18932 16992
rect 21824 16940 21876 16992
rect 22652 16983 22704 16992
rect 22652 16949 22661 16983
rect 22661 16949 22695 16983
rect 22695 16949 22704 16983
rect 22652 16940 22704 16949
rect 8379 16838 8431 16890
rect 8443 16838 8495 16890
rect 8507 16838 8559 16890
rect 8571 16838 8623 16890
rect 15776 16838 15828 16890
rect 15840 16838 15892 16890
rect 15904 16838 15956 16890
rect 15968 16838 16020 16890
rect 3148 16736 3200 16788
rect 3332 16779 3384 16788
rect 3332 16745 3341 16779
rect 3341 16745 3375 16779
rect 3375 16745 3384 16779
rect 3332 16736 3384 16745
rect 4252 16736 4304 16788
rect 5264 16736 5316 16788
rect 5448 16736 5500 16788
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 2320 16668 2372 16720
rect 2596 16668 2648 16720
rect 3976 16668 4028 16720
rect 4068 16600 4120 16652
rect 4804 16668 4856 16720
rect 7748 16668 7800 16720
rect 7932 16668 7984 16720
rect 9220 16668 9272 16720
rect 9956 16711 10008 16720
rect 9956 16677 9990 16711
rect 9990 16677 10008 16711
rect 9956 16668 10008 16677
rect 10232 16736 10284 16788
rect 10968 16736 11020 16788
rect 13084 16779 13136 16788
rect 13084 16745 13093 16779
rect 13093 16745 13127 16779
rect 13127 16745 13136 16779
rect 13084 16736 13136 16745
rect 13176 16736 13228 16788
rect 13544 16736 13596 16788
rect 4896 16600 4948 16652
rect 5448 16643 5500 16652
rect 5448 16609 5457 16643
rect 5457 16609 5491 16643
rect 5491 16609 5500 16643
rect 5448 16600 5500 16609
rect 4344 16532 4396 16584
rect 6000 16600 6052 16652
rect 6184 16600 6236 16652
rect 8944 16600 8996 16652
rect 3424 16464 3476 16516
rect 5724 16532 5776 16584
rect 6460 16396 6512 16448
rect 7472 16396 7524 16448
rect 8944 16464 8996 16516
rect 10232 16600 10284 16652
rect 11336 16600 11388 16652
rect 11888 16668 11940 16720
rect 13912 16668 13964 16720
rect 15660 16736 15712 16788
rect 14924 16668 14976 16720
rect 17960 16736 18012 16788
rect 18972 16736 19024 16788
rect 19984 16736 20036 16788
rect 22652 16736 22704 16788
rect 15384 16600 15436 16652
rect 16488 16600 16540 16652
rect 17868 16668 17920 16720
rect 19708 16668 19760 16720
rect 19892 16668 19944 16720
rect 20260 16668 20312 16720
rect 20812 16668 20864 16720
rect 21640 16711 21692 16720
rect 21640 16677 21674 16711
rect 21674 16677 21692 16711
rect 21640 16668 21692 16677
rect 19248 16600 19300 16652
rect 19340 16600 19392 16652
rect 20720 16600 20772 16652
rect 9956 16396 10008 16448
rect 10324 16396 10376 16448
rect 12900 16532 12952 16584
rect 13452 16532 13504 16584
rect 13820 16532 13872 16584
rect 15200 16532 15252 16584
rect 18788 16532 18840 16584
rect 19984 16575 20036 16584
rect 19984 16541 19993 16575
rect 19993 16541 20027 16575
rect 20027 16541 20036 16575
rect 20904 16575 20956 16584
rect 19984 16532 20036 16541
rect 20904 16541 20913 16575
rect 20913 16541 20947 16575
rect 20947 16541 20956 16575
rect 20904 16532 20956 16541
rect 11060 16507 11112 16516
rect 11060 16473 11069 16507
rect 11069 16473 11103 16507
rect 11103 16473 11112 16507
rect 11060 16464 11112 16473
rect 14280 16396 14332 16448
rect 17500 16464 17552 16516
rect 18420 16396 18472 16448
rect 20260 16396 20312 16448
rect 4680 16294 4732 16346
rect 4744 16294 4796 16346
rect 4808 16294 4860 16346
rect 4872 16294 4924 16346
rect 12078 16294 12130 16346
rect 12142 16294 12194 16346
rect 12206 16294 12258 16346
rect 12270 16294 12322 16346
rect 19475 16294 19527 16346
rect 19539 16294 19591 16346
rect 19603 16294 19655 16346
rect 19667 16294 19719 16346
rect 2780 16192 2832 16244
rect 3424 16235 3476 16244
rect 3424 16201 3433 16235
rect 3433 16201 3467 16235
rect 3467 16201 3476 16235
rect 3424 16192 3476 16201
rect 1492 16031 1544 16040
rect 1492 15997 1501 16031
rect 1501 15997 1535 16031
rect 1535 15997 1544 16031
rect 1492 15988 1544 15997
rect 1860 15988 1912 16040
rect 5908 16192 5960 16244
rect 6828 16192 6880 16244
rect 10416 16192 10468 16244
rect 10692 16192 10744 16244
rect 4252 16056 4304 16108
rect 4528 16099 4580 16108
rect 4528 16065 4540 16099
rect 4540 16065 4574 16099
rect 4574 16065 4580 16099
rect 4528 16056 4580 16065
rect 5540 16056 5592 16108
rect 5724 16056 5776 16108
rect 6276 16056 6328 16108
rect 7380 16056 7432 16108
rect 9312 16056 9364 16108
rect 10876 16056 10928 16108
rect 2688 15920 2740 15972
rect 4896 15988 4948 16040
rect 6644 15988 6696 16040
rect 6828 16031 6880 16040
rect 6828 15997 6837 16031
rect 6837 15997 6871 16031
rect 6871 15997 6880 16031
rect 6828 15988 6880 15997
rect 6736 15920 6788 15972
rect 9680 16031 9732 16040
rect 9680 15997 9689 16031
rect 9689 15997 9723 16031
rect 9723 15997 9732 16031
rect 9680 15988 9732 15997
rect 10784 15988 10836 16040
rect 11244 15988 11296 16040
rect 11612 16099 11664 16108
rect 11612 16065 11621 16099
rect 11621 16065 11655 16099
rect 11655 16065 11664 16099
rect 11980 16192 12032 16244
rect 13268 16192 13320 16244
rect 17592 16192 17644 16244
rect 16580 16124 16632 16176
rect 19800 16192 19852 16244
rect 21548 16235 21600 16244
rect 21548 16201 21557 16235
rect 21557 16201 21591 16235
rect 21591 16201 21600 16235
rect 21548 16192 21600 16201
rect 22744 16124 22796 16176
rect 11612 16056 11664 16065
rect 11796 15988 11848 16040
rect 11980 16031 12032 16040
rect 11980 15997 11989 16031
rect 11989 15997 12023 16031
rect 12023 15997 12032 16031
rect 11980 15988 12032 15997
rect 13084 16056 13136 16108
rect 13820 16099 13872 16108
rect 13820 16065 13832 16099
rect 13832 16065 13866 16099
rect 13866 16065 13872 16099
rect 13820 16056 13872 16065
rect 15200 16056 15252 16108
rect 22008 16056 22060 16108
rect 22376 16056 22428 16108
rect 14004 15988 14056 16040
rect 14096 16031 14148 16040
rect 14096 15997 14105 16031
rect 14105 15997 14139 16031
rect 14139 15997 14148 16031
rect 14096 15988 14148 15997
rect 16856 15988 16908 16040
rect 4344 15852 4396 15904
rect 4896 15852 4948 15904
rect 5172 15852 5224 15904
rect 6552 15852 6604 15904
rect 7288 15895 7340 15904
rect 7288 15861 7303 15895
rect 7303 15861 7337 15895
rect 7337 15861 7340 15895
rect 7288 15852 7340 15861
rect 8208 15852 8260 15904
rect 9312 15852 9364 15904
rect 10692 15852 10744 15904
rect 15660 15920 15712 15972
rect 11244 15852 11296 15904
rect 12072 15852 12124 15904
rect 12348 15852 12400 15904
rect 12624 15852 12676 15904
rect 12808 15895 12860 15904
rect 12808 15861 12817 15895
rect 12817 15861 12851 15895
rect 12851 15861 12860 15895
rect 12808 15852 12860 15861
rect 13452 15852 13504 15904
rect 13912 15852 13964 15904
rect 15200 15895 15252 15904
rect 15200 15861 15209 15895
rect 15209 15861 15243 15895
rect 15243 15861 15252 15895
rect 15200 15852 15252 15861
rect 16120 15852 16172 15904
rect 18696 15988 18748 16040
rect 19340 15920 19392 15972
rect 20720 15988 20772 16040
rect 20904 15988 20956 16040
rect 21824 15920 21876 15972
rect 20168 15852 20220 15904
rect 20904 15852 20956 15904
rect 21272 15895 21324 15904
rect 21272 15861 21281 15895
rect 21281 15861 21315 15895
rect 21315 15861 21324 15895
rect 21272 15852 21324 15861
rect 8379 15750 8431 15802
rect 8443 15750 8495 15802
rect 8507 15750 8559 15802
rect 8571 15750 8623 15802
rect 15776 15750 15828 15802
rect 15840 15750 15892 15802
rect 15904 15750 15956 15802
rect 15968 15750 16020 15802
rect 7196 15648 7248 15700
rect 10784 15648 10836 15700
rect 10876 15648 10928 15700
rect 12716 15648 12768 15700
rect 13084 15648 13136 15700
rect 14924 15691 14976 15700
rect 14924 15657 14933 15691
rect 14933 15657 14967 15691
rect 14967 15657 14976 15691
rect 14924 15648 14976 15657
rect 15108 15648 15160 15700
rect 19340 15691 19392 15700
rect 1860 15580 1912 15632
rect 3976 15580 4028 15632
rect 4252 15580 4304 15632
rect 2964 15512 3016 15564
rect 3148 15555 3200 15564
rect 3148 15521 3157 15555
rect 3157 15521 3191 15555
rect 3191 15521 3200 15555
rect 3148 15512 3200 15521
rect 4436 15555 4488 15564
rect 4436 15521 4445 15555
rect 4445 15521 4479 15555
rect 4479 15521 4488 15555
rect 4436 15512 4488 15521
rect 6828 15580 6880 15632
rect 7472 15580 7524 15632
rect 3332 15487 3384 15496
rect 3332 15453 3341 15487
rect 3341 15453 3375 15487
rect 3375 15453 3384 15487
rect 3332 15444 3384 15453
rect 5448 15487 5500 15496
rect 5448 15453 5460 15487
rect 5460 15453 5494 15487
rect 5494 15453 5500 15487
rect 5448 15444 5500 15453
rect 6000 15512 6052 15564
rect 8668 15512 8720 15564
rect 8944 15555 8996 15564
rect 8944 15521 8953 15555
rect 8953 15521 8987 15555
rect 8987 15521 8996 15555
rect 8944 15512 8996 15521
rect 10508 15580 10560 15632
rect 10692 15580 10744 15632
rect 9128 15512 9180 15564
rect 6460 15444 6512 15496
rect 6828 15444 6880 15496
rect 4988 15376 5040 15428
rect 10968 15555 11020 15564
rect 10968 15521 10977 15555
rect 10977 15521 11011 15555
rect 11011 15521 11020 15555
rect 10968 15512 11020 15521
rect 14004 15580 14056 15632
rect 11796 15555 11848 15564
rect 11796 15521 11805 15555
rect 11805 15521 11839 15555
rect 11839 15521 11848 15555
rect 11796 15512 11848 15521
rect 12900 15512 12952 15564
rect 13268 15512 13320 15564
rect 13912 15512 13964 15564
rect 15108 15555 15160 15564
rect 9772 15444 9824 15496
rect 10232 15487 10284 15496
rect 10232 15453 10241 15487
rect 10241 15453 10275 15487
rect 10275 15453 10284 15487
rect 10232 15444 10284 15453
rect 10416 15444 10468 15496
rect 2688 15308 2740 15360
rect 5264 15308 5316 15360
rect 5908 15308 5960 15360
rect 6736 15308 6788 15360
rect 7104 15308 7156 15360
rect 9220 15308 9272 15360
rect 9312 15308 9364 15360
rect 10600 15308 10652 15360
rect 10784 15351 10836 15360
rect 10784 15317 10793 15351
rect 10793 15317 10827 15351
rect 10827 15317 10836 15351
rect 10784 15308 10836 15317
rect 10876 15308 10928 15360
rect 12440 15444 12492 15496
rect 13084 15444 13136 15496
rect 12624 15308 12676 15360
rect 15108 15521 15117 15555
rect 15117 15521 15151 15555
rect 15151 15521 15160 15555
rect 15108 15512 15160 15521
rect 14740 15444 14792 15496
rect 17960 15580 18012 15632
rect 18788 15580 18840 15632
rect 19340 15657 19349 15691
rect 19349 15657 19383 15691
rect 19383 15657 19392 15691
rect 19340 15648 19392 15657
rect 20168 15648 20220 15700
rect 20720 15648 20772 15700
rect 19892 15580 19944 15632
rect 15844 15512 15896 15564
rect 16120 15512 16172 15564
rect 18972 15512 19024 15564
rect 20168 15555 20220 15564
rect 20168 15521 20177 15555
rect 20177 15521 20211 15555
rect 20211 15521 20220 15555
rect 20168 15512 20220 15521
rect 21272 15580 21324 15632
rect 21640 15512 21692 15564
rect 20904 15487 20956 15496
rect 17684 15376 17736 15428
rect 13544 15308 13596 15360
rect 14188 15308 14240 15360
rect 15200 15308 15252 15360
rect 15476 15308 15528 15360
rect 16120 15308 16172 15360
rect 20904 15453 20913 15487
rect 20913 15453 20947 15487
rect 20947 15453 20956 15487
rect 20904 15444 20956 15453
rect 18696 15308 18748 15360
rect 19800 15351 19852 15360
rect 19800 15317 19809 15351
rect 19809 15317 19843 15351
rect 19843 15317 19852 15351
rect 19800 15308 19852 15317
rect 21548 15308 21600 15360
rect 4680 15206 4732 15258
rect 4744 15206 4796 15258
rect 4808 15206 4860 15258
rect 4872 15206 4924 15258
rect 12078 15206 12130 15258
rect 12142 15206 12194 15258
rect 12206 15206 12258 15258
rect 12270 15206 12322 15258
rect 19475 15206 19527 15258
rect 19539 15206 19591 15258
rect 19603 15206 19655 15258
rect 19667 15206 19719 15258
rect 1860 15011 1912 15020
rect 1860 14977 1869 15011
rect 1869 14977 1903 15011
rect 1903 14977 1912 15011
rect 1860 14968 1912 14977
rect 6736 15104 6788 15156
rect 10048 15104 10100 15156
rect 11612 15104 11664 15156
rect 11888 15104 11940 15156
rect 14464 15104 14516 15156
rect 15016 15104 15068 15156
rect 17960 15104 18012 15156
rect 18972 15104 19024 15156
rect 20444 15104 20496 15156
rect 20720 15104 20772 15156
rect 11704 15036 11756 15088
rect 12716 15036 12768 15088
rect 12992 15036 13044 15088
rect 18052 15036 18104 15088
rect 19340 15036 19392 15088
rect 5356 14968 5408 15020
rect 9956 14968 10008 15020
rect 3976 14900 4028 14952
rect 4252 14900 4304 14952
rect 5172 14900 5224 14952
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 3056 14832 3108 14884
rect 7104 14875 7156 14884
rect 7104 14841 7138 14875
rect 7138 14841 7156 14875
rect 7104 14832 7156 14841
rect 9680 14900 9732 14952
rect 10232 14900 10284 14952
rect 12072 14968 12124 15020
rect 14924 14968 14976 15020
rect 18328 14968 18380 15020
rect 20168 14968 20220 15020
rect 21916 14968 21968 15020
rect 10784 14900 10836 14952
rect 9588 14832 9640 14884
rect 9956 14832 10008 14884
rect 1400 14807 1452 14816
rect 1400 14773 1409 14807
rect 1409 14773 1443 14807
rect 1443 14773 1452 14807
rect 1400 14764 1452 14773
rect 2964 14764 3016 14816
rect 3700 14764 3752 14816
rect 4988 14764 5040 14816
rect 6000 14807 6052 14816
rect 6000 14773 6009 14807
rect 6009 14773 6043 14807
rect 6043 14773 6052 14807
rect 6000 14764 6052 14773
rect 6184 14764 6236 14816
rect 8208 14807 8260 14816
rect 8208 14773 8217 14807
rect 8217 14773 8251 14807
rect 8251 14773 8260 14807
rect 8208 14764 8260 14773
rect 11796 14900 11848 14952
rect 13544 14900 13596 14952
rect 17960 14900 18012 14952
rect 18236 14943 18288 14952
rect 18236 14909 18245 14943
rect 18245 14909 18279 14943
rect 18279 14909 18288 14943
rect 18236 14900 18288 14909
rect 19248 14900 19300 14952
rect 19616 14900 19668 14952
rect 19984 14900 20036 14952
rect 20720 14900 20772 14952
rect 21732 14900 21784 14952
rect 12808 14832 12860 14884
rect 13268 14832 13320 14884
rect 14188 14832 14240 14884
rect 18788 14832 18840 14884
rect 23020 14900 23072 14952
rect 11244 14764 11296 14816
rect 11428 14764 11480 14816
rect 11612 14764 11664 14816
rect 12992 14807 13044 14816
rect 12992 14773 13001 14807
rect 13001 14773 13035 14807
rect 13035 14773 13044 14807
rect 12992 14764 13044 14773
rect 14832 14807 14884 14816
rect 14832 14773 14841 14807
rect 14841 14773 14875 14807
rect 14875 14773 14884 14807
rect 14832 14764 14884 14773
rect 15476 14764 15528 14816
rect 15568 14764 15620 14816
rect 16212 14764 16264 14816
rect 18604 14764 18656 14816
rect 19616 14764 19668 14816
rect 21456 14807 21508 14816
rect 21456 14773 21465 14807
rect 21465 14773 21499 14807
rect 21499 14773 21508 14807
rect 21456 14764 21508 14773
rect 21732 14764 21784 14816
rect 8379 14662 8431 14714
rect 8443 14662 8495 14714
rect 8507 14662 8559 14714
rect 8571 14662 8623 14714
rect 15776 14662 15828 14714
rect 15840 14662 15892 14714
rect 15904 14662 15956 14714
rect 15968 14662 16020 14714
rect 1860 14560 1912 14612
rect 3056 14603 3108 14612
rect 3056 14569 3065 14603
rect 3065 14569 3099 14603
rect 3099 14569 3108 14603
rect 3056 14560 3108 14569
rect 4068 14603 4120 14612
rect 1492 14424 1544 14476
rect 2872 14492 2924 14544
rect 4068 14569 4077 14603
rect 4077 14569 4111 14603
rect 4111 14569 4120 14603
rect 4068 14560 4120 14569
rect 9956 14560 10008 14612
rect 5264 14424 5316 14476
rect 5356 14424 5408 14476
rect 6460 14424 6512 14476
rect 8208 14424 8260 14476
rect 9864 14492 9916 14544
rect 10048 14492 10100 14544
rect 10508 14492 10560 14544
rect 11336 14560 11388 14612
rect 11980 14560 12032 14612
rect 12624 14560 12676 14612
rect 14096 14560 14148 14612
rect 14924 14603 14976 14612
rect 14924 14569 14933 14603
rect 14933 14569 14967 14603
rect 14967 14569 14976 14603
rect 14924 14560 14976 14569
rect 19156 14560 19208 14612
rect 19800 14560 19852 14612
rect 11704 14492 11756 14544
rect 3056 14356 3108 14408
rect 4712 14356 4764 14408
rect 10416 14424 10468 14476
rect 6460 14288 6512 14340
rect 4344 14220 4396 14272
rect 4988 14220 5040 14272
rect 9036 14356 9088 14408
rect 9588 14356 9640 14408
rect 10968 14356 11020 14408
rect 12532 14492 12584 14544
rect 12808 14492 12860 14544
rect 13084 14492 13136 14544
rect 19984 14492 20036 14544
rect 21640 14560 21692 14612
rect 15660 14424 15712 14476
rect 17592 14424 17644 14476
rect 17776 14467 17828 14476
rect 17776 14433 17810 14467
rect 17810 14433 17828 14467
rect 17776 14424 17828 14433
rect 19156 14467 19208 14476
rect 19156 14433 19183 14467
rect 19183 14433 19208 14467
rect 19156 14424 19208 14433
rect 19340 14467 19392 14476
rect 19340 14433 19347 14467
rect 19347 14433 19381 14467
rect 19381 14433 19392 14467
rect 19340 14424 19392 14433
rect 12440 14399 12492 14408
rect 9772 14288 9824 14340
rect 11244 14331 11296 14340
rect 11244 14297 11253 14331
rect 11253 14297 11287 14331
rect 11287 14297 11296 14331
rect 11244 14288 11296 14297
rect 11428 14288 11480 14340
rect 12440 14365 12449 14399
rect 12449 14365 12483 14399
rect 12483 14365 12492 14399
rect 12440 14356 12492 14365
rect 14648 14356 14700 14408
rect 16212 14399 16264 14408
rect 16212 14365 16221 14399
rect 16221 14365 16255 14399
rect 16255 14365 16264 14399
rect 16212 14356 16264 14365
rect 6828 14220 6880 14272
rect 7012 14220 7064 14272
rect 8668 14220 8720 14272
rect 10048 14220 10100 14272
rect 11888 14220 11940 14272
rect 13728 14220 13780 14272
rect 13912 14263 13964 14272
rect 13912 14229 13921 14263
rect 13921 14229 13955 14263
rect 13955 14229 13964 14263
rect 15752 14263 15804 14272
rect 13912 14220 13964 14229
rect 15752 14229 15761 14263
rect 15761 14229 15795 14263
rect 15795 14229 15804 14263
rect 15752 14220 15804 14229
rect 21548 14492 21600 14544
rect 18512 14288 18564 14340
rect 19616 14288 19668 14340
rect 19984 14288 20036 14340
rect 20996 14288 21048 14340
rect 17224 14220 17276 14272
rect 18880 14263 18932 14272
rect 18880 14229 18889 14263
rect 18889 14229 18923 14263
rect 18923 14229 18932 14263
rect 18880 14220 18932 14229
rect 19340 14220 19392 14272
rect 21916 14220 21968 14272
rect 4680 14118 4732 14170
rect 4744 14118 4796 14170
rect 4808 14118 4860 14170
rect 4872 14118 4924 14170
rect 12078 14118 12130 14170
rect 12142 14118 12194 14170
rect 12206 14118 12258 14170
rect 12270 14118 12322 14170
rect 19475 14118 19527 14170
rect 19539 14118 19591 14170
rect 19603 14118 19655 14170
rect 19667 14118 19719 14170
rect 2872 14059 2924 14068
rect 2872 14025 2881 14059
rect 2881 14025 2915 14059
rect 2915 14025 2924 14059
rect 2872 14016 2924 14025
rect 4252 14016 4304 14068
rect 7380 14016 7432 14068
rect 8668 14016 8720 14068
rect 9220 14016 9272 14068
rect 9680 14059 9732 14068
rect 9680 14025 9689 14059
rect 9689 14025 9723 14059
rect 9723 14025 9732 14059
rect 9680 14016 9732 14025
rect 10508 14016 10560 14068
rect 11612 14016 11664 14068
rect 11888 14016 11940 14068
rect 17776 14016 17828 14068
rect 17868 14016 17920 14068
rect 20720 14016 20772 14068
rect 6460 13948 6512 14000
rect 1492 13923 1544 13932
rect 1492 13889 1501 13923
rect 1501 13889 1535 13923
rect 1535 13889 1544 13923
rect 1492 13880 1544 13889
rect 3700 13923 3752 13932
rect 3700 13889 3709 13923
rect 3709 13889 3743 13923
rect 3743 13889 3752 13923
rect 3700 13880 3752 13889
rect 4068 13744 4120 13796
rect 4528 13744 4580 13796
rect 3148 13719 3200 13728
rect 3148 13685 3157 13719
rect 3157 13685 3191 13719
rect 3191 13685 3200 13719
rect 3148 13676 3200 13685
rect 7196 13880 7248 13932
rect 7748 13880 7800 13932
rect 9772 13880 9824 13932
rect 10692 13948 10744 14000
rect 19616 13948 19668 14000
rect 4988 13812 5040 13864
rect 5724 13812 5776 13864
rect 6276 13812 6328 13864
rect 6460 13812 6512 13864
rect 8208 13812 8260 13864
rect 6276 13719 6328 13728
rect 6276 13685 6285 13719
rect 6285 13685 6319 13719
rect 6319 13685 6328 13719
rect 6276 13676 6328 13685
rect 6736 13676 6788 13728
rect 7196 13719 7248 13728
rect 7196 13685 7205 13719
rect 7205 13685 7239 13719
rect 7239 13685 7248 13719
rect 7196 13676 7248 13685
rect 7288 13719 7340 13728
rect 7288 13685 7297 13719
rect 7297 13685 7331 13719
rect 7331 13685 7340 13719
rect 11428 13880 11480 13932
rect 11612 13923 11664 13932
rect 11612 13889 11621 13923
rect 11621 13889 11655 13923
rect 11655 13889 11664 13923
rect 11612 13880 11664 13889
rect 18880 13923 18932 13932
rect 18880 13889 18889 13923
rect 18889 13889 18923 13923
rect 18923 13889 18932 13923
rect 18880 13880 18932 13889
rect 19248 13880 19300 13932
rect 11336 13855 11388 13864
rect 9220 13744 9272 13796
rect 10048 13744 10100 13796
rect 7288 13676 7340 13685
rect 9496 13676 9548 13728
rect 11336 13821 11345 13855
rect 11345 13821 11379 13855
rect 11379 13821 11388 13855
rect 11336 13812 11388 13821
rect 11060 13744 11112 13796
rect 12440 13812 12492 13864
rect 13084 13855 13136 13864
rect 13084 13821 13118 13855
rect 13118 13821 13136 13855
rect 13084 13812 13136 13821
rect 13544 13744 13596 13796
rect 17592 13812 17644 13864
rect 19156 13812 19208 13864
rect 19800 13880 19852 13932
rect 22836 13880 22888 13932
rect 14648 13744 14700 13796
rect 14924 13744 14976 13796
rect 15016 13744 15068 13796
rect 13820 13676 13872 13728
rect 15384 13676 15436 13728
rect 17408 13744 17460 13796
rect 19340 13744 19392 13796
rect 21456 13812 21508 13864
rect 21732 13744 21784 13796
rect 18052 13676 18104 13728
rect 20996 13676 21048 13728
rect 22100 13719 22152 13728
rect 22100 13685 22109 13719
rect 22109 13685 22143 13719
rect 22143 13685 22152 13719
rect 22100 13676 22152 13685
rect 8379 13574 8431 13626
rect 8443 13574 8495 13626
rect 8507 13574 8559 13626
rect 8571 13574 8623 13626
rect 15776 13574 15828 13626
rect 15840 13574 15892 13626
rect 15904 13574 15956 13626
rect 15968 13574 16020 13626
rect 1400 13472 1452 13524
rect 3148 13472 3200 13524
rect 5356 13472 5408 13524
rect 5724 13472 5776 13524
rect 4988 13404 5040 13456
rect 6920 13472 6972 13524
rect 7380 13472 7432 13524
rect 9312 13515 9364 13524
rect 9312 13481 9321 13515
rect 9321 13481 9355 13515
rect 9355 13481 9364 13515
rect 9312 13472 9364 13481
rect 6276 13447 6328 13456
rect 6276 13413 6285 13447
rect 6285 13413 6319 13447
rect 6319 13413 6328 13447
rect 6276 13404 6328 13413
rect 7012 13447 7064 13456
rect 7012 13413 7046 13447
rect 7046 13413 7064 13447
rect 7012 13404 7064 13413
rect 7196 13404 7248 13456
rect 8944 13404 8996 13456
rect 10784 13472 10836 13524
rect 11796 13404 11848 13456
rect 1676 13379 1728 13388
rect 1676 13345 1685 13379
rect 1685 13345 1719 13379
rect 1719 13345 1728 13379
rect 1676 13336 1728 13345
rect 7288 13336 7340 13388
rect 8484 13336 8536 13388
rect 9312 13336 9364 13388
rect 11704 13336 11756 13388
rect 12164 13379 12216 13388
rect 12164 13345 12173 13379
rect 12173 13345 12207 13379
rect 12207 13345 12216 13379
rect 12164 13336 12216 13345
rect 2688 13268 2740 13320
rect 4344 13268 4396 13320
rect 6736 13311 6788 13320
rect 6736 13277 6745 13311
rect 6745 13277 6779 13311
rect 6779 13277 6788 13311
rect 6736 13268 6788 13277
rect 1860 13243 1912 13252
rect 1860 13209 1869 13243
rect 1869 13209 1903 13243
rect 1903 13209 1912 13243
rect 1860 13200 1912 13209
rect 5540 13200 5592 13252
rect 8944 13311 8996 13320
rect 8944 13277 8953 13311
rect 8953 13277 8987 13311
rect 8987 13277 8996 13311
rect 8944 13268 8996 13277
rect 10600 13268 10652 13320
rect 10692 13311 10744 13320
rect 10692 13277 10701 13311
rect 10701 13277 10735 13311
rect 10735 13277 10744 13311
rect 13728 13404 13780 13456
rect 13820 13404 13872 13456
rect 18880 13404 18932 13456
rect 19616 13472 19668 13524
rect 22100 13472 22152 13524
rect 20168 13404 20220 13456
rect 21916 13404 21968 13456
rect 13452 13336 13504 13388
rect 14188 13336 14240 13388
rect 14924 13336 14976 13388
rect 15844 13336 15896 13388
rect 16304 13336 16356 13388
rect 18512 13336 18564 13388
rect 20352 13336 20404 13388
rect 10692 13268 10744 13277
rect 3240 13132 3292 13184
rect 4344 13132 4396 13184
rect 10508 13200 10560 13252
rect 11980 13200 12032 13252
rect 8116 13175 8168 13184
rect 8116 13141 8125 13175
rect 8125 13141 8159 13175
rect 8159 13141 8168 13175
rect 8116 13132 8168 13141
rect 10048 13132 10100 13184
rect 14648 13132 14700 13184
rect 17684 13268 17736 13320
rect 16948 13200 17000 13252
rect 17868 13200 17920 13252
rect 17408 13132 17460 13184
rect 17684 13132 17736 13184
rect 19340 13243 19392 13252
rect 19340 13209 19349 13243
rect 19349 13209 19383 13243
rect 19383 13209 19392 13243
rect 20996 13268 21048 13320
rect 19340 13200 19392 13209
rect 18604 13132 18656 13184
rect 19800 13132 19852 13184
rect 22836 13132 22888 13184
rect 4680 13030 4732 13082
rect 4744 13030 4796 13082
rect 4808 13030 4860 13082
rect 4872 13030 4924 13082
rect 12078 13030 12130 13082
rect 12142 13030 12194 13082
rect 12206 13030 12258 13082
rect 12270 13030 12322 13082
rect 19475 13030 19527 13082
rect 19539 13030 19591 13082
rect 19603 13030 19655 13082
rect 19667 13030 19719 13082
rect 4344 12928 4396 12980
rect 4988 12971 5040 12980
rect 4988 12937 4997 12971
rect 4997 12937 5031 12971
rect 5031 12937 5040 12971
rect 4988 12928 5040 12937
rect 5356 12860 5408 12912
rect 9128 12928 9180 12980
rect 10324 12928 10376 12980
rect 11704 12971 11756 12980
rect 11704 12937 11713 12971
rect 11713 12937 11747 12971
rect 11747 12937 11756 12971
rect 11704 12928 11756 12937
rect 11336 12860 11388 12912
rect 8484 12792 8536 12844
rect 8944 12792 8996 12844
rect 9680 12792 9732 12844
rect 16396 12928 16448 12980
rect 20628 12928 20680 12980
rect 14004 12903 14056 12912
rect 14004 12869 14013 12903
rect 14013 12869 14047 12903
rect 14047 12869 14056 12903
rect 14004 12860 14056 12869
rect 16304 12860 16356 12912
rect 1584 12724 1636 12776
rect 4344 12724 4396 12776
rect 5540 12724 5592 12776
rect 2964 12656 3016 12708
rect 2872 12588 2924 12640
rect 4436 12656 4488 12708
rect 6828 12767 6880 12776
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 3424 12588 3476 12640
rect 7472 12656 7524 12708
rect 10508 12656 10560 12708
rect 11704 12724 11756 12776
rect 11888 12767 11940 12776
rect 11888 12733 11897 12767
rect 11897 12733 11931 12767
rect 11931 12733 11940 12767
rect 11888 12724 11940 12733
rect 11980 12724 12032 12776
rect 12440 12724 12492 12776
rect 13360 12724 13412 12776
rect 11520 12656 11572 12708
rect 7380 12588 7432 12640
rect 8852 12631 8904 12640
rect 8852 12597 8861 12631
rect 8861 12597 8895 12631
rect 8895 12597 8904 12631
rect 8852 12588 8904 12597
rect 8944 12631 8996 12640
rect 8944 12597 8953 12631
rect 8953 12597 8987 12631
rect 8987 12597 8996 12631
rect 8944 12588 8996 12597
rect 9128 12588 9180 12640
rect 9956 12631 10008 12640
rect 9956 12597 9965 12631
rect 9965 12597 9999 12631
rect 9999 12597 10008 12631
rect 9956 12588 10008 12597
rect 10324 12588 10376 12640
rect 10692 12588 10744 12640
rect 11888 12588 11940 12640
rect 11980 12588 12032 12640
rect 13268 12656 13320 12708
rect 13728 12656 13780 12708
rect 14372 12724 14424 12776
rect 14924 12724 14976 12776
rect 17868 12860 17920 12912
rect 18236 12903 18288 12912
rect 18236 12869 18245 12903
rect 18245 12869 18279 12903
rect 18279 12869 18288 12903
rect 18236 12860 18288 12869
rect 22192 12860 22244 12912
rect 16856 12792 16908 12844
rect 17132 12792 17184 12844
rect 15384 12656 15436 12708
rect 13912 12588 13964 12640
rect 14924 12588 14976 12640
rect 17868 12767 17920 12776
rect 17868 12733 17877 12767
rect 17877 12733 17911 12767
rect 17911 12733 17920 12767
rect 17868 12724 17920 12733
rect 20904 12792 20956 12844
rect 21732 12792 21784 12844
rect 22008 12792 22060 12844
rect 18604 12767 18656 12776
rect 18604 12733 18613 12767
rect 18613 12733 18647 12767
rect 18647 12733 18656 12767
rect 18604 12724 18656 12733
rect 19340 12724 19392 12776
rect 20168 12724 20220 12776
rect 16580 12588 16632 12640
rect 17224 12588 17276 12640
rect 17868 12588 17920 12640
rect 18696 12656 18748 12708
rect 19708 12656 19760 12708
rect 20996 12656 21048 12708
rect 19984 12631 20036 12640
rect 19984 12597 19993 12631
rect 19993 12597 20027 12631
rect 20027 12597 20036 12631
rect 19984 12588 20036 12597
rect 20352 12588 20404 12640
rect 22744 12588 22796 12640
rect 8379 12486 8431 12538
rect 8443 12486 8495 12538
rect 8507 12486 8559 12538
rect 8571 12486 8623 12538
rect 15776 12486 15828 12538
rect 15840 12486 15892 12538
rect 15904 12486 15956 12538
rect 15968 12486 16020 12538
rect 2964 12427 3016 12436
rect 2964 12393 2973 12427
rect 2973 12393 3007 12427
rect 3007 12393 3016 12427
rect 2964 12384 3016 12393
rect 4436 12427 4488 12436
rect 4436 12393 4445 12427
rect 4445 12393 4479 12427
rect 4479 12393 4488 12427
rect 4436 12384 4488 12393
rect 6920 12384 6972 12436
rect 5540 12316 5592 12368
rect 5816 12359 5868 12368
rect 5816 12325 5825 12359
rect 5825 12325 5859 12359
rect 5859 12325 5868 12359
rect 5816 12316 5868 12325
rect 1584 12291 1636 12300
rect 1584 12257 1593 12291
rect 1593 12257 1627 12291
rect 1627 12257 1636 12291
rect 1584 12248 1636 12257
rect 2780 12248 2832 12300
rect 5080 12248 5132 12300
rect 6644 12316 6696 12368
rect 6828 12316 6880 12368
rect 8208 12384 8260 12436
rect 9128 12384 9180 12436
rect 9312 12384 9364 12436
rect 9864 12384 9916 12436
rect 7380 12316 7432 12368
rect 7748 12316 7800 12368
rect 8024 12316 8076 12368
rect 11428 12384 11480 12436
rect 13452 12384 13504 12436
rect 14096 12384 14148 12436
rect 14740 12384 14792 12436
rect 2964 12180 3016 12232
rect 5356 12180 5408 12232
rect 6368 12180 6420 12232
rect 9220 12248 9272 12300
rect 9772 12291 9824 12300
rect 9772 12257 9781 12291
rect 9781 12257 9815 12291
rect 9815 12257 9824 12291
rect 9772 12248 9824 12257
rect 3516 12112 3568 12164
rect 10968 12248 11020 12300
rect 15292 12316 15344 12368
rect 14004 12248 14056 12300
rect 13176 12180 13228 12232
rect 4068 12087 4120 12096
rect 4068 12053 4077 12087
rect 4077 12053 4111 12087
rect 4111 12053 4120 12087
rect 4068 12044 4120 12053
rect 4436 12044 4488 12096
rect 5356 12087 5408 12096
rect 5356 12053 5365 12087
rect 5365 12053 5399 12087
rect 5399 12053 5408 12087
rect 5356 12044 5408 12053
rect 8392 12087 8444 12096
rect 8392 12053 8401 12087
rect 8401 12053 8435 12087
rect 8435 12053 8444 12087
rect 8392 12044 8444 12053
rect 8576 12044 8628 12096
rect 9680 12044 9732 12096
rect 12532 12044 12584 12096
rect 14280 12180 14332 12232
rect 15476 12291 15528 12300
rect 15476 12257 15485 12291
rect 15485 12257 15519 12291
rect 15519 12257 15528 12291
rect 15476 12248 15528 12257
rect 15660 12427 15712 12436
rect 15660 12393 15669 12427
rect 15669 12393 15703 12427
rect 15703 12393 15712 12427
rect 16396 12427 16448 12436
rect 15660 12384 15712 12393
rect 16396 12393 16405 12427
rect 16405 12393 16439 12427
rect 16439 12393 16448 12427
rect 16396 12384 16448 12393
rect 15752 12248 15804 12300
rect 17224 12248 17276 12300
rect 17868 12316 17920 12368
rect 19892 12316 19944 12368
rect 18696 12248 18748 12300
rect 19340 12248 19392 12300
rect 19800 12291 19852 12300
rect 19800 12257 19809 12291
rect 19809 12257 19843 12291
rect 19843 12257 19852 12291
rect 19800 12248 19852 12257
rect 20444 12316 20496 12368
rect 20996 12248 21048 12300
rect 21180 12291 21232 12300
rect 21180 12257 21214 12291
rect 21214 12257 21232 12291
rect 21180 12248 21232 12257
rect 15476 12112 15528 12164
rect 19892 12223 19944 12232
rect 19892 12189 19901 12223
rect 19901 12189 19935 12223
rect 19935 12189 19944 12223
rect 19892 12180 19944 12189
rect 19984 12223 20036 12232
rect 19984 12189 19993 12223
rect 19993 12189 20027 12223
rect 20027 12189 20036 12223
rect 19984 12180 20036 12189
rect 20168 12180 20220 12232
rect 22560 12223 22612 12232
rect 22560 12189 22569 12223
rect 22569 12189 22603 12223
rect 22603 12189 22612 12223
rect 22560 12180 22612 12189
rect 18788 12112 18840 12164
rect 14188 12044 14240 12096
rect 15292 12044 15344 12096
rect 21640 12044 21692 12096
rect 21824 12044 21876 12096
rect 22008 12044 22060 12096
rect 4680 11942 4732 11994
rect 4744 11942 4796 11994
rect 4808 11942 4860 11994
rect 4872 11942 4924 11994
rect 12078 11942 12130 11994
rect 12142 11942 12194 11994
rect 12206 11942 12258 11994
rect 12270 11942 12322 11994
rect 19475 11942 19527 11994
rect 19539 11942 19591 11994
rect 19603 11942 19655 11994
rect 19667 11942 19719 11994
rect 3332 11704 3384 11756
rect 4344 11772 4396 11824
rect 4436 11704 4488 11756
rect 4712 11747 4764 11756
rect 4712 11713 4721 11747
rect 4721 11713 4755 11747
rect 4755 11713 4764 11747
rect 4712 11704 4764 11713
rect 6368 11772 6420 11824
rect 10692 11840 10744 11892
rect 11704 11883 11756 11892
rect 11704 11849 11713 11883
rect 11713 11849 11747 11883
rect 11747 11849 11756 11883
rect 11704 11840 11756 11849
rect 12624 11840 12676 11892
rect 12808 11840 12860 11892
rect 13176 11840 13228 11892
rect 14004 11840 14056 11892
rect 14188 11840 14240 11892
rect 14832 11840 14884 11892
rect 14924 11840 14976 11892
rect 15200 11840 15252 11892
rect 16120 11840 16172 11892
rect 16764 11840 16816 11892
rect 17316 11840 17368 11892
rect 20904 11883 20956 11892
rect 9772 11772 9824 11824
rect 11612 11772 11664 11824
rect 12532 11772 12584 11824
rect 16396 11772 16448 11824
rect 16672 11772 16724 11824
rect 6828 11704 6880 11756
rect 8668 11704 8720 11756
rect 8852 11704 8904 11756
rect 9864 11747 9916 11756
rect 9864 11713 9873 11747
rect 9873 11713 9907 11747
rect 9907 11713 9916 11747
rect 9864 11704 9916 11713
rect 10324 11747 10376 11756
rect 10324 11713 10333 11747
rect 10333 11713 10367 11747
rect 10367 11713 10376 11747
rect 10324 11704 10376 11713
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 2964 11636 3016 11688
rect 4896 11636 4948 11688
rect 9036 11679 9088 11688
rect 9036 11645 9045 11679
rect 9045 11645 9079 11679
rect 9079 11645 9088 11679
rect 9036 11636 9088 11645
rect 10968 11636 11020 11688
rect 11980 11679 12032 11688
rect 11980 11645 11989 11679
rect 11989 11645 12023 11679
rect 12023 11645 12032 11679
rect 11980 11636 12032 11645
rect 14832 11679 14884 11688
rect 14832 11645 14841 11679
rect 14841 11645 14875 11679
rect 14875 11645 14884 11679
rect 14832 11636 14884 11645
rect 15660 11704 15712 11756
rect 16028 11704 16080 11756
rect 17500 11747 17552 11756
rect 17500 11713 17509 11747
rect 17509 11713 17543 11747
rect 17543 11713 17552 11747
rect 17500 11704 17552 11713
rect 18696 11747 18748 11756
rect 18696 11713 18705 11747
rect 18705 11713 18739 11747
rect 18739 11713 18748 11747
rect 20904 11849 20913 11883
rect 20913 11849 20947 11883
rect 20947 11849 20956 11883
rect 20904 11840 20956 11849
rect 18696 11704 18748 11713
rect 19248 11704 19300 11756
rect 19708 11704 19760 11756
rect 16764 11636 16816 11688
rect 18604 11636 18656 11688
rect 19064 11679 19116 11688
rect 19064 11645 19073 11679
rect 19073 11645 19107 11679
rect 19107 11645 19116 11679
rect 19064 11636 19116 11645
rect 19892 11636 19944 11688
rect 21272 11636 21324 11688
rect 2780 11543 2832 11552
rect 2780 11509 2789 11543
rect 2789 11509 2823 11543
rect 2823 11509 2832 11543
rect 6920 11568 6972 11620
rect 7472 11611 7524 11620
rect 7472 11577 7506 11611
rect 7506 11577 7524 11611
rect 7472 11568 7524 11577
rect 8392 11568 8444 11620
rect 11796 11568 11848 11620
rect 13176 11568 13228 11620
rect 14648 11568 14700 11620
rect 18696 11568 18748 11620
rect 22652 11568 22704 11620
rect 2780 11500 2832 11509
rect 3056 11543 3108 11552
rect 3056 11509 3065 11543
rect 3065 11509 3099 11543
rect 3099 11509 3108 11543
rect 3424 11543 3476 11552
rect 3056 11500 3108 11509
rect 3424 11509 3433 11543
rect 3433 11509 3467 11543
rect 3467 11509 3476 11543
rect 3424 11500 3476 11509
rect 3700 11500 3752 11552
rect 7840 11500 7892 11552
rect 8760 11500 8812 11552
rect 9036 11500 9088 11552
rect 11428 11500 11480 11552
rect 11612 11500 11664 11552
rect 16120 11500 16172 11552
rect 16396 11543 16448 11552
rect 16396 11509 16405 11543
rect 16405 11509 16439 11543
rect 16439 11509 16448 11543
rect 16948 11543 17000 11552
rect 16396 11500 16448 11509
rect 16948 11509 16957 11543
rect 16957 11509 16991 11543
rect 16991 11509 17000 11543
rect 16948 11500 17000 11509
rect 18052 11543 18104 11552
rect 18052 11509 18061 11543
rect 18061 11509 18095 11543
rect 18095 11509 18104 11543
rect 18052 11500 18104 11509
rect 19340 11500 19392 11552
rect 19432 11500 19484 11552
rect 20076 11500 20128 11552
rect 8379 11398 8431 11450
rect 8443 11398 8495 11450
rect 8507 11398 8559 11450
rect 8571 11398 8623 11450
rect 15776 11398 15828 11450
rect 15840 11398 15892 11450
rect 15904 11398 15956 11450
rect 15968 11398 16020 11450
rect 2964 11296 3016 11348
rect 3148 11296 3200 11348
rect 3424 11296 3476 11348
rect 4068 11296 4120 11348
rect 3148 11160 3200 11212
rect 3516 11228 3568 11280
rect 5816 11296 5868 11348
rect 7748 11296 7800 11348
rect 10416 11296 10468 11348
rect 11796 11339 11848 11348
rect 11796 11305 11805 11339
rect 11805 11305 11839 11339
rect 11839 11305 11848 11339
rect 11796 11296 11848 11305
rect 14280 11296 14332 11348
rect 15200 11296 15252 11348
rect 3424 11203 3476 11212
rect 3424 11169 3433 11203
rect 3433 11169 3467 11203
rect 3467 11169 3476 11203
rect 4436 11203 4488 11212
rect 3424 11160 3476 11169
rect 4436 11169 4445 11203
rect 4445 11169 4479 11203
rect 4479 11169 4488 11203
rect 4436 11160 4488 11169
rect 4896 11160 4948 11212
rect 6460 11160 6512 11212
rect 6644 11160 6696 11212
rect 7840 11160 7892 11212
rect 7932 11160 7984 11212
rect 11060 11228 11112 11280
rect 11704 11228 11756 11280
rect 17224 11296 17276 11348
rect 19432 11296 19484 11348
rect 19892 11296 19944 11348
rect 20260 11296 20312 11348
rect 22100 11296 22152 11348
rect 22284 11296 22336 11348
rect 22652 11339 22704 11348
rect 22652 11305 22661 11339
rect 22661 11305 22695 11339
rect 22695 11305 22704 11339
rect 22652 11296 22704 11305
rect 9680 11160 9732 11212
rect 10048 11160 10100 11212
rect 10324 11160 10376 11212
rect 11428 11160 11480 11212
rect 11520 11160 11572 11212
rect 12440 11160 12492 11212
rect 14004 11160 14056 11212
rect 14372 11160 14424 11212
rect 15936 11203 15988 11212
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 4160 11092 4212 11144
rect 4712 11135 4764 11144
rect 4712 11101 4721 11135
rect 4721 11101 4755 11135
rect 4755 11101 4764 11135
rect 4712 11092 4764 11101
rect 6828 11135 6880 11144
rect 6828 11101 6837 11135
rect 6837 11101 6871 11135
rect 6871 11101 6880 11135
rect 6828 11092 6880 11101
rect 8668 11092 8720 11144
rect 4344 11024 4396 11076
rect 3516 10956 3568 11008
rect 5540 10956 5592 11008
rect 8576 10956 8628 11008
rect 9956 11024 10008 11076
rect 10048 10956 10100 11008
rect 10232 10956 10284 11008
rect 15936 11169 15959 11203
rect 15959 11169 15988 11203
rect 15936 11160 15988 11169
rect 17224 11160 17276 11212
rect 17868 11160 17920 11212
rect 19064 11160 19116 11212
rect 19340 11160 19392 11212
rect 15200 11092 15252 11144
rect 17684 11135 17736 11144
rect 17684 11101 17693 11135
rect 17693 11101 17727 11135
rect 17727 11101 17736 11135
rect 17684 11092 17736 11101
rect 18420 11135 18472 11144
rect 18420 11101 18432 11135
rect 18432 11101 18466 11135
rect 18466 11101 18472 11135
rect 18420 11092 18472 11101
rect 18604 11092 18656 11144
rect 12992 10956 13044 11008
rect 13728 10956 13780 11008
rect 13912 10956 13964 11008
rect 14280 10956 14332 11008
rect 17224 10956 17276 11008
rect 21824 11228 21876 11280
rect 20260 11203 20312 11212
rect 20260 11169 20269 11203
rect 20269 11169 20303 11203
rect 20303 11169 20312 11203
rect 20260 11160 20312 11169
rect 20720 11092 20772 11144
rect 21272 11135 21324 11144
rect 21272 11101 21281 11135
rect 21281 11101 21315 11135
rect 21315 11101 21324 11135
rect 21272 11092 21324 11101
rect 20352 11024 20404 11076
rect 4680 10854 4732 10906
rect 4744 10854 4796 10906
rect 4808 10854 4860 10906
rect 4872 10854 4924 10906
rect 12078 10854 12130 10906
rect 12142 10854 12194 10906
rect 12206 10854 12258 10906
rect 12270 10854 12322 10906
rect 19475 10854 19527 10906
rect 19539 10854 19591 10906
rect 19603 10854 19655 10906
rect 19667 10854 19719 10906
rect 3148 10795 3200 10804
rect 3148 10761 3157 10795
rect 3157 10761 3191 10795
rect 3191 10761 3200 10795
rect 3148 10752 3200 10761
rect 4436 10752 4488 10804
rect 6460 10795 6512 10804
rect 6460 10761 6469 10795
rect 6469 10761 6503 10795
rect 6503 10761 6512 10795
rect 6460 10752 6512 10761
rect 7288 10752 7340 10804
rect 1400 10548 1452 10600
rect 3332 10548 3384 10600
rect 3516 10548 3568 10600
rect 4160 10548 4212 10600
rect 2136 10480 2188 10532
rect 5540 10480 5592 10532
rect 6276 10548 6328 10600
rect 6644 10480 6696 10532
rect 3608 10412 3660 10464
rect 8576 10752 8628 10804
rect 9496 10752 9548 10804
rect 9680 10727 9732 10736
rect 9680 10693 9689 10727
rect 9689 10693 9723 10727
rect 9723 10693 9732 10727
rect 9680 10684 9732 10693
rect 9864 10684 9916 10736
rect 10324 10752 10376 10804
rect 10692 10752 10744 10804
rect 11796 10752 11848 10804
rect 12440 10684 12492 10736
rect 15200 10684 15252 10736
rect 17684 10752 17736 10804
rect 18420 10752 18472 10804
rect 21180 10752 21232 10804
rect 19064 10684 19116 10736
rect 8760 10548 8812 10600
rect 9772 10548 9824 10600
rect 7748 10523 7800 10532
rect 7748 10489 7782 10523
rect 7782 10489 7800 10523
rect 7748 10480 7800 10489
rect 9680 10480 9732 10532
rect 11152 10548 11204 10600
rect 12440 10548 12492 10600
rect 10232 10523 10284 10532
rect 10232 10489 10266 10523
rect 10266 10489 10284 10523
rect 10232 10480 10284 10489
rect 12624 10548 12676 10600
rect 14280 10548 14332 10600
rect 18052 10616 18104 10668
rect 18880 10659 18932 10668
rect 18880 10625 18889 10659
rect 18889 10625 18923 10659
rect 18923 10625 18932 10659
rect 18880 10616 18932 10625
rect 19156 10548 19208 10600
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 19708 10548 19760 10557
rect 19984 10591 20036 10600
rect 19984 10557 20018 10591
rect 20018 10557 20036 10591
rect 19984 10548 20036 10557
rect 21640 10548 21692 10600
rect 22376 10591 22428 10600
rect 22376 10557 22385 10591
rect 22385 10557 22419 10591
rect 22419 10557 22428 10591
rect 22376 10548 22428 10557
rect 8208 10412 8260 10464
rect 9404 10412 9456 10464
rect 10508 10412 10560 10464
rect 15936 10480 15988 10532
rect 16120 10523 16172 10532
rect 16120 10489 16154 10523
rect 16154 10489 16172 10523
rect 16120 10480 16172 10489
rect 16304 10480 16356 10532
rect 16580 10480 16632 10532
rect 17592 10480 17644 10532
rect 19800 10480 19852 10532
rect 14280 10412 14332 10464
rect 17684 10455 17736 10464
rect 17684 10421 17693 10455
rect 17693 10421 17727 10455
rect 17727 10421 17736 10455
rect 17684 10412 17736 10421
rect 20536 10412 20588 10464
rect 21456 10412 21508 10464
rect 8379 10310 8431 10362
rect 8443 10310 8495 10362
rect 8507 10310 8559 10362
rect 8571 10310 8623 10362
rect 15776 10310 15828 10362
rect 15840 10310 15892 10362
rect 15904 10310 15956 10362
rect 15968 10310 16020 10362
rect 1768 10208 1820 10260
rect 4804 10208 4856 10260
rect 5540 10251 5592 10260
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 6920 10208 6972 10260
rect 9312 10208 9364 10260
rect 10232 10208 10284 10260
rect 2136 10140 2188 10192
rect 4436 10183 4488 10192
rect 4436 10149 4470 10183
rect 4470 10149 4488 10183
rect 4436 10140 4488 10149
rect 5816 10140 5868 10192
rect 7564 10140 7616 10192
rect 8300 10140 8352 10192
rect 8392 10140 8444 10192
rect 8944 10140 8996 10192
rect 9864 10140 9916 10192
rect 11704 10140 11756 10192
rect 12348 10140 12400 10192
rect 13176 10208 13228 10260
rect 14004 10208 14056 10260
rect 14556 10251 14608 10260
rect 14556 10217 14565 10251
rect 14565 10217 14599 10251
rect 14599 10217 14608 10251
rect 14556 10208 14608 10217
rect 14648 10208 14700 10260
rect 16120 10208 16172 10260
rect 17316 10208 17368 10260
rect 18420 10208 18472 10260
rect 18696 10208 18748 10260
rect 21732 10208 21784 10260
rect 22284 10251 22336 10260
rect 22284 10217 22293 10251
rect 22293 10217 22327 10251
rect 22327 10217 22336 10251
rect 22284 10208 22336 10217
rect 2780 10072 2832 10124
rect 3516 10072 3568 10124
rect 6644 10072 6696 10124
rect 6920 10072 6972 10124
rect 8208 10115 8260 10124
rect 8208 10081 8231 10115
rect 8231 10081 8260 10115
rect 8208 10072 8260 10081
rect 10232 10072 10284 10124
rect 11796 10072 11848 10124
rect 14280 10140 14332 10192
rect 9680 10047 9732 10056
rect 3332 9868 3384 9920
rect 4068 9868 4120 9920
rect 4436 9868 4488 9920
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 12440 10004 12492 10056
rect 14924 10072 14976 10124
rect 15108 10115 15160 10124
rect 15108 10081 15117 10115
rect 15117 10081 15151 10115
rect 15151 10081 15160 10115
rect 15108 10072 15160 10081
rect 16396 10140 16448 10192
rect 17040 10072 17092 10124
rect 17592 10115 17644 10124
rect 17592 10081 17601 10115
rect 17601 10081 17635 10115
rect 17635 10081 17644 10115
rect 17592 10072 17644 10081
rect 17868 10072 17920 10124
rect 18236 10115 18288 10124
rect 18236 10081 18245 10115
rect 18245 10081 18279 10115
rect 18279 10081 18288 10115
rect 18236 10072 18288 10081
rect 14648 10004 14700 10056
rect 14740 10004 14792 10056
rect 19800 10140 19852 10192
rect 20444 10140 20496 10192
rect 18788 10072 18840 10124
rect 18880 10072 18932 10124
rect 19984 10072 20036 10124
rect 21272 10115 21324 10124
rect 21272 10081 21281 10115
rect 21281 10081 21315 10115
rect 21315 10081 21324 10115
rect 21272 10072 21324 10081
rect 19708 10004 19760 10056
rect 20720 10004 20772 10056
rect 22652 10004 22704 10056
rect 8944 9868 8996 9920
rect 9496 9868 9548 9920
rect 12992 9868 13044 9920
rect 14096 9868 14148 9920
rect 14924 9911 14976 9920
rect 14924 9877 14933 9911
rect 14933 9877 14967 9911
rect 14967 9877 14976 9911
rect 14924 9868 14976 9877
rect 15200 9868 15252 9920
rect 17224 9911 17276 9920
rect 17224 9877 17233 9911
rect 17233 9877 17267 9911
rect 17267 9877 17276 9911
rect 17224 9868 17276 9877
rect 20628 9936 20680 9988
rect 19340 9868 19392 9920
rect 20904 9868 20956 9920
rect 21732 9868 21784 9920
rect 4680 9766 4732 9818
rect 4744 9766 4796 9818
rect 4808 9766 4860 9818
rect 4872 9766 4924 9818
rect 12078 9766 12130 9818
rect 12142 9766 12194 9818
rect 12206 9766 12258 9818
rect 12270 9766 12322 9818
rect 19475 9766 19527 9818
rect 19539 9766 19591 9818
rect 19603 9766 19655 9818
rect 19667 9766 19719 9818
rect 2136 9664 2188 9716
rect 2780 9639 2832 9648
rect 2780 9605 2789 9639
rect 2789 9605 2823 9639
rect 2823 9605 2832 9639
rect 2780 9596 2832 9605
rect 4160 9596 4212 9648
rect 5816 9596 5868 9648
rect 7012 9664 7064 9716
rect 7932 9664 7984 9716
rect 8392 9664 8444 9716
rect 5264 9528 5316 9580
rect 5540 9528 5592 9580
rect 8668 9596 8720 9648
rect 3332 9503 3384 9512
rect 3332 9469 3366 9503
rect 3366 9469 3384 9503
rect 1492 9392 1544 9444
rect 3332 9460 3384 9469
rect 4896 9460 4948 9512
rect 9956 9664 10008 9716
rect 10324 9664 10376 9716
rect 11796 9664 11848 9716
rect 12532 9664 12584 9716
rect 10232 9596 10284 9648
rect 11428 9596 11480 9648
rect 12992 9664 13044 9716
rect 7012 9460 7064 9512
rect 3516 9392 3568 9444
rect 6460 9392 6512 9444
rect 6644 9392 6696 9444
rect 8484 9460 8536 9512
rect 2320 9324 2372 9376
rect 4804 9324 4856 9376
rect 5264 9324 5316 9376
rect 6368 9367 6420 9376
rect 6368 9333 6377 9367
rect 6377 9333 6411 9367
rect 6411 9333 6420 9367
rect 6368 9324 6420 9333
rect 7012 9324 7064 9376
rect 7288 9324 7340 9376
rect 8576 9392 8628 9444
rect 8944 9503 8996 9512
rect 8944 9469 8978 9503
rect 8978 9469 8996 9503
rect 8944 9460 8996 9469
rect 8760 9392 8812 9444
rect 9128 9392 9180 9444
rect 9772 9324 9824 9376
rect 12624 9528 12676 9580
rect 15108 9664 15160 9716
rect 14096 9639 14148 9648
rect 14096 9605 14105 9639
rect 14105 9605 14139 9639
rect 14139 9605 14148 9639
rect 14096 9596 14148 9605
rect 16396 9596 16448 9648
rect 14740 9528 14792 9580
rect 18604 9664 18656 9716
rect 17868 9596 17920 9648
rect 17776 9528 17828 9580
rect 12440 9460 12492 9512
rect 12532 9460 12584 9512
rect 10508 9392 10560 9444
rect 13268 9460 13320 9512
rect 15016 9460 15068 9512
rect 18696 9460 18748 9512
rect 14464 9392 14516 9444
rect 14740 9392 14792 9444
rect 19156 9571 19208 9580
rect 19156 9537 19165 9571
rect 19165 9537 19199 9571
rect 19199 9537 19208 9571
rect 19156 9528 19208 9537
rect 19708 9528 19760 9580
rect 19892 9571 19944 9580
rect 19892 9537 19901 9571
rect 19901 9537 19935 9571
rect 19935 9537 19944 9571
rect 19892 9528 19944 9537
rect 20720 9528 20772 9580
rect 18972 9460 19024 9512
rect 10416 9324 10468 9376
rect 11336 9324 11388 9376
rect 15016 9367 15068 9376
rect 15016 9333 15025 9367
rect 15025 9333 15059 9367
rect 15059 9333 15068 9367
rect 15016 9324 15068 9333
rect 19064 9392 19116 9444
rect 17316 9367 17368 9376
rect 17316 9333 17325 9367
rect 17325 9333 17359 9367
rect 17359 9333 17368 9367
rect 17316 9324 17368 9333
rect 17776 9324 17828 9376
rect 18144 9367 18196 9376
rect 18144 9333 18153 9367
rect 18153 9333 18187 9367
rect 18187 9333 18196 9367
rect 18144 9324 18196 9333
rect 18236 9324 18288 9376
rect 18604 9367 18656 9376
rect 18604 9333 18613 9367
rect 18613 9333 18647 9367
rect 18647 9333 18656 9367
rect 18604 9324 18656 9333
rect 18788 9324 18840 9376
rect 22652 9392 22704 9444
rect 8379 9222 8431 9274
rect 8443 9222 8495 9274
rect 8507 9222 8559 9274
rect 8571 9222 8623 9274
rect 15776 9222 15828 9274
rect 15840 9222 15892 9274
rect 15904 9222 15956 9274
rect 15968 9222 16020 9274
rect 2320 9163 2372 9172
rect 2320 9129 2329 9163
rect 2329 9129 2363 9163
rect 2363 9129 2372 9163
rect 2320 9120 2372 9129
rect 3332 9120 3384 9172
rect 3424 9120 3476 9172
rect 4344 9120 4396 9172
rect 5080 9163 5132 9172
rect 5080 9129 5089 9163
rect 5089 9129 5123 9163
rect 5123 9129 5132 9163
rect 5080 9120 5132 9129
rect 5356 9120 5408 9172
rect 2504 9052 2556 9104
rect 2780 8984 2832 9036
rect 3976 9052 4028 9104
rect 5264 9052 5316 9104
rect 4896 8984 4948 9036
rect 5080 8984 5132 9036
rect 5356 8916 5408 8968
rect 7012 9120 7064 9172
rect 7288 9120 7340 9172
rect 8944 9163 8996 9172
rect 6368 8916 6420 8968
rect 6552 8916 6604 8968
rect 7012 8959 7064 8968
rect 7012 8925 7021 8959
rect 7021 8925 7055 8959
rect 7055 8925 7064 8959
rect 7012 8916 7064 8925
rect 8484 9052 8536 9104
rect 8944 9129 8953 9163
rect 8953 9129 8987 9163
rect 8987 9129 8996 9163
rect 8944 9120 8996 9129
rect 9496 9120 9548 9172
rect 10416 9120 10468 9172
rect 8024 8984 8076 9036
rect 8668 8984 8720 9036
rect 9128 9052 9180 9104
rect 10876 8984 10928 9036
rect 11336 8984 11388 9036
rect 7656 8848 7708 8900
rect 8760 8916 8812 8968
rect 9220 8959 9272 8968
rect 9220 8925 9229 8959
rect 9229 8925 9263 8959
rect 9263 8925 9272 8959
rect 9220 8916 9272 8925
rect 10140 8916 10192 8968
rect 8208 8848 8260 8900
rect 8392 8891 8444 8900
rect 8392 8857 8401 8891
rect 8401 8857 8435 8891
rect 8435 8857 8444 8891
rect 8392 8848 8444 8857
rect 8668 8848 8720 8900
rect 9864 8848 9916 8900
rect 11152 8848 11204 8900
rect 11428 8916 11480 8968
rect 12348 8916 12400 8968
rect 12992 9120 13044 9172
rect 13360 9120 13412 9172
rect 13636 9120 13688 9172
rect 22284 9120 22336 9172
rect 22652 9163 22704 9172
rect 22652 9129 22661 9163
rect 22661 9129 22695 9163
rect 22695 9129 22704 9163
rect 22652 9120 22704 9129
rect 13268 9052 13320 9104
rect 14924 9052 14976 9104
rect 15200 9052 15252 9104
rect 17224 9052 17276 9104
rect 17592 9052 17644 9104
rect 17868 9052 17920 9104
rect 12992 9027 13044 9036
rect 12992 8993 13001 9027
rect 13001 8993 13035 9027
rect 13035 8993 13044 9027
rect 12992 8984 13044 8993
rect 14832 8984 14884 9036
rect 16396 8984 16448 9036
rect 17500 8984 17552 9036
rect 18052 8984 18104 9036
rect 13360 8916 13412 8968
rect 16304 8916 16356 8968
rect 14740 8848 14792 8900
rect 6368 8780 6420 8832
rect 8760 8780 8812 8832
rect 9680 8780 9732 8832
rect 11612 8780 11664 8832
rect 12716 8823 12768 8832
rect 12716 8789 12725 8823
rect 12725 8789 12759 8823
rect 12759 8789 12768 8823
rect 12716 8780 12768 8789
rect 14924 8823 14976 8832
rect 14924 8789 14933 8823
rect 14933 8789 14967 8823
rect 14967 8789 14976 8823
rect 14924 8780 14976 8789
rect 15200 8780 15252 8832
rect 18236 8916 18288 8968
rect 18696 8984 18748 9036
rect 18972 8984 19024 9036
rect 19156 8984 19208 9036
rect 22100 8984 22152 9036
rect 18512 8916 18564 8968
rect 18880 8916 18932 8968
rect 19064 8959 19116 8968
rect 19064 8925 19073 8959
rect 19073 8925 19107 8959
rect 19107 8925 19116 8959
rect 19064 8916 19116 8925
rect 20720 8916 20772 8968
rect 17776 8848 17828 8900
rect 20168 8891 20220 8900
rect 17592 8780 17644 8832
rect 20168 8857 20177 8891
rect 20177 8857 20211 8891
rect 20211 8857 20220 8891
rect 20168 8848 20220 8857
rect 22192 8780 22244 8832
rect 4680 8678 4732 8730
rect 4744 8678 4796 8730
rect 4808 8678 4860 8730
rect 4872 8678 4924 8730
rect 12078 8678 12130 8730
rect 12142 8678 12194 8730
rect 12206 8678 12258 8730
rect 12270 8678 12322 8730
rect 19475 8678 19527 8730
rect 19539 8678 19591 8730
rect 19603 8678 19655 8730
rect 19667 8678 19719 8730
rect 2872 8576 2924 8628
rect 3608 8576 3660 8628
rect 3884 8576 3936 8628
rect 6736 8576 6788 8628
rect 7564 8576 7616 8628
rect 8668 8576 8720 8628
rect 4068 8508 4120 8560
rect 2596 8483 2648 8492
rect 2596 8449 2605 8483
rect 2605 8449 2639 8483
rect 2639 8449 2648 8483
rect 2596 8440 2648 8449
rect 3056 8440 3108 8492
rect 5356 8508 5408 8560
rect 8208 8508 8260 8560
rect 5172 8483 5224 8492
rect 5172 8449 5181 8483
rect 5181 8449 5215 8483
rect 5215 8449 5224 8483
rect 5172 8440 5224 8449
rect 5540 8440 5592 8492
rect 8300 8440 8352 8492
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 9404 8576 9456 8628
rect 9680 8576 9732 8628
rect 9772 8576 9824 8628
rect 12532 8576 12584 8628
rect 14004 8576 14056 8628
rect 14832 8576 14884 8628
rect 15476 8576 15528 8628
rect 16304 8576 16356 8628
rect 9220 8508 9272 8560
rect 11244 8508 11296 8560
rect 11428 8508 11480 8560
rect 14924 8508 14976 8560
rect 17500 8576 17552 8628
rect 18604 8576 18656 8628
rect 8392 8440 8444 8449
rect 3240 8372 3292 8424
rect 3700 8372 3752 8424
rect 5632 8372 5684 8424
rect 6736 8372 6788 8424
rect 7656 8372 7708 8424
rect 8484 8372 8536 8424
rect 4160 8304 4212 8356
rect 7932 8304 7984 8356
rect 8576 8304 8628 8356
rect 6736 8236 6788 8288
rect 9772 8483 9824 8492
rect 9772 8449 9781 8483
rect 9781 8449 9815 8483
rect 9815 8449 9824 8483
rect 9772 8440 9824 8449
rect 10876 8440 10928 8492
rect 12072 8440 12124 8492
rect 13360 8483 13412 8492
rect 13360 8449 13369 8483
rect 13369 8449 13403 8483
rect 13403 8449 13412 8483
rect 13360 8440 13412 8449
rect 15108 8440 15160 8492
rect 11612 8372 11664 8424
rect 12440 8415 12492 8424
rect 12440 8381 12449 8415
rect 12449 8381 12483 8415
rect 12483 8381 12492 8415
rect 13268 8415 13320 8424
rect 12440 8372 12492 8381
rect 13268 8381 13277 8415
rect 13277 8381 13311 8415
rect 13311 8381 13320 8415
rect 13268 8372 13320 8381
rect 14096 8372 14148 8424
rect 15016 8415 15068 8424
rect 15016 8381 15025 8415
rect 15025 8381 15059 8415
rect 15059 8381 15068 8415
rect 15016 8372 15068 8381
rect 15476 8372 15528 8424
rect 16856 8440 16908 8492
rect 18788 8483 18840 8492
rect 18788 8449 18797 8483
rect 18797 8449 18831 8483
rect 18831 8449 18840 8483
rect 18788 8440 18840 8449
rect 22100 8576 22152 8628
rect 17224 8415 17276 8424
rect 17224 8381 17233 8415
rect 17233 8381 17267 8415
rect 17267 8381 17276 8415
rect 17224 8372 17276 8381
rect 19156 8415 19208 8424
rect 9128 8347 9180 8356
rect 9128 8313 9137 8347
rect 9137 8313 9171 8347
rect 9171 8313 9180 8347
rect 9128 8304 9180 8313
rect 10876 8304 10928 8356
rect 12716 8304 12768 8356
rect 11612 8279 11664 8288
rect 11612 8245 11621 8279
rect 11621 8245 11655 8279
rect 11655 8245 11664 8279
rect 11612 8236 11664 8245
rect 17868 8304 17920 8356
rect 19156 8381 19165 8415
rect 19165 8381 19199 8415
rect 19199 8381 19208 8415
rect 19156 8372 19208 8381
rect 19432 8415 19484 8424
rect 19432 8381 19466 8415
rect 19466 8381 19484 8415
rect 19432 8372 19484 8381
rect 19800 8372 19852 8424
rect 20720 8372 20772 8424
rect 21364 8372 21416 8424
rect 22468 8415 22520 8424
rect 22468 8381 22477 8415
rect 22477 8381 22511 8415
rect 22511 8381 22520 8415
rect 22468 8372 22520 8381
rect 19064 8304 19116 8356
rect 19892 8304 19944 8356
rect 20444 8304 20496 8356
rect 19984 8236 20036 8288
rect 8379 8134 8431 8186
rect 8443 8134 8495 8186
rect 8507 8134 8559 8186
rect 8571 8134 8623 8186
rect 15776 8134 15828 8186
rect 15840 8134 15892 8186
rect 15904 8134 15956 8186
rect 15968 8134 16020 8186
rect 5080 8032 5132 8084
rect 7012 8032 7064 8084
rect 8944 8075 8996 8084
rect 8944 8041 8953 8075
rect 8953 8041 8987 8075
rect 8987 8041 8996 8075
rect 8944 8032 8996 8041
rect 11612 8032 11664 8084
rect 11704 8032 11756 8084
rect 12072 8032 12124 8084
rect 13912 8032 13964 8084
rect 14464 8075 14516 8084
rect 14464 8041 14473 8075
rect 14473 8041 14507 8075
rect 14507 8041 14516 8075
rect 14464 8032 14516 8041
rect 14740 8075 14792 8084
rect 14740 8041 14749 8075
rect 14749 8041 14783 8075
rect 14783 8041 14792 8075
rect 14740 8032 14792 8041
rect 17316 8032 17368 8084
rect 18328 8032 18380 8084
rect 19156 8032 19208 8084
rect 19432 8032 19484 8084
rect 19800 8032 19852 8084
rect 22192 8075 22244 8084
rect 22192 8041 22201 8075
rect 22201 8041 22235 8075
rect 22235 8041 22244 8075
rect 22192 8032 22244 8041
rect 7932 8007 7984 8016
rect 1768 7896 1820 7948
rect 3148 7939 3200 7948
rect 3148 7905 3157 7939
rect 3157 7905 3191 7939
rect 3191 7905 3200 7939
rect 3148 7896 3200 7905
rect 4344 7896 4396 7948
rect 3792 7828 3844 7880
rect 7932 7973 7941 8007
rect 7941 7973 7975 8007
rect 7975 7973 7984 8007
rect 7932 7964 7984 7973
rect 8760 7964 8812 8016
rect 9220 7964 9272 8016
rect 11244 7964 11296 8016
rect 4988 7871 5040 7880
rect 4988 7837 4997 7871
rect 4997 7837 5031 7871
rect 5031 7837 5040 7871
rect 4988 7828 5040 7837
rect 7012 7871 7064 7880
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 7932 7828 7984 7880
rect 5080 7760 5132 7812
rect 7564 7803 7616 7812
rect 5632 7692 5684 7744
rect 7564 7769 7573 7803
rect 7573 7769 7607 7803
rect 7607 7769 7616 7803
rect 7564 7760 7616 7769
rect 9680 7896 9732 7948
rect 9864 7896 9916 7948
rect 12348 7964 12400 8016
rect 20628 7964 20680 8016
rect 21272 8007 21324 8016
rect 21272 7973 21281 8007
rect 21281 7973 21315 8007
rect 21315 7973 21324 8007
rect 21272 7964 21324 7973
rect 22560 7964 22612 8016
rect 14924 7896 14976 7948
rect 16396 7896 16448 7948
rect 16672 7896 16724 7948
rect 17592 7896 17644 7948
rect 18512 7896 18564 7948
rect 19984 7939 20036 7948
rect 9588 7828 9640 7880
rect 11428 7871 11480 7880
rect 11428 7837 11437 7871
rect 11437 7837 11471 7871
rect 11471 7837 11480 7871
rect 11428 7828 11480 7837
rect 12624 7828 12676 7880
rect 9128 7760 9180 7812
rect 7196 7692 7248 7744
rect 8576 7735 8628 7744
rect 8576 7701 8585 7735
rect 8585 7701 8619 7735
rect 8619 7701 8628 7735
rect 8576 7692 8628 7701
rect 8668 7692 8720 7744
rect 9680 7760 9732 7812
rect 10876 7760 10928 7812
rect 11336 7760 11388 7812
rect 12532 7760 12584 7812
rect 14740 7828 14792 7880
rect 15476 7828 15528 7880
rect 11796 7692 11848 7744
rect 12716 7692 12768 7744
rect 13728 7692 13780 7744
rect 15660 7692 15712 7744
rect 16028 7692 16080 7744
rect 16304 7692 16356 7744
rect 19984 7905 19993 7939
rect 19993 7905 20027 7939
rect 20027 7905 20036 7939
rect 19984 7896 20036 7905
rect 20996 7939 21048 7948
rect 20996 7905 21005 7939
rect 21005 7905 21039 7939
rect 21039 7905 21048 7939
rect 20996 7896 21048 7905
rect 19156 7828 19208 7880
rect 20168 7871 20220 7880
rect 20168 7837 20177 7871
rect 20177 7837 20211 7871
rect 20211 7837 20220 7871
rect 20168 7828 20220 7837
rect 22192 7896 22244 7948
rect 22652 7828 22704 7880
rect 18328 7692 18380 7744
rect 18604 7692 18656 7744
rect 23020 7692 23072 7744
rect 4680 7590 4732 7642
rect 4744 7590 4796 7642
rect 4808 7590 4860 7642
rect 4872 7590 4924 7642
rect 12078 7590 12130 7642
rect 12142 7590 12194 7642
rect 12206 7590 12258 7642
rect 12270 7590 12322 7642
rect 19475 7590 19527 7642
rect 19539 7590 19591 7642
rect 19603 7590 19655 7642
rect 19667 7590 19719 7642
rect 5080 7488 5132 7540
rect 6644 7488 6696 7540
rect 7932 7488 7984 7540
rect 8576 7488 8628 7540
rect 12624 7488 12676 7540
rect 4988 7420 5040 7472
rect 5632 7420 5684 7472
rect 9864 7420 9916 7472
rect 10140 7420 10192 7472
rect 11428 7420 11480 7472
rect 12532 7420 12584 7472
rect 6644 7352 6696 7404
rect 8392 7352 8444 7404
rect 8576 7395 8628 7404
rect 8576 7361 8585 7395
rect 8585 7361 8619 7395
rect 8619 7361 8628 7395
rect 8576 7352 8628 7361
rect 9680 7352 9732 7404
rect 10232 7395 10284 7404
rect 10232 7361 10241 7395
rect 10241 7361 10275 7395
rect 10275 7361 10284 7395
rect 10232 7352 10284 7361
rect 6092 7284 6144 7336
rect 9864 7284 9916 7336
rect 10876 7284 10928 7336
rect 16304 7488 16356 7540
rect 19156 7488 19208 7540
rect 19892 7488 19944 7540
rect 20720 7488 20772 7540
rect 14924 7463 14976 7472
rect 14924 7429 14933 7463
rect 14933 7429 14967 7463
rect 14967 7429 14976 7463
rect 14924 7420 14976 7429
rect 15844 7395 15896 7404
rect 15844 7361 15853 7395
rect 15853 7361 15887 7395
rect 15887 7361 15896 7395
rect 15844 7352 15896 7361
rect 16120 7352 16172 7404
rect 13268 7284 13320 7336
rect 4252 7216 4304 7268
rect 7564 7216 7616 7268
rect 1952 7148 2004 7200
rect 2964 7148 3016 7200
rect 4068 7191 4120 7200
rect 4068 7157 4077 7191
rect 4077 7157 4111 7191
rect 4111 7157 4120 7191
rect 4068 7148 4120 7157
rect 5816 7148 5868 7200
rect 7196 7148 7248 7200
rect 9128 7148 9180 7200
rect 12348 7216 12400 7268
rect 15108 7284 15160 7336
rect 15292 7327 15344 7336
rect 15292 7293 15301 7327
rect 15301 7293 15335 7327
rect 15335 7293 15344 7327
rect 15292 7284 15344 7293
rect 16764 7352 16816 7404
rect 18420 7395 18472 7404
rect 18420 7361 18429 7395
rect 18429 7361 18463 7395
rect 18463 7361 18472 7395
rect 18420 7352 18472 7361
rect 19156 7395 19208 7404
rect 11612 7191 11664 7200
rect 11612 7157 11621 7191
rect 11621 7157 11655 7191
rect 11655 7157 11664 7191
rect 11612 7148 11664 7157
rect 14832 7216 14884 7268
rect 12624 7148 12676 7200
rect 15292 7148 15344 7200
rect 16856 7284 16908 7336
rect 17040 7284 17092 7336
rect 19156 7361 19165 7395
rect 19165 7361 19199 7395
rect 19199 7361 19208 7395
rect 19156 7352 19208 7361
rect 20260 7284 20312 7336
rect 20628 7284 20680 7336
rect 22744 7284 22796 7336
rect 18696 7148 18748 7200
rect 20720 7216 20772 7268
rect 22468 7259 22520 7268
rect 22468 7225 22477 7259
rect 22477 7225 22511 7259
rect 22511 7225 22520 7259
rect 22468 7216 22520 7225
rect 20996 7148 21048 7200
rect 21088 7148 21140 7200
rect 8379 7046 8431 7098
rect 8443 7046 8495 7098
rect 8507 7046 8559 7098
rect 8571 7046 8623 7098
rect 15776 7046 15828 7098
rect 15840 7046 15892 7098
rect 15904 7046 15956 7098
rect 15968 7046 16020 7098
rect 6184 6944 6236 6996
rect 6552 6987 6604 6996
rect 6552 6953 6561 6987
rect 6561 6953 6595 6987
rect 6595 6953 6604 6987
rect 6552 6944 6604 6953
rect 6920 6987 6972 6996
rect 6920 6953 6929 6987
rect 6929 6953 6963 6987
rect 6963 6953 6972 6987
rect 6920 6944 6972 6953
rect 7012 6944 7064 6996
rect 7564 6944 7616 6996
rect 7932 6987 7984 6996
rect 7932 6953 7941 6987
rect 7941 6953 7975 6987
rect 7975 6953 7984 6987
rect 7932 6944 7984 6953
rect 8668 6944 8720 6996
rect 8944 6987 8996 6996
rect 8944 6953 8953 6987
rect 8953 6953 8987 6987
rect 8987 6953 8996 6987
rect 8944 6944 8996 6953
rect 9588 6944 9640 6996
rect 11796 6944 11848 6996
rect 13268 6944 13320 6996
rect 14096 6944 14148 6996
rect 14372 6944 14424 6996
rect 14832 6944 14884 6996
rect 15292 6944 15344 6996
rect 19984 6944 20036 6996
rect 6828 6876 6880 6928
rect 7196 6876 7248 6928
rect 10416 6876 10468 6928
rect 4988 6851 5040 6860
rect 4988 6817 4997 6851
rect 4997 6817 5031 6851
rect 5031 6817 5040 6851
rect 4988 6808 5040 6817
rect 7748 6808 7800 6860
rect 5172 6783 5224 6792
rect 5172 6749 5181 6783
rect 5181 6749 5215 6783
rect 5215 6749 5224 6783
rect 5172 6740 5224 6749
rect 5632 6740 5684 6792
rect 6920 6740 6972 6792
rect 8208 6783 8260 6792
rect 4528 6715 4580 6724
rect 4528 6681 4537 6715
rect 4537 6681 4571 6715
rect 4571 6681 4580 6715
rect 4528 6672 4580 6681
rect 5448 6672 5500 6724
rect 6644 6672 6696 6724
rect 8208 6749 8217 6783
rect 8217 6749 8251 6783
rect 8251 6749 8260 6783
rect 8208 6740 8260 6749
rect 10692 6851 10744 6860
rect 10692 6817 10726 6851
rect 10726 6817 10744 6851
rect 10692 6808 10744 6817
rect 13636 6876 13688 6928
rect 13084 6808 13136 6860
rect 7932 6672 7984 6724
rect 8576 6715 8628 6724
rect 8576 6681 8585 6715
rect 8585 6681 8619 6715
rect 8619 6681 8628 6715
rect 8576 6672 8628 6681
rect 10140 6740 10192 6792
rect 10232 6740 10284 6792
rect 10416 6783 10468 6792
rect 10416 6749 10425 6783
rect 10425 6749 10459 6783
rect 10459 6749 10468 6783
rect 10416 6740 10468 6749
rect 14372 6808 14424 6860
rect 15752 6808 15804 6860
rect 16304 6808 16356 6860
rect 16396 6808 16448 6860
rect 18880 6876 18932 6928
rect 19064 6876 19116 6928
rect 18512 6808 18564 6860
rect 10048 6715 10100 6724
rect 10048 6681 10057 6715
rect 10057 6681 10091 6715
rect 10091 6681 10100 6715
rect 10048 6672 10100 6681
rect 16672 6740 16724 6792
rect 17316 6783 17368 6792
rect 17316 6749 17325 6783
rect 17325 6749 17359 6783
rect 17359 6749 17368 6783
rect 17316 6740 17368 6749
rect 18788 6740 18840 6792
rect 20444 6808 20496 6860
rect 20996 6944 21048 6996
rect 21088 6876 21140 6928
rect 20996 6808 21048 6860
rect 13268 6672 13320 6724
rect 14648 6672 14700 6724
rect 14924 6672 14976 6724
rect 6368 6604 6420 6656
rect 7012 6604 7064 6656
rect 9956 6604 10008 6656
rect 10692 6604 10744 6656
rect 11612 6604 11664 6656
rect 11796 6647 11848 6656
rect 11796 6613 11805 6647
rect 11805 6613 11839 6647
rect 11839 6613 11848 6647
rect 11796 6604 11848 6613
rect 17040 6647 17092 6656
rect 17040 6613 17049 6647
rect 17049 6613 17083 6647
rect 17083 6613 17092 6647
rect 17040 6604 17092 6613
rect 17224 6647 17276 6656
rect 17224 6613 17233 6647
rect 17233 6613 17267 6647
rect 17267 6613 17276 6647
rect 17224 6604 17276 6613
rect 18880 6672 18932 6724
rect 18696 6604 18748 6656
rect 19156 6715 19208 6724
rect 19156 6681 19165 6715
rect 19165 6681 19199 6715
rect 19199 6681 19208 6715
rect 19156 6672 19208 6681
rect 20168 6672 20220 6724
rect 22284 6808 22336 6860
rect 20444 6647 20496 6656
rect 20444 6613 20453 6647
rect 20453 6613 20487 6647
rect 20487 6613 20496 6647
rect 20444 6604 20496 6613
rect 22928 6672 22980 6724
rect 4680 6502 4732 6554
rect 4744 6502 4796 6554
rect 4808 6502 4860 6554
rect 4872 6502 4924 6554
rect 12078 6502 12130 6554
rect 12142 6502 12194 6554
rect 12206 6502 12258 6554
rect 12270 6502 12322 6554
rect 19475 6502 19527 6554
rect 19539 6502 19591 6554
rect 19603 6502 19655 6554
rect 19667 6502 19719 6554
rect 5632 6443 5684 6452
rect 5632 6409 5641 6443
rect 5641 6409 5675 6443
rect 5675 6409 5684 6443
rect 5632 6400 5684 6409
rect 8024 6400 8076 6452
rect 7932 6332 7984 6384
rect 8668 6375 8720 6384
rect 8668 6341 8677 6375
rect 8677 6341 8711 6375
rect 8711 6341 8720 6375
rect 8668 6332 8720 6341
rect 12440 6400 12492 6452
rect 10140 6332 10192 6384
rect 4068 6264 4120 6316
rect 7288 6264 7340 6316
rect 7748 6264 7800 6316
rect 8300 6264 8352 6316
rect 9680 6264 9732 6316
rect 10324 6307 10376 6316
rect 10324 6273 10333 6307
rect 10333 6273 10367 6307
rect 10367 6273 10376 6307
rect 10324 6264 10376 6273
rect 6000 6239 6052 6248
rect 6000 6205 6009 6239
rect 6009 6205 6043 6239
rect 6043 6205 6052 6239
rect 6000 6196 6052 6205
rect 8392 6196 8444 6248
rect 9404 6196 9456 6248
rect 10416 6196 10468 6248
rect 10692 6239 10744 6248
rect 10692 6205 10701 6239
rect 10701 6205 10735 6239
rect 10735 6205 10744 6239
rect 10692 6196 10744 6205
rect 9312 6128 9364 6180
rect 11336 6196 11388 6248
rect 12624 6264 12676 6316
rect 13084 6307 13136 6316
rect 13084 6273 13093 6307
rect 13093 6273 13127 6307
rect 13127 6273 13136 6307
rect 13084 6264 13136 6273
rect 15752 6332 15804 6384
rect 16580 6332 16632 6384
rect 16764 6332 16816 6384
rect 11520 6128 11572 6180
rect 11796 6128 11848 6180
rect 13636 6128 13688 6180
rect 11152 6060 11204 6112
rect 12440 6060 12492 6112
rect 14740 6239 14792 6248
rect 14740 6205 14749 6239
rect 14749 6205 14783 6239
rect 14783 6205 14792 6239
rect 14740 6196 14792 6205
rect 16672 6264 16724 6316
rect 16948 6264 17000 6316
rect 17592 6307 17644 6316
rect 17592 6273 17601 6307
rect 17601 6273 17635 6307
rect 17635 6273 17644 6307
rect 17592 6264 17644 6273
rect 16856 6196 16908 6248
rect 17684 6196 17736 6248
rect 18236 6239 18288 6248
rect 18236 6205 18245 6239
rect 18245 6205 18279 6239
rect 18279 6205 18288 6239
rect 18236 6196 18288 6205
rect 18328 6196 18380 6248
rect 20720 6332 20772 6384
rect 20444 6264 20496 6316
rect 20812 6196 20864 6248
rect 21180 6196 21232 6248
rect 14280 6060 14332 6112
rect 15292 6128 15344 6180
rect 15752 6128 15804 6180
rect 14556 6060 14608 6112
rect 18144 6128 18196 6180
rect 19156 6128 19208 6180
rect 17868 6060 17920 6112
rect 18604 6060 18656 6112
rect 18696 6060 18748 6112
rect 19340 6060 19392 6112
rect 19800 6060 19852 6112
rect 21824 6128 21876 6180
rect 22652 6060 22704 6112
rect 22744 6103 22796 6112
rect 22744 6069 22753 6103
rect 22753 6069 22787 6103
rect 22787 6069 22796 6103
rect 22744 6060 22796 6069
rect 8379 5958 8431 6010
rect 8443 5958 8495 6010
rect 8507 5958 8559 6010
rect 8571 5958 8623 6010
rect 15776 5958 15828 6010
rect 15840 5958 15892 6010
rect 15904 5958 15956 6010
rect 15968 5958 16020 6010
rect 4160 5856 4212 5908
rect 6552 5899 6604 5908
rect 6552 5865 6561 5899
rect 6561 5865 6595 5899
rect 6595 5865 6604 5899
rect 6552 5856 6604 5865
rect 7012 5899 7064 5908
rect 7012 5865 7021 5899
rect 7021 5865 7055 5899
rect 7055 5865 7064 5899
rect 7012 5856 7064 5865
rect 7656 5856 7708 5908
rect 7840 5856 7892 5908
rect 9404 5856 9456 5908
rect 13636 5899 13688 5908
rect 4436 5788 4488 5840
rect 6460 5788 6512 5840
rect 7472 5788 7524 5840
rect 9312 5788 9364 5840
rect 13636 5865 13645 5899
rect 13645 5865 13679 5899
rect 13679 5865 13688 5899
rect 13636 5856 13688 5865
rect 14280 5899 14332 5908
rect 14280 5865 14289 5899
rect 14289 5865 14323 5899
rect 14323 5865 14332 5899
rect 14280 5856 14332 5865
rect 14740 5856 14792 5908
rect 18512 5899 18564 5908
rect 12808 5788 12860 5840
rect 17868 5788 17920 5840
rect 18512 5865 18521 5899
rect 18521 5865 18555 5899
rect 18555 5865 18564 5899
rect 18512 5856 18564 5865
rect 18604 5856 18656 5908
rect 20720 5788 20772 5840
rect 9036 5720 9088 5772
rect 10692 5720 10744 5772
rect 12348 5720 12400 5772
rect 12900 5720 12952 5772
rect 5908 5652 5960 5704
rect 6276 5652 6328 5704
rect 7748 5652 7800 5704
rect 8852 5652 8904 5704
rect 9404 5652 9456 5704
rect 12256 5695 12308 5704
rect 12256 5661 12265 5695
rect 12265 5661 12299 5695
rect 12299 5661 12308 5695
rect 12256 5652 12308 5661
rect 14004 5720 14056 5772
rect 17040 5720 17092 5772
rect 17224 5720 17276 5772
rect 14372 5652 14424 5704
rect 14464 5652 14516 5704
rect 14924 5652 14976 5704
rect 16764 5695 16816 5704
rect 9588 5584 9640 5636
rect 13268 5584 13320 5636
rect 16028 5584 16080 5636
rect 16764 5661 16773 5695
rect 16773 5661 16807 5695
rect 16807 5661 16816 5695
rect 16764 5652 16816 5661
rect 20076 5720 20128 5772
rect 18788 5627 18840 5636
rect 10324 5516 10376 5568
rect 12900 5516 12952 5568
rect 14004 5516 14056 5568
rect 14372 5516 14424 5568
rect 16396 5516 16448 5568
rect 18788 5593 18797 5627
rect 18797 5593 18831 5627
rect 18831 5593 18840 5627
rect 18788 5584 18840 5593
rect 19800 5652 19852 5704
rect 21640 5720 21692 5772
rect 22284 5720 22336 5772
rect 20352 5695 20404 5704
rect 20352 5661 20361 5695
rect 20361 5661 20395 5695
rect 20395 5661 20404 5695
rect 20352 5652 20404 5661
rect 20444 5652 20496 5704
rect 22100 5695 22152 5704
rect 22100 5661 22109 5695
rect 22109 5661 22143 5695
rect 22143 5661 22152 5695
rect 22100 5652 22152 5661
rect 19340 5516 19392 5568
rect 19800 5559 19852 5568
rect 19800 5525 19809 5559
rect 19809 5525 19843 5559
rect 19843 5525 19852 5559
rect 19800 5516 19852 5525
rect 19984 5516 20036 5568
rect 20260 5516 20312 5568
rect 22744 5516 22796 5568
rect 4680 5414 4732 5466
rect 4744 5414 4796 5466
rect 4808 5414 4860 5466
rect 4872 5414 4924 5466
rect 12078 5414 12130 5466
rect 12142 5414 12194 5466
rect 12206 5414 12258 5466
rect 12270 5414 12322 5466
rect 19475 5414 19527 5466
rect 19539 5414 19591 5466
rect 19603 5414 19655 5466
rect 19667 5414 19719 5466
rect 8944 5312 8996 5364
rect 9128 5355 9180 5364
rect 9128 5321 9137 5355
rect 9137 5321 9171 5355
rect 9171 5321 9180 5355
rect 9128 5312 9180 5321
rect 9864 5312 9916 5364
rect 10692 5312 10744 5364
rect 11152 5355 11204 5364
rect 11152 5321 11161 5355
rect 11161 5321 11195 5355
rect 11195 5321 11204 5355
rect 11152 5312 11204 5321
rect 11336 5312 11388 5364
rect 13084 5312 13136 5364
rect 13360 5312 13412 5364
rect 7748 5176 7800 5228
rect 9772 5219 9824 5228
rect 9772 5185 9781 5219
rect 9781 5185 9815 5219
rect 9815 5185 9824 5219
rect 9772 5176 9824 5185
rect 7380 5108 7432 5160
rect 13452 5244 13504 5296
rect 10692 5219 10744 5228
rect 10692 5185 10701 5219
rect 10701 5185 10735 5219
rect 10735 5185 10744 5219
rect 10692 5176 10744 5185
rect 11612 5219 11664 5228
rect 11612 5185 11621 5219
rect 11621 5185 11655 5219
rect 11655 5185 11664 5219
rect 11612 5176 11664 5185
rect 11520 5151 11572 5160
rect 7932 5040 7984 5092
rect 11520 5117 11529 5151
rect 11529 5117 11563 5151
rect 11563 5117 11572 5151
rect 11520 5108 11572 5117
rect 12440 5176 12492 5228
rect 14464 5312 14516 5364
rect 14924 5312 14976 5364
rect 16856 5355 16908 5364
rect 16856 5321 16865 5355
rect 16865 5321 16899 5355
rect 16899 5321 16908 5355
rect 16856 5312 16908 5321
rect 18236 5312 18288 5364
rect 20076 5312 20128 5364
rect 21824 5312 21876 5364
rect 20720 5244 20772 5296
rect 14740 5176 14792 5228
rect 17592 5176 17644 5228
rect 17868 5176 17920 5228
rect 18144 5176 18196 5228
rect 19156 5219 19208 5228
rect 19156 5185 19165 5219
rect 19165 5185 19199 5219
rect 19199 5185 19208 5219
rect 19156 5176 19208 5185
rect 20260 5219 20312 5228
rect 20260 5185 20269 5219
rect 20269 5185 20303 5219
rect 20303 5185 20312 5219
rect 20260 5176 20312 5185
rect 20904 5176 20956 5228
rect 13360 5108 13412 5160
rect 14188 5108 14240 5160
rect 16028 5108 16080 5160
rect 9588 5015 9640 5024
rect 9588 4981 9597 5015
rect 9597 4981 9631 5015
rect 9631 4981 9640 5015
rect 9588 4972 9640 4981
rect 12624 5040 12676 5092
rect 12256 4972 12308 5024
rect 12348 4972 12400 5024
rect 12808 5015 12860 5024
rect 12808 4981 12817 5015
rect 12817 4981 12851 5015
rect 12851 4981 12860 5015
rect 12808 4972 12860 4981
rect 15568 5040 15620 5092
rect 17776 5108 17828 5160
rect 19432 5108 19484 5160
rect 20720 5108 20772 5160
rect 21180 5151 21232 5160
rect 21180 5117 21189 5151
rect 21189 5117 21223 5151
rect 21223 5117 21232 5151
rect 21180 5108 21232 5117
rect 17868 5040 17920 5092
rect 18328 5040 18380 5092
rect 17224 5015 17276 5024
rect 17224 4981 17233 5015
rect 17233 4981 17267 5015
rect 17267 4981 17276 5015
rect 17224 4972 17276 4981
rect 17500 4972 17552 5024
rect 19340 5040 19392 5092
rect 22100 5040 22152 5092
rect 8379 4870 8431 4922
rect 8443 4870 8495 4922
rect 8507 4870 8559 4922
rect 8571 4870 8623 4922
rect 15776 4870 15828 4922
rect 15840 4870 15892 4922
rect 15904 4870 15956 4922
rect 15968 4870 16020 4922
rect 9864 4811 9916 4820
rect 9864 4777 9873 4811
rect 9873 4777 9907 4811
rect 9907 4777 9916 4811
rect 9864 4768 9916 4777
rect 10784 4768 10836 4820
rect 11704 4768 11756 4820
rect 11888 4811 11940 4820
rect 11888 4777 11897 4811
rect 11897 4777 11931 4811
rect 11931 4777 11940 4811
rect 11888 4768 11940 4777
rect 11980 4768 12032 4820
rect 12992 4768 13044 4820
rect 14832 4768 14884 4820
rect 17500 4768 17552 4820
rect 17776 4811 17828 4820
rect 17776 4777 17785 4811
rect 17785 4777 17819 4811
rect 17819 4777 17828 4811
rect 17776 4768 17828 4777
rect 18236 4811 18288 4820
rect 18236 4777 18245 4811
rect 18245 4777 18279 4811
rect 18279 4777 18288 4811
rect 18236 4768 18288 4777
rect 22100 4768 22152 4820
rect 10324 4743 10376 4752
rect 10324 4709 10333 4743
rect 10333 4709 10367 4743
rect 10367 4709 10376 4743
rect 10324 4700 10376 4709
rect 13360 4743 13412 4752
rect 13360 4709 13369 4743
rect 13369 4709 13403 4743
rect 13403 4709 13412 4743
rect 13360 4700 13412 4709
rect 14556 4700 14608 4752
rect 11888 4632 11940 4684
rect 10692 4564 10744 4616
rect 11612 4564 11664 4616
rect 14188 4632 14240 4684
rect 18052 4700 18104 4752
rect 20444 4700 20496 4752
rect 15660 4632 15712 4684
rect 16672 4632 16724 4684
rect 12440 4607 12492 4616
rect 12440 4573 12449 4607
rect 12449 4573 12483 4607
rect 12483 4573 12492 4607
rect 12440 4564 12492 4573
rect 12900 4564 12952 4616
rect 14464 4607 14516 4616
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 16948 4632 17000 4684
rect 17316 4632 17368 4684
rect 19800 4632 19852 4684
rect 21180 4632 21232 4684
rect 21364 4675 21416 4684
rect 21364 4641 21398 4675
rect 21398 4641 21416 4675
rect 21364 4632 21416 4641
rect 15568 4496 15620 4548
rect 17040 4496 17092 4548
rect 18880 4496 18932 4548
rect 20076 4564 20128 4616
rect 20260 4496 20312 4548
rect 6920 4428 6972 4480
rect 11980 4428 12032 4480
rect 14924 4428 14976 4480
rect 15292 4428 15344 4480
rect 15844 4428 15896 4480
rect 16580 4428 16632 4480
rect 17684 4428 17736 4480
rect 20812 4428 20864 4480
rect 4680 4326 4732 4378
rect 4744 4326 4796 4378
rect 4808 4326 4860 4378
rect 4872 4326 4924 4378
rect 12078 4326 12130 4378
rect 12142 4326 12194 4378
rect 12206 4326 12258 4378
rect 12270 4326 12322 4378
rect 19475 4326 19527 4378
rect 19539 4326 19591 4378
rect 19603 4326 19655 4378
rect 19667 4326 19719 4378
rect 9588 4224 9640 4276
rect 13268 4224 13320 4276
rect 13636 4267 13688 4276
rect 13636 4233 13645 4267
rect 13645 4233 13679 4267
rect 13679 4233 13688 4267
rect 13636 4224 13688 4233
rect 8208 4156 8260 4208
rect 9220 4088 9272 4140
rect 11888 4131 11940 4140
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 14096 4088 14148 4140
rect 14832 4224 14884 4276
rect 18052 4267 18104 4276
rect 15660 4156 15712 4208
rect 18052 4233 18061 4267
rect 18061 4233 18095 4267
rect 18095 4233 18104 4267
rect 18052 4224 18104 4233
rect 22008 4224 22060 4276
rect 15844 4088 15896 4140
rect 17592 4088 17644 4140
rect 18880 4088 18932 4140
rect 19064 4131 19116 4140
rect 19064 4097 19073 4131
rect 19073 4097 19107 4131
rect 19107 4097 19116 4131
rect 19064 4088 19116 4097
rect 20996 4088 21048 4140
rect 21272 4088 21324 4140
rect 14004 4063 14056 4072
rect 14004 4029 14013 4063
rect 14013 4029 14047 4063
rect 14047 4029 14056 4063
rect 14004 4020 14056 4029
rect 14740 4020 14792 4072
rect 14924 4063 14976 4072
rect 14924 4029 14958 4063
rect 14958 4029 14976 4063
rect 14924 4020 14976 4029
rect 18972 4020 19024 4072
rect 20352 4020 20404 4072
rect 21180 4020 21232 4072
rect 21640 4063 21692 4072
rect 21640 4029 21674 4063
rect 21674 4029 21692 4063
rect 21640 4020 21692 4029
rect 11428 3884 11480 3936
rect 12164 3884 12216 3936
rect 16580 3995 16632 4004
rect 16580 3961 16614 3995
rect 16614 3961 16632 3995
rect 16580 3952 16632 3961
rect 19156 3952 19208 4004
rect 12624 3927 12676 3936
rect 12624 3893 12633 3927
rect 12633 3893 12667 3927
rect 12667 3893 12676 3927
rect 12992 3927 13044 3936
rect 12624 3884 12676 3893
rect 12992 3893 13001 3927
rect 13001 3893 13035 3927
rect 13035 3893 13044 3927
rect 12992 3884 13044 3893
rect 13084 3927 13136 3936
rect 13084 3893 13093 3927
rect 13093 3893 13127 3927
rect 13127 3893 13136 3927
rect 13084 3884 13136 3893
rect 14372 3884 14424 3936
rect 15016 3884 15068 3936
rect 17040 3884 17092 3936
rect 17684 3927 17736 3936
rect 17684 3893 17693 3927
rect 17693 3893 17727 3927
rect 17727 3893 17736 3927
rect 17684 3884 17736 3893
rect 18512 3927 18564 3936
rect 18512 3893 18521 3927
rect 18521 3893 18555 3927
rect 18555 3893 18564 3927
rect 18512 3884 18564 3893
rect 21272 3884 21324 3936
rect 21364 3884 21416 3936
rect 8379 3782 8431 3834
rect 8443 3782 8495 3834
rect 8507 3782 8559 3834
rect 8571 3782 8623 3834
rect 15776 3782 15828 3834
rect 15840 3782 15892 3834
rect 15904 3782 15956 3834
rect 15968 3782 16020 3834
rect 11428 3680 11480 3732
rect 13176 3680 13228 3732
rect 13544 3723 13596 3732
rect 13544 3689 13553 3723
rect 13553 3689 13587 3723
rect 13587 3689 13596 3723
rect 13544 3680 13596 3689
rect 13728 3680 13780 3732
rect 14280 3680 14332 3732
rect 16120 3723 16172 3732
rect 16120 3689 16129 3723
rect 16129 3689 16163 3723
rect 16163 3689 16172 3723
rect 16120 3680 16172 3689
rect 16948 3680 17000 3732
rect 12440 3612 12492 3664
rect 18604 3680 18656 3732
rect 20812 3680 20864 3732
rect 21640 3680 21692 3732
rect 17500 3612 17552 3664
rect 17776 3612 17828 3664
rect 20996 3612 21048 3664
rect 11612 3544 11664 3596
rect 12532 3587 12584 3596
rect 10692 3476 10744 3528
rect 11704 3519 11756 3528
rect 11704 3485 11713 3519
rect 11713 3485 11747 3519
rect 11747 3485 11756 3519
rect 11704 3476 11756 3485
rect 12532 3553 12541 3587
rect 12541 3553 12575 3587
rect 12575 3553 12584 3587
rect 12532 3544 12584 3553
rect 14004 3544 14056 3596
rect 14648 3587 14700 3596
rect 14648 3553 14657 3587
rect 14657 3553 14691 3587
rect 14691 3553 14700 3587
rect 14648 3544 14700 3553
rect 15568 3587 15620 3596
rect 15568 3553 15577 3587
rect 15577 3553 15611 3587
rect 15611 3553 15620 3587
rect 15568 3544 15620 3553
rect 18512 3544 18564 3596
rect 19248 3587 19300 3596
rect 19248 3553 19282 3587
rect 19282 3553 19300 3587
rect 19248 3544 19300 3553
rect 20352 3544 20404 3596
rect 22284 3612 22336 3664
rect 13820 3519 13872 3528
rect 13820 3485 13829 3519
rect 13829 3485 13863 3519
rect 13863 3485 13872 3519
rect 13820 3476 13872 3485
rect 14832 3519 14884 3528
rect 14832 3485 14841 3519
rect 14841 3485 14875 3519
rect 14875 3485 14884 3519
rect 14832 3476 14884 3485
rect 15108 3476 15160 3528
rect 12164 3451 12216 3460
rect 12164 3417 12173 3451
rect 12173 3417 12207 3451
rect 12207 3417 12216 3451
rect 12164 3408 12216 3417
rect 7564 3340 7616 3392
rect 13268 3340 13320 3392
rect 16304 3408 16356 3460
rect 17040 3476 17092 3528
rect 18144 3476 18196 3528
rect 18972 3519 19024 3528
rect 18972 3485 18981 3519
rect 18981 3485 19015 3519
rect 19015 3485 19024 3519
rect 18972 3476 19024 3485
rect 18420 3408 18472 3460
rect 15568 3340 15620 3392
rect 17776 3340 17828 3392
rect 19156 3340 19208 3392
rect 20444 3340 20496 3392
rect 21548 3340 21600 3392
rect 4680 3238 4732 3290
rect 4744 3238 4796 3290
rect 4808 3238 4860 3290
rect 4872 3238 4924 3290
rect 12078 3238 12130 3290
rect 12142 3238 12194 3290
rect 12206 3238 12258 3290
rect 12270 3238 12322 3290
rect 19475 3238 19527 3290
rect 19539 3238 19591 3290
rect 19603 3238 19655 3290
rect 19667 3238 19719 3290
rect 13268 3179 13320 3188
rect 13268 3145 13277 3179
rect 13277 3145 13311 3179
rect 13311 3145 13320 3179
rect 13268 3136 13320 3145
rect 14096 3179 14148 3188
rect 14096 3145 14105 3179
rect 14105 3145 14139 3179
rect 14139 3145 14148 3179
rect 14096 3136 14148 3145
rect 14188 3136 14240 3188
rect 15384 3136 15436 3188
rect 2964 3068 3016 3120
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 1768 2975 1820 2984
rect 1768 2941 1777 2975
rect 1777 2941 1811 2975
rect 1811 2941 1820 2975
rect 1768 2932 1820 2941
rect 11060 3000 11112 3052
rect 11980 3000 12032 3052
rect 14004 3000 14056 3052
rect 15016 3000 15068 3052
rect 16488 3136 16540 3188
rect 19156 3136 19208 3188
rect 19248 3136 19300 3188
rect 20352 3068 20404 3120
rect 22284 3136 22336 3188
rect 5080 2975 5132 2984
rect 5080 2941 5089 2975
rect 5089 2941 5123 2975
rect 5123 2941 5132 2975
rect 5080 2932 5132 2941
rect 17316 3000 17368 3052
rect 17684 2932 17736 2984
rect 20444 3000 20496 3052
rect 1676 2796 1728 2848
rect 14372 2796 14424 2848
rect 15108 2796 15160 2848
rect 17040 2864 17092 2916
rect 18144 2864 18196 2916
rect 21456 2932 21508 2984
rect 18328 2864 18380 2916
rect 17500 2796 17552 2848
rect 18052 2796 18104 2848
rect 20076 2796 20128 2848
rect 20904 2864 20956 2916
rect 22560 2796 22612 2848
rect 8379 2694 8431 2746
rect 8443 2694 8495 2746
rect 8507 2694 8559 2746
rect 8571 2694 8623 2746
rect 15776 2694 15828 2746
rect 15840 2694 15892 2746
rect 15904 2694 15956 2746
rect 15968 2694 16020 2746
rect 13912 2592 13964 2644
rect 15660 2592 15712 2644
rect 17500 2592 17552 2644
rect 18328 2592 18380 2644
rect 19984 2592 20036 2644
rect 20628 2592 20680 2644
rect 11704 2524 11756 2576
rect 16488 2524 16540 2576
rect 16764 2524 16816 2576
rect 14004 2456 14056 2508
rect 17408 2456 17460 2508
rect 17684 2524 17736 2576
rect 18420 2524 18472 2576
rect 18604 2567 18656 2576
rect 18604 2533 18638 2567
rect 18638 2533 18656 2567
rect 18604 2524 18656 2533
rect 20904 2524 20956 2576
rect 14372 2363 14424 2372
rect 14372 2329 14381 2363
rect 14381 2329 14415 2363
rect 14415 2329 14424 2363
rect 14372 2320 14424 2329
rect 18144 2456 18196 2508
rect 16120 2320 16172 2372
rect 17500 2320 17552 2372
rect 18052 2388 18104 2440
rect 19340 2456 19392 2508
rect 20352 2456 20404 2508
rect 21272 2456 21324 2508
rect 21088 2388 21140 2440
rect 15476 2252 15528 2304
rect 16304 2252 16356 2304
rect 17868 2252 17920 2304
rect 4680 2150 4732 2202
rect 4744 2150 4796 2202
rect 4808 2150 4860 2202
rect 4872 2150 4924 2202
rect 12078 2150 12130 2202
rect 12142 2150 12194 2202
rect 12206 2150 12258 2202
rect 12270 2150 12322 2202
rect 19475 2150 19527 2202
rect 19539 2150 19591 2202
rect 19603 2150 19655 2202
rect 19667 2150 19719 2202
rect 16764 2048 16816 2100
rect 19248 2048 19300 2100
rect 14372 1980 14424 2032
rect 17224 1980 17276 2032
rect 17408 1980 17460 2032
rect 20904 1980 20956 2032
rect 17500 1912 17552 1964
rect 21272 1912 21324 1964
rect 16304 1844 16356 1896
rect 18236 1844 18288 1896
rect 15200 1776 15252 1828
rect 19892 1776 19944 1828
rect 16396 1300 16448 1352
rect 19340 1300 19392 1352
<< metal2 >>
rect 294 23920 350 24400
rect 846 23920 902 24400
rect 1490 23920 1546 24400
rect 2134 23920 2190 24400
rect 2778 23920 2834 24400
rect 3422 23920 3478 24400
rect 4066 23920 4122 24400
rect 4710 23920 4766 24400
rect 5354 23920 5410 24400
rect 5998 23920 6054 24400
rect 6642 23920 6698 24400
rect 7286 23920 7342 24400
rect 7930 23920 7986 24400
rect 8574 23920 8630 24400
rect 9218 23920 9274 24400
rect 9862 23920 9918 24400
rect 10506 23920 10562 24400
rect 11150 23920 11206 24400
rect 11794 23920 11850 24400
rect 12438 23920 12494 24400
rect 13082 23920 13138 24400
rect 13726 23920 13782 24400
rect 14370 23920 14426 24400
rect 15014 23920 15070 24400
rect 15658 23920 15714 24400
rect 16302 23920 16358 24400
rect 16946 23920 17002 24400
rect 17590 23920 17646 24400
rect 18234 23920 18290 24400
rect 18878 23920 18934 24400
rect 19522 23920 19578 24400
rect 19798 24032 19854 24041
rect 19798 23967 19854 23976
rect 308 21146 336 23920
rect 296 21140 348 21146
rect 296 21082 348 21088
rect 860 20262 888 23920
rect 1504 21690 1532 23920
rect 1492 21684 1544 21690
rect 1492 21626 1544 21632
rect 1952 21344 2004 21350
rect 1952 21286 2004 21292
rect 1768 20936 1820 20942
rect 1768 20878 1820 20884
rect 1780 20398 1808 20878
rect 1768 20392 1820 20398
rect 1768 20334 1820 20340
rect 848 20256 900 20262
rect 848 20198 900 20204
rect 1768 19984 1820 19990
rect 1768 19926 1820 19932
rect 1400 19848 1452 19854
rect 1400 19790 1452 19796
rect 1412 19310 1440 19790
rect 1400 19304 1452 19310
rect 1400 19246 1452 19252
rect 1676 19236 1728 19242
rect 1676 19178 1728 19184
rect 1688 18970 1716 19178
rect 1676 18964 1728 18970
rect 1676 18906 1728 18912
rect 1490 18320 1546 18329
rect 1490 18255 1546 18264
rect 1400 17332 1452 17338
rect 1400 17274 1452 17280
rect 1412 16658 1440 17274
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1504 16046 1532 18255
rect 1492 16040 1544 16046
rect 1492 15982 1544 15988
rect 1400 14816 1452 14822
rect 1400 14758 1452 14764
rect 1412 13530 1440 14758
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1504 13938 1532 14418
rect 1492 13932 1544 13938
rect 1492 13874 1544 13880
rect 1400 13524 1452 13530
rect 1400 13466 1452 13472
rect 1674 13424 1730 13433
rect 1674 13359 1676 13368
rect 1728 13359 1730 13368
rect 1676 13330 1728 13336
rect 1584 12776 1636 12782
rect 1584 12718 1636 12724
rect 1596 12306 1624 12718
rect 1584 12300 1636 12306
rect 1584 12242 1636 12248
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 1412 11150 1440 11630
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10606 1440 11086
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1780 10266 1808 19926
rect 1860 16040 1912 16046
rect 1860 15982 1912 15988
rect 1872 15638 1900 15982
rect 1860 15632 1912 15638
rect 1860 15574 1912 15580
rect 1872 15026 1900 15574
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1872 14618 1900 14962
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1858 13832 1914 13841
rect 1858 13767 1914 13776
rect 1872 13258 1900 13767
rect 1860 13252 1912 13258
rect 1860 13194 1912 13200
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1492 9444 1544 9450
rect 1492 9386 1544 9392
rect 1504 9081 1532 9386
rect 1490 9072 1546 9081
rect 1490 9007 1546 9016
rect 1768 7948 1820 7954
rect 1768 7890 1820 7896
rect 1780 2990 1808 7890
rect 1964 7206 1992 21286
rect 2044 20324 2096 20330
rect 2044 20266 2096 20272
rect 2056 19718 2084 20266
rect 2148 20058 2176 23920
rect 2792 23066 2820 23920
rect 3436 23066 3464 23920
rect 4080 23066 4108 23920
rect 2792 23038 2912 23066
rect 3436 23038 3740 23066
rect 2688 21412 2740 21418
rect 2688 21354 2740 21360
rect 2412 21344 2464 21350
rect 2412 21286 2464 21292
rect 2136 20052 2188 20058
rect 2136 19994 2188 20000
rect 2044 19712 2096 19718
rect 2044 19654 2096 19660
rect 2320 19236 2372 19242
rect 2320 19178 2372 19184
rect 2332 18766 2360 19178
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2332 18086 2360 18702
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 2332 17746 2360 18022
rect 2320 17740 2372 17746
rect 2320 17682 2372 17688
rect 2228 17128 2280 17134
rect 2332 17116 2360 17682
rect 2280 17088 2360 17116
rect 2228 17070 2280 17076
rect 2332 16726 2360 17088
rect 2320 16720 2372 16726
rect 2320 16662 2372 16668
rect 2424 15473 2452 21286
rect 2596 17808 2648 17814
rect 2700 17785 2728 21354
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2792 19281 2820 19858
rect 2778 19272 2834 19281
rect 2778 19207 2834 19216
rect 2792 19174 2820 19207
rect 2780 19168 2832 19174
rect 2780 19110 2832 19116
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2596 17750 2648 17756
rect 2686 17776 2742 17785
rect 2608 17660 2636 17750
rect 2686 17711 2742 17720
rect 2792 17660 2820 17818
rect 2608 17632 2820 17660
rect 2596 16720 2648 16726
rect 2596 16662 2648 16668
rect 2502 15600 2558 15609
rect 2502 15535 2558 15544
rect 2410 15464 2466 15473
rect 2410 15399 2466 15408
rect 2136 10532 2188 10538
rect 2136 10474 2188 10480
rect 2148 10198 2176 10474
rect 2136 10192 2188 10198
rect 2136 10134 2188 10140
rect 2148 9722 2176 10134
rect 2136 9716 2188 9722
rect 2136 9658 2188 9664
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 2332 9178 2360 9318
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2516 9110 2544 15535
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2608 8498 2636 16662
rect 2884 16266 2912 23038
rect 2964 21344 3016 21350
rect 2964 21286 3016 21292
rect 3332 21344 3384 21350
rect 3332 21286 3384 21292
rect 3424 21344 3476 21350
rect 3424 21286 3476 21292
rect 2976 21078 3004 21286
rect 2964 21072 3016 21078
rect 2964 21014 3016 21020
rect 3344 20806 3372 21286
rect 3436 21010 3464 21286
rect 3424 21004 3476 21010
rect 3424 20946 3476 20952
rect 3332 20800 3384 20806
rect 3332 20742 3384 20748
rect 3344 19310 3372 20742
rect 3436 20602 3464 20946
rect 3424 20596 3476 20602
rect 3424 20538 3476 20544
rect 3424 20392 3476 20398
rect 3424 20334 3476 20340
rect 3436 19922 3464 20334
rect 3424 19916 3476 19922
rect 3424 19858 3476 19864
rect 3436 19514 3464 19858
rect 3712 19802 3740 23038
rect 3804 23038 4108 23066
rect 4724 23066 4752 23920
rect 4724 23038 5028 23066
rect 3804 19990 3832 23038
rect 4654 21788 4950 21808
rect 4710 21786 4734 21788
rect 4790 21786 4814 21788
rect 4870 21786 4894 21788
rect 4732 21734 4734 21786
rect 4796 21734 4808 21786
rect 4870 21734 4872 21786
rect 4710 21732 4734 21734
rect 4790 21732 4814 21734
rect 4870 21732 4894 21734
rect 4654 21712 4950 21732
rect 4160 21480 4212 21486
rect 4160 21422 4212 21428
rect 4068 21344 4120 21350
rect 3882 21312 3938 21321
rect 4068 21286 4120 21292
rect 3882 21247 3938 21256
rect 3896 20874 3924 21247
rect 4080 21146 4108 21286
rect 4068 21140 4120 21146
rect 4068 21082 4120 21088
rect 3884 20868 3936 20874
rect 3884 20810 3936 20816
rect 3976 20800 4028 20806
rect 3976 20742 4028 20748
rect 3792 19984 3844 19990
rect 3792 19926 3844 19932
rect 3712 19774 3924 19802
rect 3424 19508 3476 19514
rect 3424 19450 3476 19456
rect 3792 19508 3844 19514
rect 3792 19450 3844 19456
rect 3332 19304 3384 19310
rect 2962 19272 3018 19281
rect 3332 19246 3384 19252
rect 2962 19207 2964 19216
rect 3016 19207 3018 19216
rect 2964 19178 3016 19184
rect 3240 19168 3292 19174
rect 3240 19110 3292 19116
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 3160 16697 3188 16730
rect 3146 16688 3202 16697
rect 3146 16623 3202 16632
rect 2792 16250 2912 16266
rect 2780 16244 2912 16250
rect 2832 16238 2912 16244
rect 2780 16186 2832 16192
rect 2688 15972 2740 15978
rect 2688 15914 2740 15920
rect 2700 15366 2728 15914
rect 3146 15736 3202 15745
rect 3146 15671 3202 15680
rect 3160 15570 3188 15671
rect 2964 15564 3016 15570
rect 2964 15506 3016 15512
rect 3148 15564 3200 15570
rect 3148 15506 3200 15512
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2700 13326 2728 15302
rect 2976 14822 3004 15506
rect 3056 14884 3108 14890
rect 3056 14826 3108 14832
rect 2964 14816 3016 14822
rect 2964 14758 3016 14764
rect 3068 14618 3096 14826
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 2884 14385 2912 14486
rect 3068 14414 3096 14554
rect 3056 14408 3108 14414
rect 2870 14376 2926 14385
rect 3056 14350 3108 14356
rect 2870 14311 2926 14320
rect 2884 14074 2912 14311
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 3160 13530 3188 13670
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 3252 13190 3280 19110
rect 3436 18290 3464 19450
rect 3700 19304 3752 19310
rect 3700 19246 3752 19252
rect 3712 18834 3740 19246
rect 3700 18828 3752 18834
rect 3700 18770 3752 18776
rect 3712 18358 3740 18770
rect 3700 18352 3752 18358
rect 3700 18294 3752 18300
rect 3424 18284 3476 18290
rect 3424 18226 3476 18232
rect 3436 18086 3464 18226
rect 3608 18148 3660 18154
rect 3608 18090 3660 18096
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 3516 17740 3568 17746
rect 3516 17682 3568 17688
rect 3528 17338 3556 17682
rect 3620 17610 3648 18090
rect 3608 17604 3660 17610
rect 3608 17546 3660 17552
rect 3516 17332 3568 17338
rect 3516 17274 3568 17280
rect 3620 17202 3648 17546
rect 3700 17264 3752 17270
rect 3698 17232 3700 17241
rect 3752 17232 3754 17241
rect 3608 17196 3660 17202
rect 3698 17167 3754 17176
rect 3608 17138 3660 17144
rect 3332 17060 3384 17066
rect 3332 17002 3384 17008
rect 3344 16833 3372 17002
rect 3330 16824 3386 16833
rect 3330 16759 3332 16768
rect 3384 16759 3386 16768
rect 3332 16730 3384 16736
rect 3424 16516 3476 16522
rect 3424 16458 3476 16464
rect 3436 16250 3464 16458
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3332 15496 3384 15502
rect 3332 15438 3384 15444
rect 3344 15201 3372 15438
rect 3330 15192 3386 15201
rect 3330 15127 3386 15136
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3712 13938 3740 14758
rect 3700 13932 3752 13938
rect 3700 13874 3752 13880
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2792 11558 2820 12242
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2792 9654 2820 10066
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2792 9042 2820 9590
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2884 8634 2912 12582
rect 2976 12442 3004 12650
rect 3424 12640 3476 12646
rect 3252 12600 3424 12628
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 2976 12238 3004 12378
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2976 11354 3004 11630
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3068 8498 3096 11494
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 3160 11218 3188 11290
rect 3148 11212 3200 11218
rect 3148 11154 3200 11160
rect 3160 10810 3188 11154
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3146 10568 3202 10577
rect 3146 10503 3202 10512
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 3160 7954 3188 10503
rect 3252 8430 3280 12600
rect 3424 12582 3476 12588
rect 3516 12164 3568 12170
rect 3516 12106 3568 12112
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3344 10606 3372 11698
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3436 11354 3464 11494
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3528 11286 3556 12106
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3516 11280 3568 11286
rect 3516 11222 3568 11228
rect 3424 11212 3476 11218
rect 3424 11154 3476 11160
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3344 9518 3372 9862
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3344 9178 3372 9454
rect 3436 9178 3464 11154
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 3528 10606 3556 10950
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3528 10130 3556 10542
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3528 9450 3556 10066
rect 3516 9444 3568 9450
rect 3516 9386 3568 9392
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3620 8634 3648 10406
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3712 8430 3740 11494
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 3804 7886 3832 19450
rect 3896 8634 3924 19774
rect 3988 18222 4016 20742
rect 4172 20058 4200 21422
rect 4436 21344 4488 21350
rect 4436 21286 4488 21292
rect 4528 21344 4580 21350
rect 4528 21286 4580 21292
rect 4344 20936 4396 20942
rect 4344 20878 4396 20884
rect 4252 20324 4304 20330
rect 4252 20266 4304 20272
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4068 19848 4120 19854
rect 4066 19816 4068 19825
rect 4120 19816 4122 19825
rect 4066 19751 4122 19760
rect 4172 19174 4200 19994
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 4160 18828 4212 18834
rect 4160 18770 4212 18776
rect 4172 18426 4200 18770
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 4066 17776 4122 17785
rect 4066 17711 4068 17720
rect 4120 17711 4122 17720
rect 4068 17682 4120 17688
rect 4160 17672 4212 17678
rect 3988 17620 4160 17626
rect 3988 17614 4212 17620
rect 3988 17598 4200 17614
rect 3988 16726 4016 17598
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 4066 17368 4122 17377
rect 4066 17303 4122 17312
rect 4080 17270 4108 17303
rect 4068 17264 4120 17270
rect 4068 17206 4120 17212
rect 4068 17128 4120 17134
rect 4066 17096 4068 17105
rect 4120 17096 4122 17105
rect 4066 17031 4122 17040
rect 4068 16992 4120 16998
rect 4066 16960 4068 16969
rect 4120 16960 4122 16969
rect 4066 16895 4122 16904
rect 3976 16720 4028 16726
rect 3976 16662 4028 16668
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 3976 15632 4028 15638
rect 3976 15574 4028 15580
rect 3988 14958 4016 15574
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 4080 14618 4108 16594
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4080 13802 4108 14554
rect 4068 13796 4120 13802
rect 4068 13738 4120 13744
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 3974 11792 4030 11801
rect 3974 11727 4030 11736
rect 3988 9110 4016 11727
rect 4080 11354 4108 12038
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4172 11234 4200 17478
rect 4264 17241 4292 20266
rect 4356 17898 4384 20878
rect 4448 20602 4476 21286
rect 4436 20596 4488 20602
rect 4436 20538 4488 20544
rect 4448 19990 4476 20538
rect 4540 20398 4568 21286
rect 4654 20700 4950 20720
rect 4710 20698 4734 20700
rect 4790 20698 4814 20700
rect 4870 20698 4894 20700
rect 4732 20646 4734 20698
rect 4796 20646 4808 20698
rect 4870 20646 4872 20698
rect 4710 20644 4734 20646
rect 4790 20644 4814 20646
rect 4870 20644 4894 20646
rect 4654 20624 4950 20644
rect 4528 20392 4580 20398
rect 4528 20334 4580 20340
rect 4436 19984 4488 19990
rect 4436 19926 4488 19932
rect 4434 19816 4490 19825
rect 4434 19751 4490 19760
rect 4448 18057 4476 19751
rect 4540 19514 4568 20334
rect 5000 20058 5028 23038
rect 5264 21344 5316 21350
rect 5264 21286 5316 21292
rect 5172 21004 5224 21010
rect 5172 20946 5224 20952
rect 5080 20800 5132 20806
rect 5080 20742 5132 20748
rect 5092 20466 5120 20742
rect 5080 20460 5132 20466
rect 5080 20402 5132 20408
rect 4988 20052 5040 20058
rect 4988 19994 5040 20000
rect 4986 19952 5042 19961
rect 5092 19922 5120 20402
rect 4986 19887 5042 19896
rect 5080 19916 5132 19922
rect 4654 19612 4950 19632
rect 4710 19610 4734 19612
rect 4790 19610 4814 19612
rect 4870 19610 4894 19612
rect 4732 19558 4734 19610
rect 4796 19558 4808 19610
rect 4870 19558 4872 19610
rect 4710 19556 4734 19558
rect 4790 19556 4814 19558
rect 4870 19556 4894 19558
rect 4654 19536 4950 19556
rect 4528 19508 4580 19514
rect 4528 19450 4580 19456
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4724 18970 4752 19110
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4816 18850 4844 18906
rect 4632 18822 4844 18850
rect 4632 18766 4660 18822
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4654 18524 4950 18544
rect 4710 18522 4734 18524
rect 4790 18522 4814 18524
rect 4870 18522 4894 18524
rect 4732 18470 4734 18522
rect 4796 18470 4808 18522
rect 4870 18470 4872 18522
rect 4710 18468 4734 18470
rect 4790 18468 4814 18470
rect 4870 18468 4894 18470
rect 4654 18448 4950 18468
rect 4434 18048 4490 18057
rect 4434 17983 4490 17992
rect 4356 17870 4568 17898
rect 4436 17740 4488 17746
rect 4436 17682 4488 17688
rect 4448 17338 4476 17682
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4436 17332 4488 17338
rect 4436 17274 4488 17280
rect 4250 17232 4306 17241
rect 4250 17167 4306 17176
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4264 16794 4292 16934
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 4356 16590 4384 17274
rect 4540 17252 4568 17870
rect 4804 17672 4856 17678
rect 4802 17640 4804 17649
rect 4856 17640 4858 17649
rect 4802 17575 4858 17584
rect 4654 17436 4950 17456
rect 4710 17434 4734 17436
rect 4790 17434 4814 17436
rect 4870 17434 4894 17436
rect 4732 17382 4734 17434
rect 4796 17382 4808 17434
rect 4870 17382 4872 17434
rect 4710 17380 4734 17382
rect 4790 17380 4814 17382
rect 4870 17380 4894 17382
rect 4654 17360 4950 17380
rect 4620 17264 4672 17270
rect 4434 17232 4490 17241
rect 4540 17224 4620 17252
rect 4620 17206 4672 17212
rect 4434 17167 4490 17176
rect 4712 17196 4764 17202
rect 4448 16640 4476 17167
rect 4712 17138 4764 17144
rect 4724 16833 4752 17138
rect 4804 16992 4856 16998
rect 5000 16946 5028 19887
rect 5080 19858 5132 19864
rect 5080 19712 5132 19718
rect 5080 19654 5132 19660
rect 5092 19310 5120 19654
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 5080 18624 5132 18630
rect 5080 18566 5132 18572
rect 5092 17338 5120 18566
rect 5184 17338 5212 20946
rect 5276 20262 5304 21286
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 5368 19514 5396 23920
rect 6012 23066 6040 23920
rect 6012 23038 6408 23066
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5448 21072 5500 21078
rect 5448 21014 5500 21020
rect 5460 20262 5488 21014
rect 5448 20256 5500 20262
rect 5448 20198 5500 20204
rect 5448 20052 5500 20058
rect 5448 19994 5500 20000
rect 5460 19854 5488 19994
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 5356 19508 5408 19514
rect 5356 19450 5408 19456
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5264 19236 5316 19242
rect 5264 19178 5316 19184
rect 5276 18698 5304 19178
rect 5264 18692 5316 18698
rect 5264 18634 5316 18640
rect 5460 18578 5488 19450
rect 5552 19378 5580 21490
rect 6092 21412 6144 21418
rect 6092 21354 6144 21360
rect 5816 21344 5868 21350
rect 5816 21286 5868 21292
rect 5828 19990 5856 21286
rect 5816 19984 5868 19990
rect 5816 19926 5868 19932
rect 6000 19712 6052 19718
rect 6000 19654 6052 19660
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 5724 19168 5776 19174
rect 5724 19110 5776 19116
rect 5736 18902 5764 19110
rect 5724 18896 5776 18902
rect 5724 18838 5776 18844
rect 5276 18550 5488 18578
rect 5814 18592 5870 18601
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 4804 16934 4856 16940
rect 4710 16824 4766 16833
rect 4710 16759 4766 16768
rect 4816 16726 4844 16934
rect 4908 16918 5028 16946
rect 4804 16720 4856 16726
rect 4804 16662 4856 16668
rect 4908 16658 4936 16918
rect 4896 16652 4948 16658
rect 4448 16612 4568 16640
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4434 16552 4490 16561
rect 4434 16487 4490 16496
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 4264 15638 4292 16050
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4252 15632 4304 15638
rect 4252 15574 4304 15580
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 4264 14074 4292 14894
rect 4356 14278 4384 15846
rect 4448 15570 4476 16487
rect 4540 16114 4568 16612
rect 4896 16594 4948 16600
rect 4654 16348 4950 16368
rect 4710 16346 4734 16348
rect 4790 16346 4814 16348
rect 4870 16346 4894 16348
rect 4732 16294 4734 16346
rect 4796 16294 4808 16346
rect 4870 16294 4872 16346
rect 4710 16292 4734 16294
rect 4790 16292 4814 16294
rect 4870 16292 4894 16294
rect 4654 16272 4950 16292
rect 4528 16108 4580 16114
rect 4528 16050 4580 16056
rect 4896 16040 4948 16046
rect 4896 15982 4948 15988
rect 4908 15910 4936 15982
rect 4896 15904 4948 15910
rect 4948 15864 5028 15892
rect 4896 15846 4948 15852
rect 4436 15564 4488 15570
rect 4436 15506 4488 15512
rect 5000 15434 5028 15864
rect 4988 15428 5040 15434
rect 4988 15370 5040 15376
rect 4654 15260 4950 15280
rect 4710 15258 4734 15260
rect 4790 15258 4814 15260
rect 4870 15258 4894 15260
rect 4732 15206 4734 15258
rect 4796 15206 4808 15258
rect 4870 15206 4872 15258
rect 4710 15204 4734 15206
rect 4790 15204 4814 15206
rect 4870 15204 4894 15206
rect 4654 15184 4950 15204
rect 5000 14822 5028 15370
rect 4988 14816 5040 14822
rect 5092 14804 5120 17274
rect 5276 17218 5304 18550
rect 5814 18527 5870 18536
rect 5632 18148 5684 18154
rect 5632 18090 5684 18096
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 5184 17190 5304 17218
rect 5184 16674 5212 17190
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5276 16794 5304 16934
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 5184 16646 5304 16674
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5184 14958 5212 15846
rect 5276 15366 5304 16646
rect 5368 15745 5396 17274
rect 5460 16794 5488 17478
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5552 17105 5580 17274
rect 5538 17096 5594 17105
rect 5538 17031 5594 17040
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5354 15736 5410 15745
rect 5354 15671 5410 15680
rect 5460 15620 5488 16594
rect 5538 16144 5594 16153
rect 5538 16079 5540 16088
rect 5592 16079 5594 16088
rect 5540 16050 5592 16056
rect 5359 15592 5488 15620
rect 5359 15484 5387 15592
rect 5448 15496 5500 15502
rect 5359 15456 5396 15484
rect 5264 15360 5316 15366
rect 5264 15302 5316 15308
rect 5368 15026 5396 15456
rect 5448 15438 5500 15444
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 5172 14952 5224 14958
rect 5172 14894 5224 14900
rect 5092 14776 5212 14804
rect 4988 14758 5040 14764
rect 5000 14634 5028 14758
rect 5000 14606 5120 14634
rect 4434 14512 4490 14521
rect 4434 14447 4490 14456
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4252 14068 4304 14074
rect 4252 14010 4304 14016
rect 4356 13326 4384 14214
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 4356 12986 4384 13126
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4448 12866 4476 14447
rect 4712 14408 4764 14414
rect 4710 14376 4712 14385
rect 4764 14376 4766 14385
rect 4710 14311 4766 14320
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 4654 14172 4950 14192
rect 4710 14170 4734 14172
rect 4790 14170 4814 14172
rect 4870 14170 4894 14172
rect 4732 14118 4734 14170
rect 4796 14118 4808 14170
rect 4870 14118 4872 14170
rect 4710 14116 4734 14118
rect 4790 14116 4814 14118
rect 4870 14116 4894 14118
rect 4654 14096 4950 14116
rect 5000 13870 5028 14214
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 4528 13796 4580 13802
rect 4528 13738 4580 13744
rect 4540 12889 4568 13738
rect 4988 13456 5040 13462
rect 4988 13398 5040 13404
rect 4654 13084 4950 13104
rect 4710 13082 4734 13084
rect 4790 13082 4814 13084
rect 4870 13082 4894 13084
rect 4732 13030 4734 13082
rect 4796 13030 4808 13082
rect 4870 13030 4872 13082
rect 4710 13028 4734 13030
rect 4790 13028 4814 13030
rect 4870 13028 4894 13030
rect 4654 13008 4950 13028
rect 5000 12986 5028 13398
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 4080 11206 4200 11234
rect 4264 12838 4476 12866
rect 4526 12880 4582 12889
rect 4080 9926 4108 11206
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4172 10606 4200 11086
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 4172 9654 4200 10542
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 4080 7206 4108 8502
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 2976 3126 3004 7142
rect 4080 6322 4108 7142
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4172 5914 4200 8298
rect 4264 7274 4292 12838
rect 5092 12866 5120 14606
rect 4526 12815 4582 12824
rect 5000 12838 5120 12866
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 4526 12744 4582 12753
rect 4356 11830 4384 12718
rect 4436 12708 4488 12714
rect 4526 12679 4582 12688
rect 4436 12650 4488 12656
rect 4448 12442 4476 12650
rect 4436 12436 4488 12442
rect 4436 12378 4488 12384
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 4344 11824 4396 11830
rect 4344 11766 4396 11772
rect 4448 11762 4476 12038
rect 4436 11756 4488 11762
rect 4436 11698 4488 11704
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 4356 9178 4384 11018
rect 4448 10810 4476 11154
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4448 10198 4476 10746
rect 4436 10192 4488 10198
rect 4436 10134 4488 10140
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4342 8528 4398 8537
rect 4342 8463 4398 8472
rect 4356 7954 4384 8463
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4252 7268 4304 7274
rect 4252 7210 4304 7216
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4448 5846 4476 9862
rect 4540 6730 4568 12679
rect 4654 11996 4950 12016
rect 4710 11994 4734 11996
rect 4790 11994 4814 11996
rect 4870 11994 4894 11996
rect 4732 11942 4734 11994
rect 4796 11942 4808 11994
rect 4870 11942 4872 11994
rect 4710 11940 4734 11942
rect 4790 11940 4814 11942
rect 4870 11940 4894 11942
rect 4654 11920 4950 11940
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4724 11150 4752 11698
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4908 11218 4936 11630
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4712 11144 4764 11150
rect 4710 11112 4712 11121
rect 4764 11112 4766 11121
rect 4710 11047 4766 11056
rect 4654 10908 4950 10928
rect 4710 10906 4734 10908
rect 4790 10906 4814 10908
rect 4870 10906 4894 10908
rect 4732 10854 4734 10906
rect 4796 10854 4808 10906
rect 4870 10854 4872 10906
rect 4710 10852 4734 10854
rect 4790 10852 4814 10854
rect 4870 10852 4894 10854
rect 4654 10832 4950 10852
rect 4802 10296 4858 10305
rect 4802 10231 4804 10240
rect 4856 10231 4858 10240
rect 4804 10202 4856 10208
rect 4654 9820 4950 9840
rect 4710 9818 4734 9820
rect 4790 9818 4814 9820
rect 4870 9818 4894 9820
rect 4732 9766 4734 9818
rect 4796 9766 4808 9818
rect 4870 9766 4872 9818
rect 4710 9764 4734 9766
rect 4790 9764 4814 9766
rect 4870 9764 4894 9766
rect 4654 9744 4950 9764
rect 4802 9616 4858 9625
rect 4802 9551 4858 9560
rect 4816 9382 4844 9551
rect 4896 9512 4948 9518
rect 4894 9480 4896 9489
rect 4948 9480 4950 9489
rect 4894 9415 4950 9424
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4908 9042 4936 9415
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4654 8732 4950 8752
rect 4710 8730 4734 8732
rect 4790 8730 4814 8732
rect 4870 8730 4894 8732
rect 4732 8678 4734 8730
rect 4796 8678 4808 8730
rect 4870 8678 4872 8730
rect 4710 8676 4734 8678
rect 4790 8676 4814 8678
rect 4870 8676 4894 8678
rect 4654 8656 4950 8676
rect 5000 7886 5028 12838
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 5092 9178 5120 12242
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5092 8090 5120 8978
rect 5184 8498 5212 14776
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5356 14476 5408 14482
rect 5356 14418 5408 14424
rect 5276 9586 5304 14418
rect 5368 13530 5396 14418
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 5368 12238 5396 12854
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5276 9110 5304 9318
rect 5368 9178 5396 12038
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5368 8566 5396 8910
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 4654 7644 4950 7664
rect 4710 7642 4734 7644
rect 4790 7642 4814 7644
rect 4870 7642 4894 7644
rect 4732 7590 4734 7642
rect 4796 7590 4808 7642
rect 4870 7590 4872 7642
rect 4710 7588 4734 7590
rect 4790 7588 4814 7590
rect 4870 7588 4894 7590
rect 4654 7568 4950 7588
rect 5092 7546 5120 7754
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 4988 7472 5040 7478
rect 4988 7414 5040 7420
rect 5000 6866 5028 7414
rect 5170 6896 5226 6905
rect 4988 6860 5040 6866
rect 5170 6831 5226 6840
rect 4988 6802 5040 6808
rect 5184 6798 5212 6831
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5460 6730 5488 15438
rect 5538 13424 5594 13433
rect 5538 13359 5594 13368
rect 5552 13258 5580 13359
rect 5540 13252 5592 13258
rect 5540 13194 5592 13200
rect 5538 13016 5594 13025
rect 5538 12951 5594 12960
rect 5552 12782 5580 12951
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5540 12368 5592 12374
rect 5538 12336 5540 12345
rect 5592 12336 5594 12345
rect 5538 12271 5594 12280
rect 5538 11792 5594 11801
rect 5538 11727 5594 11736
rect 5552 11014 5580 11727
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5552 10266 5580 10474
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5552 9586 5580 10202
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5538 9072 5594 9081
rect 5538 9007 5594 9016
rect 5552 8498 5580 9007
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5644 8430 5672 18090
rect 5724 18080 5776 18086
rect 5828 18068 5856 18527
rect 5776 18040 5856 18068
rect 5724 18022 5776 18028
rect 5722 17640 5778 17649
rect 5722 17575 5778 17584
rect 5736 16590 5764 17575
rect 5724 16584 5776 16590
rect 5724 16526 5776 16532
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5736 15609 5764 16050
rect 5722 15600 5778 15609
rect 5722 15535 5778 15544
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5736 13530 5764 13806
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5736 13025 5764 13466
rect 5722 13016 5778 13025
rect 5722 12951 5778 12960
rect 5828 12628 5856 18040
rect 5908 18080 5960 18086
rect 5908 18022 5960 18028
rect 5920 17746 5948 18022
rect 5908 17740 5960 17746
rect 5908 17682 5960 17688
rect 6012 17202 6040 19654
rect 6104 19553 6132 21354
rect 6276 21344 6328 21350
rect 6276 21286 6328 21292
rect 6288 20398 6316 21286
rect 6276 20392 6328 20398
rect 6276 20334 6328 20340
rect 6288 19786 6316 20334
rect 6276 19780 6328 19786
rect 6276 19722 6328 19728
rect 6090 19544 6146 19553
rect 6090 19479 6146 19488
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 6000 17060 6052 17066
rect 6000 17002 6052 17008
rect 6012 16833 6040 17002
rect 5998 16824 6054 16833
rect 5920 16782 5998 16810
rect 5920 16250 5948 16782
rect 5998 16759 6054 16768
rect 6000 16652 6052 16658
rect 6000 16594 6052 16600
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 6012 15570 6040 16594
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 5908 15360 5960 15366
rect 5908 15302 5960 15308
rect 5920 12753 5948 15302
rect 6012 14822 6040 15506
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 5906 12744 5962 12753
rect 5906 12679 5962 12688
rect 5828 12600 5948 12628
rect 5816 12368 5868 12374
rect 5816 12310 5868 12316
rect 5722 12064 5778 12073
rect 5722 11999 5778 12008
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5630 7984 5686 7993
rect 5630 7919 5686 7928
rect 5644 7750 5672 7919
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5632 7472 5684 7478
rect 5736 7460 5764 11999
rect 5828 11354 5856 12310
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5828 10198 5856 11290
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5684 7432 5764 7460
rect 5632 7414 5684 7420
rect 5828 7206 5856 9590
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 4528 6724 4580 6730
rect 4528 6666 4580 6672
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 4654 6556 4950 6576
rect 4710 6554 4734 6556
rect 4790 6554 4814 6556
rect 4870 6554 4894 6556
rect 4732 6502 4734 6554
rect 4796 6502 4808 6554
rect 4870 6502 4872 6554
rect 4710 6500 4734 6502
rect 4790 6500 4814 6502
rect 4870 6500 4894 6502
rect 4654 6480 4950 6500
rect 5644 6458 5672 6734
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 4436 5840 4488 5846
rect 4436 5782 4488 5788
rect 5920 5710 5948 12600
rect 6012 6254 6040 14758
rect 6104 12481 6132 17478
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 6196 15994 6224 16594
rect 6288 16114 6316 18022
rect 6276 16108 6328 16114
rect 6276 16050 6328 16056
rect 6196 15966 6316 15994
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6090 12472 6146 12481
rect 6090 12407 6146 12416
rect 6090 12200 6146 12209
rect 6090 12135 6146 12144
rect 6104 7342 6132 12135
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6196 7002 6224 14758
rect 6288 13870 6316 15966
rect 6276 13864 6328 13870
rect 6276 13806 6328 13812
rect 6276 13728 6328 13734
rect 6276 13670 6328 13676
rect 6288 13462 6316 13670
rect 6276 13456 6328 13462
rect 6276 13398 6328 13404
rect 6380 13274 6408 23038
rect 6460 21412 6512 21418
rect 6460 21354 6512 21360
rect 6472 21010 6500 21354
rect 6460 21004 6512 21010
rect 6460 20946 6512 20952
rect 6472 20602 6500 20946
rect 6552 20800 6604 20806
rect 6552 20742 6604 20748
rect 6564 20602 6592 20742
rect 6460 20596 6512 20602
rect 6460 20538 6512 20544
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 6460 19372 6512 19378
rect 6460 19314 6512 19320
rect 6472 18630 6500 19314
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 6460 17672 6512 17678
rect 6564 17660 6592 20538
rect 6656 20330 6684 23920
rect 7300 22658 7328 23920
rect 7116 22630 7328 22658
rect 7012 21412 7064 21418
rect 7012 21354 7064 21360
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 6828 21004 6880 21010
rect 6828 20946 6880 20952
rect 6644 20324 6696 20330
rect 6644 20266 6696 20272
rect 6840 19854 6868 20946
rect 6932 20058 6960 21286
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 6840 19174 6868 19790
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6840 18970 6868 19110
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6840 18222 6868 18566
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6512 17632 6592 17660
rect 6460 17614 6512 17620
rect 6564 17134 6592 17632
rect 6828 17264 6880 17270
rect 7024 17252 7052 21354
rect 6880 17224 7052 17252
rect 6828 17206 6880 17212
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6472 15502 6500 16390
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6840 16046 6868 16186
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6458 14512 6514 14521
rect 6458 14447 6460 14456
rect 6512 14447 6514 14456
rect 6460 14418 6512 14424
rect 6460 14340 6512 14346
rect 6460 14282 6512 14288
rect 6472 14006 6500 14282
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 6288 13246 6408 13274
rect 6288 10606 6316 13246
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6380 11830 6408 12174
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 6472 11370 6500 13806
rect 6380 11342 6500 11370
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 6380 10418 6408 11342
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6472 10810 6500 11154
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6288 10390 6408 10418
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 6288 5710 6316 10390
rect 6366 9480 6422 9489
rect 6472 9450 6500 10746
rect 6366 9415 6422 9424
rect 6460 9444 6512 9450
rect 6380 9382 6408 9415
rect 6460 9386 6512 9392
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6366 9208 6422 9217
rect 6564 9160 6592 15846
rect 6656 12866 6684 15982
rect 6736 15972 6788 15978
rect 6736 15914 6788 15920
rect 6748 15366 6776 15914
rect 6840 15638 6868 15982
rect 7116 15722 7144 22630
rect 7564 22024 7616 22030
rect 7564 21966 7616 21972
rect 7576 21622 7604 21966
rect 7564 21616 7616 21622
rect 7564 21558 7616 21564
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 7380 21344 7432 21350
rect 7380 21286 7432 21292
rect 7300 21078 7328 21286
rect 7392 21146 7420 21286
rect 7380 21140 7432 21146
rect 7380 21082 7432 21088
rect 7288 21072 7340 21078
rect 7288 21014 7340 21020
rect 7392 20398 7420 21082
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 7576 20602 7604 20878
rect 7564 20596 7616 20602
rect 7564 20538 7616 20544
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 7656 19780 7708 19786
rect 7656 19722 7708 19728
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 7194 19272 7250 19281
rect 7194 19207 7250 19216
rect 7208 18358 7236 19207
rect 7576 18766 7604 19654
rect 7288 18760 7340 18766
rect 7288 18702 7340 18708
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7196 18352 7248 18358
rect 7194 18320 7196 18329
rect 7248 18320 7250 18329
rect 7194 18255 7250 18264
rect 7300 16998 7328 18702
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7576 18290 7604 18566
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 7194 16824 7250 16833
rect 7194 16759 7250 16768
rect 6932 15694 7144 15722
rect 7208 15706 7236 16759
rect 7472 16448 7524 16454
rect 7472 16390 7524 16396
rect 7380 16108 7432 16114
rect 7300 16068 7380 16096
rect 7300 15910 7328 16068
rect 7380 16050 7432 16056
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7196 15700 7248 15706
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 6736 15360 6788 15366
rect 6736 15302 6788 15308
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6748 13734 6776 15098
rect 6840 14958 6868 15438
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6840 14278 6868 14894
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 6736 13320 6788 13326
rect 6840 13308 6868 14214
rect 6932 13530 6960 15694
rect 7196 15642 7248 15648
rect 7484 15638 7512 16390
rect 7472 15632 7524 15638
rect 7472 15574 7524 15580
rect 7104 15360 7156 15366
rect 7104 15302 7156 15308
rect 7116 14890 7144 15302
rect 7104 14884 7156 14890
rect 7104 14826 7156 14832
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 7024 13462 7052 14214
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 6788 13280 6868 13308
rect 6736 13262 6788 13268
rect 6656 12838 6776 12866
rect 6644 12368 6696 12374
rect 6644 12310 6696 12316
rect 6656 12209 6684 12310
rect 6642 12200 6698 12209
rect 6642 12135 6698 12144
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6656 10538 6684 11154
rect 6644 10532 6696 10538
rect 6644 10474 6696 10480
rect 6656 10130 6684 10474
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6644 9444 6696 9450
rect 6644 9386 6696 9392
rect 6366 9143 6422 9152
rect 6380 8974 6408 9143
rect 6472 9132 6592 9160
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6380 6662 6408 8774
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 6472 5846 6500 9132
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6564 7002 6592 8910
rect 6656 7546 6684 9386
rect 6748 8634 6776 12838
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6840 12374 6868 12718
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 6828 12368 6880 12374
rect 6828 12310 6880 12316
rect 6840 11762 6868 12310
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6932 11626 6960 12378
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6734 8528 6790 8537
rect 6734 8463 6790 8472
rect 6748 8430 6776 8463
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6656 6730 6684 7346
rect 6644 6724 6696 6730
rect 6644 6666 6696 6672
rect 6748 6610 6776 8230
rect 6840 6934 6868 11086
rect 6932 10266 6960 11562
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6932 7002 6960 10066
rect 7024 9722 7052 13398
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 7010 9616 7066 9625
rect 7010 9551 7066 9560
rect 7024 9518 7052 9551
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 7024 9178 7052 9318
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 7012 8968 7064 8974
rect 7010 8936 7012 8945
rect 7064 8936 7066 8945
rect 7010 8871 7066 8880
rect 7010 8120 7066 8129
rect 7010 8055 7012 8064
rect 7064 8055 7066 8064
rect 7012 8026 7064 8032
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7024 7002 7052 7822
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 6828 6928 6880 6934
rect 7116 6882 7144 14826
rect 7380 14068 7432 14074
rect 7380 14010 7432 14016
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 7208 13841 7236 13874
rect 7194 13832 7250 13841
rect 7194 13767 7250 13776
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7288 13728 7340 13734
rect 7288 13670 7340 13676
rect 7208 13462 7236 13670
rect 7196 13456 7248 13462
rect 7196 13398 7248 13404
rect 7300 13394 7328 13670
rect 7392 13530 7420 14010
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7484 13274 7512 15574
rect 7562 14376 7618 14385
rect 7562 14311 7618 14320
rect 7208 13246 7512 13274
rect 7208 9058 7236 13246
rect 7470 13152 7526 13161
rect 7470 13087 7526 13096
rect 7286 12744 7342 12753
rect 7484 12714 7512 13087
rect 7286 12679 7342 12688
rect 7472 12708 7524 12714
rect 7300 10810 7328 12679
rect 7472 12650 7524 12656
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7392 12374 7420 12582
rect 7380 12368 7432 12374
rect 7380 12310 7432 12316
rect 7288 10804 7340 10810
rect 7288 10746 7340 10752
rect 7300 9382 7328 10746
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7286 9208 7342 9217
rect 7286 9143 7288 9152
rect 7340 9143 7342 9152
rect 7288 9114 7340 9120
rect 7208 9030 7328 9058
rect 7194 8936 7250 8945
rect 7194 8871 7250 8880
rect 7208 7886 7236 8871
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7196 7744 7248 7750
rect 7194 7712 7196 7721
rect 7248 7712 7250 7721
rect 7194 7647 7250 7656
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7208 6934 7236 7142
rect 6828 6870 6880 6876
rect 6932 6854 7144 6882
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 6932 6798 6960 6854
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 7012 6656 7064 6662
rect 6748 6582 6960 6610
rect 7012 6598 7064 6604
rect 6550 5944 6606 5953
rect 6550 5879 6552 5888
rect 6604 5879 6606 5888
rect 6552 5850 6604 5856
rect 6460 5840 6512 5846
rect 6460 5782 6512 5788
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 4654 5468 4950 5488
rect 4710 5466 4734 5468
rect 4790 5466 4814 5468
rect 4870 5466 4894 5468
rect 4732 5414 4734 5466
rect 4796 5414 4808 5466
rect 4870 5414 4872 5466
rect 4710 5412 4734 5414
rect 4790 5412 4814 5414
rect 4870 5412 4894 5414
rect 4654 5392 4950 5412
rect 6932 4486 6960 6582
rect 7024 5914 7052 6598
rect 7300 6322 7328 9030
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 7392 5166 7420 12310
rect 7472 11620 7524 11626
rect 7472 11562 7524 11568
rect 7484 5846 7512 11562
rect 7576 10198 7604 14311
rect 7564 10192 7616 10198
rect 7564 10134 7616 10140
rect 7668 9500 7696 19722
rect 7840 19440 7892 19446
rect 7840 19382 7892 19388
rect 7852 19174 7880 19382
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 7944 18902 7972 23920
rect 8588 21690 8616 23920
rect 8116 21684 8168 21690
rect 8116 21626 8168 21632
rect 8576 21684 8628 21690
rect 8576 21626 8628 21632
rect 8024 20392 8076 20398
rect 8024 20334 8076 20340
rect 8036 19922 8064 20334
rect 8128 20040 8156 21626
rect 9128 21480 9180 21486
rect 9128 21422 9180 21428
rect 8852 21412 8904 21418
rect 8852 21354 8904 21360
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8760 21344 8812 21350
rect 8760 21286 8812 21292
rect 8353 21244 8649 21264
rect 8409 21242 8433 21244
rect 8489 21242 8513 21244
rect 8569 21242 8593 21244
rect 8431 21190 8433 21242
rect 8495 21190 8507 21242
rect 8569 21190 8571 21242
rect 8409 21188 8433 21190
rect 8489 21188 8513 21190
rect 8569 21188 8593 21190
rect 8353 21168 8649 21188
rect 8680 21078 8708 21286
rect 8208 21072 8260 21078
rect 8208 21014 8260 21020
rect 8668 21072 8720 21078
rect 8668 21014 8720 21020
rect 8220 20602 8248 21014
rect 8772 20602 8800 21286
rect 8864 21146 8892 21354
rect 8852 21140 8904 21146
rect 8852 21082 8904 21088
rect 8208 20596 8260 20602
rect 8208 20538 8260 20544
rect 8760 20596 8812 20602
rect 8760 20538 8812 20544
rect 8353 20156 8649 20176
rect 8409 20154 8433 20156
rect 8489 20154 8513 20156
rect 8569 20154 8593 20156
rect 8431 20102 8433 20154
rect 8495 20102 8507 20154
rect 8569 20102 8571 20154
rect 8409 20100 8433 20102
rect 8489 20100 8513 20102
rect 8569 20100 8593 20102
rect 8353 20080 8649 20100
rect 8128 20012 8524 20040
rect 8024 19916 8076 19922
rect 8024 19858 8076 19864
rect 8208 19916 8260 19922
rect 8208 19858 8260 19864
rect 7932 18896 7984 18902
rect 7932 18838 7984 18844
rect 7932 18760 7984 18766
rect 8036 18714 8064 19858
rect 8220 19802 8248 19858
rect 8128 19774 8248 19802
rect 8128 19174 8156 19774
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8312 19310 8340 19654
rect 8300 19304 8352 19310
rect 8300 19246 8352 19252
rect 8116 19168 8168 19174
rect 8312 19156 8340 19246
rect 8496 19242 8524 20012
rect 8772 19242 8800 20538
rect 8864 20330 8892 21082
rect 8852 20324 8904 20330
rect 8852 20266 8904 20272
rect 9036 20324 9088 20330
rect 9036 20266 9088 20272
rect 9048 19825 9076 20266
rect 9034 19816 9090 19825
rect 9034 19751 9090 19760
rect 8484 19236 8536 19242
rect 8484 19178 8536 19184
rect 8668 19236 8720 19242
rect 8668 19178 8720 19184
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8116 19110 8168 19116
rect 8220 19128 8340 19156
rect 8220 18902 8248 19128
rect 8353 19068 8649 19088
rect 8409 19066 8433 19068
rect 8489 19066 8513 19068
rect 8569 19066 8593 19068
rect 8431 19014 8433 19066
rect 8495 19014 8507 19066
rect 8569 19014 8571 19066
rect 8409 19012 8433 19014
rect 8489 19012 8513 19014
rect 8569 19012 8593 19014
rect 8353 18992 8649 19012
rect 8208 18896 8260 18902
rect 8208 18838 8260 18844
rect 8300 18896 8352 18902
rect 8300 18838 8352 18844
rect 7984 18708 8064 18714
rect 7932 18702 8064 18708
rect 7944 18686 8064 18702
rect 7932 18284 7984 18290
rect 7932 18226 7984 18232
rect 7840 17536 7892 17542
rect 7838 17504 7840 17513
rect 7892 17504 7894 17513
rect 7838 17439 7894 17448
rect 7852 17134 7880 17439
rect 7840 17128 7892 17134
rect 7840 17070 7892 17076
rect 7840 16992 7892 16998
rect 7840 16934 7892 16940
rect 7748 16720 7800 16726
rect 7748 16662 7800 16668
rect 7760 13938 7788 16662
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7760 12209 7788 12310
rect 7746 12200 7802 12209
rect 7746 12135 7802 12144
rect 7852 11937 7880 16934
rect 7944 16726 7972 18226
rect 8036 18204 8064 18686
rect 8312 18358 8340 18838
rect 8680 18465 8708 19178
rect 8390 18456 8446 18465
rect 8390 18391 8446 18400
rect 8666 18456 8722 18465
rect 8666 18391 8722 18400
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 8404 18222 8432 18391
rect 8208 18216 8260 18222
rect 8036 18176 8208 18204
rect 8208 18158 8260 18164
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 8220 17796 8248 18158
rect 8944 18080 8996 18086
rect 8942 18048 8944 18057
rect 8996 18048 8998 18057
rect 8353 17980 8649 18000
rect 8942 17983 8998 17992
rect 8409 17978 8433 17980
rect 8489 17978 8513 17980
rect 8569 17978 8593 17980
rect 8431 17926 8433 17978
rect 8495 17926 8507 17978
rect 8569 17926 8571 17978
rect 8409 17924 8433 17926
rect 8489 17924 8513 17926
rect 8569 17924 8593 17926
rect 8353 17904 8649 17924
rect 8220 17768 8340 17796
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 7932 16720 7984 16726
rect 7932 16662 7984 16668
rect 8036 12374 8064 17478
rect 8312 17134 8340 17768
rect 8760 17740 8812 17746
rect 8760 17682 8812 17688
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8588 17241 8616 17614
rect 8574 17232 8630 17241
rect 8574 17167 8630 17176
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 8353 16892 8649 16912
rect 8409 16890 8433 16892
rect 8489 16890 8513 16892
rect 8569 16890 8593 16892
rect 8431 16838 8433 16890
rect 8495 16838 8507 16890
rect 8569 16838 8571 16890
rect 8409 16836 8433 16838
rect 8489 16836 8513 16838
rect 8569 16836 8593 16838
rect 8353 16816 8649 16836
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 8220 14929 8248 15846
rect 8353 15804 8649 15824
rect 8409 15802 8433 15804
rect 8489 15802 8513 15804
rect 8569 15802 8593 15804
rect 8431 15750 8433 15802
rect 8495 15750 8507 15802
rect 8569 15750 8571 15802
rect 8409 15748 8433 15750
rect 8489 15748 8513 15750
rect 8569 15748 8593 15750
rect 8353 15728 8649 15748
rect 8668 15564 8720 15570
rect 8668 15506 8720 15512
rect 8206 14920 8262 14929
rect 8206 14855 8262 14864
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8220 14482 8248 14758
rect 8353 14716 8649 14736
rect 8409 14714 8433 14716
rect 8489 14714 8513 14716
rect 8569 14714 8593 14716
rect 8431 14662 8433 14714
rect 8495 14662 8507 14714
rect 8569 14662 8571 14714
rect 8409 14660 8433 14662
rect 8489 14660 8513 14662
rect 8569 14660 8593 14662
rect 8353 14640 8649 14660
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8680 14278 8708 15506
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 8116 13184 8168 13190
rect 8114 13152 8116 13161
rect 8168 13152 8170 13161
rect 8114 13087 8170 13096
rect 8220 12442 8248 13806
rect 8353 13628 8649 13648
rect 8409 13626 8433 13628
rect 8489 13626 8513 13628
rect 8569 13626 8593 13628
rect 8431 13574 8433 13626
rect 8495 13574 8507 13626
rect 8569 13574 8571 13626
rect 8409 13572 8433 13574
rect 8489 13572 8513 13574
rect 8569 13572 8593 13574
rect 8353 13552 8649 13572
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8496 12850 8524 13330
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8353 12540 8649 12560
rect 8409 12538 8433 12540
rect 8489 12538 8513 12540
rect 8569 12538 8593 12540
rect 8431 12486 8433 12538
rect 8495 12486 8507 12538
rect 8569 12486 8571 12538
rect 8409 12484 8433 12486
rect 8489 12484 8513 12486
rect 8569 12484 8593 12486
rect 8353 12464 8649 12484
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8024 12368 8076 12374
rect 8024 12310 8076 12316
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 7838 11928 7894 11937
rect 7838 11863 7894 11872
rect 8404 11626 8432 12038
rect 8392 11620 8444 11626
rect 8392 11562 8444 11568
rect 7840 11552 7892 11558
rect 8588 11540 8616 12038
rect 8680 11762 8708 14010
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8772 11558 8800 17682
rect 9036 17672 9088 17678
rect 9036 17614 9088 17620
rect 8850 17096 8906 17105
rect 8850 17031 8906 17040
rect 8944 17060 8996 17066
rect 8864 16998 8892 17031
rect 8944 17002 8996 17008
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8850 16688 8906 16697
rect 8956 16658 8984 17002
rect 8850 16623 8906 16632
rect 8944 16652 8996 16658
rect 8864 13308 8892 16623
rect 8944 16594 8996 16600
rect 8944 16516 8996 16522
rect 8944 16458 8996 16464
rect 8956 15570 8984 16458
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 9048 15065 9076 17614
rect 9140 16153 9168 21422
rect 9232 20058 9260 23920
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9496 20528 9548 20534
rect 9416 20476 9496 20482
rect 9416 20470 9548 20476
rect 9416 20454 9536 20470
rect 9220 20052 9272 20058
rect 9220 19994 9272 20000
rect 9416 17762 9444 20454
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9586 18864 9642 18873
rect 9496 18828 9548 18834
rect 9692 18834 9720 19654
rect 9784 19242 9812 20742
rect 9876 20058 9904 23920
rect 9956 21956 10008 21962
rect 9956 21898 10008 21904
rect 9968 21690 9996 21898
rect 9956 21684 10008 21690
rect 9956 21626 10008 21632
rect 10416 21480 10468 21486
rect 10416 21422 10468 21428
rect 10048 21004 10100 21010
rect 10048 20946 10100 20952
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9772 19236 9824 19242
rect 9772 19178 9824 19184
rect 9876 18970 9904 19858
rect 10060 19310 10088 20946
rect 10428 20942 10456 21422
rect 10416 20936 10468 20942
rect 10416 20878 10468 20884
rect 10428 20398 10456 20878
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10428 19854 10456 20334
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 10138 19544 10194 19553
rect 10138 19479 10140 19488
rect 10192 19479 10194 19488
rect 10140 19450 10192 19456
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 10232 19236 10284 19242
rect 10232 19178 10284 19184
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 9586 18799 9642 18808
rect 9680 18828 9732 18834
rect 9496 18770 9548 18776
rect 9324 17734 9444 17762
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 9232 16726 9260 17478
rect 9220 16720 9272 16726
rect 9220 16662 9272 16668
rect 9324 16561 9352 17734
rect 9404 17672 9456 17678
rect 9404 17614 9456 17620
rect 9310 16552 9366 16561
rect 9310 16487 9366 16496
rect 9126 16144 9182 16153
rect 9126 16079 9182 16088
rect 9312 16108 9364 16114
rect 9140 15570 9168 16079
rect 9312 16050 9364 16056
rect 9324 15910 9352 16050
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 9416 15586 9444 17614
rect 9508 17610 9536 18770
rect 9600 18426 9628 18799
rect 9680 18770 9732 18776
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9784 18465 9812 18702
rect 9770 18456 9826 18465
rect 9588 18420 9640 18426
rect 9770 18391 9772 18400
rect 9588 18362 9640 18368
rect 9824 18391 9826 18400
rect 9772 18362 9824 18368
rect 9784 18331 9812 18362
rect 9586 18320 9642 18329
rect 9586 18255 9642 18264
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9128 15564 9180 15570
rect 9416 15558 9450 15586
rect 9422 15552 9450 15558
rect 9422 15524 9490 15552
rect 9128 15506 9180 15512
rect 9126 15464 9182 15473
rect 9462 15416 9490 15524
rect 9126 15399 9182 15408
rect 9034 15056 9090 15065
rect 8956 15014 9034 15042
rect 8956 13462 8984 15014
rect 9034 14991 9090 15000
rect 9036 14408 9088 14414
rect 9036 14350 9088 14356
rect 8944 13456 8996 13462
rect 8944 13398 8996 13404
rect 8944 13320 8996 13326
rect 8864 13280 8944 13308
rect 8944 13262 8996 13268
rect 8956 12850 8984 13262
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8864 12345 8892 12582
rect 8850 12336 8906 12345
rect 8850 12271 8906 12280
rect 8956 11801 8984 12582
rect 9048 12073 9076 14350
rect 9140 12986 9168 15399
rect 9416 15388 9490 15416
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9232 14074 9260 15302
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9126 12880 9182 12889
rect 9126 12815 9182 12824
rect 9140 12646 9168 12815
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 9034 12064 9090 12073
rect 9034 11999 9090 12008
rect 8942 11792 8998 11801
rect 8852 11756 8904 11762
rect 8942 11727 8998 11736
rect 8852 11698 8904 11704
rect 8760 11552 8812 11558
rect 8588 11512 8708 11540
rect 7840 11494 7892 11500
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7760 10538 7788 11290
rect 7852 11218 7880 11494
rect 8353 11452 8649 11472
rect 8409 11450 8433 11452
rect 8489 11450 8513 11452
rect 8569 11450 8593 11452
rect 8431 11398 8433 11450
rect 8495 11398 8507 11450
rect 8569 11398 8571 11450
rect 8409 11396 8433 11398
rect 8489 11396 8513 11398
rect 8569 11396 8593 11398
rect 8353 11376 8649 11396
rect 8680 11336 8708 11512
rect 8760 11494 8812 11500
rect 8496 11308 8708 11336
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 7748 10532 7800 10538
rect 7748 10474 7800 10480
rect 7576 9472 7696 9500
rect 7576 9466 7604 9472
rect 7567 9438 7604 9466
rect 7567 9194 7595 9438
rect 7760 9432 7788 10474
rect 7852 9602 7880 11154
rect 7944 9722 7972 11154
rect 8496 10577 8524 11308
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8588 10810 8616 10950
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8482 10568 8538 10577
rect 8482 10503 8538 10512
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8220 10130 8248 10406
rect 8353 10364 8649 10384
rect 8409 10362 8433 10364
rect 8489 10362 8513 10364
rect 8569 10362 8593 10364
rect 8431 10310 8433 10362
rect 8495 10310 8507 10362
rect 8569 10310 8571 10362
rect 8409 10308 8433 10310
rect 8489 10308 8513 10310
rect 8569 10308 8593 10310
rect 8353 10288 8649 10308
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8312 10010 8340 10134
rect 8220 9982 8340 10010
rect 7932 9716 7984 9722
rect 7932 9658 7984 9664
rect 8220 9602 8248 9982
rect 8404 9908 8432 10134
rect 8312 9880 8432 9908
rect 8312 9625 8340 9880
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 7852 9574 7972 9602
rect 7751 9404 7788 9432
rect 7751 9330 7779 9404
rect 7944 9330 7972 9574
rect 8128 9574 8248 9602
rect 8298 9616 8354 9625
rect 8128 9353 8156 9574
rect 8298 9551 8354 9560
rect 8404 9364 8432 9658
rect 8680 9654 8708 11086
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8772 9897 8800 10542
rect 8758 9888 8814 9897
rect 8758 9823 8814 9832
rect 8668 9648 8720 9654
rect 8482 9616 8538 9625
rect 8668 9590 8720 9596
rect 8482 9551 8538 9560
rect 8496 9518 8524 9551
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8576 9444 8628 9450
rect 8760 9444 8812 9450
rect 8628 9404 8708 9432
rect 8576 9386 8628 9392
rect 7668 9302 7779 9330
rect 7852 9302 7972 9330
rect 8114 9344 8170 9353
rect 7668 9194 7696 9302
rect 7567 9166 7604 9194
rect 7668 9166 7788 9194
rect 7576 8634 7604 9166
rect 7656 8900 7708 8906
rect 7656 8842 7708 8848
rect 7668 8673 7696 8842
rect 7654 8664 7710 8673
rect 7564 8628 7616 8634
rect 7654 8599 7710 8608
rect 7564 8570 7616 8576
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7562 7848 7618 7857
rect 7562 7783 7564 7792
rect 7616 7783 7618 7792
rect 7564 7754 7616 7760
rect 7562 7712 7618 7721
rect 7562 7647 7618 7656
rect 7576 7274 7604 7647
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 4654 4380 4950 4400
rect 4710 4378 4734 4380
rect 4790 4378 4814 4380
rect 4870 4378 4894 4380
rect 4732 4326 4734 4378
rect 4796 4326 4808 4378
rect 4870 4326 4872 4378
rect 4710 4324 4734 4326
rect 4790 4324 4814 4326
rect 4870 4324 4894 4326
rect 4654 4304 4950 4324
rect 7576 3398 7604 6938
rect 7668 5914 7696 8366
rect 7760 6866 7788 9166
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7760 5710 7788 6258
rect 7852 5914 7880 9302
rect 8114 9279 8170 9288
rect 8220 9336 8432 9364
rect 7930 9208 7986 9217
rect 7930 9143 7986 9152
rect 7944 8362 7972 9143
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 7932 8016 7984 8022
rect 7930 7984 7932 7993
rect 7984 7984 7986 7993
rect 7930 7919 7986 7928
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7944 7721 7972 7822
rect 7930 7712 7986 7721
rect 7930 7647 7986 7656
rect 7930 7576 7986 7585
rect 7930 7511 7932 7520
rect 7984 7511 7986 7520
rect 7932 7482 7984 7488
rect 7930 7440 7986 7449
rect 7930 7375 7986 7384
rect 7944 7002 7972 7375
rect 7932 6996 7984 7002
rect 7932 6938 7984 6944
rect 7932 6724 7984 6730
rect 7932 6666 7984 6672
rect 7944 6390 7972 6666
rect 8036 6458 8064 8978
rect 8220 8906 8248 9336
rect 8353 9276 8649 9296
rect 8409 9274 8433 9276
rect 8489 9274 8513 9276
rect 8569 9274 8593 9276
rect 8431 9222 8433 9274
rect 8495 9222 8507 9274
rect 8569 9222 8571 9274
rect 8409 9220 8433 9222
rect 8489 9220 8513 9222
rect 8569 9220 8593 9222
rect 8353 9200 8649 9220
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 8208 8560 8260 8566
rect 8404 8537 8432 8842
rect 8208 8502 8260 8508
rect 8390 8528 8446 8537
rect 8220 7970 8248 8502
rect 8300 8492 8352 8498
rect 8390 8463 8392 8472
rect 8300 8434 8352 8440
rect 8444 8463 8446 8472
rect 8392 8434 8444 8440
rect 8312 8401 8340 8434
rect 8496 8430 8524 9046
rect 8680 9042 8708 9404
rect 8760 9386 8812 9392
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8772 8974 8800 9386
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8668 8900 8720 8906
rect 8588 8860 8668 8888
rect 8484 8424 8536 8430
rect 8298 8392 8354 8401
rect 8484 8366 8536 8372
rect 8588 8362 8616 8860
rect 8668 8842 8720 8848
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8298 8327 8354 8336
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8353 8188 8649 8208
rect 8409 8186 8433 8188
rect 8489 8186 8513 8188
rect 8569 8186 8593 8188
rect 8431 8134 8433 8186
rect 8495 8134 8507 8186
rect 8569 8134 8571 8186
rect 8409 8132 8433 8134
rect 8489 8132 8513 8134
rect 8569 8132 8593 8134
rect 8353 8112 8649 8132
rect 8680 8106 8708 8570
rect 8772 8265 8800 8774
rect 8758 8256 8814 8265
rect 8758 8191 8814 8200
rect 8864 8129 8892 11698
rect 9048 11694 9076 11999
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 8942 10976 8998 10985
rect 8942 10911 8998 10920
rect 8956 10198 8984 10911
rect 8944 10192 8996 10198
rect 8944 10134 8996 10140
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 8956 9761 8984 9862
rect 8942 9752 8998 9761
rect 8942 9687 8998 9696
rect 8956 9518 8984 9687
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8942 9344 8998 9353
rect 8942 9279 8998 9288
rect 8956 9178 8984 9279
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8942 8664 8998 8673
rect 8942 8599 8998 8608
rect 8850 8120 8906 8129
rect 8680 8078 8800 8106
rect 8772 8022 8800 8078
rect 8956 8090 8984 8599
rect 8850 8055 8906 8064
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8760 8016 8812 8022
rect 8220 7942 8340 7970
rect 8760 7958 8812 7964
rect 8312 7188 8340 7942
rect 8576 7744 8628 7750
rect 8576 7686 8628 7692
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8588 7546 8616 7686
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8576 7404 8628 7410
rect 8680 7392 8708 7686
rect 8628 7364 8708 7392
rect 8576 7346 8628 7352
rect 8404 7290 8432 7346
rect 8942 7304 8998 7313
rect 8404 7262 8892 7290
rect 8220 7160 8340 7188
rect 8220 6882 8248 7160
rect 8353 7100 8649 7120
rect 8409 7098 8433 7100
rect 8489 7098 8513 7100
rect 8569 7098 8593 7100
rect 8431 7046 8433 7098
rect 8495 7046 8507 7098
rect 8569 7046 8571 7098
rect 8409 7044 8433 7046
rect 8489 7044 8513 7046
rect 8569 7044 8593 7046
rect 8353 7024 8649 7044
rect 8758 7032 8814 7041
rect 8680 7002 8758 7018
rect 8668 6996 8758 7002
rect 8720 6990 8758 6996
rect 8758 6967 8814 6976
rect 8668 6938 8720 6944
rect 8220 6854 8340 6882
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 7932 6384 7984 6390
rect 7932 6326 7984 6332
rect 7930 6216 7986 6225
rect 7930 6151 7986 6160
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7760 5234 7788 5646
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 7944 5098 7972 6151
rect 7932 5092 7984 5098
rect 7932 5034 7984 5040
rect 8220 4214 8248 6734
rect 8312 6322 8340 6854
rect 8574 6760 8630 6769
rect 8574 6695 8576 6704
rect 8628 6695 8630 6704
rect 8576 6666 8628 6672
rect 8390 6488 8446 6497
rect 8390 6423 8446 6432
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8404 6254 8432 6423
rect 8668 6384 8720 6390
rect 8666 6352 8668 6361
rect 8720 6352 8722 6361
rect 8666 6287 8722 6296
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8353 6012 8649 6032
rect 8409 6010 8433 6012
rect 8489 6010 8513 6012
rect 8569 6010 8593 6012
rect 8431 5958 8433 6010
rect 8495 5958 8507 6010
rect 8569 5958 8571 6010
rect 8409 5956 8433 5958
rect 8489 5956 8513 5958
rect 8569 5956 8593 5958
rect 8353 5936 8649 5956
rect 8864 5710 8892 7262
rect 8942 7239 8998 7248
rect 8956 7002 8984 7239
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 9048 6780 9076 11494
rect 9140 9450 9168 12378
rect 9232 12306 9260 13738
rect 9324 13530 9352 15302
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 9312 13388 9364 13394
rect 9312 13330 9364 13336
rect 9324 12442 9352 13330
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9416 12050 9444 15388
rect 9600 15348 9628 18255
rect 9876 18222 9904 18906
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9678 17232 9734 17241
rect 9678 17167 9734 17176
rect 9692 16046 9720 17167
rect 9954 16824 10010 16833
rect 9954 16759 10010 16768
rect 9968 16726 9996 16759
rect 9956 16720 10008 16726
rect 9956 16662 10008 16668
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9508 15320 9628 15348
rect 9508 13818 9536 15320
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9588 14884 9640 14890
rect 9588 14826 9640 14832
rect 9600 14414 9628 14826
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9692 14074 9720 14894
rect 9784 14346 9812 15438
rect 9968 15026 9996 16390
rect 10060 15314 10088 18566
rect 10140 18352 10192 18358
rect 10140 18294 10192 18300
rect 10152 16776 10180 18294
rect 10244 17610 10272 19178
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10336 17678 10364 18158
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10232 17604 10284 17610
rect 10232 17546 10284 17552
rect 10336 17134 10364 17614
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10232 16788 10284 16794
rect 10152 16748 10232 16776
rect 10232 16730 10284 16736
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 10244 16561 10272 16594
rect 10230 16552 10286 16561
rect 10230 16487 10286 16496
rect 10336 16454 10364 17070
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10416 16244 10468 16250
rect 10416 16186 10468 16192
rect 10428 15502 10456 16186
rect 10520 15638 10548 23920
rect 10692 19916 10744 19922
rect 10692 19858 10744 19864
rect 10704 19174 10732 19858
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10704 18970 10732 19110
rect 10692 18964 10744 18970
rect 10692 18906 10744 18912
rect 10796 18834 10824 19110
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 10782 18592 10838 18601
rect 10782 18527 10838 18536
rect 10796 18222 10824 18527
rect 10784 18216 10836 18222
rect 10784 18158 10836 18164
rect 11060 17060 11112 17066
rect 11060 17002 11112 17008
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10704 15910 10732 16186
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10704 15638 10732 15846
rect 10796 15706 10824 15982
rect 10888 15706 10916 16050
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10508 15632 10560 15638
rect 10508 15574 10560 15580
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10980 15570 11008 16730
rect 11072 16522 11100 17002
rect 11060 16516 11112 16522
rect 11060 16458 11112 16464
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10060 15286 10180 15314
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 9968 14890 9996 14962
rect 9956 14884 10008 14890
rect 9956 14826 10008 14832
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 9864 14544 9916 14550
rect 9864 14486 9916 14492
rect 9772 14340 9824 14346
rect 9772 14282 9824 14288
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 9508 13790 9628 13818
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9232 12022 9444 12050
rect 9232 9897 9260 12022
rect 9508 10810 9536 13670
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9218 9888 9274 9897
rect 9218 9823 9274 9832
rect 9218 9752 9274 9761
rect 9218 9687 9274 9696
rect 9128 9444 9180 9450
rect 9128 9386 9180 9392
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 9140 8362 9168 9046
rect 9232 8974 9260 9687
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9232 8566 9260 8910
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 9128 8356 9180 8362
rect 9128 8298 9180 8304
rect 9126 8120 9182 8129
rect 9126 8055 9182 8064
rect 9140 7818 9168 8055
rect 9220 8016 9272 8022
rect 9220 7958 9272 7964
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 8956 6752 9076 6780
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8956 5370 8984 6752
rect 9034 6624 9090 6633
rect 9034 6559 9090 6568
rect 9048 5778 9076 6559
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 9140 5370 9168 7142
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 8353 4924 8649 4944
rect 8409 4922 8433 4924
rect 8489 4922 8513 4924
rect 8569 4922 8593 4924
rect 8431 4870 8433 4922
rect 8495 4870 8507 4922
rect 8569 4870 8571 4922
rect 8409 4868 8433 4870
rect 8489 4868 8513 4870
rect 8569 4868 8593 4870
rect 8353 4848 8649 4868
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 9232 4146 9260 7958
rect 9324 6186 9352 10202
rect 9416 8634 9444 10406
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9508 9178 9536 9862
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9494 9072 9550 9081
rect 9494 9007 9550 9016
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9508 8514 9536 9007
rect 9416 8486 9536 8514
rect 9416 6254 9444 8486
rect 9600 8412 9628 13790
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9692 12753 9720 12786
rect 9678 12744 9734 12753
rect 9678 12679 9734 12688
rect 9784 12306 9812 13874
rect 9876 12442 9904 14486
rect 9968 13002 9996 14554
rect 10060 14550 10088 15098
rect 10048 14544 10100 14550
rect 10048 14486 10100 14492
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10060 13802 10088 14214
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 10060 13190 10088 13738
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 9968 12974 10088 13002
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9680 12096 9732 12102
rect 9678 12064 9680 12073
rect 9732 12064 9734 12073
rect 9678 11999 9734 12008
rect 9968 11914 9996 12582
rect 9692 11886 9996 11914
rect 9692 11218 9720 11886
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 9954 11792 10010 11801
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9692 10538 9720 10678
rect 9784 10606 9812 11766
rect 9864 11756 9916 11762
rect 9954 11727 10010 11736
rect 9864 11698 9916 11704
rect 9876 11665 9904 11698
rect 9862 11656 9918 11665
rect 9862 11591 9918 11600
rect 9876 10962 9904 11591
rect 9968 11082 9996 11727
rect 10060 11218 10088 12974
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 10048 11008 10100 11014
rect 9876 10934 9996 10962
rect 10048 10950 10100 10956
rect 9864 10736 9916 10742
rect 9864 10678 9916 10684
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9876 10418 9904 10678
rect 9692 10390 9904 10418
rect 9692 10062 9720 10390
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9692 8634 9720 8774
rect 9784 8634 9812 9318
rect 9876 8906 9904 10134
rect 9968 9722 9996 10934
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9784 8498 9812 8570
rect 9862 8528 9918 8537
rect 9772 8492 9824 8498
rect 9508 8384 9628 8412
rect 9692 8452 9772 8480
rect 9508 6769 9536 8384
rect 9692 7954 9720 8452
rect 9862 8463 9918 8472
rect 9772 8434 9824 8440
rect 9876 8378 9904 8463
rect 9784 8350 9904 8378
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9600 7002 9628 7822
rect 9692 7818 9720 7890
rect 9680 7812 9732 7818
rect 9680 7754 9732 7760
rect 9692 7410 9720 7754
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9586 6896 9642 6905
rect 9586 6831 9642 6840
rect 9494 6760 9550 6769
rect 9494 6695 9550 6704
rect 9494 6624 9550 6633
rect 9494 6559 9550 6568
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 9310 5944 9366 5953
rect 9508 5930 9536 6559
rect 9416 5914 9536 5930
rect 9310 5879 9366 5888
rect 9404 5908 9536 5914
rect 9324 5846 9352 5879
rect 9456 5902 9536 5908
rect 9404 5850 9456 5856
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9404 5704 9456 5710
rect 9402 5672 9404 5681
rect 9456 5672 9458 5681
rect 9600 5642 9628 6831
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9692 5953 9720 6258
rect 9678 5944 9734 5953
rect 9678 5879 9734 5888
rect 9402 5607 9458 5616
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 9784 5234 9812 8350
rect 9864 7948 9916 7954
rect 9864 7890 9916 7896
rect 9876 7478 9904 7890
rect 10060 7868 10088 10950
rect 10152 9217 10180 15286
rect 10244 14958 10272 15438
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10232 14952 10284 14958
rect 10232 14894 10284 14900
rect 10508 14544 10560 14550
rect 10230 14512 10286 14521
rect 10508 14486 10560 14492
rect 10230 14447 10286 14456
rect 10416 14476 10468 14482
rect 10244 11014 10272 14447
rect 10416 14418 10468 14424
rect 10322 13288 10378 13297
rect 10322 13223 10378 13232
rect 10336 12986 10364 13223
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10336 11762 10364 12582
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10336 11218 10364 11698
rect 10428 11354 10456 14418
rect 10520 14074 10548 14486
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10612 13326 10640 15302
rect 10796 14958 10824 15302
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10692 14000 10744 14006
rect 10692 13942 10744 13948
rect 10704 13326 10732 13942
rect 10796 13841 10824 14894
rect 10782 13832 10838 13841
rect 10782 13767 10838 13776
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10508 13252 10560 13258
rect 10508 13194 10560 13200
rect 10520 12714 10548 13194
rect 10508 12708 10560 12714
rect 10508 12650 10560 12656
rect 10612 12594 10640 13262
rect 10704 12646 10732 13262
rect 10520 12566 10640 12594
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10520 11665 10548 12566
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10598 11792 10654 11801
rect 10598 11727 10654 11736
rect 10506 11656 10562 11665
rect 10506 11591 10562 11600
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10336 10810 10364 11154
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10232 10532 10284 10538
rect 10232 10474 10284 10480
rect 10244 10266 10272 10474
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10244 9654 10272 10066
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10138 9208 10194 9217
rect 10138 9143 10194 9152
rect 10244 9081 10272 9590
rect 10230 9072 10286 9081
rect 10230 9007 10286 9016
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 9968 7840 10088 7868
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9876 5370 9904 7278
rect 9968 6662 9996 7840
rect 10152 7478 10180 8910
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10046 6896 10102 6905
rect 10046 6831 10102 6840
rect 10060 6730 10088 6831
rect 10244 6798 10272 7346
rect 10140 6792 10192 6798
rect 10138 6760 10140 6769
rect 10232 6792 10284 6798
rect 10192 6760 10194 6769
rect 10048 6724 10100 6730
rect 10232 6734 10284 6740
rect 10138 6695 10194 6704
rect 10048 6666 10100 6672
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 10336 6474 10364 9658
rect 10520 9450 10548 10406
rect 10508 9444 10560 9450
rect 10508 9386 10560 9392
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10428 9178 10456 9318
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10414 9072 10470 9081
rect 10414 9007 10470 9016
rect 10428 6934 10456 9007
rect 10416 6928 10468 6934
rect 10416 6870 10468 6876
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10152 6446 10364 6474
rect 10152 6390 10180 6446
rect 10140 6384 10192 6390
rect 10140 6326 10192 6332
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10336 6225 10364 6258
rect 10428 6254 10456 6734
rect 10520 6497 10548 9386
rect 10612 6905 10640 11727
rect 10704 11529 10732 11834
rect 10690 11520 10746 11529
rect 10690 11455 10746 11464
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10704 9761 10732 10746
rect 10690 9752 10746 9761
rect 10690 9687 10746 9696
rect 10796 9330 10824 13466
rect 10888 12866 10916 15302
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 10980 12968 11008 14350
rect 11060 13796 11112 13802
rect 11060 13738 11112 13744
rect 11072 13138 11100 13738
rect 11164 13682 11192 23920
rect 11808 23066 11836 23920
rect 12452 23882 12480 23920
rect 12452 23854 12572 23882
rect 11808 23038 11928 23066
rect 11796 21412 11848 21418
rect 11796 21354 11848 21360
rect 11520 21140 11572 21146
rect 11520 21082 11572 21088
rect 11348 20466 11468 20482
rect 11348 20460 11480 20466
rect 11348 20454 11428 20460
rect 11348 20330 11376 20454
rect 11428 20402 11480 20408
rect 11336 20324 11388 20330
rect 11336 20266 11388 20272
rect 11428 20324 11480 20330
rect 11428 20266 11480 20272
rect 11242 16688 11298 16697
rect 11242 16623 11298 16632
rect 11336 16652 11388 16658
rect 11256 16046 11284 16623
rect 11336 16594 11388 16600
rect 11348 16561 11376 16594
rect 11334 16552 11390 16561
rect 11334 16487 11390 16496
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11256 14822 11284 15846
rect 11440 14822 11468 20266
rect 11532 17626 11560 21082
rect 11808 20602 11836 21354
rect 11796 20596 11848 20602
rect 11796 20538 11848 20544
rect 11900 19718 11928 23038
rect 12052 21788 12348 21808
rect 12108 21786 12132 21788
rect 12188 21786 12212 21788
rect 12268 21786 12292 21788
rect 12130 21734 12132 21786
rect 12194 21734 12206 21786
rect 12268 21734 12270 21786
rect 12108 21732 12132 21734
rect 12188 21732 12212 21734
rect 12268 21732 12292 21734
rect 12052 21712 12348 21732
rect 12164 21480 12216 21486
rect 12164 21422 12216 21428
rect 12072 21344 12124 21350
rect 12072 21286 12124 21292
rect 12084 21078 12112 21286
rect 12072 21072 12124 21078
rect 12072 21014 12124 21020
rect 12176 20788 12204 21422
rect 11992 20760 12204 20788
rect 12440 20800 12492 20806
rect 11992 20398 12020 20760
rect 12440 20742 12492 20748
rect 12052 20700 12348 20720
rect 12108 20698 12132 20700
rect 12188 20698 12212 20700
rect 12268 20698 12292 20700
rect 12130 20646 12132 20698
rect 12194 20646 12206 20698
rect 12268 20646 12270 20698
rect 12108 20644 12132 20646
rect 12188 20644 12212 20646
rect 12268 20644 12292 20646
rect 12052 20624 12348 20644
rect 11980 20392 12032 20398
rect 11980 20334 12032 20340
rect 11992 20058 12020 20334
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 12176 19990 12204 20198
rect 12164 19984 12216 19990
rect 12164 19926 12216 19932
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11888 19712 11940 19718
rect 11888 19654 11940 19660
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11612 18828 11664 18834
rect 11612 18770 11664 18776
rect 11624 18426 11652 18770
rect 11612 18420 11664 18426
rect 11612 18362 11664 18368
rect 11716 18154 11744 19110
rect 11704 18148 11756 18154
rect 11704 18090 11756 18096
rect 11532 17598 11652 17626
rect 11716 17610 11744 18090
rect 11808 17814 11836 19110
rect 11992 18834 12020 19858
rect 12268 19802 12296 20198
rect 12452 19938 12480 20742
rect 12544 20330 12572 23854
rect 12900 21344 12952 21350
rect 12900 21286 12952 21292
rect 12532 20324 12584 20330
rect 12532 20266 12584 20272
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12808 20256 12860 20262
rect 12808 20198 12860 20204
rect 12360 19922 12480 19938
rect 12348 19916 12480 19922
rect 12400 19910 12480 19916
rect 12348 19858 12400 19864
rect 12084 19786 12296 19802
rect 12072 19780 12296 19786
rect 12124 19774 12296 19780
rect 12072 19722 12124 19728
rect 12728 19718 12756 20198
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12052 19612 12348 19632
rect 12108 19610 12132 19612
rect 12188 19610 12212 19612
rect 12268 19610 12292 19612
rect 12130 19558 12132 19610
rect 12194 19558 12206 19610
rect 12268 19558 12270 19610
rect 12108 19556 12132 19558
rect 12188 19556 12212 19558
rect 12268 19556 12292 19558
rect 12052 19536 12348 19556
rect 12348 19168 12400 19174
rect 12346 19136 12348 19145
rect 12400 19136 12402 19145
rect 12346 19071 12402 19080
rect 11980 18828 12032 18834
rect 11980 18770 12032 18776
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 12176 18612 12204 18770
rect 11992 18584 12204 18612
rect 11796 17808 11848 17814
rect 11796 17750 11848 17756
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11532 16998 11560 17478
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 11624 16810 11652 17598
rect 11704 17604 11756 17610
rect 11704 17546 11756 17552
rect 11992 17338 12020 18584
rect 12052 18524 12348 18544
rect 12108 18522 12132 18524
rect 12188 18522 12212 18524
rect 12268 18522 12292 18524
rect 12130 18470 12132 18522
rect 12194 18470 12206 18522
rect 12268 18470 12270 18522
rect 12108 18468 12132 18470
rect 12188 18468 12212 18470
rect 12268 18468 12292 18470
rect 12052 18448 12348 18468
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 12084 17814 12112 18226
rect 12452 18222 12480 19654
rect 12530 19544 12586 19553
rect 12530 19479 12532 19488
rect 12584 19479 12586 19488
rect 12532 19450 12584 19456
rect 12544 19332 12756 19360
rect 12544 18970 12572 19332
rect 12622 19272 12678 19281
rect 12622 19207 12678 19216
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12636 18834 12664 19207
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12348 18148 12400 18154
rect 12348 18090 12400 18096
rect 12072 17808 12124 17814
rect 12072 17750 12124 17756
rect 12360 17746 12388 18090
rect 12532 18080 12584 18086
rect 12532 18022 12584 18028
rect 12440 17808 12492 17814
rect 12440 17750 12492 17756
rect 12348 17740 12400 17746
rect 12348 17682 12400 17688
rect 12452 17649 12480 17750
rect 12438 17640 12494 17649
rect 12438 17575 12494 17584
rect 12052 17436 12348 17456
rect 12108 17434 12132 17436
rect 12188 17434 12212 17436
rect 12268 17434 12292 17436
rect 12130 17382 12132 17434
rect 12194 17382 12206 17434
rect 12268 17382 12270 17434
rect 12108 17380 12132 17382
rect 12188 17380 12212 17382
rect 12268 17380 12292 17382
rect 12052 17360 12348 17380
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 12256 17264 12308 17270
rect 12256 17206 12308 17212
rect 12268 17105 12296 17206
rect 12254 17096 12310 17105
rect 12254 17031 12310 17040
rect 11532 16782 11652 16810
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11256 14346 11284 14758
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 11348 13870 11376 14554
rect 11428 14340 11480 14346
rect 11428 14282 11480 14288
rect 11440 13938 11468 14282
rect 11428 13932 11480 13938
rect 11428 13874 11480 13880
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11164 13654 11468 13682
rect 11072 13110 11284 13138
rect 10980 12940 11100 12968
rect 10888 12838 11008 12866
rect 10980 12306 11008 12838
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10874 12200 10930 12209
rect 10874 12135 10930 12144
rect 10704 9302 10824 9330
rect 10704 7041 10732 9302
rect 10888 9160 10916 12135
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10796 9132 10916 9160
rect 10690 7032 10746 7041
rect 10690 6967 10746 6976
rect 10598 6896 10654 6905
rect 10598 6831 10654 6840
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10704 6662 10732 6802
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10506 6488 10562 6497
rect 10506 6423 10562 6432
rect 10416 6248 10468 6254
rect 10322 6216 10378 6225
rect 10416 6190 10468 6196
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10322 6151 10378 6160
rect 10336 5574 10364 6151
rect 10704 5778 10732 6190
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 9862 5264 9918 5273
rect 9772 5228 9824 5234
rect 10704 5234 10732 5306
rect 9862 5199 9918 5208
rect 10692 5228 10744 5234
rect 9772 5170 9824 5176
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9600 4282 9628 4966
rect 9876 4826 9904 5199
rect 10692 5170 10744 5176
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 10324 4752 10376 4758
rect 10322 4720 10324 4729
rect 10376 4720 10378 4729
rect 10322 4655 10378 4664
rect 10704 4622 10732 5170
rect 10796 4826 10824 9132
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10888 8498 10916 8978
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 10888 8362 10916 8434
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 10876 7812 10928 7818
rect 10876 7754 10928 7760
rect 10888 7342 10916 7754
rect 10980 7585 11008 11630
rect 11072 11286 11100 12940
rect 11150 12880 11206 12889
rect 11150 12815 11206 12824
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 11164 11132 11192 12815
rect 11072 11104 11192 11132
rect 11072 8786 11100 11104
rect 11152 10600 11204 10606
rect 11256 10588 11284 13110
rect 11336 12912 11388 12918
rect 11336 12854 11388 12860
rect 11204 10560 11284 10588
rect 11152 10542 11204 10548
rect 11164 8906 11192 10542
rect 11348 9382 11376 12854
rect 11440 12442 11468 13654
rect 11532 12714 11560 16782
rect 11888 16720 11940 16726
rect 11888 16662 11940 16668
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11624 15162 11652 16050
rect 11796 16040 11848 16046
rect 11796 15982 11848 15988
rect 11808 15570 11836 15982
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11900 15162 11928 16662
rect 12052 16348 12348 16368
rect 12108 16346 12132 16348
rect 12188 16346 12212 16348
rect 12268 16346 12292 16348
rect 12130 16294 12132 16346
rect 12194 16294 12206 16346
rect 12268 16294 12270 16346
rect 12108 16292 12132 16294
rect 12188 16292 12212 16294
rect 12268 16292 12292 16294
rect 12052 16272 12348 16292
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11992 16130 12020 16186
rect 11992 16102 12112 16130
rect 11980 16040 12032 16046
rect 11980 15982 12032 15988
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11704 15088 11756 15094
rect 11704 15030 11756 15036
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11624 14074 11652 14758
rect 11716 14550 11744 15030
rect 11796 14952 11848 14958
rect 11796 14894 11848 14900
rect 11704 14544 11756 14550
rect 11704 14486 11756 14492
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11520 12708 11572 12714
rect 11520 12650 11572 12656
rect 11518 12608 11574 12617
rect 11518 12543 11574 12552
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11428 11552 11480 11558
rect 11428 11494 11480 11500
rect 11440 11218 11468 11494
rect 11532 11218 11560 12543
rect 11624 11830 11652 13874
rect 11808 13462 11836 14894
rect 11900 14278 11928 15098
rect 11992 14618 12020 15982
rect 12084 15910 12112 16102
rect 12072 15904 12124 15910
rect 12072 15846 12124 15852
rect 12348 15904 12400 15910
rect 12400 15864 12480 15892
rect 12348 15846 12400 15852
rect 12452 15502 12480 15864
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 12052 15260 12348 15280
rect 12108 15258 12132 15260
rect 12188 15258 12212 15260
rect 12268 15258 12292 15260
rect 12130 15206 12132 15258
rect 12194 15206 12206 15258
rect 12268 15206 12270 15258
rect 12108 15204 12132 15206
rect 12188 15204 12212 15206
rect 12268 15204 12292 15206
rect 12052 15184 12348 15204
rect 12070 15056 12126 15065
rect 12070 14991 12072 15000
rect 12124 14991 12126 15000
rect 12072 14962 12124 14968
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 12544 14550 12572 18022
rect 12728 17882 12756 19332
rect 12820 18222 12848 20198
rect 12912 19242 12940 21286
rect 13096 20534 13124 23920
rect 13740 23882 13768 23920
rect 13464 23854 13768 23882
rect 13176 21004 13228 21010
rect 13176 20946 13228 20952
rect 13084 20528 13136 20534
rect 13084 20470 13136 20476
rect 13188 20398 13216 20946
rect 13176 20392 13228 20398
rect 13176 20334 13228 20340
rect 13188 20262 13216 20334
rect 13360 20324 13412 20330
rect 13360 20266 13412 20272
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 13082 19408 13138 19417
rect 13082 19343 13084 19352
rect 13136 19343 13138 19352
rect 13084 19314 13136 19320
rect 12900 19236 12952 19242
rect 12900 19178 12952 19184
rect 13268 18828 13320 18834
rect 13268 18770 13320 18776
rect 13280 18630 13308 18770
rect 13084 18624 13136 18630
rect 13268 18624 13320 18630
rect 13136 18572 13216 18578
rect 13084 18566 13216 18572
rect 13268 18566 13320 18572
rect 13096 18550 13216 18566
rect 12808 18216 12860 18222
rect 12808 18158 12860 18164
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 12820 17746 12848 18158
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 12820 17490 12848 17682
rect 12900 17604 12952 17610
rect 12900 17546 12952 17552
rect 12636 17462 12848 17490
rect 12636 17202 12664 17462
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 12912 16590 12940 17546
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 13096 16794 13124 16934
rect 13188 16794 13216 18550
rect 13280 17134 13308 18566
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 13176 16788 13228 16794
rect 13176 16730 13228 16736
rect 12900 16584 12952 16590
rect 12900 16526 12952 16532
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 12622 16144 12678 16153
rect 12622 16079 12678 16088
rect 12990 16144 13046 16153
rect 12990 16079 13046 16088
rect 13084 16108 13136 16114
rect 12636 15910 12664 16079
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12714 15736 12770 15745
rect 12714 15671 12716 15680
rect 12768 15671 12770 15680
rect 12716 15642 12768 15648
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12636 14618 12664 15302
rect 12716 15088 12768 15094
rect 12716 15030 12768 15036
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12532 14544 12584 14550
rect 12532 14486 12584 14492
rect 12440 14408 12492 14414
rect 12636 14385 12664 14554
rect 12440 14350 12492 14356
rect 12622 14376 12678 14385
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 12052 14172 12348 14192
rect 12108 14170 12132 14172
rect 12188 14170 12212 14172
rect 12268 14170 12292 14172
rect 12130 14118 12132 14170
rect 12194 14118 12206 14170
rect 12268 14118 12270 14170
rect 12108 14116 12132 14118
rect 12188 14116 12212 14118
rect 12268 14116 12292 14118
rect 12052 14096 12348 14116
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11796 13456 11848 13462
rect 11796 13398 11848 13404
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11716 12986 11744 13330
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11900 12782 11928 14010
rect 12452 13870 12480 14350
rect 12622 14311 12678 14320
rect 12440 13864 12492 13870
rect 12162 13832 12218 13841
rect 12440 13806 12492 13812
rect 12162 13767 12218 13776
rect 12176 13394 12204 13767
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 11980 13252 12032 13258
rect 11980 13194 12032 13200
rect 11992 12782 12020 13194
rect 12052 13084 12348 13104
rect 12108 13082 12132 13084
rect 12188 13082 12212 13084
rect 12268 13082 12292 13084
rect 12130 13030 12132 13082
rect 12194 13030 12206 13082
rect 12268 13030 12270 13082
rect 12108 13028 12132 13030
rect 12188 13028 12212 13030
rect 12268 13028 12292 13030
rect 12052 13008 12348 13028
rect 12728 12889 12756 15030
rect 12820 14890 12848 15846
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12808 14884 12860 14890
rect 12808 14826 12860 14832
rect 12808 14544 12860 14550
rect 12808 14486 12860 14492
rect 12714 12880 12770 12889
rect 12714 12815 12770 12824
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12714 12744 12770 12753
rect 11716 11898 11744 12718
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11612 11824 11664 11830
rect 11612 11766 11664 11772
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11428 11212 11480 11218
rect 11428 11154 11480 11160
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11440 9654 11468 11154
rect 11518 11112 11574 11121
rect 11518 11047 11574 11056
rect 11428 9648 11480 9654
rect 11428 9590 11480 9596
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11256 9132 11468 9160
rect 11152 8900 11204 8906
rect 11152 8842 11204 8848
rect 11072 8758 11192 8786
rect 10966 7576 11022 7585
rect 10966 7511 11022 7520
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 11164 6202 11192 8758
rect 11256 8566 11284 9132
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11244 8560 11296 8566
rect 11244 8502 11296 8508
rect 11256 8022 11284 8502
rect 11244 8016 11296 8022
rect 11244 7958 11296 7964
rect 11348 7818 11376 8978
rect 11440 8974 11468 9132
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 11426 8664 11482 8673
rect 11426 8599 11482 8608
rect 11440 8566 11468 8599
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 11440 7478 11468 7822
rect 11428 7472 11480 7478
rect 11428 7414 11480 7420
rect 11532 7290 11560 11047
rect 11624 9353 11652 11494
rect 11808 11354 11836 11562
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 11716 10985 11744 11222
rect 11702 10976 11758 10985
rect 11702 10911 11758 10920
rect 11794 10840 11850 10849
rect 11794 10775 11796 10784
rect 11848 10775 11850 10784
rect 11796 10746 11848 10752
rect 11704 10192 11756 10198
rect 11704 10134 11756 10140
rect 11610 9344 11666 9353
rect 11610 9279 11666 9288
rect 11612 8832 11664 8838
rect 11612 8774 11664 8780
rect 11624 8430 11652 8774
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11624 8090 11652 8230
rect 11716 8090 11744 10134
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 11808 9722 11836 10066
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 11794 8392 11850 8401
rect 11794 8327 11850 8336
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11610 7984 11666 7993
rect 11610 7919 11666 7928
rect 11624 7721 11652 7919
rect 11808 7750 11836 8327
rect 11796 7744 11848 7750
rect 11610 7712 11666 7721
rect 11796 7686 11848 7692
rect 11610 7647 11666 7656
rect 11532 7262 11744 7290
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11624 6662 11652 7142
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11072 6174 11192 6202
rect 11336 6248 11388 6254
rect 11336 6190 11388 6196
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 9588 4276 9640 4282
rect 9588 4218 9640 4224
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 8353 3836 8649 3856
rect 8409 3834 8433 3836
rect 8489 3834 8513 3836
rect 8569 3834 8593 3836
rect 8431 3782 8433 3834
rect 8495 3782 8507 3834
rect 8569 3782 8571 3834
rect 8409 3780 8433 3782
rect 8489 3780 8513 3782
rect 8569 3780 8593 3782
rect 8353 3760 8649 3780
rect 10704 3534 10732 4558
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 4654 3292 4950 3312
rect 4710 3290 4734 3292
rect 4790 3290 4814 3292
rect 4870 3290 4894 3292
rect 4732 3238 4734 3290
rect 4796 3238 4808 3290
rect 4870 3238 4872 3290
rect 4710 3236 4734 3238
rect 4790 3236 4814 3238
rect 4870 3236 4894 3238
rect 4654 3216 4950 3236
rect 2964 3120 3016 3126
rect 1950 3088 2006 3097
rect 2964 3062 3016 3068
rect 11072 3058 11100 6174
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11164 5370 11192 6054
rect 11348 5370 11376 6190
rect 11520 6180 11572 6186
rect 11520 6122 11572 6128
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11532 5166 11560 6122
rect 11624 5234 11652 6598
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11520 5160 11572 5166
rect 11716 5137 11744 7262
rect 11794 7032 11850 7041
rect 11794 6967 11796 6976
rect 11848 6967 11850 6976
rect 11796 6938 11848 6944
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11808 6186 11836 6598
rect 11796 6180 11848 6186
rect 11796 6122 11848 6128
rect 11520 5102 11572 5108
rect 11702 5128 11758 5137
rect 11702 5063 11758 5072
rect 11702 4856 11758 4865
rect 11900 4826 11928 12582
rect 11992 11694 12020 12582
rect 12052 11996 12348 12016
rect 12108 11994 12132 11996
rect 12188 11994 12212 11996
rect 12268 11994 12292 11996
rect 12130 11942 12132 11994
rect 12194 11942 12206 11994
rect 12268 11942 12270 11994
rect 12108 11940 12132 11942
rect 12188 11940 12212 11942
rect 12268 11940 12292 11942
rect 12052 11920 12348 11940
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 12452 11218 12480 12718
rect 12820 12730 12848 14486
rect 12770 12702 12848 12730
rect 12714 12679 12770 12688
rect 12728 12458 12756 12679
rect 12912 12617 12940 15506
rect 13004 15094 13032 16079
rect 13084 16050 13136 16056
rect 13096 15706 13124 16050
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 13280 15570 13308 16186
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 12992 15088 13044 15094
rect 12992 15030 13044 15036
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 12898 12608 12954 12617
rect 12898 12543 12954 12552
rect 12636 12430 12756 12458
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12544 11937 12572 12038
rect 12530 11928 12586 11937
rect 12636 11898 12664 12430
rect 12714 12200 12770 12209
rect 12714 12135 12770 12144
rect 12530 11863 12586 11872
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12052 10908 12348 10928
rect 12108 10906 12132 10908
rect 12188 10906 12212 10908
rect 12268 10906 12292 10908
rect 12130 10854 12132 10906
rect 12194 10854 12206 10906
rect 12268 10854 12270 10906
rect 12108 10852 12132 10854
rect 12188 10852 12212 10854
rect 12268 10852 12292 10854
rect 12052 10832 12348 10852
rect 12452 10742 12480 11154
rect 12440 10736 12492 10742
rect 12360 10696 12440 10724
rect 11978 10296 12034 10305
rect 11978 10231 12034 10240
rect 11992 4826 12020 10231
rect 12360 10198 12388 10696
rect 12440 10678 12492 10684
rect 12440 10600 12492 10606
rect 12544 10577 12572 11766
rect 12624 10600 12676 10606
rect 12440 10542 12492 10548
rect 12530 10568 12586 10577
rect 12348 10192 12400 10198
rect 12348 10134 12400 10140
rect 12452 10146 12480 10542
rect 12624 10542 12676 10548
rect 12530 10503 12586 10512
rect 12452 10118 12572 10146
rect 12440 10056 12492 10062
rect 12544 10033 12572 10118
rect 12440 9998 12492 10004
rect 12530 10024 12586 10033
rect 12052 9820 12348 9840
rect 12108 9818 12132 9820
rect 12188 9818 12212 9820
rect 12268 9818 12292 9820
rect 12130 9766 12132 9818
rect 12194 9766 12206 9818
rect 12268 9766 12270 9818
rect 12108 9764 12132 9766
rect 12188 9764 12212 9766
rect 12268 9764 12292 9766
rect 12052 9744 12348 9764
rect 12452 9602 12480 9998
rect 12530 9959 12586 9968
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12360 9574 12480 9602
rect 12360 8974 12388 9574
rect 12544 9518 12572 9658
rect 12636 9586 12664 10542
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12452 9330 12480 9454
rect 12452 9302 12572 9330
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12052 8732 12348 8752
rect 12108 8730 12132 8732
rect 12188 8730 12212 8732
rect 12268 8730 12292 8732
rect 12130 8678 12132 8730
rect 12194 8678 12206 8730
rect 12268 8678 12270 8730
rect 12108 8676 12132 8678
rect 12188 8676 12212 8678
rect 12268 8676 12292 8678
rect 12052 8656 12348 8676
rect 12544 8634 12572 9302
rect 12728 8945 12756 12135
rect 13004 12050 13032 14758
rect 13096 14550 13124 15438
rect 13268 14884 13320 14890
rect 13268 14826 13320 14832
rect 13280 14793 13308 14826
rect 13266 14784 13322 14793
rect 13266 14719 13322 14728
rect 13084 14544 13136 14550
rect 13084 14486 13136 14492
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 13096 12345 13124 13806
rect 13372 12866 13400 20266
rect 13464 17105 13492 23854
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13740 21078 13768 21286
rect 13728 21072 13780 21078
rect 13728 21014 13780 21020
rect 13740 20058 13768 21014
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 13832 20058 13860 20946
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 14200 19854 14228 21490
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 13544 19712 13596 19718
rect 13544 19654 13596 19660
rect 13556 19310 13584 19654
rect 14200 19514 14228 19790
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 13910 19408 13966 19417
rect 13910 19343 13966 19352
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13636 19304 13688 19310
rect 13924 19292 13952 19343
rect 13636 19246 13688 19252
rect 13832 19264 13952 19292
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13450 17096 13506 17105
rect 13450 17031 13506 17040
rect 13556 16794 13584 18566
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13464 15910 13492 16526
rect 13452 15904 13504 15910
rect 13452 15846 13504 15852
rect 13464 13512 13492 15846
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13556 14958 13584 15302
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13556 13802 13584 14894
rect 13544 13796 13596 13802
rect 13544 13738 13596 13744
rect 13464 13484 13584 13512
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13280 12838 13400 12866
rect 13280 12714 13308 12838
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13268 12708 13320 12714
rect 13268 12650 13320 12656
rect 13082 12336 13138 12345
rect 13082 12271 13138 12280
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 12912 12022 13032 12050
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12714 8936 12770 8945
rect 12714 8871 12770 8880
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12162 8528 12218 8537
rect 12072 8492 12124 8498
rect 12162 8463 12218 8472
rect 12072 8434 12124 8440
rect 12084 8090 12112 8434
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12176 8004 12204 8463
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12348 8016 12400 8022
rect 12176 7976 12348 8004
rect 12348 7958 12400 7964
rect 12052 7644 12348 7664
rect 12108 7642 12132 7644
rect 12188 7642 12212 7644
rect 12268 7642 12292 7644
rect 12130 7590 12132 7642
rect 12194 7590 12206 7642
rect 12268 7590 12270 7642
rect 12108 7588 12132 7590
rect 12188 7588 12212 7590
rect 12268 7588 12292 7590
rect 12052 7568 12348 7588
rect 12348 7268 12400 7274
rect 12348 7210 12400 7216
rect 12360 6905 12388 7210
rect 12346 6896 12402 6905
rect 12346 6831 12402 6840
rect 12052 6556 12348 6576
rect 12108 6554 12132 6556
rect 12188 6554 12212 6556
rect 12268 6554 12292 6556
rect 12130 6502 12132 6554
rect 12194 6502 12206 6554
rect 12268 6502 12270 6554
rect 12108 6500 12132 6502
rect 12188 6500 12212 6502
rect 12268 6500 12292 6502
rect 12052 6480 12348 6500
rect 12452 6458 12480 8366
rect 12728 8362 12756 8774
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12532 7812 12584 7818
rect 12532 7754 12584 7760
rect 12544 7478 12572 7754
rect 12636 7546 12664 7822
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12544 6304 12572 7414
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12636 6497 12664 7142
rect 12622 6488 12678 6497
rect 12622 6423 12678 6432
rect 12624 6316 12676 6322
rect 12268 6276 12624 6304
rect 12268 5710 12296 6276
rect 12624 6258 12676 6264
rect 12440 6112 12492 6118
rect 12728 6066 12756 7686
rect 12440 6054 12492 6060
rect 12348 5772 12400 5778
rect 12452 5760 12480 6054
rect 12400 5732 12480 5760
rect 12348 5714 12400 5720
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12052 5468 12348 5488
rect 12108 5466 12132 5468
rect 12188 5466 12212 5468
rect 12268 5466 12292 5468
rect 12130 5414 12132 5466
rect 12194 5414 12206 5466
rect 12268 5414 12270 5466
rect 12108 5412 12132 5414
rect 12188 5412 12212 5414
rect 12268 5412 12292 5414
rect 12052 5392 12348 5412
rect 12452 5234 12480 5732
rect 12544 6038 12756 6066
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12438 5128 12494 5137
rect 12438 5063 12494 5072
rect 12256 5024 12308 5030
rect 12254 4992 12256 5001
rect 12348 5024 12400 5030
rect 12308 4992 12310 5001
rect 12348 4966 12400 4972
rect 12254 4927 12310 4936
rect 12360 4865 12388 4966
rect 12346 4856 12402 4865
rect 11702 4791 11704 4800
rect 11756 4791 11758 4800
rect 11888 4820 11940 4826
rect 11704 4762 11756 4768
rect 11888 4762 11940 4768
rect 11980 4820 12032 4826
rect 12346 4791 12402 4800
rect 11980 4762 12032 4768
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11900 4570 11928 4626
rect 12452 4622 12480 5063
rect 12440 4616 12492 4622
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11440 3738 11468 3878
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11624 3602 11652 4558
rect 11900 4542 12020 4570
rect 12440 4558 12492 4564
rect 11992 4486 12020 4542
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 12052 4380 12348 4400
rect 12108 4378 12132 4380
rect 12188 4378 12212 4380
rect 12268 4378 12292 4380
rect 12130 4326 12132 4378
rect 12194 4326 12206 4378
rect 12268 4326 12270 4378
rect 12108 4324 12132 4326
rect 12188 4324 12212 4326
rect 12268 4324 12292 4326
rect 12052 4304 12348 4324
rect 11886 4176 11942 4185
rect 11886 4111 11888 4120
rect 11940 4111 11942 4120
rect 11888 4082 11940 4088
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 1950 3023 1952 3032
rect 2004 3023 2006 3032
rect 11060 3052 11112 3058
rect 1952 2994 2004 3000
rect 11060 2994 11112 3000
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1688 480 1716 2790
rect 4654 2204 4950 2224
rect 4710 2202 4734 2204
rect 4790 2202 4814 2204
rect 4870 2202 4894 2204
rect 4732 2150 4734 2202
rect 4796 2150 4808 2202
rect 4870 2150 4872 2202
rect 4710 2148 4734 2150
rect 4790 2148 4814 2150
rect 4870 2148 4894 2150
rect 4654 2128 4950 2148
rect 5092 480 5120 2926
rect 8353 2748 8649 2768
rect 8409 2746 8433 2748
rect 8489 2746 8513 2748
rect 8569 2746 8593 2748
rect 8431 2694 8433 2746
rect 8495 2694 8507 2746
rect 8569 2694 8571 2746
rect 8409 2692 8433 2694
rect 8489 2692 8513 2694
rect 8569 2692 8593 2694
rect 8353 2672 8649 2692
rect 11716 2582 11744 3470
rect 12176 3466 12204 3878
rect 12544 3754 12572 6038
rect 12820 5930 12848 11834
rect 12912 11529 12940 12022
rect 13188 11898 13216 12174
rect 13266 11928 13322 11937
rect 13176 11892 13228 11898
rect 13266 11863 13322 11872
rect 13176 11834 13228 11840
rect 13174 11656 13230 11665
rect 13174 11591 13176 11600
rect 13228 11591 13230 11600
rect 13176 11562 13228 11568
rect 12898 11520 12954 11529
rect 12898 11455 12954 11464
rect 12898 11248 12954 11257
rect 12898 11183 12954 11192
rect 12636 5902 12848 5930
rect 12636 5098 12664 5902
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12820 5030 12848 5782
rect 12912 5778 12940 11183
rect 12992 11008 13044 11014
rect 12990 10976 12992 10985
rect 13044 10976 13046 10985
rect 12990 10911 13046 10920
rect 12990 10840 13046 10849
rect 12990 10775 13046 10784
rect 13004 10169 13032 10775
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 12990 10160 13046 10169
rect 12990 10095 13046 10104
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 13004 9722 13032 9862
rect 12992 9716 13044 9722
rect 12992 9658 13044 9664
rect 13004 9178 13032 9658
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12912 4622 12940 5510
rect 13004 4826 13032 8978
rect 13082 7576 13138 7585
rect 13082 7511 13138 7520
rect 13096 6866 13124 7511
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 13096 5370 13124 6258
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 12990 4312 13046 4321
rect 12990 4247 13046 4256
rect 13004 3942 13032 4247
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12992 3936 13044 3942
rect 13084 3936 13136 3942
rect 12992 3878 13044 3884
rect 13082 3904 13084 3913
rect 13136 3904 13138 3913
rect 12452 3726 12572 3754
rect 12452 3670 12480 3726
rect 12440 3664 12492 3670
rect 12440 3606 12492 3612
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12164 3460 12216 3466
rect 12164 3402 12216 3408
rect 12052 3292 12348 3312
rect 12108 3290 12132 3292
rect 12188 3290 12212 3292
rect 12268 3290 12292 3292
rect 12130 3238 12132 3290
rect 12194 3238 12206 3290
rect 12268 3238 12270 3290
rect 12108 3236 12132 3238
rect 12188 3236 12212 3238
rect 12268 3236 12292 3238
rect 12052 3216 12348 3236
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 11704 2576 11756 2582
rect 8574 2544 8630 2553
rect 11704 2518 11756 2524
rect 8574 2479 8630 2488
rect 8588 480 8616 2479
rect 11992 2088 12020 2994
rect 12544 2553 12572 3538
rect 12636 3369 12664 3878
rect 13082 3839 13138 3848
rect 13188 3738 13216 10202
rect 13280 9518 13308 11863
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 13372 9178 13400 12718
rect 13464 12442 13492 13330
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 13280 8430 13308 9046
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13372 8498 13400 8910
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13358 8392 13414 8401
rect 13358 8327 13414 8336
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13280 7002 13308 7278
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13268 6724 13320 6730
rect 13268 6666 13320 6672
rect 13280 5642 13308 6666
rect 13268 5636 13320 5642
rect 13268 5578 13320 5584
rect 13372 5522 13400 8327
rect 13280 5494 13400 5522
rect 13280 4282 13308 5494
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13372 5166 13400 5306
rect 13464 5302 13492 12378
rect 13452 5296 13504 5302
rect 13452 5238 13504 5244
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 13358 4856 13414 4865
rect 13358 4791 13414 4800
rect 13372 4758 13400 4791
rect 13360 4752 13412 4758
rect 13360 4694 13412 4700
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13556 3738 13584 13484
rect 13648 11257 13676 19246
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13740 14362 13768 17818
rect 13832 17066 13860 19264
rect 14096 18352 14148 18358
rect 14096 18294 14148 18300
rect 13912 18080 13964 18086
rect 13912 18022 13964 18028
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 13832 16590 13860 17002
rect 13924 16726 13952 18022
rect 14004 17672 14056 17678
rect 14004 17614 14056 17620
rect 14016 17338 14044 17614
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 14108 16833 14136 18294
rect 14280 18148 14332 18154
rect 14280 18090 14332 18096
rect 14292 17882 14320 18090
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 14384 17134 14412 23920
rect 14740 21684 14792 21690
rect 14740 21626 14792 21632
rect 14464 21412 14516 21418
rect 14464 21354 14516 21360
rect 14476 20806 14504 21354
rect 14648 21004 14700 21010
rect 14648 20946 14700 20952
rect 14464 20800 14516 20806
rect 14464 20742 14516 20748
rect 14556 20800 14608 20806
rect 14556 20742 14608 20748
rect 14476 20398 14504 20742
rect 14464 20392 14516 20398
rect 14464 20334 14516 20340
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 14094 16824 14150 16833
rect 14094 16759 14150 16768
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 14280 16448 14332 16454
rect 14476 16436 14504 17070
rect 14332 16408 14504 16436
rect 14280 16390 14332 16396
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13832 15337 13860 16050
rect 14004 16040 14056 16046
rect 14004 15982 14056 15988
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13924 15570 13952 15846
rect 14016 15638 14044 15982
rect 14004 15632 14056 15638
rect 14004 15574 14056 15580
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 13818 15328 13874 15337
rect 13818 15263 13874 15272
rect 14108 14618 14136 15982
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14200 14890 14228 15302
rect 14188 14884 14240 14890
rect 14188 14826 14240 14832
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 14292 14396 14320 16390
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 14292 14368 14412 14396
rect 13740 14334 13952 14362
rect 13924 14278 13952 14334
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13740 13462 13768 14214
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13832 13462 13860 13670
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13634 11248 13690 11257
rect 13634 11183 13690 11192
rect 13740 11098 13768 12650
rect 13648 11070 13768 11098
rect 13648 9178 13676 11070
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13740 10849 13768 10950
rect 13726 10840 13782 10849
rect 13726 10775 13782 10784
rect 13832 10441 13860 13398
rect 14188 13388 14240 13394
rect 14188 13330 14240 13336
rect 14004 12912 14056 12918
rect 14004 12854 14056 12860
rect 14016 12753 14044 12854
rect 14002 12744 14058 12753
rect 14002 12679 14058 12688
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13924 11014 13952 12582
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 14108 12345 14136 12378
rect 14094 12336 14150 12345
rect 14004 12300 14056 12306
rect 14094 12271 14150 12280
rect 14004 12242 14056 12248
rect 14016 11898 14044 12242
rect 14200 12102 14228 13330
rect 14384 12889 14412 14368
rect 14370 12880 14426 12889
rect 14370 12815 14426 12824
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 14384 12481 14412 12718
rect 14370 12472 14426 12481
rect 14370 12407 14426 12416
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14094 11928 14150 11937
rect 14004 11892 14056 11898
rect 14094 11863 14150 11872
rect 14188 11892 14240 11898
rect 14004 11834 14056 11840
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13818 10432 13874 10441
rect 13818 10367 13874 10376
rect 13924 10282 13952 10950
rect 13740 10254 13952 10282
rect 14016 10266 14044 11154
rect 14004 10260 14056 10266
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13634 8392 13690 8401
rect 13634 8327 13690 8336
rect 13648 7041 13676 8327
rect 13740 7750 13768 10254
rect 14004 10202 14056 10208
rect 13818 10160 13874 10169
rect 13818 10095 13874 10104
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13832 7154 13860 10095
rect 14108 10010 14136 11863
rect 14188 11834 14240 11840
rect 13924 9982 14136 10010
rect 13924 8090 13952 9982
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14108 9654 14136 9862
rect 14096 9648 14148 9654
rect 14096 9590 14148 9596
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 13832 7126 13952 7154
rect 13634 7032 13690 7041
rect 13634 6967 13690 6976
rect 13636 6928 13688 6934
rect 13688 6888 13768 6916
rect 13636 6870 13688 6876
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13648 5914 13676 6122
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13634 5808 13690 5817
rect 13634 5743 13690 5752
rect 13648 4282 13676 5743
rect 13740 5409 13768 6888
rect 13818 6080 13874 6089
rect 13818 6015 13874 6024
rect 13726 5400 13782 5409
rect 13726 5335 13782 5344
rect 13832 5250 13860 6015
rect 13740 5222 13860 5250
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13740 3738 13768 5222
rect 13818 5128 13874 5137
rect 13818 5063 13874 5072
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13832 3534 13860 5063
rect 13924 5001 13952 7126
rect 14016 5778 14044 8570
rect 14108 8430 14136 9590
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14004 5772 14056 5778
rect 14004 5714 14056 5720
rect 14004 5568 14056 5574
rect 14004 5510 14056 5516
rect 13910 4992 13966 5001
rect 13910 4927 13966 4936
rect 14016 4865 14044 5510
rect 14002 4856 14058 4865
rect 14002 4791 14058 4800
rect 13910 4584 13966 4593
rect 13910 4519 13966 4528
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13268 3392 13320 3398
rect 12622 3360 12678 3369
rect 13268 3334 13320 3340
rect 12622 3295 12678 3304
rect 13280 3194 13308 3334
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13924 2650 13952 4519
rect 14108 4146 14136 6938
rect 14200 5953 14228 11834
rect 14292 11354 14320 12174
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14292 10606 14320 10950
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 14292 10198 14320 10406
rect 14280 10192 14332 10198
rect 14280 10134 14332 10140
rect 14384 7002 14412 11154
rect 14476 11121 14504 15098
rect 14462 11112 14518 11121
rect 14462 11047 14518 11056
rect 14568 10266 14596 20742
rect 14660 20602 14688 20946
rect 14648 20596 14700 20602
rect 14648 20538 14700 20544
rect 14660 19378 14688 20538
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14752 18222 14780 21626
rect 15028 19922 15056 23920
rect 15568 21480 15620 21486
rect 15568 21422 15620 21428
rect 15108 21344 15160 21350
rect 15108 21286 15160 21292
rect 15120 20806 15148 21286
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 15108 20800 15160 20806
rect 15108 20742 15160 20748
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 15212 20398 15240 20742
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 15016 19916 15068 19922
rect 15016 19858 15068 19864
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14844 18426 14872 19790
rect 14924 19780 14976 19786
rect 14924 19722 14976 19728
rect 14936 19378 14964 19722
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 14936 18766 14964 19314
rect 15014 19272 15070 19281
rect 15014 19207 15070 19216
rect 14924 18760 14976 18766
rect 14924 18702 14976 18708
rect 14832 18420 14884 18426
rect 14832 18362 14884 18368
rect 14936 18290 14964 18702
rect 15028 18698 15056 19207
rect 15212 19174 15240 20334
rect 15304 20262 15332 20878
rect 15476 20324 15528 20330
rect 15476 20266 15528 20272
rect 15292 20256 15344 20262
rect 15292 20198 15344 20204
rect 15304 19854 15332 20198
rect 15292 19848 15344 19854
rect 15344 19808 15424 19836
rect 15292 19790 15344 19796
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 15108 18828 15160 18834
rect 15108 18770 15160 18776
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 15120 18737 15148 18770
rect 15106 18728 15162 18737
rect 15016 18692 15068 18698
rect 15106 18663 15162 18672
rect 15016 18634 15068 18640
rect 14924 18284 14976 18290
rect 14924 18226 14976 18232
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 14832 17604 14884 17610
rect 14832 17546 14884 17552
rect 14844 17270 14872 17546
rect 14936 17338 14964 18022
rect 15212 17864 15240 18770
rect 15120 17836 15240 17864
rect 15120 17610 15148 17836
rect 15304 17814 15332 19110
rect 15396 18834 15424 19808
rect 15488 19514 15516 20266
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 15384 18828 15436 18834
rect 15384 18770 15436 18776
rect 15476 18828 15528 18834
rect 15476 18770 15528 18776
rect 15488 18329 15516 18770
rect 15474 18320 15530 18329
rect 15474 18255 15530 18264
rect 15384 18148 15436 18154
rect 15384 18090 15436 18096
rect 15292 17808 15344 17814
rect 15292 17750 15344 17756
rect 15108 17604 15160 17610
rect 15108 17546 15160 17552
rect 15120 17490 15148 17546
rect 15120 17462 15240 17490
rect 14924 17332 14976 17338
rect 14924 17274 14976 17280
rect 14832 17264 14884 17270
rect 14832 17206 14884 17212
rect 15212 17134 15240 17462
rect 15200 17128 15252 17134
rect 14922 17096 14978 17105
rect 15200 17070 15252 17076
rect 14922 17031 14978 17040
rect 14936 16998 14964 17031
rect 14924 16992 14976 16998
rect 14924 16934 14976 16940
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 14924 16720 14976 16726
rect 14924 16662 14976 16668
rect 14936 15706 14964 16662
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14660 13977 14688 14350
rect 14646 13968 14702 13977
rect 14646 13903 14702 13912
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14660 13190 14688 13738
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14660 11744 14688 13126
rect 14752 12442 14780 15438
rect 15028 15162 15056 16934
rect 15212 16590 15240 17070
rect 15396 16658 15424 18090
rect 15476 17808 15528 17814
rect 15476 17750 15528 17756
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 15212 16114 15240 16526
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15200 15904 15252 15910
rect 15198 15872 15200 15881
rect 15252 15872 15254 15881
rect 15198 15807 15254 15816
rect 15106 15736 15162 15745
rect 15106 15671 15108 15680
rect 15160 15671 15162 15680
rect 15108 15642 15160 15648
rect 15108 15564 15160 15570
rect 15108 15506 15160 15512
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14844 11898 14872 14758
rect 14936 14618 14964 14962
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14936 14113 14964 14554
rect 14922 14104 14978 14113
rect 14922 14039 14978 14048
rect 14924 13796 14976 13802
rect 14924 13738 14976 13744
rect 15016 13796 15068 13802
rect 15016 13738 15068 13744
rect 14936 13394 14964 13738
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14936 12782 14964 13330
rect 14924 12776 14976 12782
rect 14924 12718 14976 12724
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14936 11898 14964 12582
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 14660 11716 14780 11744
rect 14648 11620 14700 11626
rect 14648 11562 14700 11568
rect 14660 10266 14688 11562
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14648 10260 14700 10266
rect 14648 10202 14700 10208
rect 14752 10146 14780 11716
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14568 10118 14780 10146
rect 14464 9444 14516 9450
rect 14464 9386 14516 9392
rect 14476 8090 14504 9386
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14462 7712 14518 7721
rect 14462 7647 14518 7656
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 14372 6860 14424 6866
rect 14372 6802 14424 6808
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14186 5944 14242 5953
rect 14292 5914 14320 6054
rect 14384 5930 14412 6802
rect 14476 6089 14504 7647
rect 14568 6202 14596 10118
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14660 6730 14688 9998
rect 14752 9586 14780 9998
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14740 9444 14792 9450
rect 14740 9386 14792 9392
rect 14752 9081 14780 9386
rect 14738 9072 14794 9081
rect 14844 9042 14872 11630
rect 14922 10976 14978 10985
rect 14922 10911 14978 10920
rect 14936 10130 14964 10911
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 14936 9110 14964 9862
rect 15028 9518 15056 13738
rect 15120 10130 15148 15506
rect 15488 15366 15516 17750
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 15212 12220 15240 15302
rect 15580 15008 15608 21422
rect 15672 19961 15700 23920
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 16488 21548 16540 21554
rect 16488 21490 16540 21496
rect 15750 21244 16046 21264
rect 15806 21242 15830 21244
rect 15886 21242 15910 21244
rect 15966 21242 15990 21244
rect 15828 21190 15830 21242
rect 15892 21190 15904 21242
rect 15966 21190 15968 21242
rect 15806 21188 15830 21190
rect 15886 21188 15910 21190
rect 15966 21188 15990 21190
rect 15750 21168 16046 21188
rect 16132 20466 16160 21490
rect 16304 21344 16356 21350
rect 16304 21286 16356 21292
rect 16212 20528 16264 20534
rect 16212 20470 16264 20476
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 15750 20156 16046 20176
rect 15806 20154 15830 20156
rect 15886 20154 15910 20156
rect 15966 20154 15990 20156
rect 15828 20102 15830 20154
rect 15892 20102 15904 20154
rect 15966 20102 15968 20154
rect 15806 20100 15830 20102
rect 15886 20100 15910 20102
rect 15966 20100 15990 20102
rect 15750 20080 16046 20100
rect 15658 19952 15714 19961
rect 15658 19887 15714 19896
rect 16224 19768 16252 20470
rect 16316 20369 16344 21286
rect 16302 20360 16358 20369
rect 16302 20295 16358 20304
rect 16304 20256 16356 20262
rect 16304 20198 16356 20204
rect 16316 19990 16344 20198
rect 16304 19984 16356 19990
rect 16304 19926 16356 19932
rect 16132 19740 16252 19768
rect 16132 19417 16160 19740
rect 16396 19712 16448 19718
rect 16224 19672 16396 19700
rect 16118 19408 16174 19417
rect 15936 19372 15988 19378
rect 16118 19343 16174 19352
rect 15936 19314 15988 19320
rect 15948 19258 15976 19314
rect 16132 19310 16160 19343
rect 15672 19230 15976 19258
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 15672 17105 15700 19230
rect 15750 19068 16046 19088
rect 15806 19066 15830 19068
rect 15886 19066 15910 19068
rect 15966 19066 15990 19068
rect 15828 19014 15830 19066
rect 15892 19014 15904 19066
rect 15966 19014 15968 19066
rect 15806 19012 15830 19014
rect 15886 19012 15910 19014
rect 15966 19012 15990 19014
rect 15750 18992 16046 19012
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 15750 17980 16046 18000
rect 15806 17978 15830 17980
rect 15886 17978 15910 17980
rect 15966 17978 15990 17980
rect 15828 17926 15830 17978
rect 15892 17926 15904 17978
rect 15966 17926 15968 17978
rect 15806 17924 15830 17926
rect 15886 17924 15910 17926
rect 15966 17924 15990 17926
rect 15750 17904 16046 17924
rect 16132 17814 16160 18906
rect 16224 18902 16252 19672
rect 16396 19654 16448 19660
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16212 18896 16264 18902
rect 16212 18838 16264 18844
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 16224 17882 16252 18226
rect 16316 18154 16344 19110
rect 16396 18420 16448 18426
rect 16396 18362 16448 18368
rect 16304 18148 16356 18154
rect 16304 18090 16356 18096
rect 16212 17876 16264 17882
rect 16212 17818 16264 17824
rect 16120 17808 16172 17814
rect 16120 17750 16172 17756
rect 16304 17808 16356 17814
rect 16304 17750 16356 17756
rect 15658 17096 15714 17105
rect 15658 17031 15714 17040
rect 15750 16892 16046 16912
rect 15806 16890 15830 16892
rect 15886 16890 15910 16892
rect 15966 16890 15990 16892
rect 15828 16838 15830 16890
rect 15892 16838 15904 16890
rect 15966 16838 15968 16890
rect 15806 16836 15830 16838
rect 15886 16836 15910 16838
rect 15966 16836 15990 16838
rect 15750 16816 16046 16836
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15672 15978 15700 16730
rect 16316 16425 16344 17750
rect 16302 16416 16358 16425
rect 16408 16402 16436 18362
rect 16500 17338 16528 21490
rect 16580 20460 16632 20466
rect 16580 20402 16632 20408
rect 16592 19378 16620 20402
rect 16684 19718 16712 21966
rect 16960 21962 16988 23920
rect 16948 21956 17000 21962
rect 16948 21898 17000 21904
rect 16764 21616 16816 21622
rect 16764 21558 16816 21564
rect 16776 20466 16804 21558
rect 16856 21344 16908 21350
rect 16856 21286 16908 21292
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16580 19372 16632 19378
rect 16580 19314 16632 19320
rect 16672 19304 16724 19310
rect 16672 19246 16724 19252
rect 16578 18728 16634 18737
rect 16578 18663 16634 18672
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 16500 16658 16528 17274
rect 16488 16652 16540 16658
rect 16488 16594 16540 16600
rect 16408 16374 16528 16402
rect 16302 16351 16358 16360
rect 15660 15972 15712 15978
rect 15660 15914 15712 15920
rect 15672 15473 15700 15914
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 15750 15804 16046 15824
rect 15806 15802 15830 15804
rect 15886 15802 15910 15804
rect 15966 15802 15990 15804
rect 15828 15750 15830 15802
rect 15892 15750 15904 15802
rect 15966 15750 15968 15802
rect 15806 15748 15830 15750
rect 15886 15748 15910 15750
rect 15966 15748 15990 15750
rect 15750 15728 16046 15748
rect 16132 15570 16160 15846
rect 15844 15564 15896 15570
rect 15844 15506 15896 15512
rect 16120 15564 16172 15570
rect 16120 15506 16172 15512
rect 15658 15464 15714 15473
rect 15658 15399 15714 15408
rect 15304 14980 15608 15008
rect 15304 12374 15332 14980
rect 15856 14929 15884 15506
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 15842 14920 15898 14929
rect 15842 14855 15898 14864
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15396 12714 15424 13670
rect 15384 12708 15436 12714
rect 15384 12650 15436 12656
rect 15292 12368 15344 12374
rect 15396 12345 15424 12650
rect 15292 12310 15344 12316
rect 15382 12336 15438 12345
rect 15488 12306 15516 14758
rect 15382 12271 15438 12280
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15212 12192 15424 12220
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15212 11354 15240 11834
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15212 10742 15240 11086
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15120 9722 15148 10066
rect 15198 10024 15254 10033
rect 15198 9959 15254 9968
rect 15212 9926 15240 9959
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 15108 9716 15160 9722
rect 15108 9658 15160 9664
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 14924 9104 14976 9110
rect 14924 9046 14976 9052
rect 14738 9007 14794 9016
rect 14832 9036 14884 9042
rect 14832 8978 14884 8984
rect 14740 8900 14792 8906
rect 14740 8842 14792 8848
rect 14752 8090 14780 8842
rect 14844 8634 14872 8978
rect 14922 8936 14978 8945
rect 14922 8871 14978 8880
rect 14936 8838 14964 8871
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 14832 8628 14884 8634
rect 14832 8570 14884 8576
rect 14936 8566 14964 8774
rect 14924 8560 14976 8566
rect 14924 8502 14976 8508
rect 15028 8430 15056 9318
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 15212 8838 15240 9046
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15016 8424 15068 8430
rect 15016 8366 15068 8372
rect 15014 8120 15070 8129
rect 14740 8084 14792 8090
rect 15014 8055 15070 8064
rect 14740 8026 14792 8032
rect 14924 7948 14976 7954
rect 14924 7890 14976 7896
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 14752 6254 14780 7822
rect 14936 7478 14964 7890
rect 15028 7721 15056 8055
rect 15014 7712 15070 7721
rect 15014 7647 15070 7656
rect 14924 7472 14976 7478
rect 15120 7426 15148 8434
rect 14924 7414 14976 7420
rect 15028 7398 15148 7426
rect 14832 7268 14884 7274
rect 14832 7210 14884 7216
rect 14844 7002 14872 7210
rect 15028 7177 15056 7398
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 15014 7168 15070 7177
rect 15014 7103 15070 7112
rect 14832 6996 14884 7002
rect 14832 6938 14884 6944
rect 14740 6248 14792 6254
rect 14568 6174 14688 6202
rect 14740 6190 14792 6196
rect 14556 6112 14608 6118
rect 14462 6080 14518 6089
rect 14556 6054 14608 6060
rect 14462 6015 14518 6024
rect 14568 5930 14596 6054
rect 14186 5879 14242 5888
rect 14280 5908 14332 5914
rect 14200 5166 14228 5879
rect 14384 5902 14596 5930
rect 14280 5850 14332 5856
rect 14370 5808 14426 5817
rect 14292 5766 14370 5794
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14188 4684 14240 4690
rect 14188 4626 14240 4632
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14004 4072 14056 4078
rect 14002 4040 14004 4049
rect 14056 4040 14058 4049
rect 14002 3975 14058 3984
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 14016 3058 14044 3538
rect 14094 3224 14150 3233
rect 14200 3194 14228 4626
rect 14292 3738 14320 5766
rect 14370 5743 14426 5752
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14384 5574 14412 5646
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14476 5370 14504 5646
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14476 4622 14504 5306
rect 14568 4758 14596 5902
rect 14556 4752 14608 4758
rect 14660 4729 14688 6174
rect 14752 5914 14780 6190
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14752 5234 14780 5850
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14556 4694 14608 4700
rect 14646 4720 14702 4729
rect 14646 4655 14702 4664
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14370 4176 14426 4185
rect 14370 4111 14426 4120
rect 14384 3942 14412 4111
rect 14752 4078 14780 5170
rect 14844 4826 14872 6938
rect 14924 6724 14976 6730
rect 14924 6666 14976 6672
rect 14936 5710 14964 6666
rect 15014 6352 15070 6361
rect 15014 6287 15070 6296
rect 14924 5704 14976 5710
rect 14924 5646 14976 5652
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14936 4486 14964 5306
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 14740 4072 14792 4078
rect 14646 4040 14702 4049
rect 14740 4014 14792 4020
rect 14646 3975 14702 3984
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14660 3602 14688 3975
rect 14648 3596 14700 3602
rect 14648 3538 14700 3544
rect 14844 3534 14872 4218
rect 14936 4078 14964 4422
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 15028 3942 15056 6287
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14094 3159 14096 3168
rect 14148 3159 14150 3168
rect 14188 3188 14240 3194
rect 14096 3130 14148 3136
rect 14188 3130 14240 3136
rect 15028 3058 15056 3878
rect 15120 3534 15148 7278
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 15106 3088 15162 3097
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 15016 3052 15068 3058
rect 15106 3023 15162 3032
rect 15016 2994 15068 3000
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 12530 2544 12586 2553
rect 14016 2514 14044 2994
rect 14370 2952 14426 2961
rect 14370 2887 14426 2896
rect 14384 2854 14412 2887
rect 15120 2854 15148 3023
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 12530 2479 12586 2488
rect 14004 2508 14056 2514
rect 14004 2450 14056 2456
rect 14372 2372 14424 2378
rect 14372 2314 14424 2320
rect 12052 2204 12348 2224
rect 12108 2202 12132 2204
rect 12188 2202 12212 2204
rect 12268 2202 12292 2204
rect 12130 2150 12132 2202
rect 12194 2150 12206 2202
rect 12268 2150 12270 2202
rect 12108 2148 12132 2150
rect 12188 2148 12212 2150
rect 12268 2148 12292 2150
rect 12052 2128 12348 2148
rect 11992 2060 12112 2088
rect 12084 480 12112 2060
rect 14384 2038 14412 2314
rect 14372 2032 14424 2038
rect 14372 1974 14424 1980
rect 15212 1834 15240 8774
rect 15304 7342 15332 12038
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15304 7002 15332 7142
rect 15292 6996 15344 7002
rect 15292 6938 15344 6944
rect 15292 6180 15344 6186
rect 15292 6122 15344 6128
rect 15304 4486 15332 6122
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 15396 3194 15424 12192
rect 15476 12164 15528 12170
rect 15476 12106 15528 12112
rect 15488 8634 15516 12106
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15488 7886 15516 8366
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15580 7392 15608 14758
rect 15750 14716 16046 14736
rect 15806 14714 15830 14716
rect 15886 14714 15910 14716
rect 15966 14714 15990 14716
rect 15828 14662 15830 14714
rect 15892 14662 15904 14714
rect 15966 14662 15968 14714
rect 15806 14660 15830 14662
rect 15886 14660 15910 14662
rect 15966 14660 15990 14662
rect 15750 14640 16046 14660
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15672 12442 15700 14418
rect 15752 14272 15804 14278
rect 15750 14240 15752 14249
rect 15804 14240 15806 14249
rect 15750 14175 15806 14184
rect 15750 13628 16046 13648
rect 15806 13626 15830 13628
rect 15886 13626 15910 13628
rect 15966 13626 15990 13628
rect 15828 13574 15830 13626
rect 15892 13574 15904 13626
rect 15966 13574 15968 13626
rect 15806 13572 15830 13574
rect 15886 13572 15910 13574
rect 15966 13572 15990 13574
rect 15750 13552 16046 13572
rect 16132 13433 16160 15302
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16224 14657 16252 14758
rect 16210 14648 16266 14657
rect 16210 14583 16266 14592
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16118 13424 16174 13433
rect 15844 13388 15896 13394
rect 16118 13359 16174 13368
rect 15844 13330 15896 13336
rect 15856 13161 15884 13330
rect 15842 13152 15898 13161
rect 15842 13087 15898 13096
rect 15750 12540 16046 12560
rect 15806 12538 15830 12540
rect 15886 12538 15910 12540
rect 15966 12538 15990 12540
rect 15828 12486 15830 12538
rect 15892 12486 15904 12538
rect 15966 12486 15968 12538
rect 15806 12484 15830 12486
rect 15886 12484 15910 12486
rect 15966 12484 15990 12486
rect 15750 12464 16046 12484
rect 15660 12436 15712 12442
rect 16132 12424 16160 13359
rect 15660 12378 15712 12384
rect 16040 12396 16160 12424
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15764 11937 15792 12242
rect 15750 11928 15806 11937
rect 15750 11863 15806 11872
rect 16040 11762 16068 12396
rect 16224 12356 16252 14350
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16316 12918 16344 13330
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 16132 12328 16252 12356
rect 16132 11898 16160 12328
rect 16316 12220 16344 12854
rect 16408 12442 16436 12922
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16224 12192 16344 12220
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 15672 10985 15700 11698
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 15750 11452 16046 11472
rect 15806 11450 15830 11452
rect 15886 11450 15910 11452
rect 15966 11450 15990 11452
rect 15828 11398 15830 11450
rect 15892 11398 15904 11450
rect 15966 11398 15968 11450
rect 15806 11396 15830 11398
rect 15886 11396 15910 11398
rect 15966 11396 15990 11398
rect 15750 11376 16046 11396
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 15658 10976 15714 10985
rect 15658 10911 15714 10920
rect 15658 10840 15714 10849
rect 15658 10775 15714 10784
rect 15672 7834 15700 10775
rect 15948 10538 15976 11154
rect 16132 10538 16160 11494
rect 15936 10532 15988 10538
rect 15936 10474 15988 10480
rect 16120 10532 16172 10538
rect 16120 10474 16172 10480
rect 15750 10364 16046 10384
rect 15806 10362 15830 10364
rect 15886 10362 15910 10364
rect 15966 10362 15990 10364
rect 15828 10310 15830 10362
rect 15892 10310 15904 10362
rect 15966 10310 15968 10362
rect 15806 10308 15830 10310
rect 15886 10308 15910 10310
rect 15966 10308 15990 10310
rect 15750 10288 16046 10308
rect 16132 10266 16160 10474
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16118 10160 16174 10169
rect 16118 10095 16174 10104
rect 15750 9276 16046 9296
rect 15806 9274 15830 9276
rect 15886 9274 15910 9276
rect 15966 9274 15990 9276
rect 15828 9222 15830 9274
rect 15892 9222 15904 9274
rect 15966 9222 15968 9274
rect 15806 9220 15830 9222
rect 15886 9220 15910 9222
rect 15966 9220 15990 9222
rect 15750 9200 16046 9220
rect 15750 8188 16046 8208
rect 15806 8186 15830 8188
rect 15886 8186 15910 8188
rect 15966 8186 15990 8188
rect 15828 8134 15830 8186
rect 15892 8134 15904 8186
rect 15966 8134 15968 8186
rect 15806 8132 15830 8134
rect 15886 8132 15910 8134
rect 15966 8132 15990 8134
rect 15750 8112 16046 8132
rect 16132 7834 16160 10095
rect 15672 7806 15792 7834
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15488 7364 15608 7392
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15488 2310 15516 7364
rect 15672 7324 15700 7686
rect 15580 7296 15700 7324
rect 15580 5273 15608 7296
rect 15764 7188 15792 7806
rect 16040 7806 16160 7834
rect 16040 7750 16068 7806
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 15842 7440 15898 7449
rect 15842 7375 15844 7384
rect 15896 7375 15898 7384
rect 16120 7404 16172 7410
rect 15844 7346 15896 7352
rect 16120 7346 16172 7352
rect 15672 7160 15792 7188
rect 15566 5264 15622 5273
rect 15566 5199 15622 5208
rect 15672 5137 15700 7160
rect 15750 7100 16046 7120
rect 15806 7098 15830 7100
rect 15886 7098 15910 7100
rect 15966 7098 15990 7100
rect 15828 7046 15830 7098
rect 15892 7046 15904 7098
rect 15966 7046 15968 7098
rect 15806 7044 15830 7046
rect 15886 7044 15910 7046
rect 15966 7044 15990 7046
rect 15750 7024 16046 7044
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15764 6390 15792 6802
rect 15752 6384 15804 6390
rect 15752 6326 15804 6332
rect 15764 6186 15792 6326
rect 15752 6180 15804 6186
rect 15752 6122 15804 6128
rect 15750 6012 16046 6032
rect 15806 6010 15830 6012
rect 15886 6010 15910 6012
rect 15966 6010 15990 6012
rect 15828 5958 15830 6010
rect 15892 5958 15904 6010
rect 15966 5958 15968 6010
rect 15806 5956 15830 5958
rect 15886 5956 15910 5958
rect 15966 5956 15990 5958
rect 15750 5936 16046 5956
rect 16028 5636 16080 5642
rect 16028 5578 16080 5584
rect 16040 5166 16068 5578
rect 16028 5160 16080 5166
rect 15658 5128 15714 5137
rect 15568 5092 15620 5098
rect 16028 5102 16080 5108
rect 15658 5063 15714 5072
rect 15568 5034 15620 5040
rect 15580 4554 15608 5034
rect 15750 4924 16046 4944
rect 15806 4922 15830 4924
rect 15886 4922 15910 4924
rect 15966 4922 15990 4924
rect 15828 4870 15830 4922
rect 15892 4870 15904 4922
rect 15966 4870 15968 4922
rect 15806 4868 15830 4870
rect 15886 4868 15910 4870
rect 15966 4868 15990 4870
rect 15750 4848 16046 4868
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15568 4548 15620 4554
rect 15568 4490 15620 4496
rect 15672 4214 15700 4626
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 15660 4208 15712 4214
rect 15660 4150 15712 4156
rect 15566 3632 15622 3641
rect 15566 3567 15568 3576
rect 15620 3567 15622 3576
rect 15568 3538 15620 3544
rect 15568 3392 15620 3398
rect 15568 3334 15620 3340
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 15200 1828 15252 1834
rect 15200 1770 15252 1776
rect 15580 480 15608 3334
rect 15672 2650 15700 4150
rect 15856 4146 15884 4422
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 15750 3836 16046 3856
rect 15806 3834 15830 3836
rect 15886 3834 15910 3836
rect 15966 3834 15990 3836
rect 15828 3782 15830 3834
rect 15892 3782 15904 3834
rect 15966 3782 15968 3834
rect 15806 3780 15830 3782
rect 15886 3780 15910 3782
rect 15966 3780 15990 3782
rect 15750 3760 16046 3780
rect 16132 3738 16160 7346
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16224 3618 16252 12192
rect 16408 11830 16436 12378
rect 16396 11824 16448 11830
rect 16396 11766 16448 11772
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16304 10532 16356 10538
rect 16304 10474 16356 10480
rect 16316 10033 16344 10474
rect 16408 10198 16436 11494
rect 16396 10192 16448 10198
rect 16396 10134 16448 10140
rect 16302 10024 16358 10033
rect 16302 9959 16358 9968
rect 16316 9330 16344 9959
rect 16408 9654 16436 10134
rect 16396 9648 16448 9654
rect 16396 9590 16448 9596
rect 16316 9302 16436 9330
rect 16408 9042 16436 9302
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16316 8634 16344 8910
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16316 7546 16344 7686
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16316 6866 16344 7482
rect 16408 6866 16436 7890
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 16302 6760 16358 6769
rect 16302 6695 16358 6704
rect 16132 3590 16252 3618
rect 15750 2748 16046 2768
rect 15806 2746 15830 2748
rect 15886 2746 15910 2748
rect 15966 2746 15990 2748
rect 15828 2694 15830 2746
rect 15892 2694 15904 2746
rect 15966 2694 15968 2746
rect 15806 2692 15830 2694
rect 15886 2692 15910 2694
rect 15966 2692 15990 2694
rect 15750 2672 16046 2692
rect 15660 2644 15712 2650
rect 15660 2586 15712 2592
rect 16132 2378 16160 3590
rect 16316 3466 16344 6695
rect 16396 5568 16448 5574
rect 16396 5510 16448 5516
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 16304 2304 16356 2310
rect 16304 2246 16356 2252
rect 16316 1902 16344 2246
rect 16304 1896 16356 1902
rect 16304 1838 16356 1844
rect 16408 1358 16436 5510
rect 16500 3194 16528 16374
rect 16592 16266 16620 18663
rect 16684 17649 16712 19246
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16776 18873 16804 19110
rect 16868 18970 16896 21286
rect 16960 21146 16988 21286
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 16856 18964 16908 18970
rect 16856 18906 16908 18912
rect 16762 18864 16818 18873
rect 16762 18799 16818 18808
rect 16856 18216 16908 18222
rect 16856 18158 16908 18164
rect 16670 17640 16726 17649
rect 16670 17575 16726 17584
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16684 16998 16712 17478
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16868 16697 16896 18158
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16854 16688 16910 16697
rect 16854 16623 16910 16632
rect 16592 16238 16804 16266
rect 16580 16176 16632 16182
rect 16578 16144 16580 16153
rect 16632 16144 16634 16153
rect 16578 16079 16634 16088
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16592 11257 16620 12582
rect 16776 11898 16804 16238
rect 16856 16040 16908 16046
rect 16856 15982 16908 15988
rect 16868 13025 16896 15982
rect 16960 13258 16988 18022
rect 16948 13252 17000 13258
rect 16948 13194 17000 13200
rect 16854 13016 16910 13025
rect 16854 12951 16910 12960
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16672 11824 16724 11830
rect 16672 11766 16724 11772
rect 16578 11248 16634 11257
rect 16578 11183 16634 11192
rect 16580 10532 16632 10538
rect 16580 10474 16632 10480
rect 16592 7993 16620 10474
rect 16578 7984 16634 7993
rect 16684 7954 16712 11766
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16578 7919 16634 7928
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 16776 7410 16804 11630
rect 16868 8498 16896 12786
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16684 6610 16712 6734
rect 16592 6582 16712 6610
rect 16592 6390 16620 6582
rect 16868 6497 16896 7278
rect 16854 6488 16910 6497
rect 16854 6423 16910 6432
rect 16580 6384 16632 6390
rect 16580 6326 16632 6332
rect 16764 6384 16816 6390
rect 16764 6326 16816 6332
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 16684 4690 16712 6258
rect 16776 5710 16804 6326
rect 16960 6322 16988 11494
rect 17052 10130 17080 20198
rect 17236 19786 17264 20198
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17224 19780 17276 19786
rect 17224 19722 17276 19728
rect 17132 19712 17184 19718
rect 17132 19654 17184 19660
rect 17144 17746 17172 19654
rect 17420 19394 17448 19994
rect 17236 19366 17448 19394
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 17144 14521 17172 17206
rect 17130 14512 17186 14521
rect 17130 14447 17186 14456
rect 17236 14362 17264 19366
rect 17408 19304 17460 19310
rect 17408 19246 17460 19252
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17144 14334 17264 14362
rect 17144 12850 17172 14334
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 17236 12646 17264 14214
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17328 12458 17356 19110
rect 17420 18057 17448 19246
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17512 18358 17540 18702
rect 17500 18352 17552 18358
rect 17500 18294 17552 18300
rect 17500 18080 17552 18086
rect 17406 18048 17462 18057
rect 17500 18022 17552 18028
rect 17406 17983 17462 17992
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17420 17134 17448 17478
rect 17512 17241 17540 18022
rect 17498 17232 17554 17241
rect 17498 17167 17554 17176
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17500 16516 17552 16522
rect 17500 16458 17552 16464
rect 17408 13796 17460 13802
rect 17408 13738 17460 13744
rect 17420 13190 17448 13738
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 17144 12430 17356 12458
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 17038 9752 17094 9761
rect 17038 9687 17094 9696
rect 17052 7342 17080 9687
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 17038 6896 17094 6905
rect 17038 6831 17094 6840
rect 17052 6662 17080 6831
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 16868 5370 16896 6190
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 16948 4684 17000 4690
rect 16948 4626 17000 4632
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16592 4010 16620 4422
rect 16580 4004 16632 4010
rect 16580 3946 16632 3952
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16488 2576 16540 2582
rect 16592 2564 16620 3946
rect 16960 3738 16988 4626
rect 17052 4554 17080 5714
rect 17040 4548 17092 4554
rect 17040 4490 17092 4496
rect 17144 4049 17172 12430
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 17236 11354 17264 12242
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 17224 11212 17276 11218
rect 17224 11154 17276 11160
rect 17236 11121 17264 11154
rect 17222 11112 17278 11121
rect 17222 11047 17278 11056
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 17236 10713 17264 10950
rect 17222 10704 17278 10713
rect 17222 10639 17278 10648
rect 17328 10266 17356 11834
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17236 9110 17264 9862
rect 17314 9480 17370 9489
rect 17314 9415 17370 9424
rect 17328 9382 17356 9415
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17236 7993 17264 8366
rect 17328 8090 17356 9318
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17222 7984 17278 7993
rect 17222 7919 17278 7928
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17236 5778 17264 6598
rect 17224 5772 17276 5778
rect 17224 5714 17276 5720
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17130 4040 17186 4049
rect 17130 3975 17186 3984
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 17052 3534 17080 3878
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17052 2922 17080 3470
rect 17040 2916 17092 2922
rect 17040 2858 17092 2864
rect 16540 2536 16620 2564
rect 16764 2576 16816 2582
rect 16488 2518 16540 2524
rect 16764 2518 16816 2524
rect 16776 2106 16804 2518
rect 16764 2100 16816 2106
rect 16764 2042 16816 2048
rect 17236 2038 17264 4966
rect 17328 4690 17356 6734
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17420 4593 17448 13126
rect 17512 11880 17540 16458
rect 17604 16250 17632 23920
rect 17684 21616 17736 21622
rect 17684 21558 17736 21564
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 17696 15609 17724 21558
rect 18052 21072 18104 21078
rect 18052 21014 18104 21020
rect 17776 20800 17828 20806
rect 17776 20742 17828 20748
rect 17682 15600 17738 15609
rect 17682 15535 17738 15544
rect 17684 15428 17736 15434
rect 17684 15370 17736 15376
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17604 13870 17632 14418
rect 17592 13864 17644 13870
rect 17696 13852 17724 15370
rect 17788 14657 17816 20742
rect 18064 20398 18092 21014
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 17868 19916 17920 19922
rect 18064 19904 18092 20334
rect 17920 19876 18092 19904
rect 17868 19858 17920 19864
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 17972 19281 18000 19654
rect 18064 19310 18092 19876
rect 18052 19304 18104 19310
rect 17958 19272 18014 19281
rect 18052 19246 18104 19252
rect 17958 19207 18014 19216
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17868 18216 17920 18222
rect 17868 18158 17920 18164
rect 17880 16726 17908 18158
rect 17972 17785 18000 19110
rect 18064 18290 18092 19246
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 18064 17814 18092 18226
rect 18052 17808 18104 17814
rect 17958 17776 18014 17785
rect 18052 17750 18104 17756
rect 17958 17711 18014 17720
rect 18064 17082 18092 17750
rect 17972 17054 18092 17082
rect 17972 16794 18000 17054
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 17868 16720 17920 16726
rect 17868 16662 17920 16668
rect 17774 14648 17830 14657
rect 17774 14583 17830 14592
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17788 14074 17816 14418
rect 17880 14074 17908 16662
rect 17960 15632 18012 15638
rect 17960 15574 18012 15580
rect 17972 15162 18000 15574
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 18064 15094 18092 16934
rect 18052 15088 18104 15094
rect 18052 15030 18104 15036
rect 18248 14958 18276 23920
rect 18892 23882 18920 23920
rect 18800 23854 18920 23882
rect 18696 21956 18748 21962
rect 18696 21898 18748 21904
rect 18328 21888 18380 21894
rect 18328 21830 18380 21836
rect 18340 21486 18368 21830
rect 18604 21548 18656 21554
rect 18604 21490 18656 21496
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 18512 18624 18564 18630
rect 18512 18566 18564 18572
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 18340 15201 18368 16934
rect 18432 16454 18460 17614
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18326 15192 18382 15201
rect 18326 15127 18382 15136
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 17696 13824 17816 13852
rect 17592 13806 17644 13812
rect 17604 13716 17632 13806
rect 17604 13688 17724 13716
rect 17696 13326 17724 13688
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17684 13184 17736 13190
rect 17684 13126 17736 13132
rect 17512 11852 17632 11880
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17512 9042 17540 11698
rect 17604 10538 17632 11852
rect 17696 11150 17724 13126
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 17682 10976 17738 10985
rect 17682 10911 17738 10920
rect 17696 10810 17724 10911
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17592 10532 17644 10538
rect 17592 10474 17644 10480
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 17604 9110 17632 10066
rect 17592 9104 17644 9110
rect 17592 9046 17644 9052
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 17512 8634 17540 8978
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17604 7954 17632 8774
rect 17592 7948 17644 7954
rect 17592 7890 17644 7896
rect 17604 6322 17632 7890
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 17696 6254 17724 10406
rect 17788 9761 17816 13824
rect 17868 13252 17920 13258
rect 17868 13194 17920 13200
rect 17880 12918 17908 13194
rect 17868 12912 17920 12918
rect 17868 12854 17920 12860
rect 17868 12776 17920 12782
rect 17866 12744 17868 12753
rect 17920 12744 17922 12753
rect 17866 12679 17922 12688
rect 17868 12640 17920 12646
rect 17868 12582 17920 12588
rect 17880 12374 17908 12582
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17866 11248 17922 11257
rect 17866 11183 17868 11192
rect 17920 11183 17922 11192
rect 17868 11154 17920 11160
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17774 9752 17830 9761
rect 17774 9687 17830 9696
rect 17880 9654 17908 10066
rect 17868 9648 17920 9654
rect 17868 9590 17920 9596
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17788 9466 17816 9522
rect 17788 9438 17908 9466
rect 17776 9376 17828 9382
rect 17880 9353 17908 9438
rect 17776 9318 17828 9324
rect 17866 9344 17922 9353
rect 17788 8906 17816 9318
rect 17866 9279 17922 9288
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 17776 8900 17828 8906
rect 17776 8842 17828 8848
rect 17880 8362 17908 9046
rect 17868 8356 17920 8362
rect 17868 8298 17920 8304
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 17880 6118 17908 8298
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 17868 5840 17920 5846
rect 17868 5782 17920 5788
rect 17682 5400 17738 5409
rect 17682 5335 17738 5344
rect 17592 5228 17644 5234
rect 17592 5170 17644 5176
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 17512 4826 17540 4966
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 17406 4584 17462 4593
rect 17406 4519 17462 4528
rect 17604 4146 17632 5170
rect 17696 4486 17724 5335
rect 17880 5234 17908 5782
rect 17868 5228 17920 5234
rect 17868 5170 17920 5176
rect 17776 5160 17828 5166
rect 17776 5102 17828 5108
rect 17788 4826 17816 5102
rect 17868 5092 17920 5098
rect 17868 5034 17920 5040
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17500 3664 17552 3670
rect 17500 3606 17552 3612
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 17328 2961 17356 2994
rect 17314 2952 17370 2961
rect 17314 2887 17370 2896
rect 17512 2854 17540 3606
rect 17696 2990 17724 3878
rect 17776 3664 17828 3670
rect 17776 3606 17828 3612
rect 17788 3398 17816 3606
rect 17776 3392 17828 3398
rect 17776 3334 17828 3340
rect 17684 2984 17736 2990
rect 17684 2926 17736 2932
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17512 2650 17724 2666
rect 17500 2644 17724 2650
rect 17552 2638 17724 2644
rect 17500 2586 17552 2592
rect 17696 2582 17724 2638
rect 17684 2576 17736 2582
rect 17684 2518 17736 2524
rect 17408 2508 17460 2514
rect 17408 2450 17460 2456
rect 17420 2038 17448 2450
rect 17500 2372 17552 2378
rect 17500 2314 17552 2320
rect 17224 2032 17276 2038
rect 17224 1974 17276 1980
rect 17408 2032 17460 2038
rect 17408 1974 17460 1980
rect 17512 1970 17540 2314
rect 17880 2310 17908 5034
rect 17972 3641 18000 14894
rect 18052 13728 18104 13734
rect 18052 13670 18104 13676
rect 18064 11642 18092 13670
rect 18234 13288 18290 13297
rect 18234 13223 18290 13232
rect 18248 12918 18276 13223
rect 18236 12912 18288 12918
rect 18236 12854 18288 12860
rect 18340 11665 18368 14962
rect 18524 14521 18552 18566
rect 18616 14822 18644 21490
rect 18708 19990 18736 21898
rect 18800 20058 18828 23854
rect 19246 23352 19302 23361
rect 19246 23287 19302 23296
rect 19154 22672 19210 22681
rect 19154 22607 19210 22616
rect 18880 21480 18932 21486
rect 18880 21422 18932 21428
rect 18892 21078 18920 21422
rect 19062 21312 19118 21321
rect 19062 21247 19118 21256
rect 18880 21072 18932 21078
rect 18880 21014 18932 21020
rect 19076 20602 19104 21247
rect 19168 21146 19196 22607
rect 19260 21350 19288 23287
rect 19536 21962 19564 23920
rect 19524 21956 19576 21962
rect 19524 21898 19576 21904
rect 19449 21788 19745 21808
rect 19505 21786 19529 21788
rect 19585 21786 19609 21788
rect 19665 21786 19689 21788
rect 19527 21734 19529 21786
rect 19591 21734 19603 21786
rect 19665 21734 19667 21786
rect 19505 21732 19529 21734
rect 19585 21732 19609 21734
rect 19665 21732 19689 21734
rect 19449 21712 19745 21732
rect 19812 21690 19840 23967
rect 20166 23920 20222 24400
rect 20810 23920 20866 24400
rect 21454 23920 21510 24400
rect 22098 23920 22154 24400
rect 22742 23920 22798 24400
rect 23386 23920 23442 24400
rect 24030 23920 24086 24400
rect 20180 23882 20208 23920
rect 19996 23854 20208 23882
rect 19890 21992 19946 22001
rect 19890 21927 19946 21936
rect 19800 21684 19852 21690
rect 19800 21626 19852 21632
rect 19904 21486 19932 21927
rect 19892 21480 19944 21486
rect 19892 21422 19944 21428
rect 19340 21412 19392 21418
rect 19340 21354 19392 21360
rect 19248 21344 19300 21350
rect 19248 21286 19300 21292
rect 19156 21140 19208 21146
rect 19156 21082 19208 21088
rect 19352 20806 19380 21354
rect 19800 21004 19852 21010
rect 19800 20946 19852 20952
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19449 20700 19745 20720
rect 19505 20698 19529 20700
rect 19585 20698 19609 20700
rect 19665 20698 19689 20700
rect 19527 20646 19529 20698
rect 19591 20646 19603 20698
rect 19665 20646 19667 20698
rect 19505 20644 19529 20646
rect 19585 20644 19609 20646
rect 19665 20644 19689 20646
rect 19449 20624 19745 20644
rect 19812 20602 19840 20946
rect 19890 20632 19946 20641
rect 19064 20596 19116 20602
rect 19064 20538 19116 20544
rect 19800 20596 19852 20602
rect 19890 20567 19946 20576
rect 19800 20538 19852 20544
rect 19156 20324 19208 20330
rect 19156 20266 19208 20272
rect 19168 20058 19196 20266
rect 19338 20088 19394 20097
rect 18788 20052 18840 20058
rect 18788 19994 18840 20000
rect 19156 20052 19208 20058
rect 19338 20023 19394 20032
rect 19156 19994 19208 20000
rect 18696 19984 18748 19990
rect 18696 19926 18748 19932
rect 18880 19916 18932 19922
rect 18880 19858 18932 19864
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18800 19553 18828 19790
rect 18786 19544 18842 19553
rect 18786 19479 18842 19488
rect 18696 19304 18748 19310
rect 18696 19246 18748 19252
rect 18708 18426 18736 19246
rect 18892 18970 18920 19858
rect 19248 19712 19300 19718
rect 19246 19680 19248 19689
rect 19300 19680 19302 19689
rect 19246 19615 19302 19624
rect 19352 19514 19380 20023
rect 19812 19990 19840 20538
rect 19800 19984 19852 19990
rect 19800 19926 19852 19932
rect 19800 19848 19852 19854
rect 19800 19790 19852 19796
rect 19449 19612 19745 19632
rect 19505 19610 19529 19612
rect 19585 19610 19609 19612
rect 19665 19610 19689 19612
rect 19527 19558 19529 19610
rect 19591 19558 19603 19610
rect 19665 19558 19667 19610
rect 19505 19556 19529 19558
rect 19585 19556 19609 19558
rect 19665 19556 19689 19558
rect 19449 19536 19745 19556
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19432 19440 19484 19446
rect 19432 19382 19484 19388
rect 19248 19236 19300 19242
rect 19248 19178 19300 19184
rect 19260 19122 19288 19178
rect 19260 19094 19380 19122
rect 18880 18964 18932 18970
rect 18880 18906 18932 18912
rect 19352 18426 19380 19094
rect 19444 18902 19472 19382
rect 19432 18896 19484 18902
rect 19432 18838 19484 18844
rect 19812 18766 19840 19790
rect 19904 19786 19932 20567
rect 19996 20330 20024 23854
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 19984 20324 20036 20330
rect 19984 20266 20036 20272
rect 19892 19780 19944 19786
rect 19892 19722 19944 19728
rect 19892 19372 19944 19378
rect 19892 19314 19944 19320
rect 19800 18760 19852 18766
rect 19800 18702 19852 18708
rect 19449 18524 19745 18544
rect 19505 18522 19529 18524
rect 19585 18522 19609 18524
rect 19665 18522 19689 18524
rect 19527 18470 19529 18522
rect 19591 18470 19603 18522
rect 19665 18470 19667 18522
rect 19505 18468 19529 18470
rect 19585 18468 19609 18470
rect 19665 18468 19689 18470
rect 19449 18448 19745 18468
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 18788 18148 18840 18154
rect 18788 18090 18840 18096
rect 18800 17882 18828 18090
rect 18788 17876 18840 17882
rect 18788 17818 18840 17824
rect 19352 17814 19380 18362
rect 19340 17808 19392 17814
rect 19340 17750 19392 17756
rect 18972 17740 19024 17746
rect 18972 17682 19024 17688
rect 19248 17740 19300 17746
rect 19248 17682 19300 17688
rect 18984 17134 19012 17682
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18708 15366 18736 15982
rect 18800 15638 18828 16526
rect 18788 15632 18840 15638
rect 18788 15574 18840 15580
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 18510 14512 18566 14521
rect 18510 14447 18566 14456
rect 18512 14340 18564 14346
rect 18512 14282 18564 14288
rect 18524 13394 18552 14282
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18694 13152 18750 13161
rect 18616 12782 18644 13126
rect 18694 13087 18750 13096
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 18708 12714 18736 13087
rect 18696 12708 18748 12714
rect 18696 12650 18748 12656
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18708 11762 18736 12242
rect 18800 12170 18828 14826
rect 18892 14770 18920 16934
rect 18984 16794 19012 17070
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 18972 15564 19024 15570
rect 18972 15506 19024 15512
rect 18984 15162 19012 15506
rect 18972 15156 19024 15162
rect 18972 15098 19024 15104
rect 18892 14742 19012 14770
rect 18880 14272 18932 14278
rect 18880 14214 18932 14220
rect 18892 13938 18920 14214
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 18892 13462 18920 13874
rect 18880 13456 18932 13462
rect 18880 13398 18932 13404
rect 18788 12164 18840 12170
rect 18840 12124 18920 12152
rect 18788 12106 18840 12112
rect 18786 11928 18842 11937
rect 18786 11863 18842 11872
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18604 11688 18656 11694
rect 18326 11656 18382 11665
rect 18064 11614 18184 11642
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 18064 10674 18092 11494
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 18156 9625 18184 11614
rect 18604 11630 18656 11636
rect 18326 11591 18382 11600
rect 18616 11150 18644 11630
rect 18696 11620 18748 11626
rect 18696 11562 18748 11568
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18432 10810 18460 11086
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18236 10124 18288 10130
rect 18288 10084 18368 10112
rect 18236 10066 18288 10072
rect 18340 10033 18368 10084
rect 18326 10024 18382 10033
rect 18326 9959 18382 9968
rect 18142 9616 18198 9625
rect 18142 9551 18198 9560
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18156 9081 18184 9318
rect 18142 9072 18198 9081
rect 18052 9036 18104 9042
rect 18142 9007 18198 9016
rect 18052 8978 18104 8984
rect 18064 7449 18092 8978
rect 18248 8974 18276 9318
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18340 8090 18368 9959
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18340 7750 18368 8026
rect 18432 7936 18460 10202
rect 18616 9722 18644 11086
rect 18708 10266 18736 11562
rect 18696 10260 18748 10266
rect 18800 10248 18828 11863
rect 18892 10674 18920 12124
rect 18984 11937 19012 14742
rect 19076 12073 19104 17478
rect 19260 16658 19288 17682
rect 19812 17678 19840 18702
rect 19904 17746 19932 19314
rect 20088 18358 20116 21830
rect 20536 21480 20588 21486
rect 20536 21422 20588 21428
rect 20260 21344 20312 21350
rect 20260 21286 20312 21292
rect 20272 21078 20300 21286
rect 20260 21072 20312 21078
rect 20260 21014 20312 21020
rect 20168 20800 20220 20806
rect 20168 20742 20220 20748
rect 20180 20466 20208 20742
rect 20168 20460 20220 20466
rect 20168 20402 20220 20408
rect 20272 20330 20300 21014
rect 20548 20913 20576 21422
rect 20534 20904 20590 20913
rect 20534 20839 20590 20848
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 20260 20324 20312 20330
rect 20260 20266 20312 20272
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 20076 18352 20128 18358
rect 20076 18294 20128 18300
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19892 17740 19944 17746
rect 19892 17682 19944 17688
rect 19800 17672 19852 17678
rect 19800 17614 19852 17620
rect 19449 17436 19745 17456
rect 19505 17434 19529 17436
rect 19585 17434 19609 17436
rect 19665 17434 19689 17436
rect 19527 17382 19529 17434
rect 19591 17382 19603 17434
rect 19665 17382 19667 17434
rect 19505 17380 19529 17382
rect 19585 17380 19609 17382
rect 19665 17380 19689 17382
rect 19449 17360 19745 17380
rect 19812 17270 19840 17614
rect 19800 17264 19852 17270
rect 19852 17212 19932 17218
rect 19800 17206 19932 17212
rect 19812 17190 19932 17206
rect 19996 17202 20024 18022
rect 19800 17128 19852 17134
rect 19800 17070 19852 17076
rect 19904 17082 19932 17190
rect 19984 17196 20036 17202
rect 19984 17138 20036 17144
rect 19708 16720 19760 16726
rect 19812 16674 19840 17070
rect 19904 17054 20024 17082
rect 19996 16794 20024 17054
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 19760 16668 19840 16674
rect 19708 16662 19840 16668
rect 19892 16720 19944 16726
rect 19892 16662 19944 16668
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19340 16652 19392 16658
rect 19720 16646 19840 16662
rect 19340 16594 19392 16600
rect 19352 15978 19380 16594
rect 19449 16348 19745 16368
rect 19505 16346 19529 16348
rect 19585 16346 19609 16348
rect 19665 16346 19689 16348
rect 19527 16294 19529 16346
rect 19591 16294 19603 16346
rect 19665 16294 19667 16346
rect 19505 16292 19529 16294
rect 19585 16292 19609 16294
rect 19665 16292 19689 16294
rect 19449 16272 19745 16292
rect 19812 16250 19840 16646
rect 19800 16244 19852 16250
rect 19800 16186 19852 16192
rect 19340 15972 19392 15978
rect 19340 15914 19392 15920
rect 19352 15706 19380 15914
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19904 15638 19932 16662
rect 19996 16590 20024 16730
rect 19984 16584 20036 16590
rect 19984 16526 20036 16532
rect 19892 15632 19944 15638
rect 19892 15574 19944 15580
rect 19338 15464 19394 15473
rect 19338 15399 19394 15408
rect 19352 15314 19380 15399
rect 19168 15286 19380 15314
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19168 14618 19196 15286
rect 19449 15260 19745 15280
rect 19505 15258 19529 15260
rect 19585 15258 19609 15260
rect 19665 15258 19689 15260
rect 19527 15206 19529 15258
rect 19591 15206 19603 15258
rect 19665 15206 19667 15258
rect 19505 15204 19529 15206
rect 19585 15204 19609 15206
rect 19665 15204 19689 15206
rect 19449 15184 19745 15204
rect 19340 15088 19392 15094
rect 19338 15056 19340 15065
rect 19392 15056 19394 15065
rect 19338 14991 19394 15000
rect 19248 14952 19300 14958
rect 19616 14952 19668 14958
rect 19248 14894 19300 14900
rect 19614 14920 19616 14929
rect 19668 14920 19670 14929
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 19154 14512 19210 14521
rect 19154 14447 19156 14456
rect 19208 14447 19210 14456
rect 19156 14418 19208 14424
rect 19260 13938 19288 14894
rect 19670 14878 19748 14906
rect 19614 14855 19670 14864
rect 19616 14816 19668 14822
rect 19616 14758 19668 14764
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 19352 14278 19380 14418
rect 19628 14346 19656 14758
rect 19616 14340 19668 14346
rect 19616 14282 19668 14288
rect 19340 14272 19392 14278
rect 19720 14260 19748 14878
rect 19812 14618 19840 15302
rect 19982 15056 20038 15065
rect 19982 14991 20038 15000
rect 19996 14958 20024 14991
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 19982 14784 20038 14793
rect 19982 14719 20038 14728
rect 19800 14612 19852 14618
rect 19800 14554 19852 14560
rect 19996 14550 20024 14719
rect 19984 14544 20036 14550
rect 19984 14486 20036 14492
rect 19984 14340 20036 14346
rect 19984 14282 20036 14288
rect 19720 14232 19840 14260
rect 19340 14214 19392 14220
rect 19449 14172 19745 14192
rect 19505 14170 19529 14172
rect 19585 14170 19609 14172
rect 19665 14170 19689 14172
rect 19527 14118 19529 14170
rect 19591 14118 19603 14170
rect 19665 14118 19667 14170
rect 19505 14116 19529 14118
rect 19585 14116 19609 14118
rect 19665 14116 19689 14118
rect 19449 14096 19745 14116
rect 19616 14000 19668 14006
rect 19616 13942 19668 13948
rect 19248 13932 19300 13938
rect 19248 13874 19300 13880
rect 19156 13864 19208 13870
rect 19156 13806 19208 13812
rect 19062 12064 19118 12073
rect 19062 11999 19118 12008
rect 18970 11928 19026 11937
rect 18970 11863 19026 11872
rect 19168 11778 19196 13806
rect 18984 11750 19196 11778
rect 19260 11762 19288 13874
rect 19340 13796 19392 13802
rect 19340 13738 19392 13744
rect 19352 13433 19380 13738
rect 19628 13530 19656 13942
rect 19812 13938 19840 14232
rect 19800 13932 19852 13938
rect 19852 13892 19932 13920
rect 19800 13874 19852 13880
rect 19616 13524 19668 13530
rect 19616 13466 19668 13472
rect 19338 13424 19394 13433
rect 19338 13359 19394 13368
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19352 12782 19380 13194
rect 19800 13184 19852 13190
rect 19800 13126 19852 13132
rect 19449 13084 19745 13104
rect 19505 13082 19529 13084
rect 19585 13082 19609 13084
rect 19665 13082 19689 13084
rect 19527 13030 19529 13082
rect 19591 13030 19603 13082
rect 19665 13030 19667 13082
rect 19505 13028 19529 13030
rect 19585 13028 19609 13030
rect 19665 13028 19689 13030
rect 19449 13008 19745 13028
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 19708 12708 19760 12714
rect 19708 12650 19760 12656
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19248 11756 19300 11762
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 18800 10220 18920 10248
rect 18696 10202 18748 10208
rect 18892 10130 18920 10220
rect 18788 10124 18840 10130
rect 18788 10066 18840 10072
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18604 9716 18656 9722
rect 18604 9658 18656 9664
rect 18694 9616 18750 9625
rect 18694 9551 18750 9560
rect 18708 9518 18736 9551
rect 18696 9512 18748 9518
rect 18696 9454 18748 9460
rect 18800 9382 18828 10066
rect 18984 9897 19012 11750
rect 19248 11698 19300 11704
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 19076 11218 19104 11630
rect 19352 11558 19380 12242
rect 19720 12186 19748 12650
rect 19812 12306 19840 13126
rect 19904 12889 19932 13892
rect 19890 12880 19946 12889
rect 19890 12815 19946 12824
rect 19996 12730 20024 14282
rect 19904 12702 20024 12730
rect 19904 12374 19932 12702
rect 19984 12640 20036 12646
rect 20088 12617 20116 18158
rect 20180 17649 20208 20198
rect 20364 19854 20392 20402
rect 20442 20360 20498 20369
rect 20442 20295 20498 20304
rect 20456 20262 20484 20295
rect 20444 20256 20496 20262
rect 20444 20198 20496 20204
rect 20824 19922 20852 23920
rect 21088 21344 21140 21350
rect 21088 21286 21140 21292
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 20916 20398 20944 20878
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 20626 19408 20682 19417
rect 20626 19343 20682 19352
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20166 17640 20222 17649
rect 20166 17575 20222 17584
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 20180 17134 20208 17478
rect 20168 17128 20220 17134
rect 20168 17070 20220 17076
rect 20272 16726 20300 19110
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20364 18193 20392 18566
rect 20350 18184 20406 18193
rect 20350 18119 20406 18128
rect 20352 18080 20404 18086
rect 20350 18048 20352 18057
rect 20444 18080 20496 18086
rect 20404 18048 20406 18057
rect 20444 18022 20496 18028
rect 20350 17983 20406 17992
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20260 16720 20312 16726
rect 20260 16662 20312 16668
rect 20260 16448 20312 16454
rect 20260 16390 20312 16396
rect 20168 15904 20220 15910
rect 20168 15846 20220 15852
rect 20180 15706 20208 15846
rect 20168 15700 20220 15706
rect 20168 15642 20220 15648
rect 20168 15564 20220 15570
rect 20168 15506 20220 15512
rect 20180 15026 20208 15506
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 20168 13456 20220 13462
rect 20168 13398 20220 13404
rect 20180 12782 20208 13398
rect 20168 12776 20220 12782
rect 20168 12718 20220 12724
rect 19984 12582 20036 12588
rect 20074 12608 20130 12617
rect 19892 12368 19944 12374
rect 19892 12310 19944 12316
rect 19800 12300 19852 12306
rect 19800 12242 19852 12248
rect 19996 12238 20024 12582
rect 20074 12543 20130 12552
rect 20074 12472 20130 12481
rect 20272 12458 20300 16390
rect 20364 13394 20392 17614
rect 20456 17338 20484 18022
rect 20536 17740 20588 17746
rect 20536 17682 20588 17688
rect 20444 17332 20496 17338
rect 20444 17274 20496 17280
rect 20444 15156 20496 15162
rect 20444 15098 20496 15104
rect 20456 14113 20484 15098
rect 20442 14104 20498 14113
rect 20442 14039 20498 14048
rect 20352 13388 20404 13394
rect 20352 13330 20404 13336
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20074 12407 20130 12416
rect 20180 12430 20300 12458
rect 19892 12232 19944 12238
rect 19720 12158 19840 12186
rect 19892 12174 19944 12180
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 19449 11996 19745 12016
rect 19505 11994 19529 11996
rect 19585 11994 19609 11996
rect 19665 11994 19689 11996
rect 19527 11942 19529 11994
rect 19591 11942 19603 11994
rect 19665 11942 19667 11994
rect 19505 11940 19529 11942
rect 19585 11940 19609 11942
rect 19665 11940 19689 11942
rect 19449 11920 19745 11940
rect 19706 11792 19762 11801
rect 19706 11727 19708 11736
rect 19760 11727 19762 11736
rect 19708 11698 19760 11704
rect 19340 11552 19392 11558
rect 19154 11520 19210 11529
rect 19340 11494 19392 11500
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19154 11455 19210 11464
rect 19064 11212 19116 11218
rect 19064 11154 19116 11160
rect 19062 11112 19118 11121
rect 19062 11047 19118 11056
rect 19076 10742 19104 11047
rect 19064 10736 19116 10742
rect 19064 10678 19116 10684
rect 19168 10606 19196 11455
rect 19444 11354 19472 11494
rect 19432 11348 19484 11354
rect 19260 11308 19432 11336
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19260 10112 19288 11308
rect 19432 11290 19484 11296
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19076 10084 19288 10112
rect 18970 9888 19026 9897
rect 18970 9823 19026 9832
rect 19076 9602 19104 10084
rect 19352 10010 19380 11154
rect 19449 10908 19745 10928
rect 19505 10906 19529 10908
rect 19585 10906 19609 10908
rect 19665 10906 19689 10908
rect 19527 10854 19529 10906
rect 19591 10854 19603 10906
rect 19665 10854 19667 10906
rect 19505 10852 19529 10854
rect 19585 10852 19609 10854
rect 19665 10852 19689 10854
rect 19449 10832 19745 10852
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19720 10062 19748 10542
rect 19812 10538 19840 12158
rect 19904 11694 19932 12174
rect 19892 11688 19944 11694
rect 19892 11630 19944 11636
rect 19904 11354 19932 11630
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 19996 10606 20024 12174
rect 20088 11558 20116 12407
rect 20180 12322 20208 12430
rect 20180 12294 20300 12322
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 20074 11384 20130 11393
rect 20074 11319 20130 11328
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19800 10532 19852 10538
rect 19800 10474 19852 10480
rect 19800 10192 19852 10198
rect 19800 10134 19852 10140
rect 19708 10056 19760 10062
rect 18984 9574 19104 9602
rect 19260 9982 19380 10010
rect 19706 10024 19708 10033
rect 19760 10024 19762 10033
rect 19156 9580 19208 9586
rect 18984 9518 19012 9574
rect 19260 9568 19288 9982
rect 19706 9959 19762 9968
rect 19720 9933 19748 9959
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19352 9625 19380 9862
rect 19449 9820 19745 9840
rect 19505 9818 19529 9820
rect 19585 9818 19609 9820
rect 19665 9818 19689 9820
rect 19527 9766 19529 9818
rect 19591 9766 19603 9818
rect 19665 9766 19667 9818
rect 19505 9764 19529 9766
rect 19585 9764 19609 9766
rect 19665 9764 19689 9766
rect 19449 9744 19745 9764
rect 19208 9540 19288 9568
rect 19338 9616 19394 9625
rect 19338 9551 19394 9560
rect 19708 9580 19760 9586
rect 19156 9522 19208 9528
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 18510 9208 18566 9217
rect 18510 9143 18566 9152
rect 18524 8974 18552 9143
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18616 8634 18644 9318
rect 18696 9036 18748 9042
rect 18696 8978 18748 8984
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18512 7948 18564 7954
rect 18432 7908 18512 7936
rect 18512 7890 18564 7896
rect 18328 7744 18380 7750
rect 18604 7744 18656 7750
rect 18328 7686 18380 7692
rect 18602 7712 18604 7721
rect 18656 7712 18658 7721
rect 18050 7440 18106 7449
rect 18050 7375 18106 7384
rect 18340 6254 18368 7686
rect 18602 7647 18658 7656
rect 18418 7440 18474 7449
rect 18418 7375 18420 7384
rect 18472 7375 18474 7384
rect 18420 7346 18472 7352
rect 18708 7206 18736 8978
rect 18800 8498 18828 9318
rect 18878 9072 18934 9081
rect 18984 9042 19012 9454
rect 19064 9444 19116 9450
rect 19064 9386 19116 9392
rect 19076 9081 19104 9386
rect 19154 9344 19210 9353
rect 19154 9279 19210 9288
rect 19062 9072 19118 9081
rect 18878 9007 18934 9016
rect 18972 9036 19024 9042
rect 18892 8974 18920 9007
rect 19168 9042 19196 9279
rect 19260 9217 19288 9540
rect 19708 9522 19760 9528
rect 19720 9489 19748 9522
rect 19706 9480 19762 9489
rect 19706 9415 19762 9424
rect 19246 9208 19302 9217
rect 19246 9143 19302 9152
rect 19062 9007 19118 9016
rect 19156 9036 19208 9042
rect 18972 8978 19024 8984
rect 19156 8978 19208 8984
rect 18880 8968 18932 8974
rect 18880 8910 18932 8916
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 19338 8936 19394 8945
rect 18878 8664 18934 8673
rect 18878 8599 18934 8608
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18892 7018 18920 8599
rect 19076 8362 19104 8910
rect 19338 8871 19394 8880
rect 19246 8800 19302 8809
rect 19246 8735 19302 8744
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 19064 8356 19116 8362
rect 19064 8298 19116 8304
rect 19168 8090 19196 8366
rect 19156 8084 19208 8090
rect 19156 8026 19208 8032
rect 19156 7880 19208 7886
rect 19156 7822 19208 7828
rect 19168 7546 19196 7822
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19168 7410 19196 7482
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19260 7313 19288 8735
rect 19246 7304 19302 7313
rect 19246 7239 19302 7248
rect 18432 6990 18920 7018
rect 18236 6248 18288 6254
rect 18236 6190 18288 6196
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 18144 6180 18196 6186
rect 18144 6122 18196 6128
rect 18156 5234 18184 6122
rect 18248 5370 18276 6190
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 18248 4826 18276 5306
rect 18328 5092 18380 5098
rect 18328 5034 18380 5040
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 18052 4752 18104 4758
rect 18052 4694 18104 4700
rect 18064 4282 18092 4694
rect 18052 4276 18104 4282
rect 18052 4218 18104 4224
rect 18340 3890 18368 5034
rect 18432 4185 18460 6990
rect 18880 6928 18932 6934
rect 18880 6870 18932 6876
rect 19064 6928 19116 6934
rect 19064 6870 19116 6876
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 18524 5914 18552 6802
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18708 6118 18736 6598
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18616 5914 18644 6054
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18800 5642 18828 6734
rect 18892 6730 18920 6870
rect 18880 6724 18932 6730
rect 18880 6666 18932 6672
rect 18788 5636 18840 5642
rect 18788 5578 18840 5584
rect 18880 4548 18932 4554
rect 18880 4490 18932 4496
rect 18418 4176 18474 4185
rect 18892 4146 18920 4490
rect 19076 4146 19104 6870
rect 19156 6724 19208 6730
rect 19156 6666 19208 6672
rect 19168 6186 19196 6666
rect 19352 6202 19380 8871
rect 19449 8732 19745 8752
rect 19505 8730 19529 8732
rect 19585 8730 19609 8732
rect 19665 8730 19689 8732
rect 19527 8678 19529 8730
rect 19591 8678 19603 8730
rect 19665 8678 19667 8730
rect 19505 8676 19529 8678
rect 19585 8676 19609 8678
rect 19665 8676 19689 8678
rect 19449 8656 19745 8676
rect 19812 8430 19840 10134
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19904 9081 19932 9522
rect 19890 9072 19946 9081
rect 19890 9007 19946 9016
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19800 8424 19852 8430
rect 19800 8366 19852 8372
rect 19444 8090 19472 8366
rect 19892 8356 19944 8362
rect 19892 8298 19944 8304
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19800 8084 19852 8090
rect 19800 8026 19852 8032
rect 19449 7644 19745 7664
rect 19505 7642 19529 7644
rect 19585 7642 19609 7644
rect 19665 7642 19689 7644
rect 19527 7590 19529 7642
rect 19591 7590 19603 7642
rect 19665 7590 19667 7642
rect 19505 7588 19529 7590
rect 19585 7588 19609 7590
rect 19665 7588 19689 7590
rect 19449 7568 19745 7588
rect 19449 6556 19745 6576
rect 19505 6554 19529 6556
rect 19585 6554 19609 6556
rect 19665 6554 19689 6556
rect 19527 6502 19529 6554
rect 19591 6502 19603 6554
rect 19665 6502 19667 6554
rect 19505 6500 19529 6502
rect 19585 6500 19609 6502
rect 19665 6500 19689 6502
rect 19449 6480 19745 6500
rect 19156 6180 19208 6186
rect 19156 6122 19208 6128
rect 19260 6174 19380 6202
rect 19154 5672 19210 5681
rect 19154 5607 19210 5616
rect 19168 5234 19196 5607
rect 19156 5228 19208 5234
rect 19156 5170 19208 5176
rect 19260 4321 19288 6174
rect 19812 6118 19840 8026
rect 19904 7546 19932 8298
rect 19996 8294 20024 10066
rect 19984 8288 20036 8294
rect 19984 8230 20036 8236
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 19892 7540 19944 7546
rect 19892 7482 19944 7488
rect 19996 7002 20024 7890
rect 19984 6996 20036 7002
rect 19984 6938 20036 6944
rect 20088 6882 20116 11319
rect 20180 10044 20208 12174
rect 20272 11354 20300 12294
rect 20364 11801 20392 12582
rect 20548 12481 20576 17682
rect 20640 12986 20668 19343
rect 20916 19310 20944 20334
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20732 16658 20760 18226
rect 20812 18216 20864 18222
rect 20812 18158 20864 18164
rect 20824 17678 20852 18158
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20824 17134 20852 17614
rect 20812 17128 20864 17134
rect 20812 17070 20864 17076
rect 20824 16726 20852 17070
rect 20812 16720 20864 16726
rect 20812 16662 20864 16668
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 20732 16046 20760 16594
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 20916 16046 20944 16526
rect 20994 16144 21050 16153
rect 20994 16079 21050 16088
rect 20720 16040 20772 16046
rect 20720 15982 20772 15988
rect 20904 16040 20956 16046
rect 20904 15982 20956 15988
rect 20904 15904 20956 15910
rect 20904 15846 20956 15852
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 20732 15162 20760 15642
rect 20916 15502 20944 15846
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20732 14074 20760 14894
rect 20810 14648 20866 14657
rect 20810 14583 20866 14592
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20628 12980 20680 12986
rect 20628 12922 20680 12928
rect 20534 12472 20590 12481
rect 20534 12407 20590 12416
rect 20444 12368 20496 12374
rect 20444 12310 20496 12316
rect 20350 11792 20406 11801
rect 20350 11727 20406 11736
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20260 11212 20312 11218
rect 20260 11154 20312 11160
rect 20272 10169 20300 11154
rect 20352 11076 20404 11082
rect 20352 11018 20404 11024
rect 20258 10160 20314 10169
rect 20258 10095 20314 10104
rect 20180 10016 20300 10044
rect 20166 9072 20222 9081
rect 20166 9007 20222 9016
rect 20180 8906 20208 9007
rect 20168 8900 20220 8906
rect 20168 8842 20220 8848
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 19904 6854 20116 6882
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19800 6112 19852 6118
rect 19800 6054 19852 6060
rect 19352 5574 19380 6054
rect 19800 5704 19852 5710
rect 19800 5646 19852 5652
rect 19812 5574 19840 5646
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19800 5568 19852 5574
rect 19800 5510 19852 5516
rect 19449 5468 19745 5488
rect 19505 5466 19529 5468
rect 19585 5466 19609 5468
rect 19665 5466 19689 5468
rect 19527 5414 19529 5466
rect 19591 5414 19603 5466
rect 19665 5414 19667 5466
rect 19505 5412 19529 5414
rect 19585 5412 19609 5414
rect 19665 5412 19689 5414
rect 19449 5392 19745 5412
rect 19432 5160 19484 5166
rect 19430 5128 19432 5137
rect 19484 5128 19486 5137
rect 19340 5092 19392 5098
rect 19430 5063 19486 5072
rect 19340 5034 19392 5040
rect 19246 4312 19302 4321
rect 19246 4247 19302 4256
rect 18418 4111 18474 4120
rect 18880 4140 18932 4146
rect 18880 4082 18932 4088
rect 19064 4140 19116 4146
rect 19064 4082 19116 4088
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 18248 3862 18368 3890
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 17958 3632 18014 3641
rect 17958 3567 18014 3576
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 18156 2922 18184 3470
rect 18144 2916 18196 2922
rect 18144 2858 18196 2864
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 18064 2446 18092 2790
rect 18156 2514 18184 2858
rect 18144 2508 18196 2514
rect 18144 2450 18196 2456
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 17868 2304 17920 2310
rect 17868 2246 17920 2252
rect 17500 1964 17552 1970
rect 17500 1906 17552 1912
rect 18248 1902 18276 3862
rect 18524 3602 18552 3878
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 18512 3596 18564 3602
rect 18512 3538 18564 3544
rect 18420 3460 18472 3466
rect 18420 3402 18472 3408
rect 18328 2916 18380 2922
rect 18328 2858 18380 2864
rect 18340 2650 18368 2858
rect 18328 2644 18380 2650
rect 18328 2586 18380 2592
rect 18340 2553 18368 2586
rect 18432 2582 18460 3402
rect 18616 2582 18644 3674
rect 18984 3534 19012 4014
rect 19156 4004 19208 4010
rect 19156 3946 19208 3952
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 19168 3398 19196 3946
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19156 3392 19208 3398
rect 19156 3334 19208 3340
rect 19260 3194 19288 3538
rect 19156 3188 19208 3194
rect 19156 3130 19208 3136
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 18420 2576 18472 2582
rect 18326 2544 18382 2553
rect 18420 2518 18472 2524
rect 18604 2576 18656 2582
rect 18604 2518 18656 2524
rect 18326 2479 18382 2488
rect 18236 1896 18288 1902
rect 18236 1838 18288 1844
rect 19168 1442 19196 3130
rect 19260 2106 19288 3130
rect 19352 2514 19380 5034
rect 19812 4690 19840 5510
rect 19904 4865 19932 6854
rect 20074 6760 20130 6769
rect 20180 6730 20208 7822
rect 20272 7449 20300 10016
rect 20258 7440 20314 7449
rect 20258 7375 20314 7384
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 20074 6695 20130 6704
rect 20168 6724 20220 6730
rect 20088 6610 20116 6695
rect 20168 6666 20220 6672
rect 20088 6582 20208 6610
rect 20076 5772 20128 5778
rect 20076 5714 20128 5720
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19890 4856 19946 4865
rect 19890 4791 19946 4800
rect 19800 4684 19852 4690
rect 19800 4626 19852 4632
rect 19449 4380 19745 4400
rect 19505 4378 19529 4380
rect 19585 4378 19609 4380
rect 19665 4378 19689 4380
rect 19527 4326 19529 4378
rect 19591 4326 19603 4378
rect 19665 4326 19667 4378
rect 19505 4324 19529 4326
rect 19585 4324 19609 4326
rect 19665 4324 19689 4326
rect 19449 4304 19745 4324
rect 19449 3292 19745 3312
rect 19505 3290 19529 3292
rect 19585 3290 19609 3292
rect 19665 3290 19689 3292
rect 19527 3238 19529 3290
rect 19591 3238 19603 3290
rect 19665 3238 19667 3290
rect 19505 3236 19529 3238
rect 19585 3236 19609 3238
rect 19665 3236 19689 3238
rect 19449 3216 19745 3236
rect 19996 2650 20024 5510
rect 20088 5370 20116 5714
rect 20076 5364 20128 5370
rect 20076 5306 20128 5312
rect 20074 5264 20130 5273
rect 20074 5199 20130 5208
rect 20088 4622 20116 5199
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 20088 2854 20116 4558
rect 20180 4321 20208 6582
rect 20272 5574 20300 7278
rect 20364 5710 20392 11018
rect 20456 10198 20484 12310
rect 20824 11914 20852 14583
rect 20916 14328 20944 15438
rect 21008 14521 21036 16079
rect 20994 14512 21050 14521
rect 20994 14447 21050 14456
rect 20996 14340 21048 14346
rect 20916 14300 20996 14328
rect 20996 14282 21048 14288
rect 21008 13734 21036 14282
rect 20996 13728 21048 13734
rect 20996 13670 21048 13676
rect 21008 13326 21036 13670
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 20904 12844 20956 12850
rect 20904 12786 20956 12792
rect 20548 11886 20852 11914
rect 20916 11898 20944 12786
rect 21008 12714 21036 13262
rect 20996 12708 21048 12714
rect 20996 12650 21048 12656
rect 21008 12306 21036 12650
rect 20996 12300 21048 12306
rect 20996 12242 21048 12248
rect 20904 11892 20956 11898
rect 20548 10470 20576 11886
rect 20904 11834 20956 11840
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20626 10704 20682 10713
rect 20626 10639 20682 10648
rect 20536 10464 20588 10470
rect 20536 10406 20588 10412
rect 20444 10192 20496 10198
rect 20444 10134 20496 10140
rect 20444 8356 20496 8362
rect 20444 8298 20496 8304
rect 20456 6866 20484 8298
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20444 6656 20496 6662
rect 20444 6598 20496 6604
rect 20456 6322 20484 6598
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20352 5704 20404 5710
rect 20350 5672 20352 5681
rect 20444 5704 20496 5710
rect 20404 5672 20406 5681
rect 20444 5646 20496 5652
rect 20350 5607 20406 5616
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 20272 4554 20300 5170
rect 20456 4758 20484 5646
rect 20444 4752 20496 4758
rect 20444 4694 20496 4700
rect 20260 4548 20312 4554
rect 20260 4490 20312 4496
rect 20166 4312 20222 4321
rect 20166 4247 20222 4256
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20364 3602 20392 4014
rect 20548 3641 20576 10406
rect 20640 9994 20668 10639
rect 20732 10062 20760 11086
rect 20810 10840 20866 10849
rect 20810 10775 20866 10784
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20628 9988 20680 9994
rect 20628 9930 20680 9936
rect 20732 9586 20760 9998
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20732 8974 20760 9522
rect 20720 8968 20772 8974
rect 20720 8910 20772 8916
rect 20732 8430 20760 8910
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20628 8016 20680 8022
rect 20628 7958 20680 7964
rect 20640 7342 20668 7958
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 20732 7449 20760 7482
rect 20718 7440 20774 7449
rect 20718 7375 20774 7384
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20720 7268 20772 7274
rect 20720 7210 20772 7216
rect 20626 7168 20682 7177
rect 20626 7103 20682 7112
rect 20534 3632 20590 3641
rect 20352 3596 20404 3602
rect 20534 3567 20590 3576
rect 20352 3538 20404 3544
rect 20364 3126 20392 3538
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 20352 3120 20404 3126
rect 20352 3062 20404 3068
rect 20076 2848 20128 2854
rect 20076 2790 20128 2796
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 20364 2514 20392 3062
rect 20456 3058 20484 3334
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 20640 2650 20668 7103
rect 20732 6390 20760 7210
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 20824 6254 20852 10775
rect 20904 9920 20956 9926
rect 20904 9862 20956 9868
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 20720 5840 20772 5846
rect 20720 5782 20772 5788
rect 20732 5302 20760 5782
rect 20720 5296 20772 5302
rect 20720 5238 20772 5244
rect 20916 5234 20944 9862
rect 20994 7984 21050 7993
rect 20994 7919 20996 7928
rect 21048 7919 21050 7928
rect 20996 7890 21048 7896
rect 21008 7585 21036 7890
rect 20994 7576 21050 7585
rect 20994 7511 21050 7520
rect 21100 7290 21128 21286
rect 21468 20330 21496 23920
rect 21916 21616 21968 21622
rect 21916 21558 21968 21564
rect 21824 21548 21876 21554
rect 21824 21490 21876 21496
rect 21548 21344 21600 21350
rect 21548 21286 21600 21292
rect 21640 21344 21692 21350
rect 21640 21286 21692 21292
rect 21560 20806 21588 21286
rect 21652 21078 21680 21286
rect 21640 21072 21692 21078
rect 21640 21014 21692 21020
rect 21548 20800 21600 20806
rect 21548 20742 21600 20748
rect 21560 20398 21588 20742
rect 21836 20602 21864 21490
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 21548 20392 21600 20398
rect 21548 20334 21600 20340
rect 21456 20324 21508 20330
rect 21456 20266 21508 20272
rect 21732 20256 21784 20262
rect 21732 20198 21784 20204
rect 21640 19916 21692 19922
rect 21640 19858 21692 19864
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21284 18766 21312 19110
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 21284 18222 21312 18702
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 21192 17814 21220 18022
rect 21180 17808 21232 17814
rect 21180 17750 21232 17756
rect 21192 17338 21220 17750
rect 21180 17332 21232 17338
rect 21180 17274 21232 17280
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21284 15638 21312 15846
rect 21272 15632 21324 15638
rect 21272 15574 21324 15580
rect 21376 13716 21404 19654
rect 21652 19174 21680 19858
rect 21744 19854 21772 20198
rect 21836 19854 21864 20538
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 21824 19848 21876 19854
rect 21824 19790 21876 19796
rect 21744 19310 21772 19790
rect 21732 19304 21784 19310
rect 21732 19246 21784 19252
rect 21640 19168 21692 19174
rect 21640 19110 21692 19116
rect 21652 18902 21680 19110
rect 21640 18896 21692 18902
rect 21640 18838 21692 18844
rect 21548 17536 21600 17542
rect 21548 17478 21600 17484
rect 21560 16250 21588 17478
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 21652 16726 21680 17002
rect 21824 16992 21876 16998
rect 21824 16934 21876 16940
rect 21640 16720 21692 16726
rect 21640 16662 21692 16668
rect 21548 16244 21600 16250
rect 21600 16204 21772 16232
rect 21548 16186 21600 16192
rect 21640 15564 21692 15570
rect 21640 15506 21692 15512
rect 21548 15360 21600 15366
rect 21548 15302 21600 15308
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21468 13870 21496 14758
rect 21560 14550 21588 15302
rect 21652 14618 21680 15506
rect 21744 14958 21772 16204
rect 21836 15978 21864 16934
rect 21824 15972 21876 15978
rect 21824 15914 21876 15920
rect 21928 15144 21956 21558
rect 22008 19916 22060 19922
rect 22008 19858 22060 19864
rect 22020 18737 22048 19858
rect 22112 18834 22140 23920
rect 22192 21480 22244 21486
rect 22192 21422 22244 21428
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 22006 18728 22062 18737
rect 22006 18663 22062 18672
rect 22204 18057 22232 21422
rect 22284 21344 22336 21350
rect 22284 21286 22336 21292
rect 22190 18048 22246 18057
rect 22190 17983 22246 17992
rect 22008 17536 22060 17542
rect 22008 17478 22060 17484
rect 22020 17134 22048 17478
rect 22008 17128 22060 17134
rect 22008 17070 22060 17076
rect 22020 16114 22048 17070
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 21836 15116 21956 15144
rect 21732 14952 21784 14958
rect 21732 14894 21784 14900
rect 21732 14816 21784 14822
rect 21732 14758 21784 14764
rect 21640 14612 21692 14618
rect 21640 14554 21692 14560
rect 21548 14544 21600 14550
rect 21548 14486 21600 14492
rect 21456 13864 21508 13870
rect 21456 13806 21508 13812
rect 21744 13802 21772 14758
rect 21732 13796 21784 13802
rect 21732 13738 21784 13744
rect 21376 13688 21496 13716
rect 21468 12356 21496 13688
rect 21744 12850 21772 13738
rect 21732 12844 21784 12850
rect 21732 12786 21784 12792
rect 21836 12458 21864 15116
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 21928 14278 21956 14962
rect 21916 14272 21968 14278
rect 21916 14214 21968 14220
rect 21928 13462 21956 14214
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22112 13530 22140 13670
rect 22100 13524 22152 13530
rect 22100 13466 22152 13472
rect 21916 13456 21968 13462
rect 21916 13398 21968 13404
rect 22192 12912 22244 12918
rect 22192 12854 22244 12860
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 21744 12430 21864 12458
rect 21744 12356 21772 12430
rect 21468 12328 21588 12356
rect 21744 12328 21956 12356
rect 21180 12300 21232 12306
rect 21180 12242 21232 12248
rect 21192 10810 21220 12242
rect 21272 11688 21324 11694
rect 21272 11630 21324 11636
rect 21284 11150 21312 11630
rect 21272 11144 21324 11150
rect 21272 11086 21324 11092
rect 21180 10804 21232 10810
rect 21180 10746 21232 10752
rect 21454 10568 21510 10577
rect 21454 10503 21510 10512
rect 21468 10470 21496 10503
rect 21456 10464 21508 10470
rect 21456 10406 21508 10412
rect 21272 10124 21324 10130
rect 21272 10066 21324 10072
rect 21284 9489 21312 10066
rect 21270 9480 21326 9489
rect 21270 9415 21326 9424
rect 21364 8424 21416 8430
rect 21364 8366 21416 8372
rect 21270 8256 21326 8265
rect 21270 8191 21326 8200
rect 21284 8022 21312 8191
rect 21272 8016 21324 8022
rect 21272 7958 21324 7964
rect 21100 7262 21312 7290
rect 20996 7200 21048 7206
rect 20996 7142 21048 7148
rect 21088 7200 21140 7206
rect 21088 7142 21140 7148
rect 21008 7002 21036 7142
rect 20996 6996 21048 7002
rect 20996 6938 21048 6944
rect 21100 6934 21128 7142
rect 21088 6928 21140 6934
rect 21088 6870 21140 6876
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 21008 6361 21036 6802
rect 20994 6352 21050 6361
rect 20994 6287 21050 6296
rect 20904 5228 20956 5234
rect 20904 5170 20956 5176
rect 20720 5160 20772 5166
rect 20718 5128 20720 5137
rect 20772 5128 20774 5137
rect 20718 5063 20774 5072
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 20824 3738 20852 4422
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 21008 3670 21036 4082
rect 20996 3664 21048 3670
rect 20996 3606 21048 3612
rect 20904 2916 20956 2922
rect 20904 2858 20956 2864
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 20916 2582 20944 2858
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 19340 2508 19392 2514
rect 19340 2450 19392 2456
rect 20352 2508 20404 2514
rect 20352 2450 20404 2456
rect 19890 2272 19946 2281
rect 19449 2204 19745 2224
rect 19890 2207 19946 2216
rect 19505 2202 19529 2204
rect 19585 2202 19609 2204
rect 19665 2202 19689 2204
rect 19527 2150 19529 2202
rect 19591 2150 19603 2202
rect 19665 2150 19667 2202
rect 19505 2148 19529 2150
rect 19585 2148 19609 2150
rect 19665 2148 19689 2150
rect 19449 2128 19745 2148
rect 19248 2100 19300 2106
rect 19248 2042 19300 2048
rect 19904 1834 19932 2207
rect 20916 2038 20944 2518
rect 21100 2446 21128 6870
rect 21180 6248 21232 6254
rect 21180 6190 21232 6196
rect 21192 5166 21220 6190
rect 21180 5160 21232 5166
rect 21180 5102 21232 5108
rect 21192 4690 21220 5102
rect 21180 4684 21232 4690
rect 21180 4626 21232 4632
rect 21192 4078 21220 4626
rect 21284 4146 21312 7262
rect 21376 5273 21404 8366
rect 21454 7576 21510 7585
rect 21454 7511 21510 7520
rect 21362 5264 21418 5273
rect 21362 5199 21418 5208
rect 21364 4684 21416 4690
rect 21364 4626 21416 4632
rect 21272 4140 21324 4146
rect 21272 4082 21324 4088
rect 21180 4072 21232 4078
rect 21180 4014 21232 4020
rect 21376 3942 21404 4626
rect 21272 3936 21324 3942
rect 21272 3878 21324 3884
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 21284 2514 21312 3878
rect 21468 2990 21496 7511
rect 21560 3398 21588 12328
rect 21730 12200 21786 12209
rect 21730 12135 21786 12144
rect 21640 12096 21692 12102
rect 21640 12038 21692 12044
rect 21652 10606 21680 12038
rect 21640 10600 21692 10606
rect 21640 10542 21692 10548
rect 21744 10266 21772 12135
rect 21824 12096 21876 12102
rect 21824 12038 21876 12044
rect 21836 11286 21864 12038
rect 21824 11280 21876 11286
rect 21824 11222 21876 11228
rect 21732 10260 21784 10266
rect 21732 10202 21784 10208
rect 21732 9920 21784 9926
rect 21732 9862 21784 9868
rect 21640 5772 21692 5778
rect 21640 5714 21692 5720
rect 21652 4078 21680 5714
rect 21640 4072 21692 4078
rect 21640 4014 21692 4020
rect 21652 3738 21680 4014
rect 21640 3732 21692 3738
rect 21640 3674 21692 3680
rect 21548 3392 21600 3398
rect 21548 3334 21600 3340
rect 21456 2984 21508 2990
rect 21744 2961 21772 9862
rect 21824 6180 21876 6186
rect 21824 6122 21876 6128
rect 21836 5370 21864 6122
rect 21824 5364 21876 5370
rect 21824 5306 21876 5312
rect 21928 4468 21956 12328
rect 22020 12102 22048 12786
rect 22008 12096 22060 12102
rect 22008 12038 22060 12044
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22112 9330 22140 11290
rect 22204 11234 22232 12854
rect 22296 11354 22324 21286
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22468 19916 22520 19922
rect 22468 19858 22520 19864
rect 22480 18970 22508 19858
rect 22468 18964 22520 18970
rect 22468 18906 22520 18912
rect 22480 18222 22508 18906
rect 22468 18216 22520 18222
rect 22468 18158 22520 18164
rect 22376 18148 22428 18154
rect 22376 18090 22428 18096
rect 22388 16114 22416 18090
rect 22572 17377 22600 20334
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 22664 17882 22692 19654
rect 22652 17876 22704 17882
rect 22652 17818 22704 17824
rect 22558 17368 22614 17377
rect 22558 17303 22614 17312
rect 22468 17128 22520 17134
rect 22468 17070 22520 17076
rect 22480 16697 22508 17070
rect 22652 16992 22704 16998
rect 22652 16934 22704 16940
rect 22664 16794 22692 16934
rect 22652 16788 22704 16794
rect 22652 16730 22704 16736
rect 22466 16688 22522 16697
rect 22466 16623 22522 16632
rect 22756 16182 22784 23920
rect 22928 20256 22980 20262
rect 22928 20198 22980 20204
rect 22744 16176 22796 16182
rect 22744 16118 22796 16124
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22836 13932 22888 13938
rect 22836 13874 22888 13880
rect 22848 13190 22876 13874
rect 22836 13184 22888 13190
rect 22836 13126 22888 13132
rect 22374 12744 22430 12753
rect 22374 12679 22430 12688
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22204 11206 22324 11234
rect 22296 10266 22324 11206
rect 22388 10606 22416 12679
rect 22744 12640 22796 12646
rect 22744 12582 22796 12588
rect 22560 12232 22612 12238
rect 22560 12174 22612 12180
rect 22376 10600 22428 10606
rect 22376 10542 22428 10548
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22112 9302 22416 9330
rect 22284 9172 22336 9178
rect 22284 9114 22336 9120
rect 22100 9036 22152 9042
rect 22100 8978 22152 8984
rect 22112 8634 22140 8978
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 22100 8628 22152 8634
rect 22100 8570 22152 8576
rect 22204 8090 22232 8774
rect 22192 8084 22244 8090
rect 22192 8026 22244 8032
rect 22192 7948 22244 7954
rect 22192 7890 22244 7896
rect 22100 5704 22152 5710
rect 22100 5646 22152 5652
rect 22112 5273 22140 5646
rect 22098 5264 22154 5273
rect 22098 5199 22154 5208
rect 22100 5092 22152 5098
rect 22100 5034 22152 5040
rect 22112 4826 22140 5034
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 22204 4706 22232 7890
rect 22296 6866 22324 9114
rect 22284 6860 22336 6866
rect 22284 6802 22336 6808
rect 22284 5772 22336 5778
rect 22284 5714 22336 5720
rect 21836 4440 21956 4468
rect 22112 4678 22232 4706
rect 21836 3097 21864 4440
rect 22008 4276 22060 4282
rect 22008 4218 22060 4224
rect 22020 4185 22048 4218
rect 22006 4176 22062 4185
rect 22006 4111 22062 4120
rect 21822 3088 21878 3097
rect 21822 3023 21878 3032
rect 21456 2926 21508 2932
rect 21730 2952 21786 2961
rect 21730 2887 21786 2896
rect 21272 2508 21324 2514
rect 21272 2450 21324 2456
rect 21088 2440 21140 2446
rect 21088 2382 21140 2388
rect 20904 2032 20956 2038
rect 20904 1974 20956 1980
rect 21284 1970 21312 2450
rect 21272 1964 21324 1970
rect 21272 1906 21324 1912
rect 19892 1828 19944 1834
rect 19892 1770 19944 1776
rect 22112 1601 22140 4678
rect 22296 3670 22324 5714
rect 22388 4185 22416 9302
rect 22466 8800 22522 8809
rect 22466 8735 22522 8744
rect 22480 8430 22508 8735
rect 22468 8424 22520 8430
rect 22468 8366 22520 8372
rect 22572 8022 22600 12174
rect 22652 11620 22704 11626
rect 22652 11562 22704 11568
rect 22664 11354 22692 11562
rect 22652 11348 22704 11354
rect 22652 11290 22704 11296
rect 22664 10062 22692 11290
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22652 9444 22704 9450
rect 22652 9386 22704 9392
rect 22664 9178 22692 9386
rect 22652 9172 22704 9178
rect 22652 9114 22704 9120
rect 22560 8016 22612 8022
rect 22560 7958 22612 7964
rect 22664 7886 22692 9114
rect 22652 7880 22704 7886
rect 22652 7822 22704 7828
rect 22756 7426 22784 12582
rect 22664 7398 22784 7426
rect 22468 7268 22520 7274
rect 22468 7210 22520 7216
rect 22480 6225 22508 7210
rect 22466 6216 22522 6225
rect 22466 6151 22522 6160
rect 22664 6118 22692 7398
rect 22744 7336 22796 7342
rect 22744 7278 22796 7284
rect 22756 6905 22784 7278
rect 22742 6896 22798 6905
rect 22742 6831 22798 6840
rect 22652 6112 22704 6118
rect 22652 6054 22704 6060
rect 22744 6112 22796 6118
rect 22744 6054 22796 6060
rect 22374 4176 22430 4185
rect 22374 4111 22430 4120
rect 22284 3664 22336 3670
rect 22284 3606 22336 3612
rect 22296 3194 22324 3606
rect 22284 3188 22336 3194
rect 22284 3130 22336 3136
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 22098 1592 22154 1601
rect 22098 1527 22154 1536
rect 19076 1414 19196 1442
rect 16396 1352 16448 1358
rect 16396 1294 16448 1300
rect 19076 480 19104 1414
rect 19340 1352 19392 1358
rect 19340 1294 19392 1300
rect 19352 921 19380 1294
rect 19338 912 19394 921
rect 19338 847 19394 856
rect 22572 480 22600 2790
rect 1674 0 1730 480
rect 5078 0 5134 480
rect 8574 0 8630 480
rect 12070 0 12126 480
rect 15566 0 15622 480
rect 19062 0 19118 480
rect 22558 0 22614 480
rect 22664 377 22692 6054
rect 22756 5574 22784 6054
rect 22744 5568 22796 5574
rect 22848 5545 22876 13126
rect 22940 6730 22968 20198
rect 23020 14952 23072 14958
rect 23020 14894 23072 14900
rect 23032 7750 23060 14894
rect 23400 11121 23428 23920
rect 24044 20330 24072 23920
rect 24032 20324 24084 20330
rect 24032 20266 24084 20272
rect 23386 11112 23442 11121
rect 23386 11047 23442 11056
rect 23020 7744 23072 7750
rect 23020 7686 23072 7692
rect 22928 6724 22980 6730
rect 22928 6666 22980 6672
rect 22744 5510 22796 5516
rect 22834 5536 22890 5545
rect 22834 5471 22890 5480
rect 22650 368 22706 377
rect 22650 303 22706 312
<< via2 >>
rect 19798 23976 19854 24032
rect 1490 18264 1546 18320
rect 1674 13388 1730 13424
rect 1674 13368 1676 13388
rect 1676 13368 1728 13388
rect 1728 13368 1730 13388
rect 1858 13776 1914 13832
rect 1490 9016 1546 9072
rect 2778 19216 2834 19272
rect 2686 17720 2742 17776
rect 2502 15544 2558 15600
rect 2410 15408 2466 15464
rect 4654 21786 4710 21788
rect 4734 21786 4790 21788
rect 4814 21786 4870 21788
rect 4894 21786 4950 21788
rect 4654 21734 4680 21786
rect 4680 21734 4710 21786
rect 4734 21734 4744 21786
rect 4744 21734 4790 21786
rect 4814 21734 4860 21786
rect 4860 21734 4870 21786
rect 4894 21734 4924 21786
rect 4924 21734 4950 21786
rect 4654 21732 4710 21734
rect 4734 21732 4790 21734
rect 4814 21732 4870 21734
rect 4894 21732 4950 21734
rect 3882 21256 3938 21312
rect 2962 19236 3018 19272
rect 2962 19216 2964 19236
rect 2964 19216 3016 19236
rect 3016 19216 3018 19236
rect 3146 16632 3202 16688
rect 3146 15680 3202 15736
rect 2870 14320 2926 14376
rect 3698 17212 3700 17232
rect 3700 17212 3752 17232
rect 3752 17212 3754 17232
rect 3698 17176 3754 17212
rect 3330 16788 3386 16824
rect 3330 16768 3332 16788
rect 3332 16768 3384 16788
rect 3384 16768 3386 16788
rect 3330 15136 3386 15192
rect 3146 10512 3202 10568
rect 4066 19796 4068 19816
rect 4068 19796 4120 19816
rect 4120 19796 4122 19816
rect 4066 19760 4122 19796
rect 4066 17740 4122 17776
rect 4066 17720 4068 17740
rect 4068 17720 4120 17740
rect 4120 17720 4122 17740
rect 4066 17312 4122 17368
rect 4066 17076 4068 17096
rect 4068 17076 4120 17096
rect 4120 17076 4122 17096
rect 4066 17040 4122 17076
rect 4066 16940 4068 16960
rect 4068 16940 4120 16960
rect 4120 16940 4122 16960
rect 4066 16904 4122 16940
rect 3974 11736 4030 11792
rect 4654 20698 4710 20700
rect 4734 20698 4790 20700
rect 4814 20698 4870 20700
rect 4894 20698 4950 20700
rect 4654 20646 4680 20698
rect 4680 20646 4710 20698
rect 4734 20646 4744 20698
rect 4744 20646 4790 20698
rect 4814 20646 4860 20698
rect 4860 20646 4870 20698
rect 4894 20646 4924 20698
rect 4924 20646 4950 20698
rect 4654 20644 4710 20646
rect 4734 20644 4790 20646
rect 4814 20644 4870 20646
rect 4894 20644 4950 20646
rect 4434 19760 4490 19816
rect 4986 19896 5042 19952
rect 4654 19610 4710 19612
rect 4734 19610 4790 19612
rect 4814 19610 4870 19612
rect 4894 19610 4950 19612
rect 4654 19558 4680 19610
rect 4680 19558 4710 19610
rect 4734 19558 4744 19610
rect 4744 19558 4790 19610
rect 4814 19558 4860 19610
rect 4860 19558 4870 19610
rect 4894 19558 4924 19610
rect 4924 19558 4950 19610
rect 4654 19556 4710 19558
rect 4734 19556 4790 19558
rect 4814 19556 4870 19558
rect 4894 19556 4950 19558
rect 4654 18522 4710 18524
rect 4734 18522 4790 18524
rect 4814 18522 4870 18524
rect 4894 18522 4950 18524
rect 4654 18470 4680 18522
rect 4680 18470 4710 18522
rect 4734 18470 4744 18522
rect 4744 18470 4790 18522
rect 4814 18470 4860 18522
rect 4860 18470 4870 18522
rect 4894 18470 4924 18522
rect 4924 18470 4950 18522
rect 4654 18468 4710 18470
rect 4734 18468 4790 18470
rect 4814 18468 4870 18470
rect 4894 18468 4950 18470
rect 4434 17992 4490 18048
rect 4250 17176 4306 17232
rect 4802 17620 4804 17640
rect 4804 17620 4856 17640
rect 4856 17620 4858 17640
rect 4802 17584 4858 17620
rect 4654 17434 4710 17436
rect 4734 17434 4790 17436
rect 4814 17434 4870 17436
rect 4894 17434 4950 17436
rect 4654 17382 4680 17434
rect 4680 17382 4710 17434
rect 4734 17382 4744 17434
rect 4744 17382 4790 17434
rect 4814 17382 4860 17434
rect 4860 17382 4870 17434
rect 4894 17382 4924 17434
rect 4924 17382 4950 17434
rect 4654 17380 4710 17382
rect 4734 17380 4790 17382
rect 4814 17380 4870 17382
rect 4894 17380 4950 17382
rect 4434 17176 4490 17232
rect 4710 16768 4766 16824
rect 4434 16496 4490 16552
rect 4654 16346 4710 16348
rect 4734 16346 4790 16348
rect 4814 16346 4870 16348
rect 4894 16346 4950 16348
rect 4654 16294 4680 16346
rect 4680 16294 4710 16346
rect 4734 16294 4744 16346
rect 4744 16294 4790 16346
rect 4814 16294 4860 16346
rect 4860 16294 4870 16346
rect 4894 16294 4924 16346
rect 4924 16294 4950 16346
rect 4654 16292 4710 16294
rect 4734 16292 4790 16294
rect 4814 16292 4870 16294
rect 4894 16292 4950 16294
rect 4654 15258 4710 15260
rect 4734 15258 4790 15260
rect 4814 15258 4870 15260
rect 4894 15258 4950 15260
rect 4654 15206 4680 15258
rect 4680 15206 4710 15258
rect 4734 15206 4744 15258
rect 4744 15206 4790 15258
rect 4814 15206 4860 15258
rect 4860 15206 4870 15258
rect 4894 15206 4924 15258
rect 4924 15206 4950 15258
rect 4654 15204 4710 15206
rect 4734 15204 4790 15206
rect 4814 15204 4870 15206
rect 4894 15204 4950 15206
rect 5814 18536 5870 18592
rect 5538 17040 5594 17096
rect 5354 15680 5410 15736
rect 5538 16108 5594 16144
rect 5538 16088 5540 16108
rect 5540 16088 5592 16108
rect 5592 16088 5594 16108
rect 4434 14456 4490 14512
rect 4710 14356 4712 14376
rect 4712 14356 4764 14376
rect 4764 14356 4766 14376
rect 4710 14320 4766 14356
rect 4654 14170 4710 14172
rect 4734 14170 4790 14172
rect 4814 14170 4870 14172
rect 4894 14170 4950 14172
rect 4654 14118 4680 14170
rect 4680 14118 4710 14170
rect 4734 14118 4744 14170
rect 4744 14118 4790 14170
rect 4814 14118 4860 14170
rect 4860 14118 4870 14170
rect 4894 14118 4924 14170
rect 4924 14118 4950 14170
rect 4654 14116 4710 14118
rect 4734 14116 4790 14118
rect 4814 14116 4870 14118
rect 4894 14116 4950 14118
rect 4654 13082 4710 13084
rect 4734 13082 4790 13084
rect 4814 13082 4870 13084
rect 4894 13082 4950 13084
rect 4654 13030 4680 13082
rect 4680 13030 4710 13082
rect 4734 13030 4744 13082
rect 4744 13030 4790 13082
rect 4814 13030 4860 13082
rect 4860 13030 4870 13082
rect 4894 13030 4924 13082
rect 4924 13030 4950 13082
rect 4654 13028 4710 13030
rect 4734 13028 4790 13030
rect 4814 13028 4870 13030
rect 4894 13028 4950 13030
rect 4526 12824 4582 12880
rect 4526 12688 4582 12744
rect 4342 8472 4398 8528
rect 4654 11994 4710 11996
rect 4734 11994 4790 11996
rect 4814 11994 4870 11996
rect 4894 11994 4950 11996
rect 4654 11942 4680 11994
rect 4680 11942 4710 11994
rect 4734 11942 4744 11994
rect 4744 11942 4790 11994
rect 4814 11942 4860 11994
rect 4860 11942 4870 11994
rect 4894 11942 4924 11994
rect 4924 11942 4950 11994
rect 4654 11940 4710 11942
rect 4734 11940 4790 11942
rect 4814 11940 4870 11942
rect 4894 11940 4950 11942
rect 4710 11092 4712 11112
rect 4712 11092 4764 11112
rect 4764 11092 4766 11112
rect 4710 11056 4766 11092
rect 4654 10906 4710 10908
rect 4734 10906 4790 10908
rect 4814 10906 4870 10908
rect 4894 10906 4950 10908
rect 4654 10854 4680 10906
rect 4680 10854 4710 10906
rect 4734 10854 4744 10906
rect 4744 10854 4790 10906
rect 4814 10854 4860 10906
rect 4860 10854 4870 10906
rect 4894 10854 4924 10906
rect 4924 10854 4950 10906
rect 4654 10852 4710 10854
rect 4734 10852 4790 10854
rect 4814 10852 4870 10854
rect 4894 10852 4950 10854
rect 4802 10260 4858 10296
rect 4802 10240 4804 10260
rect 4804 10240 4856 10260
rect 4856 10240 4858 10260
rect 4654 9818 4710 9820
rect 4734 9818 4790 9820
rect 4814 9818 4870 9820
rect 4894 9818 4950 9820
rect 4654 9766 4680 9818
rect 4680 9766 4710 9818
rect 4734 9766 4744 9818
rect 4744 9766 4790 9818
rect 4814 9766 4860 9818
rect 4860 9766 4870 9818
rect 4894 9766 4924 9818
rect 4924 9766 4950 9818
rect 4654 9764 4710 9766
rect 4734 9764 4790 9766
rect 4814 9764 4870 9766
rect 4894 9764 4950 9766
rect 4802 9560 4858 9616
rect 4894 9460 4896 9480
rect 4896 9460 4948 9480
rect 4948 9460 4950 9480
rect 4894 9424 4950 9460
rect 4654 8730 4710 8732
rect 4734 8730 4790 8732
rect 4814 8730 4870 8732
rect 4894 8730 4950 8732
rect 4654 8678 4680 8730
rect 4680 8678 4710 8730
rect 4734 8678 4744 8730
rect 4744 8678 4790 8730
rect 4814 8678 4860 8730
rect 4860 8678 4870 8730
rect 4894 8678 4924 8730
rect 4924 8678 4950 8730
rect 4654 8676 4710 8678
rect 4734 8676 4790 8678
rect 4814 8676 4870 8678
rect 4894 8676 4950 8678
rect 4654 7642 4710 7644
rect 4734 7642 4790 7644
rect 4814 7642 4870 7644
rect 4894 7642 4950 7644
rect 4654 7590 4680 7642
rect 4680 7590 4710 7642
rect 4734 7590 4744 7642
rect 4744 7590 4790 7642
rect 4814 7590 4860 7642
rect 4860 7590 4870 7642
rect 4894 7590 4924 7642
rect 4924 7590 4950 7642
rect 4654 7588 4710 7590
rect 4734 7588 4790 7590
rect 4814 7588 4870 7590
rect 4894 7588 4950 7590
rect 5170 6840 5226 6896
rect 5538 13368 5594 13424
rect 5538 12960 5594 13016
rect 5538 12316 5540 12336
rect 5540 12316 5592 12336
rect 5592 12316 5594 12336
rect 5538 12280 5594 12316
rect 5538 11736 5594 11792
rect 5538 9016 5594 9072
rect 5722 17584 5778 17640
rect 5722 15544 5778 15600
rect 5722 12960 5778 13016
rect 6090 19488 6146 19544
rect 5998 16768 6054 16824
rect 5906 12688 5962 12744
rect 5722 12008 5778 12064
rect 5630 7928 5686 7984
rect 4654 6554 4710 6556
rect 4734 6554 4790 6556
rect 4814 6554 4870 6556
rect 4894 6554 4950 6556
rect 4654 6502 4680 6554
rect 4680 6502 4710 6554
rect 4734 6502 4744 6554
rect 4744 6502 4790 6554
rect 4814 6502 4860 6554
rect 4860 6502 4870 6554
rect 4894 6502 4924 6554
rect 4924 6502 4950 6554
rect 4654 6500 4710 6502
rect 4734 6500 4790 6502
rect 4814 6500 4870 6502
rect 4894 6500 4950 6502
rect 6090 12416 6146 12472
rect 6090 12144 6146 12200
rect 6458 14476 6514 14512
rect 6458 14456 6460 14476
rect 6460 14456 6512 14476
rect 6512 14456 6514 14476
rect 6366 9424 6422 9480
rect 6366 9152 6422 9208
rect 7194 19216 7250 19272
rect 7194 18300 7196 18320
rect 7196 18300 7248 18320
rect 7248 18300 7250 18320
rect 7194 18264 7250 18300
rect 7194 16768 7250 16824
rect 6642 12144 6698 12200
rect 6734 8472 6790 8528
rect 7010 9560 7066 9616
rect 7010 8916 7012 8936
rect 7012 8916 7064 8936
rect 7064 8916 7066 8936
rect 7010 8880 7066 8916
rect 7010 8084 7066 8120
rect 7010 8064 7012 8084
rect 7012 8064 7064 8084
rect 7064 8064 7066 8084
rect 7194 13776 7250 13832
rect 7562 14320 7618 14376
rect 7470 13096 7526 13152
rect 7286 12688 7342 12744
rect 7286 9172 7342 9208
rect 7286 9152 7288 9172
rect 7288 9152 7340 9172
rect 7340 9152 7342 9172
rect 7194 8880 7250 8936
rect 7194 7692 7196 7712
rect 7196 7692 7248 7712
rect 7248 7692 7250 7712
rect 7194 7656 7250 7692
rect 6550 5908 6606 5944
rect 6550 5888 6552 5908
rect 6552 5888 6604 5908
rect 6604 5888 6606 5908
rect 4654 5466 4710 5468
rect 4734 5466 4790 5468
rect 4814 5466 4870 5468
rect 4894 5466 4950 5468
rect 4654 5414 4680 5466
rect 4680 5414 4710 5466
rect 4734 5414 4744 5466
rect 4744 5414 4790 5466
rect 4814 5414 4860 5466
rect 4860 5414 4870 5466
rect 4894 5414 4924 5466
rect 4924 5414 4950 5466
rect 4654 5412 4710 5414
rect 4734 5412 4790 5414
rect 4814 5412 4870 5414
rect 4894 5412 4950 5414
rect 8353 21242 8409 21244
rect 8433 21242 8489 21244
rect 8513 21242 8569 21244
rect 8593 21242 8649 21244
rect 8353 21190 8379 21242
rect 8379 21190 8409 21242
rect 8433 21190 8443 21242
rect 8443 21190 8489 21242
rect 8513 21190 8559 21242
rect 8559 21190 8569 21242
rect 8593 21190 8623 21242
rect 8623 21190 8649 21242
rect 8353 21188 8409 21190
rect 8433 21188 8489 21190
rect 8513 21188 8569 21190
rect 8593 21188 8649 21190
rect 8353 20154 8409 20156
rect 8433 20154 8489 20156
rect 8513 20154 8569 20156
rect 8593 20154 8649 20156
rect 8353 20102 8379 20154
rect 8379 20102 8409 20154
rect 8433 20102 8443 20154
rect 8443 20102 8489 20154
rect 8513 20102 8559 20154
rect 8559 20102 8569 20154
rect 8593 20102 8623 20154
rect 8623 20102 8649 20154
rect 8353 20100 8409 20102
rect 8433 20100 8489 20102
rect 8513 20100 8569 20102
rect 8593 20100 8649 20102
rect 9034 19760 9090 19816
rect 8353 19066 8409 19068
rect 8433 19066 8489 19068
rect 8513 19066 8569 19068
rect 8593 19066 8649 19068
rect 8353 19014 8379 19066
rect 8379 19014 8409 19066
rect 8433 19014 8443 19066
rect 8443 19014 8489 19066
rect 8513 19014 8559 19066
rect 8559 19014 8569 19066
rect 8593 19014 8623 19066
rect 8623 19014 8649 19066
rect 8353 19012 8409 19014
rect 8433 19012 8489 19014
rect 8513 19012 8569 19014
rect 8593 19012 8649 19014
rect 7838 17484 7840 17504
rect 7840 17484 7892 17504
rect 7892 17484 7894 17504
rect 7838 17448 7894 17484
rect 7746 12144 7802 12200
rect 8390 18400 8446 18456
rect 8666 18400 8722 18456
rect 8942 18028 8944 18048
rect 8944 18028 8996 18048
rect 8996 18028 8998 18048
rect 8942 17992 8998 18028
rect 8353 17978 8409 17980
rect 8433 17978 8489 17980
rect 8513 17978 8569 17980
rect 8593 17978 8649 17980
rect 8353 17926 8379 17978
rect 8379 17926 8409 17978
rect 8433 17926 8443 17978
rect 8443 17926 8489 17978
rect 8513 17926 8559 17978
rect 8559 17926 8569 17978
rect 8593 17926 8623 17978
rect 8623 17926 8649 17978
rect 8353 17924 8409 17926
rect 8433 17924 8489 17926
rect 8513 17924 8569 17926
rect 8593 17924 8649 17926
rect 8574 17176 8630 17232
rect 8353 16890 8409 16892
rect 8433 16890 8489 16892
rect 8513 16890 8569 16892
rect 8593 16890 8649 16892
rect 8353 16838 8379 16890
rect 8379 16838 8409 16890
rect 8433 16838 8443 16890
rect 8443 16838 8489 16890
rect 8513 16838 8559 16890
rect 8559 16838 8569 16890
rect 8593 16838 8623 16890
rect 8623 16838 8649 16890
rect 8353 16836 8409 16838
rect 8433 16836 8489 16838
rect 8513 16836 8569 16838
rect 8593 16836 8649 16838
rect 8353 15802 8409 15804
rect 8433 15802 8489 15804
rect 8513 15802 8569 15804
rect 8593 15802 8649 15804
rect 8353 15750 8379 15802
rect 8379 15750 8409 15802
rect 8433 15750 8443 15802
rect 8443 15750 8489 15802
rect 8513 15750 8559 15802
rect 8559 15750 8569 15802
rect 8593 15750 8623 15802
rect 8623 15750 8649 15802
rect 8353 15748 8409 15750
rect 8433 15748 8489 15750
rect 8513 15748 8569 15750
rect 8593 15748 8649 15750
rect 8206 14864 8262 14920
rect 8353 14714 8409 14716
rect 8433 14714 8489 14716
rect 8513 14714 8569 14716
rect 8593 14714 8649 14716
rect 8353 14662 8379 14714
rect 8379 14662 8409 14714
rect 8433 14662 8443 14714
rect 8443 14662 8489 14714
rect 8513 14662 8559 14714
rect 8559 14662 8569 14714
rect 8593 14662 8623 14714
rect 8623 14662 8649 14714
rect 8353 14660 8409 14662
rect 8433 14660 8489 14662
rect 8513 14660 8569 14662
rect 8593 14660 8649 14662
rect 8114 13132 8116 13152
rect 8116 13132 8168 13152
rect 8168 13132 8170 13152
rect 8114 13096 8170 13132
rect 8353 13626 8409 13628
rect 8433 13626 8489 13628
rect 8513 13626 8569 13628
rect 8593 13626 8649 13628
rect 8353 13574 8379 13626
rect 8379 13574 8409 13626
rect 8433 13574 8443 13626
rect 8443 13574 8489 13626
rect 8513 13574 8559 13626
rect 8559 13574 8569 13626
rect 8593 13574 8623 13626
rect 8623 13574 8649 13626
rect 8353 13572 8409 13574
rect 8433 13572 8489 13574
rect 8513 13572 8569 13574
rect 8593 13572 8649 13574
rect 8353 12538 8409 12540
rect 8433 12538 8489 12540
rect 8513 12538 8569 12540
rect 8593 12538 8649 12540
rect 8353 12486 8379 12538
rect 8379 12486 8409 12538
rect 8433 12486 8443 12538
rect 8443 12486 8489 12538
rect 8513 12486 8559 12538
rect 8559 12486 8569 12538
rect 8593 12486 8623 12538
rect 8623 12486 8649 12538
rect 8353 12484 8409 12486
rect 8433 12484 8489 12486
rect 8513 12484 8569 12486
rect 8593 12484 8649 12486
rect 7838 11872 7894 11928
rect 8850 17040 8906 17096
rect 8850 16632 8906 16688
rect 9586 18808 9642 18864
rect 10138 19508 10194 19544
rect 10138 19488 10140 19508
rect 10140 19488 10192 19508
rect 10192 19488 10194 19508
rect 9310 16496 9366 16552
rect 9126 16088 9182 16144
rect 9770 18420 9826 18456
rect 9770 18400 9772 18420
rect 9772 18400 9824 18420
rect 9824 18400 9826 18420
rect 9586 18264 9642 18320
rect 9126 15408 9182 15464
rect 9034 15000 9090 15056
rect 8850 12280 8906 12336
rect 9126 12824 9182 12880
rect 9034 12008 9090 12064
rect 8942 11736 8998 11792
rect 8353 11450 8409 11452
rect 8433 11450 8489 11452
rect 8513 11450 8569 11452
rect 8593 11450 8649 11452
rect 8353 11398 8379 11450
rect 8379 11398 8409 11450
rect 8433 11398 8443 11450
rect 8443 11398 8489 11450
rect 8513 11398 8559 11450
rect 8559 11398 8569 11450
rect 8593 11398 8623 11450
rect 8623 11398 8649 11450
rect 8353 11396 8409 11398
rect 8433 11396 8489 11398
rect 8513 11396 8569 11398
rect 8593 11396 8649 11398
rect 8482 10512 8538 10568
rect 8353 10362 8409 10364
rect 8433 10362 8489 10364
rect 8513 10362 8569 10364
rect 8593 10362 8649 10364
rect 8353 10310 8379 10362
rect 8379 10310 8409 10362
rect 8433 10310 8443 10362
rect 8443 10310 8489 10362
rect 8513 10310 8559 10362
rect 8559 10310 8569 10362
rect 8593 10310 8623 10362
rect 8623 10310 8649 10362
rect 8353 10308 8409 10310
rect 8433 10308 8489 10310
rect 8513 10308 8569 10310
rect 8593 10308 8649 10310
rect 8298 9560 8354 9616
rect 8758 9832 8814 9888
rect 8482 9560 8538 9616
rect 7654 8608 7710 8664
rect 7562 7812 7618 7848
rect 7562 7792 7564 7812
rect 7564 7792 7616 7812
rect 7616 7792 7618 7812
rect 7562 7656 7618 7712
rect 4654 4378 4710 4380
rect 4734 4378 4790 4380
rect 4814 4378 4870 4380
rect 4894 4378 4950 4380
rect 4654 4326 4680 4378
rect 4680 4326 4710 4378
rect 4734 4326 4744 4378
rect 4744 4326 4790 4378
rect 4814 4326 4860 4378
rect 4860 4326 4870 4378
rect 4894 4326 4924 4378
rect 4924 4326 4950 4378
rect 4654 4324 4710 4326
rect 4734 4324 4790 4326
rect 4814 4324 4870 4326
rect 4894 4324 4950 4326
rect 8114 9288 8170 9344
rect 7930 9152 7986 9208
rect 7930 7964 7932 7984
rect 7932 7964 7984 7984
rect 7984 7964 7986 7984
rect 7930 7928 7986 7964
rect 7930 7656 7986 7712
rect 7930 7540 7986 7576
rect 7930 7520 7932 7540
rect 7932 7520 7984 7540
rect 7984 7520 7986 7540
rect 7930 7384 7986 7440
rect 8353 9274 8409 9276
rect 8433 9274 8489 9276
rect 8513 9274 8569 9276
rect 8593 9274 8649 9276
rect 8353 9222 8379 9274
rect 8379 9222 8409 9274
rect 8433 9222 8443 9274
rect 8443 9222 8489 9274
rect 8513 9222 8559 9274
rect 8559 9222 8569 9274
rect 8593 9222 8623 9274
rect 8623 9222 8649 9274
rect 8353 9220 8409 9222
rect 8433 9220 8489 9222
rect 8513 9220 8569 9222
rect 8593 9220 8649 9222
rect 8390 8492 8446 8528
rect 8390 8472 8392 8492
rect 8392 8472 8444 8492
rect 8444 8472 8446 8492
rect 8298 8336 8354 8392
rect 8353 8186 8409 8188
rect 8433 8186 8489 8188
rect 8513 8186 8569 8188
rect 8593 8186 8649 8188
rect 8353 8134 8379 8186
rect 8379 8134 8409 8186
rect 8433 8134 8443 8186
rect 8443 8134 8489 8186
rect 8513 8134 8559 8186
rect 8559 8134 8569 8186
rect 8593 8134 8623 8186
rect 8623 8134 8649 8186
rect 8353 8132 8409 8134
rect 8433 8132 8489 8134
rect 8513 8132 8569 8134
rect 8593 8132 8649 8134
rect 8758 8200 8814 8256
rect 8942 10920 8998 10976
rect 8942 9696 8998 9752
rect 8942 9288 8998 9344
rect 8942 8608 8998 8664
rect 8850 8064 8906 8120
rect 8353 7098 8409 7100
rect 8433 7098 8489 7100
rect 8513 7098 8569 7100
rect 8593 7098 8649 7100
rect 8353 7046 8379 7098
rect 8379 7046 8409 7098
rect 8433 7046 8443 7098
rect 8443 7046 8489 7098
rect 8513 7046 8559 7098
rect 8559 7046 8569 7098
rect 8593 7046 8623 7098
rect 8623 7046 8649 7098
rect 8353 7044 8409 7046
rect 8433 7044 8489 7046
rect 8513 7044 8569 7046
rect 8593 7044 8649 7046
rect 8758 6976 8814 7032
rect 7930 6160 7986 6216
rect 8574 6724 8630 6760
rect 8574 6704 8576 6724
rect 8576 6704 8628 6724
rect 8628 6704 8630 6724
rect 8390 6432 8446 6488
rect 8666 6332 8668 6352
rect 8668 6332 8720 6352
rect 8720 6332 8722 6352
rect 8666 6296 8722 6332
rect 8353 6010 8409 6012
rect 8433 6010 8489 6012
rect 8513 6010 8569 6012
rect 8593 6010 8649 6012
rect 8353 5958 8379 6010
rect 8379 5958 8409 6010
rect 8433 5958 8443 6010
rect 8443 5958 8489 6010
rect 8513 5958 8559 6010
rect 8559 5958 8569 6010
rect 8593 5958 8623 6010
rect 8623 5958 8649 6010
rect 8353 5956 8409 5958
rect 8433 5956 8489 5958
rect 8513 5956 8569 5958
rect 8593 5956 8649 5958
rect 8942 7248 8998 7304
rect 9678 17176 9734 17232
rect 9954 16768 10010 16824
rect 10230 16496 10286 16552
rect 10782 18536 10838 18592
rect 9218 9832 9274 9888
rect 9218 9696 9274 9752
rect 9126 8064 9182 8120
rect 9034 6568 9090 6624
rect 8353 4922 8409 4924
rect 8433 4922 8489 4924
rect 8513 4922 8569 4924
rect 8593 4922 8649 4924
rect 8353 4870 8379 4922
rect 8379 4870 8409 4922
rect 8433 4870 8443 4922
rect 8443 4870 8489 4922
rect 8513 4870 8559 4922
rect 8559 4870 8569 4922
rect 8593 4870 8623 4922
rect 8623 4870 8649 4922
rect 8353 4868 8409 4870
rect 8433 4868 8489 4870
rect 8513 4868 8569 4870
rect 8593 4868 8649 4870
rect 9494 9016 9550 9072
rect 9678 12688 9734 12744
rect 9678 12044 9680 12064
rect 9680 12044 9732 12064
rect 9732 12044 9734 12064
rect 9678 12008 9734 12044
rect 9954 11736 10010 11792
rect 9862 11600 9918 11656
rect 9862 8472 9918 8528
rect 9586 6840 9642 6896
rect 9494 6704 9550 6760
rect 9494 6568 9550 6624
rect 9310 5888 9366 5944
rect 9402 5652 9404 5672
rect 9404 5652 9456 5672
rect 9456 5652 9458 5672
rect 9402 5616 9458 5652
rect 9678 5888 9734 5944
rect 10230 14456 10286 14512
rect 10322 13232 10378 13288
rect 10782 13776 10838 13832
rect 10598 11736 10654 11792
rect 10506 11600 10562 11656
rect 10138 9152 10194 9208
rect 10230 9016 10286 9072
rect 10046 6840 10102 6896
rect 10138 6740 10140 6760
rect 10140 6740 10192 6760
rect 10192 6740 10194 6760
rect 10138 6704 10194 6740
rect 10414 9016 10470 9072
rect 10690 11464 10746 11520
rect 10690 9696 10746 9752
rect 11242 16632 11298 16688
rect 11334 16496 11390 16552
rect 12052 21786 12108 21788
rect 12132 21786 12188 21788
rect 12212 21786 12268 21788
rect 12292 21786 12348 21788
rect 12052 21734 12078 21786
rect 12078 21734 12108 21786
rect 12132 21734 12142 21786
rect 12142 21734 12188 21786
rect 12212 21734 12258 21786
rect 12258 21734 12268 21786
rect 12292 21734 12322 21786
rect 12322 21734 12348 21786
rect 12052 21732 12108 21734
rect 12132 21732 12188 21734
rect 12212 21732 12268 21734
rect 12292 21732 12348 21734
rect 12052 20698 12108 20700
rect 12132 20698 12188 20700
rect 12212 20698 12268 20700
rect 12292 20698 12348 20700
rect 12052 20646 12078 20698
rect 12078 20646 12108 20698
rect 12132 20646 12142 20698
rect 12142 20646 12188 20698
rect 12212 20646 12258 20698
rect 12258 20646 12268 20698
rect 12292 20646 12322 20698
rect 12322 20646 12348 20698
rect 12052 20644 12108 20646
rect 12132 20644 12188 20646
rect 12212 20644 12268 20646
rect 12292 20644 12348 20646
rect 12052 19610 12108 19612
rect 12132 19610 12188 19612
rect 12212 19610 12268 19612
rect 12292 19610 12348 19612
rect 12052 19558 12078 19610
rect 12078 19558 12108 19610
rect 12132 19558 12142 19610
rect 12142 19558 12188 19610
rect 12212 19558 12258 19610
rect 12258 19558 12268 19610
rect 12292 19558 12322 19610
rect 12322 19558 12348 19610
rect 12052 19556 12108 19558
rect 12132 19556 12188 19558
rect 12212 19556 12268 19558
rect 12292 19556 12348 19558
rect 12346 19116 12348 19136
rect 12348 19116 12400 19136
rect 12400 19116 12402 19136
rect 12346 19080 12402 19116
rect 12052 18522 12108 18524
rect 12132 18522 12188 18524
rect 12212 18522 12268 18524
rect 12292 18522 12348 18524
rect 12052 18470 12078 18522
rect 12078 18470 12108 18522
rect 12132 18470 12142 18522
rect 12142 18470 12188 18522
rect 12212 18470 12258 18522
rect 12258 18470 12268 18522
rect 12292 18470 12322 18522
rect 12322 18470 12348 18522
rect 12052 18468 12108 18470
rect 12132 18468 12188 18470
rect 12212 18468 12268 18470
rect 12292 18468 12348 18470
rect 12530 19508 12586 19544
rect 12530 19488 12532 19508
rect 12532 19488 12584 19508
rect 12584 19488 12586 19508
rect 12622 19216 12678 19272
rect 12438 17584 12494 17640
rect 12052 17434 12108 17436
rect 12132 17434 12188 17436
rect 12212 17434 12268 17436
rect 12292 17434 12348 17436
rect 12052 17382 12078 17434
rect 12078 17382 12108 17434
rect 12132 17382 12142 17434
rect 12142 17382 12188 17434
rect 12212 17382 12258 17434
rect 12258 17382 12268 17434
rect 12292 17382 12322 17434
rect 12322 17382 12348 17434
rect 12052 17380 12108 17382
rect 12132 17380 12188 17382
rect 12212 17380 12268 17382
rect 12292 17380 12348 17382
rect 12254 17040 12310 17096
rect 10874 12144 10930 12200
rect 10690 6976 10746 7032
rect 10598 6840 10654 6896
rect 10506 6432 10562 6488
rect 10322 6160 10378 6216
rect 9862 5208 9918 5264
rect 10322 4700 10324 4720
rect 10324 4700 10376 4720
rect 10376 4700 10378 4720
rect 10322 4664 10378 4700
rect 11150 12824 11206 12880
rect 12052 16346 12108 16348
rect 12132 16346 12188 16348
rect 12212 16346 12268 16348
rect 12292 16346 12348 16348
rect 12052 16294 12078 16346
rect 12078 16294 12108 16346
rect 12132 16294 12142 16346
rect 12142 16294 12188 16346
rect 12212 16294 12258 16346
rect 12258 16294 12268 16346
rect 12292 16294 12322 16346
rect 12322 16294 12348 16346
rect 12052 16292 12108 16294
rect 12132 16292 12188 16294
rect 12212 16292 12268 16294
rect 12292 16292 12348 16294
rect 11518 12552 11574 12608
rect 12052 15258 12108 15260
rect 12132 15258 12188 15260
rect 12212 15258 12268 15260
rect 12292 15258 12348 15260
rect 12052 15206 12078 15258
rect 12078 15206 12108 15258
rect 12132 15206 12142 15258
rect 12142 15206 12188 15258
rect 12212 15206 12258 15258
rect 12258 15206 12268 15258
rect 12292 15206 12322 15258
rect 12322 15206 12348 15258
rect 12052 15204 12108 15206
rect 12132 15204 12188 15206
rect 12212 15204 12268 15206
rect 12292 15204 12348 15206
rect 12070 15020 12126 15056
rect 12070 15000 12072 15020
rect 12072 15000 12124 15020
rect 12124 15000 12126 15020
rect 13082 19372 13138 19408
rect 13082 19352 13084 19372
rect 13084 19352 13136 19372
rect 13136 19352 13138 19372
rect 12622 16088 12678 16144
rect 12990 16088 13046 16144
rect 12714 15700 12770 15736
rect 12714 15680 12716 15700
rect 12716 15680 12768 15700
rect 12768 15680 12770 15700
rect 12052 14170 12108 14172
rect 12132 14170 12188 14172
rect 12212 14170 12268 14172
rect 12292 14170 12348 14172
rect 12052 14118 12078 14170
rect 12078 14118 12108 14170
rect 12132 14118 12142 14170
rect 12142 14118 12188 14170
rect 12212 14118 12258 14170
rect 12258 14118 12268 14170
rect 12292 14118 12322 14170
rect 12322 14118 12348 14170
rect 12052 14116 12108 14118
rect 12132 14116 12188 14118
rect 12212 14116 12268 14118
rect 12292 14116 12348 14118
rect 12622 14320 12678 14376
rect 12162 13776 12218 13832
rect 12052 13082 12108 13084
rect 12132 13082 12188 13084
rect 12212 13082 12268 13084
rect 12292 13082 12348 13084
rect 12052 13030 12078 13082
rect 12078 13030 12108 13082
rect 12132 13030 12142 13082
rect 12142 13030 12188 13082
rect 12212 13030 12258 13082
rect 12258 13030 12268 13082
rect 12292 13030 12322 13082
rect 12322 13030 12348 13082
rect 12052 13028 12108 13030
rect 12132 13028 12188 13030
rect 12212 13028 12268 13030
rect 12292 13028 12348 13030
rect 12714 12824 12770 12880
rect 11518 11056 11574 11112
rect 10966 7520 11022 7576
rect 11426 8608 11482 8664
rect 11702 10920 11758 10976
rect 11794 10804 11850 10840
rect 11794 10784 11796 10804
rect 11796 10784 11848 10804
rect 11848 10784 11850 10804
rect 11610 9288 11666 9344
rect 11794 8336 11850 8392
rect 11610 7928 11666 7984
rect 11610 7656 11666 7712
rect 8353 3834 8409 3836
rect 8433 3834 8489 3836
rect 8513 3834 8569 3836
rect 8593 3834 8649 3836
rect 8353 3782 8379 3834
rect 8379 3782 8409 3834
rect 8433 3782 8443 3834
rect 8443 3782 8489 3834
rect 8513 3782 8559 3834
rect 8559 3782 8569 3834
rect 8593 3782 8623 3834
rect 8623 3782 8649 3834
rect 8353 3780 8409 3782
rect 8433 3780 8489 3782
rect 8513 3780 8569 3782
rect 8593 3780 8649 3782
rect 4654 3290 4710 3292
rect 4734 3290 4790 3292
rect 4814 3290 4870 3292
rect 4894 3290 4950 3292
rect 4654 3238 4680 3290
rect 4680 3238 4710 3290
rect 4734 3238 4744 3290
rect 4744 3238 4790 3290
rect 4814 3238 4860 3290
rect 4860 3238 4870 3290
rect 4894 3238 4924 3290
rect 4924 3238 4950 3290
rect 4654 3236 4710 3238
rect 4734 3236 4790 3238
rect 4814 3236 4870 3238
rect 4894 3236 4950 3238
rect 1950 3052 2006 3088
rect 11794 6996 11850 7032
rect 11794 6976 11796 6996
rect 11796 6976 11848 6996
rect 11848 6976 11850 6996
rect 11702 5072 11758 5128
rect 11702 4820 11758 4856
rect 12052 11994 12108 11996
rect 12132 11994 12188 11996
rect 12212 11994 12268 11996
rect 12292 11994 12348 11996
rect 12052 11942 12078 11994
rect 12078 11942 12108 11994
rect 12132 11942 12142 11994
rect 12142 11942 12188 11994
rect 12212 11942 12258 11994
rect 12258 11942 12268 11994
rect 12292 11942 12322 11994
rect 12322 11942 12348 11994
rect 12052 11940 12108 11942
rect 12132 11940 12188 11942
rect 12212 11940 12268 11942
rect 12292 11940 12348 11942
rect 12714 12688 12770 12744
rect 12898 12552 12954 12608
rect 12530 11872 12586 11928
rect 12714 12144 12770 12200
rect 12052 10906 12108 10908
rect 12132 10906 12188 10908
rect 12212 10906 12268 10908
rect 12292 10906 12348 10908
rect 12052 10854 12078 10906
rect 12078 10854 12108 10906
rect 12132 10854 12142 10906
rect 12142 10854 12188 10906
rect 12212 10854 12258 10906
rect 12258 10854 12268 10906
rect 12292 10854 12322 10906
rect 12322 10854 12348 10906
rect 12052 10852 12108 10854
rect 12132 10852 12188 10854
rect 12212 10852 12268 10854
rect 12292 10852 12348 10854
rect 11978 10240 12034 10296
rect 12530 10512 12586 10568
rect 12052 9818 12108 9820
rect 12132 9818 12188 9820
rect 12212 9818 12268 9820
rect 12292 9818 12348 9820
rect 12052 9766 12078 9818
rect 12078 9766 12108 9818
rect 12132 9766 12142 9818
rect 12142 9766 12188 9818
rect 12212 9766 12258 9818
rect 12258 9766 12268 9818
rect 12292 9766 12322 9818
rect 12322 9766 12348 9818
rect 12052 9764 12108 9766
rect 12132 9764 12188 9766
rect 12212 9764 12268 9766
rect 12292 9764 12348 9766
rect 12530 9968 12586 10024
rect 12052 8730 12108 8732
rect 12132 8730 12188 8732
rect 12212 8730 12268 8732
rect 12292 8730 12348 8732
rect 12052 8678 12078 8730
rect 12078 8678 12108 8730
rect 12132 8678 12142 8730
rect 12142 8678 12188 8730
rect 12212 8678 12258 8730
rect 12258 8678 12268 8730
rect 12292 8678 12322 8730
rect 12322 8678 12348 8730
rect 12052 8676 12108 8678
rect 12132 8676 12188 8678
rect 12212 8676 12268 8678
rect 12292 8676 12348 8678
rect 13266 14728 13322 14784
rect 13910 19352 13966 19408
rect 13450 17040 13506 17096
rect 13082 12280 13138 12336
rect 12714 8880 12770 8936
rect 12162 8472 12218 8528
rect 12052 7642 12108 7644
rect 12132 7642 12188 7644
rect 12212 7642 12268 7644
rect 12292 7642 12348 7644
rect 12052 7590 12078 7642
rect 12078 7590 12108 7642
rect 12132 7590 12142 7642
rect 12142 7590 12188 7642
rect 12212 7590 12258 7642
rect 12258 7590 12268 7642
rect 12292 7590 12322 7642
rect 12322 7590 12348 7642
rect 12052 7588 12108 7590
rect 12132 7588 12188 7590
rect 12212 7588 12268 7590
rect 12292 7588 12348 7590
rect 12346 6840 12402 6896
rect 12052 6554 12108 6556
rect 12132 6554 12188 6556
rect 12212 6554 12268 6556
rect 12292 6554 12348 6556
rect 12052 6502 12078 6554
rect 12078 6502 12108 6554
rect 12132 6502 12142 6554
rect 12142 6502 12188 6554
rect 12212 6502 12258 6554
rect 12258 6502 12268 6554
rect 12292 6502 12322 6554
rect 12322 6502 12348 6554
rect 12052 6500 12108 6502
rect 12132 6500 12188 6502
rect 12212 6500 12268 6502
rect 12292 6500 12348 6502
rect 12622 6432 12678 6488
rect 12052 5466 12108 5468
rect 12132 5466 12188 5468
rect 12212 5466 12268 5468
rect 12292 5466 12348 5468
rect 12052 5414 12078 5466
rect 12078 5414 12108 5466
rect 12132 5414 12142 5466
rect 12142 5414 12188 5466
rect 12212 5414 12258 5466
rect 12258 5414 12268 5466
rect 12292 5414 12322 5466
rect 12322 5414 12348 5466
rect 12052 5412 12108 5414
rect 12132 5412 12188 5414
rect 12212 5412 12268 5414
rect 12292 5412 12348 5414
rect 12438 5072 12494 5128
rect 12254 4972 12256 4992
rect 12256 4972 12308 4992
rect 12308 4972 12310 4992
rect 12254 4936 12310 4972
rect 11702 4800 11704 4820
rect 11704 4800 11756 4820
rect 11756 4800 11758 4820
rect 12346 4800 12402 4856
rect 12052 4378 12108 4380
rect 12132 4378 12188 4380
rect 12212 4378 12268 4380
rect 12292 4378 12348 4380
rect 12052 4326 12078 4378
rect 12078 4326 12108 4378
rect 12132 4326 12142 4378
rect 12142 4326 12188 4378
rect 12212 4326 12258 4378
rect 12258 4326 12268 4378
rect 12292 4326 12322 4378
rect 12322 4326 12348 4378
rect 12052 4324 12108 4326
rect 12132 4324 12188 4326
rect 12212 4324 12268 4326
rect 12292 4324 12348 4326
rect 11886 4140 11942 4176
rect 11886 4120 11888 4140
rect 11888 4120 11940 4140
rect 11940 4120 11942 4140
rect 1950 3032 1952 3052
rect 1952 3032 2004 3052
rect 2004 3032 2006 3052
rect 4654 2202 4710 2204
rect 4734 2202 4790 2204
rect 4814 2202 4870 2204
rect 4894 2202 4950 2204
rect 4654 2150 4680 2202
rect 4680 2150 4710 2202
rect 4734 2150 4744 2202
rect 4744 2150 4790 2202
rect 4814 2150 4860 2202
rect 4860 2150 4870 2202
rect 4894 2150 4924 2202
rect 4924 2150 4950 2202
rect 4654 2148 4710 2150
rect 4734 2148 4790 2150
rect 4814 2148 4870 2150
rect 4894 2148 4950 2150
rect 8353 2746 8409 2748
rect 8433 2746 8489 2748
rect 8513 2746 8569 2748
rect 8593 2746 8649 2748
rect 8353 2694 8379 2746
rect 8379 2694 8409 2746
rect 8433 2694 8443 2746
rect 8443 2694 8489 2746
rect 8513 2694 8559 2746
rect 8559 2694 8569 2746
rect 8593 2694 8623 2746
rect 8623 2694 8649 2746
rect 8353 2692 8409 2694
rect 8433 2692 8489 2694
rect 8513 2692 8569 2694
rect 8593 2692 8649 2694
rect 13266 11872 13322 11928
rect 13174 11620 13230 11656
rect 13174 11600 13176 11620
rect 13176 11600 13228 11620
rect 13228 11600 13230 11620
rect 12898 11464 12954 11520
rect 12898 11192 12954 11248
rect 12990 10956 12992 10976
rect 12992 10956 13044 10976
rect 13044 10956 13046 10976
rect 12990 10920 13046 10956
rect 12990 10784 13046 10840
rect 12990 10104 13046 10160
rect 13082 7520 13138 7576
rect 12990 4256 13046 4312
rect 13082 3884 13084 3904
rect 13084 3884 13136 3904
rect 13136 3884 13138 3904
rect 12052 3290 12108 3292
rect 12132 3290 12188 3292
rect 12212 3290 12268 3292
rect 12292 3290 12348 3292
rect 12052 3238 12078 3290
rect 12078 3238 12108 3290
rect 12132 3238 12142 3290
rect 12142 3238 12188 3290
rect 12212 3238 12258 3290
rect 12258 3238 12268 3290
rect 12292 3238 12322 3290
rect 12322 3238 12348 3290
rect 12052 3236 12108 3238
rect 12132 3236 12188 3238
rect 12212 3236 12268 3238
rect 12292 3236 12348 3238
rect 8574 2488 8630 2544
rect 13082 3848 13138 3884
rect 13358 8336 13414 8392
rect 13358 4800 13414 4856
rect 14094 16768 14150 16824
rect 13818 15272 13874 15328
rect 13634 11192 13690 11248
rect 13726 10784 13782 10840
rect 14002 12688 14058 12744
rect 14094 12280 14150 12336
rect 14370 12824 14426 12880
rect 14370 12416 14426 12472
rect 14094 11872 14150 11928
rect 13818 10376 13874 10432
rect 13634 8336 13690 8392
rect 13818 10104 13874 10160
rect 13634 6976 13690 7032
rect 13634 5752 13690 5808
rect 13818 6024 13874 6080
rect 13726 5344 13782 5400
rect 13818 5072 13874 5128
rect 13910 4936 13966 4992
rect 14002 4800 14058 4856
rect 13910 4528 13966 4584
rect 12622 3304 12678 3360
rect 14462 11056 14518 11112
rect 15014 19216 15070 19272
rect 15106 18672 15162 18728
rect 15474 18264 15530 18320
rect 14922 17040 14978 17096
rect 14646 13912 14702 13968
rect 15198 15852 15200 15872
rect 15200 15852 15252 15872
rect 15252 15852 15254 15872
rect 15198 15816 15254 15852
rect 15106 15700 15162 15736
rect 15106 15680 15108 15700
rect 15108 15680 15160 15700
rect 15160 15680 15162 15700
rect 14922 14048 14978 14104
rect 14462 7656 14518 7712
rect 14186 5888 14242 5944
rect 14738 9016 14794 9072
rect 14922 10920 14978 10976
rect 15750 21242 15806 21244
rect 15830 21242 15886 21244
rect 15910 21242 15966 21244
rect 15990 21242 16046 21244
rect 15750 21190 15776 21242
rect 15776 21190 15806 21242
rect 15830 21190 15840 21242
rect 15840 21190 15886 21242
rect 15910 21190 15956 21242
rect 15956 21190 15966 21242
rect 15990 21190 16020 21242
rect 16020 21190 16046 21242
rect 15750 21188 15806 21190
rect 15830 21188 15886 21190
rect 15910 21188 15966 21190
rect 15990 21188 16046 21190
rect 15750 20154 15806 20156
rect 15830 20154 15886 20156
rect 15910 20154 15966 20156
rect 15990 20154 16046 20156
rect 15750 20102 15776 20154
rect 15776 20102 15806 20154
rect 15830 20102 15840 20154
rect 15840 20102 15886 20154
rect 15910 20102 15956 20154
rect 15956 20102 15966 20154
rect 15990 20102 16020 20154
rect 16020 20102 16046 20154
rect 15750 20100 15806 20102
rect 15830 20100 15886 20102
rect 15910 20100 15966 20102
rect 15990 20100 16046 20102
rect 15658 19896 15714 19952
rect 16302 20304 16358 20360
rect 16118 19352 16174 19408
rect 15750 19066 15806 19068
rect 15830 19066 15886 19068
rect 15910 19066 15966 19068
rect 15990 19066 16046 19068
rect 15750 19014 15776 19066
rect 15776 19014 15806 19066
rect 15830 19014 15840 19066
rect 15840 19014 15886 19066
rect 15910 19014 15956 19066
rect 15956 19014 15966 19066
rect 15990 19014 16020 19066
rect 16020 19014 16046 19066
rect 15750 19012 15806 19014
rect 15830 19012 15886 19014
rect 15910 19012 15966 19014
rect 15990 19012 16046 19014
rect 15750 17978 15806 17980
rect 15830 17978 15886 17980
rect 15910 17978 15966 17980
rect 15990 17978 16046 17980
rect 15750 17926 15776 17978
rect 15776 17926 15806 17978
rect 15830 17926 15840 17978
rect 15840 17926 15886 17978
rect 15910 17926 15956 17978
rect 15956 17926 15966 17978
rect 15990 17926 16020 17978
rect 16020 17926 16046 17978
rect 15750 17924 15806 17926
rect 15830 17924 15886 17926
rect 15910 17924 15966 17926
rect 15990 17924 16046 17926
rect 15658 17040 15714 17096
rect 15750 16890 15806 16892
rect 15830 16890 15886 16892
rect 15910 16890 15966 16892
rect 15990 16890 16046 16892
rect 15750 16838 15776 16890
rect 15776 16838 15806 16890
rect 15830 16838 15840 16890
rect 15840 16838 15886 16890
rect 15910 16838 15956 16890
rect 15956 16838 15966 16890
rect 15990 16838 16020 16890
rect 16020 16838 16046 16890
rect 15750 16836 15806 16838
rect 15830 16836 15886 16838
rect 15910 16836 15966 16838
rect 15990 16836 16046 16838
rect 16302 16360 16358 16416
rect 16578 18672 16634 18728
rect 15750 15802 15806 15804
rect 15830 15802 15886 15804
rect 15910 15802 15966 15804
rect 15990 15802 16046 15804
rect 15750 15750 15776 15802
rect 15776 15750 15806 15802
rect 15830 15750 15840 15802
rect 15840 15750 15886 15802
rect 15910 15750 15956 15802
rect 15956 15750 15966 15802
rect 15990 15750 16020 15802
rect 16020 15750 16046 15802
rect 15750 15748 15806 15750
rect 15830 15748 15886 15750
rect 15910 15748 15966 15750
rect 15990 15748 16046 15750
rect 15658 15408 15714 15464
rect 15842 14864 15898 14920
rect 15382 12280 15438 12336
rect 15198 9968 15254 10024
rect 14922 8880 14978 8936
rect 15014 8064 15070 8120
rect 15014 7656 15070 7712
rect 15014 7112 15070 7168
rect 14462 6024 14518 6080
rect 14002 4020 14004 4040
rect 14004 4020 14056 4040
rect 14056 4020 14058 4040
rect 14002 3984 14058 4020
rect 14094 3188 14150 3224
rect 14370 5752 14426 5808
rect 14646 4664 14702 4720
rect 14370 4120 14426 4176
rect 15014 6296 15070 6352
rect 14646 3984 14702 4040
rect 14094 3168 14096 3188
rect 14096 3168 14148 3188
rect 14148 3168 14150 3188
rect 15106 3032 15162 3088
rect 12530 2488 12586 2544
rect 14370 2896 14426 2952
rect 12052 2202 12108 2204
rect 12132 2202 12188 2204
rect 12212 2202 12268 2204
rect 12292 2202 12348 2204
rect 12052 2150 12078 2202
rect 12078 2150 12108 2202
rect 12132 2150 12142 2202
rect 12142 2150 12188 2202
rect 12212 2150 12258 2202
rect 12258 2150 12268 2202
rect 12292 2150 12322 2202
rect 12322 2150 12348 2202
rect 12052 2148 12108 2150
rect 12132 2148 12188 2150
rect 12212 2148 12268 2150
rect 12292 2148 12348 2150
rect 15750 14714 15806 14716
rect 15830 14714 15886 14716
rect 15910 14714 15966 14716
rect 15990 14714 16046 14716
rect 15750 14662 15776 14714
rect 15776 14662 15806 14714
rect 15830 14662 15840 14714
rect 15840 14662 15886 14714
rect 15910 14662 15956 14714
rect 15956 14662 15966 14714
rect 15990 14662 16020 14714
rect 16020 14662 16046 14714
rect 15750 14660 15806 14662
rect 15830 14660 15886 14662
rect 15910 14660 15966 14662
rect 15990 14660 16046 14662
rect 15750 14220 15752 14240
rect 15752 14220 15804 14240
rect 15804 14220 15806 14240
rect 15750 14184 15806 14220
rect 15750 13626 15806 13628
rect 15830 13626 15886 13628
rect 15910 13626 15966 13628
rect 15990 13626 16046 13628
rect 15750 13574 15776 13626
rect 15776 13574 15806 13626
rect 15830 13574 15840 13626
rect 15840 13574 15886 13626
rect 15910 13574 15956 13626
rect 15956 13574 15966 13626
rect 15990 13574 16020 13626
rect 16020 13574 16046 13626
rect 15750 13572 15806 13574
rect 15830 13572 15886 13574
rect 15910 13572 15966 13574
rect 15990 13572 16046 13574
rect 16210 14592 16266 14648
rect 16118 13368 16174 13424
rect 15842 13096 15898 13152
rect 15750 12538 15806 12540
rect 15830 12538 15886 12540
rect 15910 12538 15966 12540
rect 15990 12538 16046 12540
rect 15750 12486 15776 12538
rect 15776 12486 15806 12538
rect 15830 12486 15840 12538
rect 15840 12486 15886 12538
rect 15910 12486 15956 12538
rect 15956 12486 15966 12538
rect 15990 12486 16020 12538
rect 16020 12486 16046 12538
rect 15750 12484 15806 12486
rect 15830 12484 15886 12486
rect 15910 12484 15966 12486
rect 15990 12484 16046 12486
rect 15750 11872 15806 11928
rect 15750 11450 15806 11452
rect 15830 11450 15886 11452
rect 15910 11450 15966 11452
rect 15990 11450 16046 11452
rect 15750 11398 15776 11450
rect 15776 11398 15806 11450
rect 15830 11398 15840 11450
rect 15840 11398 15886 11450
rect 15910 11398 15956 11450
rect 15956 11398 15966 11450
rect 15990 11398 16020 11450
rect 16020 11398 16046 11450
rect 15750 11396 15806 11398
rect 15830 11396 15886 11398
rect 15910 11396 15966 11398
rect 15990 11396 16046 11398
rect 15658 10920 15714 10976
rect 15658 10784 15714 10840
rect 15750 10362 15806 10364
rect 15830 10362 15886 10364
rect 15910 10362 15966 10364
rect 15990 10362 16046 10364
rect 15750 10310 15776 10362
rect 15776 10310 15806 10362
rect 15830 10310 15840 10362
rect 15840 10310 15886 10362
rect 15910 10310 15956 10362
rect 15956 10310 15966 10362
rect 15990 10310 16020 10362
rect 16020 10310 16046 10362
rect 15750 10308 15806 10310
rect 15830 10308 15886 10310
rect 15910 10308 15966 10310
rect 15990 10308 16046 10310
rect 16118 10104 16174 10160
rect 15750 9274 15806 9276
rect 15830 9274 15886 9276
rect 15910 9274 15966 9276
rect 15990 9274 16046 9276
rect 15750 9222 15776 9274
rect 15776 9222 15806 9274
rect 15830 9222 15840 9274
rect 15840 9222 15886 9274
rect 15910 9222 15956 9274
rect 15956 9222 15966 9274
rect 15990 9222 16020 9274
rect 16020 9222 16046 9274
rect 15750 9220 15806 9222
rect 15830 9220 15886 9222
rect 15910 9220 15966 9222
rect 15990 9220 16046 9222
rect 15750 8186 15806 8188
rect 15830 8186 15886 8188
rect 15910 8186 15966 8188
rect 15990 8186 16046 8188
rect 15750 8134 15776 8186
rect 15776 8134 15806 8186
rect 15830 8134 15840 8186
rect 15840 8134 15886 8186
rect 15910 8134 15956 8186
rect 15956 8134 15966 8186
rect 15990 8134 16020 8186
rect 16020 8134 16046 8186
rect 15750 8132 15806 8134
rect 15830 8132 15886 8134
rect 15910 8132 15966 8134
rect 15990 8132 16046 8134
rect 15842 7404 15898 7440
rect 15842 7384 15844 7404
rect 15844 7384 15896 7404
rect 15896 7384 15898 7404
rect 15566 5208 15622 5264
rect 15750 7098 15806 7100
rect 15830 7098 15886 7100
rect 15910 7098 15966 7100
rect 15990 7098 16046 7100
rect 15750 7046 15776 7098
rect 15776 7046 15806 7098
rect 15830 7046 15840 7098
rect 15840 7046 15886 7098
rect 15910 7046 15956 7098
rect 15956 7046 15966 7098
rect 15990 7046 16020 7098
rect 16020 7046 16046 7098
rect 15750 7044 15806 7046
rect 15830 7044 15886 7046
rect 15910 7044 15966 7046
rect 15990 7044 16046 7046
rect 15750 6010 15806 6012
rect 15830 6010 15886 6012
rect 15910 6010 15966 6012
rect 15990 6010 16046 6012
rect 15750 5958 15776 6010
rect 15776 5958 15806 6010
rect 15830 5958 15840 6010
rect 15840 5958 15886 6010
rect 15910 5958 15956 6010
rect 15956 5958 15966 6010
rect 15990 5958 16020 6010
rect 16020 5958 16046 6010
rect 15750 5956 15806 5958
rect 15830 5956 15886 5958
rect 15910 5956 15966 5958
rect 15990 5956 16046 5958
rect 15658 5072 15714 5128
rect 15750 4922 15806 4924
rect 15830 4922 15886 4924
rect 15910 4922 15966 4924
rect 15990 4922 16046 4924
rect 15750 4870 15776 4922
rect 15776 4870 15806 4922
rect 15830 4870 15840 4922
rect 15840 4870 15886 4922
rect 15910 4870 15956 4922
rect 15956 4870 15966 4922
rect 15990 4870 16020 4922
rect 16020 4870 16046 4922
rect 15750 4868 15806 4870
rect 15830 4868 15886 4870
rect 15910 4868 15966 4870
rect 15990 4868 16046 4870
rect 15566 3596 15622 3632
rect 15566 3576 15568 3596
rect 15568 3576 15620 3596
rect 15620 3576 15622 3596
rect 15750 3834 15806 3836
rect 15830 3834 15886 3836
rect 15910 3834 15966 3836
rect 15990 3834 16046 3836
rect 15750 3782 15776 3834
rect 15776 3782 15806 3834
rect 15830 3782 15840 3834
rect 15840 3782 15886 3834
rect 15910 3782 15956 3834
rect 15956 3782 15966 3834
rect 15990 3782 16020 3834
rect 16020 3782 16046 3834
rect 15750 3780 15806 3782
rect 15830 3780 15886 3782
rect 15910 3780 15966 3782
rect 15990 3780 16046 3782
rect 16302 9968 16358 10024
rect 16302 6704 16358 6760
rect 15750 2746 15806 2748
rect 15830 2746 15886 2748
rect 15910 2746 15966 2748
rect 15990 2746 16046 2748
rect 15750 2694 15776 2746
rect 15776 2694 15806 2746
rect 15830 2694 15840 2746
rect 15840 2694 15886 2746
rect 15910 2694 15956 2746
rect 15956 2694 15966 2746
rect 15990 2694 16020 2746
rect 16020 2694 16046 2746
rect 15750 2692 15806 2694
rect 15830 2692 15886 2694
rect 15910 2692 15966 2694
rect 15990 2692 16046 2694
rect 16762 18808 16818 18864
rect 16670 17584 16726 17640
rect 16854 16632 16910 16688
rect 16578 16124 16580 16144
rect 16580 16124 16632 16144
rect 16632 16124 16634 16144
rect 16578 16088 16634 16124
rect 16854 12960 16910 13016
rect 16578 11192 16634 11248
rect 16578 7928 16634 7984
rect 16854 6432 16910 6488
rect 17130 14456 17186 14512
rect 17406 17992 17462 18048
rect 17498 17176 17554 17232
rect 17038 9696 17094 9752
rect 17038 6840 17094 6896
rect 17222 11056 17278 11112
rect 17222 10648 17278 10704
rect 17314 9424 17370 9480
rect 17222 7928 17278 7984
rect 17130 3984 17186 4040
rect 17682 15544 17738 15600
rect 17958 19216 18014 19272
rect 17958 17720 18014 17776
rect 17774 14592 17830 14648
rect 18326 15136 18382 15192
rect 17682 10920 17738 10976
rect 17866 12724 17868 12744
rect 17868 12724 17920 12744
rect 17920 12724 17922 12744
rect 17866 12688 17922 12724
rect 17866 11212 17922 11248
rect 17866 11192 17868 11212
rect 17868 11192 17920 11212
rect 17920 11192 17922 11212
rect 17774 9696 17830 9752
rect 17866 9288 17922 9344
rect 17682 5344 17738 5400
rect 17406 4528 17462 4584
rect 17314 2896 17370 2952
rect 18234 13232 18290 13288
rect 19246 23296 19302 23352
rect 19154 22616 19210 22672
rect 19062 21256 19118 21312
rect 19449 21786 19505 21788
rect 19529 21786 19585 21788
rect 19609 21786 19665 21788
rect 19689 21786 19745 21788
rect 19449 21734 19475 21786
rect 19475 21734 19505 21786
rect 19529 21734 19539 21786
rect 19539 21734 19585 21786
rect 19609 21734 19655 21786
rect 19655 21734 19665 21786
rect 19689 21734 19719 21786
rect 19719 21734 19745 21786
rect 19449 21732 19505 21734
rect 19529 21732 19585 21734
rect 19609 21732 19665 21734
rect 19689 21732 19745 21734
rect 19890 21936 19946 21992
rect 19449 20698 19505 20700
rect 19529 20698 19585 20700
rect 19609 20698 19665 20700
rect 19689 20698 19745 20700
rect 19449 20646 19475 20698
rect 19475 20646 19505 20698
rect 19529 20646 19539 20698
rect 19539 20646 19585 20698
rect 19609 20646 19655 20698
rect 19655 20646 19665 20698
rect 19689 20646 19719 20698
rect 19719 20646 19745 20698
rect 19449 20644 19505 20646
rect 19529 20644 19585 20646
rect 19609 20644 19665 20646
rect 19689 20644 19745 20646
rect 19890 20576 19946 20632
rect 19338 20032 19394 20088
rect 18786 19488 18842 19544
rect 19246 19660 19248 19680
rect 19248 19660 19300 19680
rect 19300 19660 19302 19680
rect 19246 19624 19302 19660
rect 19449 19610 19505 19612
rect 19529 19610 19585 19612
rect 19609 19610 19665 19612
rect 19689 19610 19745 19612
rect 19449 19558 19475 19610
rect 19475 19558 19505 19610
rect 19529 19558 19539 19610
rect 19539 19558 19585 19610
rect 19609 19558 19655 19610
rect 19655 19558 19665 19610
rect 19689 19558 19719 19610
rect 19719 19558 19745 19610
rect 19449 19556 19505 19558
rect 19529 19556 19585 19558
rect 19609 19556 19665 19558
rect 19689 19556 19745 19558
rect 19449 18522 19505 18524
rect 19529 18522 19585 18524
rect 19609 18522 19665 18524
rect 19689 18522 19745 18524
rect 19449 18470 19475 18522
rect 19475 18470 19505 18522
rect 19529 18470 19539 18522
rect 19539 18470 19585 18522
rect 19609 18470 19655 18522
rect 19655 18470 19665 18522
rect 19689 18470 19719 18522
rect 19719 18470 19745 18522
rect 19449 18468 19505 18470
rect 19529 18468 19585 18470
rect 19609 18468 19665 18470
rect 19689 18468 19745 18470
rect 18510 14456 18566 14512
rect 18694 13096 18750 13152
rect 18786 11872 18842 11928
rect 18326 11600 18382 11656
rect 18326 9968 18382 10024
rect 18142 9560 18198 9616
rect 18142 9016 18198 9072
rect 20534 20848 20590 20904
rect 19449 17434 19505 17436
rect 19529 17434 19585 17436
rect 19609 17434 19665 17436
rect 19689 17434 19745 17436
rect 19449 17382 19475 17434
rect 19475 17382 19505 17434
rect 19529 17382 19539 17434
rect 19539 17382 19585 17434
rect 19609 17382 19655 17434
rect 19655 17382 19665 17434
rect 19689 17382 19719 17434
rect 19719 17382 19745 17434
rect 19449 17380 19505 17382
rect 19529 17380 19585 17382
rect 19609 17380 19665 17382
rect 19689 17380 19745 17382
rect 19449 16346 19505 16348
rect 19529 16346 19585 16348
rect 19609 16346 19665 16348
rect 19689 16346 19745 16348
rect 19449 16294 19475 16346
rect 19475 16294 19505 16346
rect 19529 16294 19539 16346
rect 19539 16294 19585 16346
rect 19609 16294 19655 16346
rect 19655 16294 19665 16346
rect 19689 16294 19719 16346
rect 19719 16294 19745 16346
rect 19449 16292 19505 16294
rect 19529 16292 19585 16294
rect 19609 16292 19665 16294
rect 19689 16292 19745 16294
rect 19338 15408 19394 15464
rect 19449 15258 19505 15260
rect 19529 15258 19585 15260
rect 19609 15258 19665 15260
rect 19689 15258 19745 15260
rect 19449 15206 19475 15258
rect 19475 15206 19505 15258
rect 19529 15206 19539 15258
rect 19539 15206 19585 15258
rect 19609 15206 19655 15258
rect 19655 15206 19665 15258
rect 19689 15206 19719 15258
rect 19719 15206 19745 15258
rect 19449 15204 19505 15206
rect 19529 15204 19585 15206
rect 19609 15204 19665 15206
rect 19689 15204 19745 15206
rect 19338 15036 19340 15056
rect 19340 15036 19392 15056
rect 19392 15036 19394 15056
rect 19338 15000 19394 15036
rect 19614 14900 19616 14920
rect 19616 14900 19668 14920
rect 19668 14900 19670 14920
rect 19154 14476 19210 14512
rect 19154 14456 19156 14476
rect 19156 14456 19208 14476
rect 19208 14456 19210 14476
rect 19614 14864 19670 14900
rect 19982 15000 20038 15056
rect 19982 14728 20038 14784
rect 19449 14170 19505 14172
rect 19529 14170 19585 14172
rect 19609 14170 19665 14172
rect 19689 14170 19745 14172
rect 19449 14118 19475 14170
rect 19475 14118 19505 14170
rect 19529 14118 19539 14170
rect 19539 14118 19585 14170
rect 19609 14118 19655 14170
rect 19655 14118 19665 14170
rect 19689 14118 19719 14170
rect 19719 14118 19745 14170
rect 19449 14116 19505 14118
rect 19529 14116 19585 14118
rect 19609 14116 19665 14118
rect 19689 14116 19745 14118
rect 19062 12008 19118 12064
rect 18970 11872 19026 11928
rect 19338 13368 19394 13424
rect 19449 13082 19505 13084
rect 19529 13082 19585 13084
rect 19609 13082 19665 13084
rect 19689 13082 19745 13084
rect 19449 13030 19475 13082
rect 19475 13030 19505 13082
rect 19529 13030 19539 13082
rect 19539 13030 19585 13082
rect 19609 13030 19655 13082
rect 19655 13030 19665 13082
rect 19689 13030 19719 13082
rect 19719 13030 19745 13082
rect 19449 13028 19505 13030
rect 19529 13028 19585 13030
rect 19609 13028 19665 13030
rect 19689 13028 19745 13030
rect 18694 9560 18750 9616
rect 19890 12824 19946 12880
rect 20442 20304 20498 20360
rect 20626 19352 20682 19408
rect 20166 17584 20222 17640
rect 20350 18128 20406 18184
rect 20350 18028 20352 18048
rect 20352 18028 20404 18048
rect 20404 18028 20406 18048
rect 20350 17992 20406 18028
rect 20074 12552 20130 12608
rect 20074 12416 20130 12472
rect 20442 14048 20498 14104
rect 19449 11994 19505 11996
rect 19529 11994 19585 11996
rect 19609 11994 19665 11996
rect 19689 11994 19745 11996
rect 19449 11942 19475 11994
rect 19475 11942 19505 11994
rect 19529 11942 19539 11994
rect 19539 11942 19585 11994
rect 19609 11942 19655 11994
rect 19655 11942 19665 11994
rect 19689 11942 19719 11994
rect 19719 11942 19745 11994
rect 19449 11940 19505 11942
rect 19529 11940 19585 11942
rect 19609 11940 19665 11942
rect 19689 11940 19745 11942
rect 19706 11756 19762 11792
rect 19706 11736 19708 11756
rect 19708 11736 19760 11756
rect 19760 11736 19762 11756
rect 19154 11464 19210 11520
rect 19062 11056 19118 11112
rect 18970 9832 19026 9888
rect 19449 10906 19505 10908
rect 19529 10906 19585 10908
rect 19609 10906 19665 10908
rect 19689 10906 19745 10908
rect 19449 10854 19475 10906
rect 19475 10854 19505 10906
rect 19529 10854 19539 10906
rect 19539 10854 19585 10906
rect 19609 10854 19655 10906
rect 19655 10854 19665 10906
rect 19689 10854 19719 10906
rect 19719 10854 19745 10906
rect 19449 10852 19505 10854
rect 19529 10852 19585 10854
rect 19609 10852 19665 10854
rect 19689 10852 19745 10854
rect 20074 11328 20130 11384
rect 19706 10004 19708 10024
rect 19708 10004 19760 10024
rect 19760 10004 19762 10024
rect 19706 9968 19762 10004
rect 19449 9818 19505 9820
rect 19529 9818 19585 9820
rect 19609 9818 19665 9820
rect 19689 9818 19745 9820
rect 19449 9766 19475 9818
rect 19475 9766 19505 9818
rect 19529 9766 19539 9818
rect 19539 9766 19585 9818
rect 19609 9766 19655 9818
rect 19655 9766 19665 9818
rect 19689 9766 19719 9818
rect 19719 9766 19745 9818
rect 19449 9764 19505 9766
rect 19529 9764 19585 9766
rect 19609 9764 19665 9766
rect 19689 9764 19745 9766
rect 19338 9560 19394 9616
rect 18510 9152 18566 9208
rect 18602 7692 18604 7712
rect 18604 7692 18656 7712
rect 18656 7692 18658 7712
rect 18050 7384 18106 7440
rect 18602 7656 18658 7692
rect 18418 7404 18474 7440
rect 18418 7384 18420 7404
rect 18420 7384 18472 7404
rect 18472 7384 18474 7404
rect 18878 9016 18934 9072
rect 19154 9288 19210 9344
rect 19062 9016 19118 9072
rect 19706 9424 19762 9480
rect 19246 9152 19302 9208
rect 18878 8608 18934 8664
rect 19338 8880 19394 8936
rect 19246 8744 19302 8800
rect 19246 7248 19302 7304
rect 18418 4120 18474 4176
rect 19449 8730 19505 8732
rect 19529 8730 19585 8732
rect 19609 8730 19665 8732
rect 19689 8730 19745 8732
rect 19449 8678 19475 8730
rect 19475 8678 19505 8730
rect 19529 8678 19539 8730
rect 19539 8678 19585 8730
rect 19609 8678 19655 8730
rect 19655 8678 19665 8730
rect 19689 8678 19719 8730
rect 19719 8678 19745 8730
rect 19449 8676 19505 8678
rect 19529 8676 19585 8678
rect 19609 8676 19665 8678
rect 19689 8676 19745 8678
rect 19890 9016 19946 9072
rect 19449 7642 19505 7644
rect 19529 7642 19585 7644
rect 19609 7642 19665 7644
rect 19689 7642 19745 7644
rect 19449 7590 19475 7642
rect 19475 7590 19505 7642
rect 19529 7590 19539 7642
rect 19539 7590 19585 7642
rect 19609 7590 19655 7642
rect 19655 7590 19665 7642
rect 19689 7590 19719 7642
rect 19719 7590 19745 7642
rect 19449 7588 19505 7590
rect 19529 7588 19585 7590
rect 19609 7588 19665 7590
rect 19689 7588 19745 7590
rect 19449 6554 19505 6556
rect 19529 6554 19585 6556
rect 19609 6554 19665 6556
rect 19689 6554 19745 6556
rect 19449 6502 19475 6554
rect 19475 6502 19505 6554
rect 19529 6502 19539 6554
rect 19539 6502 19585 6554
rect 19609 6502 19655 6554
rect 19655 6502 19665 6554
rect 19689 6502 19719 6554
rect 19719 6502 19745 6554
rect 19449 6500 19505 6502
rect 19529 6500 19585 6502
rect 19609 6500 19665 6502
rect 19689 6500 19745 6502
rect 19154 5616 19210 5672
rect 20994 16088 21050 16144
rect 20810 14592 20866 14648
rect 20534 12416 20590 12472
rect 20350 11736 20406 11792
rect 20258 10104 20314 10160
rect 20166 9016 20222 9072
rect 19449 5466 19505 5468
rect 19529 5466 19585 5468
rect 19609 5466 19665 5468
rect 19689 5466 19745 5468
rect 19449 5414 19475 5466
rect 19475 5414 19505 5466
rect 19529 5414 19539 5466
rect 19539 5414 19585 5466
rect 19609 5414 19655 5466
rect 19655 5414 19665 5466
rect 19689 5414 19719 5466
rect 19719 5414 19745 5466
rect 19449 5412 19505 5414
rect 19529 5412 19585 5414
rect 19609 5412 19665 5414
rect 19689 5412 19745 5414
rect 19430 5108 19432 5128
rect 19432 5108 19484 5128
rect 19484 5108 19486 5128
rect 19430 5072 19486 5108
rect 19246 4256 19302 4312
rect 17958 3576 18014 3632
rect 18326 2488 18382 2544
rect 20074 6704 20130 6760
rect 20258 7384 20314 7440
rect 19890 4800 19946 4856
rect 19449 4378 19505 4380
rect 19529 4378 19585 4380
rect 19609 4378 19665 4380
rect 19689 4378 19745 4380
rect 19449 4326 19475 4378
rect 19475 4326 19505 4378
rect 19529 4326 19539 4378
rect 19539 4326 19585 4378
rect 19609 4326 19655 4378
rect 19655 4326 19665 4378
rect 19689 4326 19719 4378
rect 19719 4326 19745 4378
rect 19449 4324 19505 4326
rect 19529 4324 19585 4326
rect 19609 4324 19665 4326
rect 19689 4324 19745 4326
rect 19449 3290 19505 3292
rect 19529 3290 19585 3292
rect 19609 3290 19665 3292
rect 19689 3290 19745 3292
rect 19449 3238 19475 3290
rect 19475 3238 19505 3290
rect 19529 3238 19539 3290
rect 19539 3238 19585 3290
rect 19609 3238 19655 3290
rect 19655 3238 19665 3290
rect 19689 3238 19719 3290
rect 19719 3238 19745 3290
rect 19449 3236 19505 3238
rect 19529 3236 19585 3238
rect 19609 3236 19665 3238
rect 19689 3236 19745 3238
rect 20074 5208 20130 5264
rect 20994 14456 21050 14512
rect 20626 10648 20682 10704
rect 20350 5652 20352 5672
rect 20352 5652 20404 5672
rect 20404 5652 20406 5672
rect 20350 5616 20406 5652
rect 20166 4256 20222 4312
rect 20810 10784 20866 10840
rect 20718 7384 20774 7440
rect 20626 7112 20682 7168
rect 20534 3576 20590 3632
rect 20994 7948 21050 7984
rect 20994 7928 20996 7948
rect 20996 7928 21048 7948
rect 21048 7928 21050 7948
rect 20994 7520 21050 7576
rect 22006 18672 22062 18728
rect 22190 17992 22246 18048
rect 21454 10512 21510 10568
rect 21270 9424 21326 9480
rect 21270 8200 21326 8256
rect 20994 6296 21050 6352
rect 20718 5108 20720 5128
rect 20720 5108 20772 5128
rect 20772 5108 20774 5128
rect 20718 5072 20774 5108
rect 19890 2216 19946 2272
rect 19449 2202 19505 2204
rect 19529 2202 19585 2204
rect 19609 2202 19665 2204
rect 19689 2202 19745 2204
rect 19449 2150 19475 2202
rect 19475 2150 19505 2202
rect 19529 2150 19539 2202
rect 19539 2150 19585 2202
rect 19609 2150 19655 2202
rect 19655 2150 19665 2202
rect 19689 2150 19719 2202
rect 19719 2150 19745 2202
rect 19449 2148 19505 2150
rect 19529 2148 19585 2150
rect 19609 2148 19665 2150
rect 19689 2148 19745 2150
rect 21454 7520 21510 7576
rect 21362 5208 21418 5264
rect 21730 12144 21786 12200
rect 22558 17312 22614 17368
rect 22466 16632 22522 16688
rect 22374 12688 22430 12744
rect 22098 5208 22154 5264
rect 22006 4120 22062 4176
rect 21822 3032 21878 3088
rect 21730 2896 21786 2952
rect 22466 8744 22522 8800
rect 22466 6160 22522 6216
rect 22742 6840 22798 6896
rect 22374 4120 22430 4176
rect 22098 1536 22154 1592
rect 19338 856 19394 912
rect 23386 11056 23442 11112
rect 22834 5480 22890 5536
rect 22650 312 22706 368
<< metal3 >>
rect 19793 24034 19859 24037
rect 23920 24034 24400 24064
rect 19793 24032 24400 24034
rect 19793 23976 19798 24032
rect 19854 23976 24400 24032
rect 19793 23974 24400 23976
rect 19793 23971 19859 23974
rect 23920 23944 24400 23974
rect 19241 23354 19307 23357
rect 23920 23354 24400 23384
rect 19241 23352 24400 23354
rect 19241 23296 19246 23352
rect 19302 23296 24400 23352
rect 19241 23294 24400 23296
rect 19241 23291 19307 23294
rect 23920 23264 24400 23294
rect 19149 22674 19215 22677
rect 23920 22674 24400 22704
rect 19149 22672 24400 22674
rect 19149 22616 19154 22672
rect 19210 22616 24400 22672
rect 19149 22614 24400 22616
rect 19149 22611 19215 22614
rect 23920 22584 24400 22614
rect 19885 21994 19951 21997
rect 23920 21994 24400 22024
rect 19885 21992 24400 21994
rect 19885 21936 19890 21992
rect 19946 21936 24400 21992
rect 19885 21934 24400 21936
rect 19885 21931 19951 21934
rect 23920 21904 24400 21934
rect 4642 21792 4962 21793
rect 4642 21728 4650 21792
rect 4714 21728 4730 21792
rect 4794 21728 4810 21792
rect 4874 21728 4890 21792
rect 4954 21728 4962 21792
rect 4642 21727 4962 21728
rect 12040 21792 12360 21793
rect 12040 21728 12048 21792
rect 12112 21728 12128 21792
rect 12192 21728 12208 21792
rect 12272 21728 12288 21792
rect 12352 21728 12360 21792
rect 12040 21727 12360 21728
rect 19437 21792 19757 21793
rect 19437 21728 19445 21792
rect 19509 21728 19525 21792
rect 19589 21728 19605 21792
rect 19669 21728 19685 21792
rect 19749 21728 19757 21792
rect 19437 21727 19757 21728
rect 0 21314 480 21344
rect 3877 21314 3943 21317
rect 0 21312 3943 21314
rect 0 21256 3882 21312
rect 3938 21256 3943 21312
rect 0 21254 3943 21256
rect 0 21224 480 21254
rect 3877 21251 3943 21254
rect 19057 21314 19123 21317
rect 23920 21314 24400 21344
rect 19057 21312 24400 21314
rect 19057 21256 19062 21312
rect 19118 21256 24400 21312
rect 19057 21254 24400 21256
rect 19057 21251 19123 21254
rect 8341 21248 8661 21249
rect 8341 21184 8349 21248
rect 8413 21184 8429 21248
rect 8493 21184 8509 21248
rect 8573 21184 8589 21248
rect 8653 21184 8661 21248
rect 8341 21183 8661 21184
rect 15738 21248 16058 21249
rect 15738 21184 15746 21248
rect 15810 21184 15826 21248
rect 15890 21184 15906 21248
rect 15970 21184 15986 21248
rect 16050 21184 16058 21248
rect 23920 21224 24400 21254
rect 15738 21183 16058 21184
rect 14222 20844 14228 20908
rect 14292 20906 14298 20908
rect 20529 20906 20595 20909
rect 14292 20904 20595 20906
rect 14292 20848 20534 20904
rect 20590 20848 20595 20904
rect 14292 20846 20595 20848
rect 14292 20844 14298 20846
rect 20529 20843 20595 20846
rect 4642 20704 4962 20705
rect 4642 20640 4650 20704
rect 4714 20640 4730 20704
rect 4794 20640 4810 20704
rect 4874 20640 4890 20704
rect 4954 20640 4962 20704
rect 4642 20639 4962 20640
rect 12040 20704 12360 20705
rect 12040 20640 12048 20704
rect 12112 20640 12128 20704
rect 12192 20640 12208 20704
rect 12272 20640 12288 20704
rect 12352 20640 12360 20704
rect 12040 20639 12360 20640
rect 19437 20704 19757 20705
rect 19437 20640 19445 20704
rect 19509 20640 19525 20704
rect 19589 20640 19605 20704
rect 19669 20640 19685 20704
rect 19749 20640 19757 20704
rect 19437 20639 19757 20640
rect 19885 20634 19951 20637
rect 23920 20634 24400 20664
rect 19885 20632 24400 20634
rect 19885 20576 19890 20632
rect 19946 20576 24400 20632
rect 19885 20574 24400 20576
rect 19885 20571 19951 20574
rect 23920 20544 24400 20574
rect 15326 20300 15332 20364
rect 15396 20362 15402 20364
rect 16297 20362 16363 20365
rect 20437 20362 20503 20365
rect 15396 20360 20503 20362
rect 15396 20304 16302 20360
rect 16358 20304 20442 20360
rect 20498 20304 20503 20360
rect 15396 20302 20503 20304
rect 15396 20300 15402 20302
rect 16297 20299 16363 20302
rect 20437 20299 20503 20302
rect 8341 20160 8661 20161
rect 8341 20096 8349 20160
rect 8413 20096 8429 20160
rect 8493 20096 8509 20160
rect 8573 20096 8589 20160
rect 8653 20096 8661 20160
rect 8341 20095 8661 20096
rect 15738 20160 16058 20161
rect 15738 20096 15746 20160
rect 15810 20096 15826 20160
rect 15890 20096 15906 20160
rect 15970 20096 15986 20160
rect 16050 20096 16058 20160
rect 15738 20095 16058 20096
rect 19333 20090 19399 20093
rect 23920 20090 24400 20120
rect 19333 20088 24400 20090
rect 19333 20032 19338 20088
rect 19394 20032 24400 20088
rect 19333 20030 24400 20032
rect 19333 20027 19399 20030
rect 23920 20000 24400 20030
rect 4981 19954 5047 19957
rect 15653 19954 15719 19957
rect 4981 19952 15719 19954
rect 4981 19896 4986 19952
rect 5042 19896 15658 19952
rect 15714 19896 15719 19952
rect 4981 19894 15719 19896
rect 4981 19891 5047 19894
rect 15653 19891 15719 19894
rect 4061 19818 4127 19821
rect 4429 19818 4495 19821
rect 9029 19818 9095 19821
rect 4061 19816 9095 19818
rect 4061 19760 4066 19816
rect 4122 19760 4434 19816
rect 4490 19760 9034 19816
rect 9090 19760 9095 19816
rect 4061 19758 9095 19760
rect 4061 19755 4127 19758
rect 4429 19755 4495 19758
rect 9029 19755 9095 19758
rect 14406 19620 14412 19684
rect 14476 19682 14482 19684
rect 19241 19682 19307 19685
rect 14476 19680 19307 19682
rect 14476 19624 19246 19680
rect 19302 19624 19307 19680
rect 14476 19622 19307 19624
rect 14476 19620 14482 19622
rect 19241 19619 19307 19622
rect 4642 19616 4962 19617
rect 4642 19552 4650 19616
rect 4714 19552 4730 19616
rect 4794 19552 4810 19616
rect 4874 19552 4890 19616
rect 4954 19552 4962 19616
rect 4642 19551 4962 19552
rect 12040 19616 12360 19617
rect 12040 19552 12048 19616
rect 12112 19552 12128 19616
rect 12192 19552 12208 19616
rect 12272 19552 12288 19616
rect 12352 19552 12360 19616
rect 12040 19551 12360 19552
rect 19437 19616 19757 19617
rect 19437 19552 19445 19616
rect 19509 19552 19525 19616
rect 19589 19552 19605 19616
rect 19669 19552 19685 19616
rect 19749 19552 19757 19616
rect 19437 19551 19757 19552
rect 6085 19546 6151 19549
rect 6678 19546 6684 19548
rect 6085 19544 6684 19546
rect 6085 19488 6090 19544
rect 6146 19488 6684 19544
rect 6085 19486 6684 19488
rect 6085 19483 6151 19486
rect 6678 19484 6684 19486
rect 6748 19546 6754 19548
rect 10133 19546 10199 19549
rect 6748 19544 10199 19546
rect 6748 19488 10138 19544
rect 10194 19488 10199 19544
rect 6748 19486 10199 19488
rect 6748 19484 6754 19486
rect 10133 19483 10199 19486
rect 12525 19546 12591 19549
rect 18781 19546 18847 19549
rect 12525 19544 18847 19546
rect 12525 19488 12530 19544
rect 12586 19488 18786 19544
rect 18842 19488 18847 19544
rect 12525 19486 18847 19488
rect 12525 19483 12591 19486
rect 18781 19483 18847 19486
rect 13077 19410 13143 19413
rect 13905 19410 13971 19413
rect 16113 19410 16179 19413
rect 13077 19408 16179 19410
rect 13077 19352 13082 19408
rect 13138 19352 13910 19408
rect 13966 19352 16118 19408
rect 16174 19352 16179 19408
rect 13077 19350 16179 19352
rect 13077 19347 13143 19350
rect 13905 19347 13971 19350
rect 16113 19347 16179 19350
rect 20621 19410 20687 19413
rect 23920 19410 24400 19440
rect 20621 19408 24400 19410
rect 20621 19352 20626 19408
rect 20682 19352 24400 19408
rect 20621 19350 24400 19352
rect 20621 19347 20687 19350
rect 23920 19320 24400 19350
rect 2773 19274 2839 19277
rect 2957 19274 3023 19277
rect 2773 19272 3023 19274
rect 2773 19216 2778 19272
rect 2834 19216 2962 19272
rect 3018 19216 3023 19272
rect 2773 19214 3023 19216
rect 2773 19211 2839 19214
rect 2957 19211 3023 19214
rect 7189 19274 7255 19277
rect 12617 19274 12683 19277
rect 7189 19272 12683 19274
rect 7189 19216 7194 19272
rect 7250 19216 12622 19272
rect 12678 19216 12683 19272
rect 7189 19214 12683 19216
rect 7189 19211 7255 19214
rect 12617 19211 12683 19214
rect 15009 19274 15075 19277
rect 17953 19274 18019 19277
rect 15009 19272 18019 19274
rect 15009 19216 15014 19272
rect 15070 19216 17958 19272
rect 18014 19216 18019 19272
rect 15009 19214 18019 19216
rect 15009 19211 15075 19214
rect 17953 19211 18019 19214
rect 11646 19076 11652 19140
rect 11716 19138 11722 19140
rect 12341 19138 12407 19141
rect 11716 19136 12407 19138
rect 11716 19080 12346 19136
rect 12402 19080 12407 19136
rect 11716 19078 12407 19080
rect 11716 19076 11722 19078
rect 12341 19075 12407 19078
rect 8341 19072 8661 19073
rect 8341 19008 8349 19072
rect 8413 19008 8429 19072
rect 8493 19008 8509 19072
rect 8573 19008 8589 19072
rect 8653 19008 8661 19072
rect 8341 19007 8661 19008
rect 15738 19072 16058 19073
rect 15738 19008 15746 19072
rect 15810 19008 15826 19072
rect 15890 19008 15906 19072
rect 15970 19008 15986 19072
rect 16050 19008 16058 19072
rect 15738 19007 16058 19008
rect 9581 18866 9647 18869
rect 16757 18866 16823 18869
rect 9581 18864 16823 18866
rect 9581 18808 9586 18864
rect 9642 18808 16762 18864
rect 16818 18808 16823 18864
rect 9581 18806 16823 18808
rect 9581 18803 9647 18806
rect 16757 18803 16823 18806
rect 15101 18730 15167 18733
rect 16573 18730 16639 18733
rect 15101 18728 16639 18730
rect 15101 18672 15106 18728
rect 15162 18672 16578 18728
rect 16634 18672 16639 18728
rect 15101 18670 16639 18672
rect 15101 18667 15167 18670
rect 16573 18667 16639 18670
rect 22001 18730 22067 18733
rect 23920 18730 24400 18760
rect 22001 18728 24400 18730
rect 22001 18672 22006 18728
rect 22062 18672 24400 18728
rect 22001 18670 24400 18672
rect 22001 18667 22067 18670
rect 23920 18640 24400 18670
rect 5809 18594 5875 18597
rect 10777 18594 10843 18597
rect 5809 18592 10843 18594
rect 5809 18536 5814 18592
rect 5870 18536 10782 18592
rect 10838 18536 10843 18592
rect 5809 18534 10843 18536
rect 5809 18531 5875 18534
rect 10777 18531 10843 18534
rect 4642 18528 4962 18529
rect 4642 18464 4650 18528
rect 4714 18464 4730 18528
rect 4794 18464 4810 18528
rect 4874 18464 4890 18528
rect 4954 18464 4962 18528
rect 4642 18463 4962 18464
rect 12040 18528 12360 18529
rect 12040 18464 12048 18528
rect 12112 18464 12128 18528
rect 12192 18464 12208 18528
rect 12272 18464 12288 18528
rect 12352 18464 12360 18528
rect 12040 18463 12360 18464
rect 19437 18528 19757 18529
rect 19437 18464 19445 18528
rect 19509 18464 19525 18528
rect 19589 18464 19605 18528
rect 19669 18464 19685 18528
rect 19749 18464 19757 18528
rect 19437 18463 19757 18464
rect 8385 18458 8451 18461
rect 8661 18458 8727 18461
rect 9765 18458 9831 18461
rect 8385 18456 9831 18458
rect 8385 18400 8390 18456
rect 8446 18400 8666 18456
rect 8722 18400 9770 18456
rect 9826 18400 9831 18456
rect 8385 18398 9831 18400
rect 8385 18395 8451 18398
rect 8661 18395 8727 18398
rect 9765 18395 9831 18398
rect 1485 18322 1551 18325
rect 7189 18322 7255 18325
rect 1485 18320 7255 18322
rect 1485 18264 1490 18320
rect 1546 18264 7194 18320
rect 7250 18264 7255 18320
rect 1485 18262 7255 18264
rect 1485 18259 1551 18262
rect 7189 18259 7255 18262
rect 9581 18322 9647 18325
rect 15469 18322 15535 18325
rect 9581 18320 15535 18322
rect 9581 18264 9586 18320
rect 9642 18264 15474 18320
rect 15530 18264 15535 18320
rect 9581 18262 15535 18264
rect 9581 18259 9647 18262
rect 15469 18259 15535 18262
rect 14038 18124 14044 18188
rect 14108 18186 14114 18188
rect 20345 18186 20411 18189
rect 14108 18184 20411 18186
rect 14108 18128 20350 18184
rect 20406 18128 20411 18184
rect 14108 18126 20411 18128
rect 14108 18124 14114 18126
rect 20345 18123 20411 18126
rect 4429 18052 4495 18053
rect 4429 18048 4476 18052
rect 4540 18050 4546 18052
rect 8937 18050 9003 18053
rect 17401 18050 17467 18053
rect 20345 18052 20411 18053
rect 17534 18050 17540 18052
rect 4429 17992 4434 18048
rect 4429 17988 4476 17992
rect 4540 17990 4586 18050
rect 8937 18048 9736 18050
rect 8937 17992 8942 18048
rect 8998 17992 9736 18048
rect 8937 17990 9736 17992
rect 4540 17988 4546 17990
rect 4429 17987 4495 17988
rect 8937 17987 9003 17990
rect 8341 17984 8661 17985
rect 8341 17920 8349 17984
rect 8413 17920 8429 17984
rect 8493 17920 8509 17984
rect 8573 17920 8589 17984
rect 8653 17920 8661 17984
rect 8341 17919 8661 17920
rect 2681 17778 2747 17781
rect 4061 17778 4127 17781
rect 2681 17776 4127 17778
rect 2681 17720 2686 17776
rect 2742 17720 4066 17776
rect 4122 17720 4127 17776
rect 2681 17718 4127 17720
rect 9676 17778 9736 17990
rect 17401 18048 17540 18050
rect 17401 17992 17406 18048
rect 17462 17992 17540 18048
rect 17401 17990 17540 17992
rect 17401 17987 17467 17990
rect 17534 17988 17540 17990
rect 17604 17988 17610 18052
rect 20294 17988 20300 18052
rect 20364 18050 20411 18052
rect 22185 18050 22251 18053
rect 23920 18050 24400 18080
rect 20364 18048 20456 18050
rect 20406 17992 20456 18048
rect 20364 17990 20456 17992
rect 22185 18048 24400 18050
rect 22185 17992 22190 18048
rect 22246 17992 24400 18048
rect 22185 17990 24400 17992
rect 20364 17988 20411 17990
rect 20345 17987 20411 17988
rect 22185 17987 22251 17990
rect 15738 17984 16058 17985
rect 15738 17920 15746 17984
rect 15810 17920 15826 17984
rect 15890 17920 15906 17984
rect 15970 17920 15986 17984
rect 16050 17920 16058 17984
rect 23920 17960 24400 17990
rect 15738 17919 16058 17920
rect 17953 17778 18019 17781
rect 9676 17776 18019 17778
rect 9676 17720 17958 17776
rect 18014 17720 18019 17776
rect 9676 17718 18019 17720
rect 2681 17715 2747 17718
rect 4061 17715 4127 17718
rect 17953 17715 18019 17718
rect 4797 17642 4863 17645
rect 5717 17642 5783 17645
rect 4797 17640 5783 17642
rect 4797 17584 4802 17640
rect 4858 17584 5722 17640
rect 5778 17584 5783 17640
rect 4797 17582 5783 17584
rect 4797 17579 4863 17582
rect 5717 17579 5783 17582
rect 12433 17642 12499 17645
rect 16665 17642 16731 17645
rect 12433 17640 16731 17642
rect 12433 17584 12438 17640
rect 12494 17584 16670 17640
rect 16726 17584 16731 17640
rect 12433 17582 16731 17584
rect 12433 17579 12499 17582
rect 16665 17579 16731 17582
rect 19190 17580 19196 17644
rect 19260 17642 19266 17644
rect 20161 17642 20227 17645
rect 19260 17640 20227 17642
rect 19260 17584 20166 17640
rect 20222 17584 20227 17640
rect 19260 17582 20227 17584
rect 19260 17580 19266 17582
rect 20161 17579 20227 17582
rect 7833 17506 7899 17509
rect 7966 17506 7972 17508
rect 7833 17504 7972 17506
rect 7833 17448 7838 17504
rect 7894 17448 7972 17504
rect 7833 17446 7972 17448
rect 7833 17443 7899 17446
rect 7966 17444 7972 17446
rect 8036 17444 8042 17508
rect 4642 17440 4962 17441
rect 4642 17376 4650 17440
rect 4714 17376 4730 17440
rect 4794 17376 4810 17440
rect 4874 17376 4890 17440
rect 4954 17376 4962 17440
rect 4642 17375 4962 17376
rect 12040 17440 12360 17441
rect 12040 17376 12048 17440
rect 12112 17376 12128 17440
rect 12192 17376 12208 17440
rect 12272 17376 12288 17440
rect 12352 17376 12360 17440
rect 12040 17375 12360 17376
rect 19437 17440 19757 17441
rect 19437 17376 19445 17440
rect 19509 17376 19525 17440
rect 19589 17376 19605 17440
rect 19669 17376 19685 17440
rect 19749 17376 19757 17440
rect 19437 17375 19757 17376
rect 4061 17370 4127 17373
rect 22553 17370 22619 17373
rect 23920 17370 24400 17400
rect 4061 17368 4492 17370
rect 4061 17312 4066 17368
rect 4122 17312 4492 17368
rect 4061 17310 4492 17312
rect 4061 17307 4127 17310
rect 4432 17237 4492 17310
rect 22553 17368 24400 17370
rect 22553 17312 22558 17368
rect 22614 17312 24400 17368
rect 22553 17310 24400 17312
rect 22553 17307 22619 17310
rect 23920 17280 24400 17310
rect 3693 17234 3759 17237
rect 4245 17234 4311 17237
rect 3693 17232 4311 17234
rect 3693 17176 3698 17232
rect 3754 17176 4250 17232
rect 4306 17176 4311 17232
rect 3693 17174 4311 17176
rect 3693 17171 3759 17174
rect 4245 17171 4311 17174
rect 4429 17232 4495 17237
rect 4429 17176 4434 17232
rect 4490 17176 4495 17232
rect 4429 17171 4495 17176
rect 8569 17234 8635 17237
rect 8886 17234 8892 17236
rect 8569 17232 8892 17234
rect 8569 17176 8574 17232
rect 8630 17176 8892 17232
rect 8569 17174 8892 17176
rect 8569 17171 8635 17174
rect 8886 17172 8892 17174
rect 8956 17172 8962 17236
rect 9673 17234 9739 17237
rect 17493 17234 17559 17237
rect 9673 17232 17559 17234
rect 9673 17176 9678 17232
rect 9734 17176 17498 17232
rect 17554 17176 17559 17232
rect 9673 17174 17559 17176
rect 9673 17171 9739 17174
rect 17493 17171 17559 17174
rect 4061 17098 4127 17101
rect 5533 17098 5599 17101
rect 8845 17098 8911 17101
rect 4061 17096 5599 17098
rect 4061 17040 4066 17096
rect 4122 17040 5538 17096
rect 5594 17040 5599 17096
rect 4061 17038 5599 17040
rect 4061 17035 4127 17038
rect 5533 17035 5599 17038
rect 8204 17096 8911 17098
rect 8204 17040 8850 17096
rect 8906 17040 8911 17096
rect 8204 17038 8911 17040
rect 4061 16962 4127 16965
rect 8204 16962 8264 17038
rect 8845 17035 8911 17038
rect 12249 17098 12315 17101
rect 13445 17098 13511 17101
rect 12249 17096 13511 17098
rect 12249 17040 12254 17096
rect 12310 17040 13450 17096
rect 13506 17040 13511 17096
rect 12249 17038 13511 17040
rect 12249 17035 12315 17038
rect 13445 17035 13511 17038
rect 14917 17098 14983 17101
rect 15653 17098 15719 17101
rect 14917 17096 15719 17098
rect 14917 17040 14922 17096
rect 14978 17040 15658 17096
rect 15714 17040 15719 17096
rect 14917 17038 15719 17040
rect 14917 17035 14983 17038
rect 15653 17035 15719 17038
rect 4061 16960 8264 16962
rect 4061 16904 4066 16960
rect 4122 16904 8264 16960
rect 4061 16902 8264 16904
rect 4061 16899 4127 16902
rect 8341 16896 8661 16897
rect 8341 16832 8349 16896
rect 8413 16832 8429 16896
rect 8493 16832 8509 16896
rect 8573 16832 8589 16896
rect 8653 16832 8661 16896
rect 8341 16831 8661 16832
rect 15738 16896 16058 16897
rect 15738 16832 15746 16896
rect 15810 16832 15826 16896
rect 15890 16832 15906 16896
rect 15970 16832 15986 16896
rect 16050 16832 16058 16896
rect 15738 16831 16058 16832
rect 3325 16826 3391 16829
rect 4705 16826 4771 16829
rect 3325 16824 4771 16826
rect 3325 16768 3330 16824
rect 3386 16768 4710 16824
rect 4766 16768 4771 16824
rect 3325 16766 4771 16768
rect 3325 16763 3391 16766
rect 4705 16763 4771 16766
rect 5993 16826 6059 16829
rect 7189 16826 7255 16829
rect 5993 16824 7255 16826
rect 5993 16768 5998 16824
rect 6054 16768 7194 16824
rect 7250 16768 7255 16824
rect 5993 16766 7255 16768
rect 5993 16763 6059 16766
rect 7189 16763 7255 16766
rect 9949 16826 10015 16829
rect 14089 16826 14155 16829
rect 9949 16824 14155 16826
rect 9949 16768 9954 16824
rect 10010 16768 14094 16824
rect 14150 16768 14155 16824
rect 9949 16766 14155 16768
rect 9949 16763 10015 16766
rect 14089 16763 14155 16766
rect 3141 16690 3207 16693
rect 8845 16690 8911 16693
rect 3141 16688 8911 16690
rect 3141 16632 3146 16688
rect 3202 16632 8850 16688
rect 8906 16632 8911 16688
rect 3141 16630 8911 16632
rect 3141 16627 3207 16630
rect 8845 16627 8911 16630
rect 11237 16690 11303 16693
rect 16849 16690 16915 16693
rect 11237 16688 16915 16690
rect 11237 16632 11242 16688
rect 11298 16632 16854 16688
rect 16910 16632 16915 16688
rect 11237 16630 16915 16632
rect 11237 16627 11303 16630
rect 16849 16627 16915 16630
rect 22461 16690 22527 16693
rect 23920 16690 24400 16720
rect 22461 16688 24400 16690
rect 22461 16632 22466 16688
rect 22522 16632 24400 16688
rect 22461 16630 24400 16632
rect 22461 16627 22527 16630
rect 23920 16600 24400 16630
rect 4429 16554 4495 16557
rect 9305 16554 9371 16557
rect 4429 16552 9371 16554
rect 4429 16496 4434 16552
rect 4490 16496 9310 16552
rect 9366 16496 9371 16552
rect 4429 16494 9371 16496
rect 4429 16491 4495 16494
rect 9305 16491 9371 16494
rect 10225 16554 10291 16557
rect 11329 16554 11395 16557
rect 10225 16552 11395 16554
rect 10225 16496 10230 16552
rect 10286 16496 11334 16552
rect 11390 16496 11395 16552
rect 10225 16494 11395 16496
rect 10225 16491 10291 16494
rect 11329 16491 11395 16494
rect 16297 16416 16363 16421
rect 16297 16360 16302 16416
rect 16358 16360 16363 16416
rect 16297 16355 16363 16360
rect 4642 16352 4962 16353
rect 4642 16288 4650 16352
rect 4714 16288 4730 16352
rect 4794 16288 4810 16352
rect 4874 16288 4890 16352
rect 4954 16288 4962 16352
rect 4642 16287 4962 16288
rect 12040 16352 12360 16353
rect 12040 16288 12048 16352
rect 12112 16288 12128 16352
rect 12192 16288 12208 16352
rect 12272 16288 12288 16352
rect 12352 16288 12360 16352
rect 12040 16287 12360 16288
rect 16300 16282 16360 16355
rect 19437 16352 19757 16353
rect 19437 16288 19445 16352
rect 19509 16288 19525 16352
rect 19589 16288 19605 16352
rect 19669 16288 19685 16352
rect 19749 16288 19757 16352
rect 19437 16287 19757 16288
rect 12436 16222 16360 16282
rect 5533 16146 5599 16149
rect 9121 16146 9187 16149
rect 5533 16144 9187 16146
rect 5533 16088 5538 16144
rect 5594 16088 9126 16144
rect 9182 16088 9187 16144
rect 5533 16086 9187 16088
rect 5533 16083 5599 16086
rect 9121 16083 9187 16086
rect 11830 16084 11836 16148
rect 11900 16146 11906 16148
rect 12436 16146 12496 16222
rect 11900 16086 12496 16146
rect 12617 16146 12683 16149
rect 12985 16146 13051 16149
rect 16573 16146 16639 16149
rect 12617 16144 16639 16146
rect 12617 16088 12622 16144
rect 12678 16088 12990 16144
rect 13046 16088 16578 16144
rect 16634 16088 16639 16144
rect 12617 16086 16639 16088
rect 11900 16084 11906 16086
rect 12617 16083 12683 16086
rect 12985 16083 13051 16086
rect 16573 16083 16639 16086
rect 20989 16146 21055 16149
rect 23920 16146 24400 16176
rect 20989 16144 24400 16146
rect 20989 16088 20994 16144
rect 21050 16088 24400 16144
rect 20989 16086 24400 16088
rect 20989 16083 21055 16086
rect 23920 16056 24400 16086
rect 13670 15812 13676 15876
rect 13740 15874 13746 15876
rect 15193 15874 15259 15877
rect 13740 15872 15259 15874
rect 13740 15816 15198 15872
rect 15254 15816 15259 15872
rect 13740 15814 15259 15816
rect 13740 15812 13746 15814
rect 15193 15811 15259 15814
rect 8341 15808 8661 15809
rect 8341 15744 8349 15808
rect 8413 15744 8429 15808
rect 8493 15744 8509 15808
rect 8573 15744 8589 15808
rect 8653 15744 8661 15808
rect 8341 15743 8661 15744
rect 15738 15808 16058 15809
rect 15738 15744 15746 15808
rect 15810 15744 15826 15808
rect 15890 15744 15906 15808
rect 15970 15744 15986 15808
rect 16050 15744 16058 15808
rect 15738 15743 16058 15744
rect 3141 15738 3207 15741
rect 5349 15740 5415 15741
rect 5349 15738 5396 15740
rect 3141 15736 5396 15738
rect 3141 15680 3146 15736
rect 3202 15680 5354 15736
rect 3141 15678 5396 15680
rect 3141 15675 3207 15678
rect 5349 15676 5396 15678
rect 5460 15676 5466 15740
rect 12709 15738 12775 15741
rect 15101 15738 15167 15741
rect 12709 15736 15167 15738
rect 12709 15680 12714 15736
rect 12770 15680 15106 15736
rect 15162 15680 15167 15736
rect 12709 15678 15167 15680
rect 5349 15675 5415 15676
rect 12709 15675 12775 15678
rect 15101 15675 15167 15678
rect 2497 15602 2563 15605
rect 5717 15602 5783 15605
rect 2497 15600 5783 15602
rect 2497 15544 2502 15600
rect 2558 15544 5722 15600
rect 5778 15544 5783 15600
rect 2497 15542 5783 15544
rect 2497 15539 2563 15542
rect 5717 15539 5783 15542
rect 17677 15602 17743 15605
rect 19926 15602 19932 15604
rect 17677 15600 19932 15602
rect 17677 15544 17682 15600
rect 17738 15544 19932 15600
rect 17677 15542 19932 15544
rect 17677 15539 17743 15542
rect 19926 15540 19932 15542
rect 19996 15540 20002 15604
rect 2405 15466 2471 15469
rect 9121 15466 9187 15469
rect 2405 15464 9187 15466
rect 2405 15408 2410 15464
rect 2466 15408 9126 15464
rect 9182 15408 9187 15464
rect 2405 15406 9187 15408
rect 2405 15403 2471 15406
rect 9121 15403 9187 15406
rect 15510 15404 15516 15468
rect 15580 15466 15586 15468
rect 15653 15466 15719 15469
rect 15580 15464 15719 15466
rect 15580 15408 15658 15464
rect 15714 15408 15719 15464
rect 15580 15406 15719 15408
rect 15580 15404 15586 15406
rect 15653 15403 15719 15406
rect 19333 15466 19399 15469
rect 23920 15466 24400 15496
rect 19333 15464 24400 15466
rect 19333 15408 19338 15464
rect 19394 15408 24400 15464
rect 19333 15406 24400 15408
rect 19333 15403 19399 15406
rect 23920 15376 24400 15406
rect 13813 15332 13879 15333
rect 13813 15328 13860 15332
rect 13924 15330 13930 15332
rect 13813 15272 13818 15328
rect 13813 15268 13860 15272
rect 13924 15270 13970 15330
rect 13924 15268 13930 15270
rect 13813 15267 13879 15268
rect 4642 15264 4962 15265
rect 0 15194 480 15224
rect 4642 15200 4650 15264
rect 4714 15200 4730 15264
rect 4794 15200 4810 15264
rect 4874 15200 4890 15264
rect 4954 15200 4962 15264
rect 4642 15199 4962 15200
rect 12040 15264 12360 15265
rect 12040 15200 12048 15264
rect 12112 15200 12128 15264
rect 12192 15200 12208 15264
rect 12272 15200 12288 15264
rect 12352 15200 12360 15264
rect 12040 15199 12360 15200
rect 19437 15264 19757 15265
rect 19437 15200 19445 15264
rect 19509 15200 19525 15264
rect 19589 15200 19605 15264
rect 19669 15200 19685 15264
rect 19749 15200 19757 15264
rect 19437 15199 19757 15200
rect 3325 15194 3391 15197
rect 0 15192 3391 15194
rect 0 15136 3330 15192
rect 3386 15136 3391 15192
rect 0 15134 3391 15136
rect 0 15104 480 15134
rect 3325 15131 3391 15134
rect 18321 15194 18387 15197
rect 18454 15194 18460 15196
rect 18321 15192 18460 15194
rect 18321 15136 18326 15192
rect 18382 15136 18460 15192
rect 18321 15134 18460 15136
rect 18321 15131 18387 15134
rect 18454 15132 18460 15134
rect 18524 15132 18530 15196
rect 9029 15058 9095 15061
rect 12065 15058 12131 15061
rect 9029 15056 12131 15058
rect 9029 15000 9034 15056
rect 9090 15000 12070 15056
rect 12126 15000 12131 15056
rect 9029 14998 12131 15000
rect 9029 14995 9095 14998
rect 12065 14995 12131 14998
rect 19333 15058 19399 15061
rect 19977 15058 20043 15061
rect 19333 15056 20043 15058
rect 19333 15000 19338 15056
rect 19394 15000 19982 15056
rect 20038 15000 20043 15056
rect 19333 14998 20043 15000
rect 19333 14995 19399 14998
rect 19977 14995 20043 14998
rect 7046 14860 7052 14924
rect 7116 14922 7122 14924
rect 8201 14922 8267 14925
rect 7116 14920 8267 14922
rect 7116 14864 8206 14920
rect 8262 14864 8267 14920
rect 7116 14862 8267 14864
rect 7116 14860 7122 14862
rect 8201 14859 8267 14862
rect 15837 14922 15903 14925
rect 19609 14922 19675 14925
rect 15837 14920 19675 14922
rect 15837 14864 15842 14920
rect 15898 14864 19614 14920
rect 19670 14864 19675 14920
rect 15837 14862 19675 14864
rect 15837 14859 15903 14862
rect 19609 14859 19675 14862
rect 9990 14724 9996 14788
rect 10060 14786 10066 14788
rect 13261 14786 13327 14789
rect 10060 14784 13327 14786
rect 10060 14728 13266 14784
rect 13322 14728 13327 14784
rect 10060 14726 13327 14728
rect 10060 14724 10066 14726
rect 13261 14723 13327 14726
rect 19977 14786 20043 14789
rect 23920 14786 24400 14816
rect 19977 14784 24400 14786
rect 19977 14728 19982 14784
rect 20038 14728 24400 14784
rect 19977 14726 24400 14728
rect 19977 14723 20043 14726
rect 8341 14720 8661 14721
rect 8341 14656 8349 14720
rect 8413 14656 8429 14720
rect 8493 14656 8509 14720
rect 8573 14656 8589 14720
rect 8653 14656 8661 14720
rect 8341 14655 8661 14656
rect 15738 14720 16058 14721
rect 15738 14656 15746 14720
rect 15810 14656 15826 14720
rect 15890 14656 15906 14720
rect 15970 14656 15986 14720
rect 16050 14656 16058 14720
rect 23920 14696 24400 14726
rect 15738 14655 16058 14656
rect 16205 14652 16271 14653
rect 16205 14648 16252 14652
rect 16316 14650 16322 14652
rect 17769 14650 17835 14653
rect 20805 14650 20871 14653
rect 16205 14592 16210 14648
rect 16205 14588 16252 14592
rect 16316 14590 16362 14650
rect 17769 14648 20871 14650
rect 17769 14592 17774 14648
rect 17830 14592 20810 14648
rect 20866 14592 20871 14648
rect 17769 14590 20871 14592
rect 16316 14588 16322 14590
rect 16205 14587 16271 14588
rect 17769 14587 17835 14590
rect 20805 14587 20871 14590
rect 4429 14514 4495 14517
rect 6453 14514 6519 14517
rect 4429 14512 6519 14514
rect 4429 14456 4434 14512
rect 4490 14456 6458 14512
rect 6514 14456 6519 14512
rect 4429 14454 6519 14456
rect 4429 14451 4495 14454
rect 6453 14451 6519 14454
rect 10225 14514 10291 14517
rect 17125 14514 17191 14517
rect 10225 14512 17191 14514
rect 10225 14456 10230 14512
rect 10286 14456 17130 14512
rect 17186 14456 17191 14512
rect 10225 14454 17191 14456
rect 10225 14451 10291 14454
rect 17125 14451 17191 14454
rect 18505 14514 18571 14517
rect 18638 14514 18644 14516
rect 18505 14512 18644 14514
rect 18505 14456 18510 14512
rect 18566 14456 18644 14512
rect 18505 14454 18644 14456
rect 18505 14451 18571 14454
rect 18638 14452 18644 14454
rect 18708 14452 18714 14516
rect 19149 14514 19215 14517
rect 20989 14514 21055 14517
rect 19149 14512 21055 14514
rect 19149 14456 19154 14512
rect 19210 14456 20994 14512
rect 21050 14456 21055 14512
rect 19149 14454 21055 14456
rect 19149 14451 19215 14454
rect 20989 14451 21055 14454
rect 2865 14378 2931 14381
rect 4705 14378 4771 14381
rect 2865 14376 4771 14378
rect 2865 14320 2870 14376
rect 2926 14320 4710 14376
rect 4766 14320 4771 14376
rect 2865 14318 4771 14320
rect 2865 14315 2931 14318
rect 4705 14315 4771 14318
rect 7557 14378 7623 14381
rect 12617 14378 12683 14381
rect 7557 14376 12683 14378
rect 7557 14320 7562 14376
rect 7618 14320 12622 14376
rect 12678 14320 12683 14376
rect 7557 14318 12683 14320
rect 7557 14315 7623 14318
rect 12617 14315 12683 14318
rect 15142 14180 15148 14244
rect 15212 14242 15218 14244
rect 15745 14242 15811 14245
rect 15212 14240 15811 14242
rect 15212 14184 15750 14240
rect 15806 14184 15811 14240
rect 15212 14182 15811 14184
rect 15212 14180 15218 14182
rect 15745 14179 15811 14182
rect 4642 14176 4962 14177
rect 4642 14112 4650 14176
rect 4714 14112 4730 14176
rect 4794 14112 4810 14176
rect 4874 14112 4890 14176
rect 4954 14112 4962 14176
rect 4642 14111 4962 14112
rect 12040 14176 12360 14177
rect 12040 14112 12048 14176
rect 12112 14112 12128 14176
rect 12192 14112 12208 14176
rect 12272 14112 12288 14176
rect 12352 14112 12360 14176
rect 12040 14111 12360 14112
rect 19437 14176 19757 14177
rect 19437 14112 19445 14176
rect 19509 14112 19525 14176
rect 19589 14112 19605 14176
rect 19669 14112 19685 14176
rect 19749 14112 19757 14176
rect 19437 14111 19757 14112
rect 12566 14044 12572 14108
rect 12636 14106 12642 14108
rect 14917 14106 14983 14109
rect 12636 14104 14983 14106
rect 12636 14048 14922 14104
rect 14978 14048 14983 14104
rect 12636 14046 14983 14048
rect 12636 14044 12642 14046
rect 14917 14043 14983 14046
rect 20437 14106 20503 14109
rect 23920 14106 24400 14136
rect 20437 14104 24400 14106
rect 20437 14048 20442 14104
rect 20498 14048 24400 14104
rect 20437 14046 24400 14048
rect 20437 14043 20503 14046
rect 23920 14016 24400 14046
rect 9622 13908 9628 13972
rect 9692 13970 9698 13972
rect 14641 13970 14707 13973
rect 9692 13968 14707 13970
rect 9692 13912 14646 13968
rect 14702 13912 14707 13968
rect 9692 13910 14707 13912
rect 9692 13908 9698 13910
rect 14641 13907 14707 13910
rect 1853 13834 1919 13837
rect 7189 13834 7255 13837
rect 1853 13832 7255 13834
rect 1853 13776 1858 13832
rect 1914 13776 7194 13832
rect 7250 13776 7255 13832
rect 1853 13774 7255 13776
rect 1853 13771 1919 13774
rect 7189 13771 7255 13774
rect 10777 13834 10843 13837
rect 12157 13834 12223 13837
rect 10777 13832 12223 13834
rect 10777 13776 10782 13832
rect 10838 13776 12162 13832
rect 12218 13776 12223 13832
rect 10777 13774 12223 13776
rect 10777 13771 10843 13774
rect 12157 13771 12223 13774
rect 8341 13632 8661 13633
rect 8341 13568 8349 13632
rect 8413 13568 8429 13632
rect 8493 13568 8509 13632
rect 8573 13568 8589 13632
rect 8653 13568 8661 13632
rect 8341 13567 8661 13568
rect 15738 13632 16058 13633
rect 15738 13568 15746 13632
rect 15810 13568 15826 13632
rect 15890 13568 15906 13632
rect 15970 13568 15986 13632
rect 16050 13568 16058 13632
rect 15738 13567 16058 13568
rect 1669 13426 1735 13429
rect 5533 13426 5599 13429
rect 1669 13424 5599 13426
rect 1669 13368 1674 13424
rect 1730 13368 5538 13424
rect 5594 13368 5599 13424
rect 1669 13366 5599 13368
rect 1669 13363 1735 13366
rect 5533 13363 5599 13366
rect 10358 13364 10364 13428
rect 10428 13426 10434 13428
rect 16113 13426 16179 13429
rect 10428 13424 16179 13426
rect 10428 13368 16118 13424
rect 16174 13368 16179 13424
rect 10428 13366 16179 13368
rect 10428 13364 10434 13366
rect 16113 13363 16179 13366
rect 19333 13426 19399 13429
rect 23920 13426 24400 13456
rect 19333 13424 24400 13426
rect 19333 13368 19338 13424
rect 19394 13368 24400 13424
rect 19333 13366 24400 13368
rect 19333 13363 19399 13366
rect 23920 13336 24400 13366
rect 10317 13290 10383 13293
rect 18229 13290 18295 13293
rect 10317 13288 18295 13290
rect 10317 13232 10322 13288
rect 10378 13232 18234 13288
rect 18290 13232 18295 13288
rect 10317 13230 18295 13232
rect 10317 13227 10383 13230
rect 18229 13227 18295 13230
rect 6494 13092 6500 13156
rect 6564 13154 6570 13156
rect 7465 13154 7531 13157
rect 8109 13154 8175 13157
rect 6564 13152 8175 13154
rect 6564 13096 7470 13152
rect 7526 13096 8114 13152
rect 8170 13096 8175 13152
rect 6564 13094 8175 13096
rect 6564 13092 6570 13094
rect 7465 13091 7531 13094
rect 8109 13091 8175 13094
rect 15837 13154 15903 13157
rect 18689 13154 18755 13157
rect 15837 13152 18755 13154
rect 15837 13096 15842 13152
rect 15898 13096 18694 13152
rect 18750 13096 18755 13152
rect 15837 13094 18755 13096
rect 15837 13091 15903 13094
rect 18689 13091 18755 13094
rect 4642 13088 4962 13089
rect 4642 13024 4650 13088
rect 4714 13024 4730 13088
rect 4794 13024 4810 13088
rect 4874 13024 4890 13088
rect 4954 13024 4962 13088
rect 4642 13023 4962 13024
rect 12040 13088 12360 13089
rect 12040 13024 12048 13088
rect 12112 13024 12128 13088
rect 12192 13024 12208 13088
rect 12272 13024 12288 13088
rect 12352 13024 12360 13088
rect 12040 13023 12360 13024
rect 19437 13088 19757 13089
rect 19437 13024 19445 13088
rect 19509 13024 19525 13088
rect 19589 13024 19605 13088
rect 19669 13024 19685 13088
rect 19749 13024 19757 13088
rect 19437 13023 19757 13024
rect 5533 13018 5599 13021
rect 5717 13018 5783 13021
rect 16849 13018 16915 13021
rect 5533 13016 5783 13018
rect 5533 12960 5538 13016
rect 5594 12960 5722 13016
rect 5778 12960 5783 13016
rect 5533 12958 5783 12960
rect 5533 12955 5599 12958
rect 5717 12955 5783 12958
rect 12436 13016 16915 13018
rect 12436 12960 16854 13016
rect 16910 12960 16915 13016
rect 12436 12958 16915 12960
rect 4521 12882 4587 12885
rect 9121 12882 9187 12885
rect 4521 12880 9187 12882
rect 4521 12824 4526 12880
rect 4582 12824 9126 12880
rect 9182 12824 9187 12880
rect 4521 12822 9187 12824
rect 4521 12819 4587 12822
rect 9121 12819 9187 12822
rect 11145 12882 11211 12885
rect 12436 12882 12496 12958
rect 16849 12955 16915 12958
rect 12709 12882 12775 12885
rect 11145 12880 12496 12882
rect 11145 12824 11150 12880
rect 11206 12824 12496 12880
rect 11145 12822 12496 12824
rect 12574 12880 12775 12882
rect 12574 12824 12714 12880
rect 12770 12824 12775 12880
rect 12574 12822 12775 12824
rect 11145 12819 11211 12822
rect 4521 12748 4587 12749
rect 4470 12684 4476 12748
rect 4540 12746 4587 12748
rect 4540 12744 4632 12746
rect 4582 12688 4632 12744
rect 4540 12686 4632 12688
rect 4540 12684 4587 12686
rect 5758 12684 5764 12748
rect 5828 12746 5834 12748
rect 5901 12746 5967 12749
rect 5828 12744 5967 12746
rect 5828 12688 5906 12744
rect 5962 12688 5967 12744
rect 5828 12686 5967 12688
rect 5828 12684 5834 12686
rect 4521 12683 4587 12684
rect 5901 12683 5967 12686
rect 7281 12746 7347 12749
rect 9673 12746 9739 12749
rect 7281 12744 9739 12746
rect 7281 12688 7286 12744
rect 7342 12688 9678 12744
rect 9734 12688 9739 12744
rect 7281 12686 9739 12688
rect 7281 12683 7347 12686
rect 9673 12683 9739 12686
rect 11513 12610 11579 12613
rect 11646 12610 11652 12612
rect 11513 12608 11652 12610
rect 11513 12552 11518 12608
rect 11574 12552 11652 12608
rect 11513 12550 11652 12552
rect 11513 12547 11579 12550
rect 11646 12548 11652 12550
rect 11716 12548 11722 12612
rect 8341 12544 8661 12545
rect 8341 12480 8349 12544
rect 8413 12480 8429 12544
rect 8493 12480 8509 12544
rect 8573 12480 8589 12544
rect 8653 12480 8661 12544
rect 8341 12479 8661 12480
rect 6085 12474 6151 12477
rect 6310 12474 6316 12476
rect 6085 12472 6316 12474
rect 6085 12416 6090 12472
rect 6146 12416 6316 12472
rect 6085 12414 6316 12416
rect 6085 12411 6151 12414
rect 6310 12412 6316 12414
rect 6380 12412 6386 12476
rect 5533 12338 5599 12341
rect 8845 12338 8911 12341
rect 12574 12338 12634 12822
rect 12709 12819 12775 12822
rect 14365 12882 14431 12885
rect 19885 12882 19951 12885
rect 14365 12880 17924 12882
rect 14365 12824 14370 12880
rect 14426 12824 17924 12880
rect 14365 12822 17924 12824
rect 14365 12819 14431 12822
rect 17864 12749 17924 12822
rect 19885 12880 19994 12882
rect 19885 12824 19890 12880
rect 19946 12824 19994 12880
rect 19885 12819 19994 12824
rect 12709 12746 12775 12749
rect 13997 12746 14063 12749
rect 12709 12744 14063 12746
rect 12709 12688 12714 12744
rect 12770 12688 14002 12744
rect 14058 12688 14063 12744
rect 12709 12686 14063 12688
rect 12709 12683 12775 12686
rect 13997 12683 14063 12686
rect 17861 12744 17927 12749
rect 17861 12688 17866 12744
rect 17922 12688 17927 12744
rect 17861 12683 17927 12688
rect 12750 12548 12756 12612
rect 12820 12610 12826 12612
rect 12893 12610 12959 12613
rect 12820 12608 12959 12610
rect 12820 12552 12898 12608
rect 12954 12552 12959 12608
rect 12820 12550 12959 12552
rect 12820 12548 12826 12550
rect 12893 12547 12959 12550
rect 15738 12544 16058 12545
rect 15738 12480 15746 12544
rect 15810 12480 15826 12544
rect 15890 12480 15906 12544
rect 15970 12480 15986 12544
rect 16050 12480 16058 12544
rect 15738 12479 16058 12480
rect 12934 12412 12940 12476
rect 13004 12474 13010 12476
rect 14365 12474 14431 12477
rect 13004 12472 14431 12474
rect 13004 12416 14370 12472
rect 14426 12416 14431 12472
rect 13004 12414 14431 12416
rect 19934 12474 19994 12819
rect 22369 12746 22435 12749
rect 23920 12746 24400 12776
rect 22369 12744 24400 12746
rect 22369 12688 22374 12744
rect 22430 12688 24400 12744
rect 22369 12686 24400 12688
rect 22369 12683 22435 12686
rect 23920 12656 24400 12686
rect 20069 12612 20135 12613
rect 20069 12608 20116 12612
rect 20180 12610 20186 12612
rect 20069 12552 20074 12608
rect 20069 12548 20116 12552
rect 20180 12550 20226 12610
rect 20180 12548 20186 12550
rect 20069 12547 20135 12548
rect 20069 12474 20135 12477
rect 20529 12476 20595 12477
rect 20478 12474 20484 12476
rect 19934 12472 20135 12474
rect 19934 12416 20074 12472
rect 20130 12416 20135 12472
rect 19934 12414 20135 12416
rect 20438 12414 20484 12474
rect 20548 12472 20595 12476
rect 20590 12416 20595 12472
rect 13004 12412 13010 12414
rect 14365 12411 14431 12414
rect 20069 12411 20135 12414
rect 20478 12412 20484 12414
rect 20548 12412 20595 12416
rect 20529 12411 20595 12412
rect 5533 12336 8911 12338
rect 5533 12280 5538 12336
rect 5594 12280 8850 12336
rect 8906 12280 8911 12336
rect 5533 12278 8911 12280
rect 5533 12275 5599 12278
rect 8845 12275 8911 12278
rect 9998 12278 12634 12338
rect 13077 12338 13143 12341
rect 13302 12338 13308 12340
rect 13077 12336 13308 12338
rect 13077 12280 13082 12336
rect 13138 12280 13308 12336
rect 13077 12278 13308 12280
rect 5758 12140 5764 12204
rect 5828 12202 5834 12204
rect 6085 12202 6151 12205
rect 5828 12200 6151 12202
rect 5828 12144 6090 12200
rect 6146 12144 6151 12200
rect 5828 12142 6151 12144
rect 5828 12140 5834 12142
rect 6085 12139 6151 12142
rect 6637 12202 6703 12205
rect 7741 12202 7807 12205
rect 6637 12200 7807 12202
rect 6637 12144 6642 12200
rect 6698 12144 7746 12200
rect 7802 12144 7807 12200
rect 6637 12142 7807 12144
rect 6637 12139 6703 12142
rect 7741 12139 7807 12142
rect 5717 12066 5783 12069
rect 6310 12066 6316 12068
rect 5717 12064 6316 12066
rect 5717 12008 5722 12064
rect 5778 12008 6316 12064
rect 5717 12006 6316 12008
rect 5717 12003 5783 12006
rect 6310 12004 6316 12006
rect 6380 12004 6386 12068
rect 9029 12066 9095 12069
rect 9673 12066 9739 12069
rect 9029 12064 9739 12066
rect 9029 12008 9034 12064
rect 9090 12008 9678 12064
rect 9734 12008 9739 12064
rect 9029 12006 9739 12008
rect 9029 12003 9095 12006
rect 9673 12003 9739 12006
rect 4642 12000 4962 12001
rect 4642 11936 4650 12000
rect 4714 11936 4730 12000
rect 4794 11936 4810 12000
rect 4874 11936 4890 12000
rect 4954 11936 4962 12000
rect 4642 11935 4962 11936
rect 7833 11930 7899 11933
rect 5030 11928 7899 11930
rect 5030 11872 7838 11928
rect 7894 11872 7899 11928
rect 5030 11870 7899 11872
rect 3969 11794 4035 11797
rect 5030 11794 5090 11870
rect 7833 11867 7899 11870
rect 9998 11797 10058 12278
rect 13077 12275 13143 12278
rect 13302 12276 13308 12278
rect 13372 12338 13378 12340
rect 14089 12338 14155 12341
rect 13372 12336 14155 12338
rect 13372 12280 14094 12336
rect 14150 12280 14155 12336
rect 13372 12278 14155 12280
rect 13372 12276 13378 12278
rect 14089 12275 14155 12278
rect 15377 12336 15443 12341
rect 15377 12280 15382 12336
rect 15438 12280 15443 12336
rect 15377 12275 15443 12280
rect 10869 12202 10935 12205
rect 12709 12204 12775 12205
rect 12709 12202 12756 12204
rect 10869 12200 12588 12202
rect 10869 12144 10874 12200
rect 10930 12144 12588 12200
rect 10869 12142 12588 12144
rect 12664 12200 12756 12202
rect 12664 12144 12714 12200
rect 12664 12142 12756 12144
rect 10869 12139 10935 12142
rect 12528 12066 12588 12142
rect 12709 12140 12756 12142
rect 12820 12140 12826 12204
rect 12709 12139 12775 12140
rect 15380 12066 15440 12275
rect 21725 12202 21791 12205
rect 23920 12202 24400 12232
rect 21725 12200 24400 12202
rect 21725 12144 21730 12200
rect 21786 12144 24400 12200
rect 21725 12142 24400 12144
rect 21725 12139 21791 12142
rect 23920 12112 24400 12142
rect 12528 12006 15440 12066
rect 18822 12004 18828 12068
rect 18892 12066 18898 12068
rect 19057 12066 19123 12069
rect 18892 12064 19123 12066
rect 18892 12008 19062 12064
rect 19118 12008 19123 12064
rect 18892 12006 19123 12008
rect 18892 12004 18898 12006
rect 19057 12003 19123 12006
rect 12040 12000 12360 12001
rect 12040 11936 12048 12000
rect 12112 11936 12128 12000
rect 12192 11936 12208 12000
rect 12272 11936 12288 12000
rect 12352 11936 12360 12000
rect 12040 11935 12360 11936
rect 19437 12000 19757 12001
rect 19437 11936 19445 12000
rect 19509 11936 19525 12000
rect 19589 11936 19605 12000
rect 19669 11936 19685 12000
rect 19749 11936 19757 12000
rect 19437 11935 19757 11936
rect 12525 11930 12591 11933
rect 13261 11930 13327 11933
rect 12525 11928 13327 11930
rect 12525 11872 12530 11928
rect 12586 11872 13266 11928
rect 13322 11872 13327 11928
rect 12525 11870 13327 11872
rect 12525 11867 12591 11870
rect 13261 11867 13327 11870
rect 14089 11930 14155 11933
rect 15745 11930 15811 11933
rect 18781 11930 18847 11933
rect 14089 11928 18847 11930
rect 14089 11872 14094 11928
rect 14150 11872 15750 11928
rect 15806 11872 18786 11928
rect 18842 11872 18847 11928
rect 14089 11870 18847 11872
rect 14089 11867 14155 11870
rect 15745 11867 15811 11870
rect 18781 11867 18847 11870
rect 18965 11932 19031 11933
rect 18965 11928 19012 11932
rect 19076 11930 19082 11932
rect 18965 11872 18970 11928
rect 18965 11868 19012 11872
rect 19076 11870 19122 11930
rect 19076 11868 19082 11870
rect 18965 11867 19031 11868
rect 3969 11792 5090 11794
rect 3969 11736 3974 11792
rect 4030 11736 5090 11792
rect 3969 11734 5090 11736
rect 5533 11794 5599 11797
rect 8937 11794 9003 11797
rect 5533 11792 9003 11794
rect 5533 11736 5538 11792
rect 5594 11736 8942 11792
rect 8998 11736 9003 11792
rect 5533 11734 9003 11736
rect 3969 11731 4035 11734
rect 5533 11731 5599 11734
rect 8937 11731 9003 11734
rect 9949 11792 10058 11797
rect 9949 11736 9954 11792
rect 10010 11736 10058 11792
rect 9949 11734 10058 11736
rect 10593 11794 10659 11797
rect 19701 11794 19767 11797
rect 20345 11794 20411 11797
rect 10593 11792 20411 11794
rect 10593 11736 10598 11792
rect 10654 11736 19706 11792
rect 19762 11736 20350 11792
rect 20406 11736 20411 11792
rect 10593 11734 20411 11736
rect 9949 11731 10015 11734
rect 10593 11731 10659 11734
rect 19701 11731 19767 11734
rect 20345 11731 20411 11734
rect 9857 11658 9923 11661
rect 10501 11658 10567 11661
rect 9857 11656 10567 11658
rect 9857 11600 9862 11656
rect 9918 11600 10506 11656
rect 10562 11600 10567 11656
rect 9857 11598 10567 11600
rect 9857 11595 9923 11598
rect 10501 11595 10567 11598
rect 13169 11658 13235 11661
rect 18321 11658 18387 11661
rect 13169 11656 18387 11658
rect 13169 11600 13174 11656
rect 13230 11600 18326 11656
rect 18382 11600 18387 11656
rect 13169 11598 18387 11600
rect 13169 11595 13235 11598
rect 18321 11595 18387 11598
rect 10685 11522 10751 11525
rect 12893 11522 12959 11525
rect 10685 11520 12959 11522
rect 10685 11464 10690 11520
rect 10746 11464 12898 11520
rect 12954 11464 12959 11520
rect 10685 11462 12959 11464
rect 10685 11459 10751 11462
rect 12893 11459 12959 11462
rect 19149 11522 19215 11525
rect 23920 11522 24400 11552
rect 19149 11520 24400 11522
rect 19149 11464 19154 11520
rect 19210 11464 24400 11520
rect 19149 11462 24400 11464
rect 19149 11459 19215 11462
rect 8341 11456 8661 11457
rect 8341 11392 8349 11456
rect 8413 11392 8429 11456
rect 8493 11392 8509 11456
rect 8573 11392 8589 11456
rect 8653 11392 8661 11456
rect 8341 11391 8661 11392
rect 15738 11456 16058 11457
rect 15738 11392 15746 11456
rect 15810 11392 15826 11456
rect 15890 11392 15906 11456
rect 15970 11392 15986 11456
rect 16050 11392 16058 11456
rect 23920 11432 24400 11462
rect 15738 11391 16058 11392
rect 15326 11386 15332 11388
rect 9630 11326 15332 11386
rect 8150 11188 8156 11252
rect 8220 11250 8226 11252
rect 9630 11250 9690 11326
rect 15326 11324 15332 11326
rect 15396 11324 15402 11388
rect 20069 11386 20135 11389
rect 20294 11386 20300 11388
rect 20069 11384 20300 11386
rect 20069 11328 20074 11384
rect 20130 11328 20300 11384
rect 20069 11326 20300 11328
rect 20069 11323 20135 11326
rect 20294 11324 20300 11326
rect 20364 11324 20370 11388
rect 8220 11190 9690 11250
rect 12893 11250 12959 11253
rect 13629 11250 13695 11253
rect 16573 11250 16639 11253
rect 17861 11250 17927 11253
rect 12893 11248 13695 11250
rect 12893 11192 12898 11248
rect 12954 11192 13634 11248
rect 13690 11192 13695 11248
rect 12893 11190 13695 11192
rect 8220 11188 8226 11190
rect 12893 11187 12959 11190
rect 13629 11187 13695 11190
rect 14598 11248 17927 11250
rect 14598 11192 16578 11248
rect 16634 11192 17866 11248
rect 17922 11192 17927 11248
rect 14598 11190 17927 11192
rect 4705 11114 4771 11117
rect 5022 11114 5028 11116
rect 4705 11112 5028 11114
rect 4705 11056 4710 11112
rect 4766 11056 5028 11112
rect 4705 11054 5028 11056
rect 4705 11051 4771 11054
rect 5022 11052 5028 11054
rect 5092 11052 5098 11116
rect 11513 11114 11579 11117
rect 14457 11114 14523 11117
rect 11513 11112 14523 11114
rect 11513 11056 11518 11112
rect 11574 11056 14462 11112
rect 14518 11056 14523 11112
rect 11513 11054 14523 11056
rect 11513 11051 11579 11054
rect 14457 11051 14523 11054
rect 8937 10978 9003 10981
rect 11697 10978 11763 10981
rect 8937 10976 11763 10978
rect 8937 10920 8942 10976
rect 8998 10920 11702 10976
rect 11758 10920 11763 10976
rect 8937 10918 11763 10920
rect 8937 10915 9003 10918
rect 11697 10915 11763 10918
rect 12985 10978 13051 10981
rect 14598 10978 14658 11190
rect 16573 11187 16639 11190
rect 17861 11187 17927 11190
rect 15142 11052 15148 11116
rect 15212 11114 15218 11116
rect 17217 11114 17283 11117
rect 15212 11112 17283 11114
rect 15212 11056 17222 11112
rect 17278 11056 17283 11112
rect 15212 11054 17283 11056
rect 15212 11052 15218 11054
rect 17217 11051 17283 11054
rect 19057 11114 19123 11117
rect 23381 11114 23447 11117
rect 19057 11112 23447 11114
rect 19057 11056 19062 11112
rect 19118 11056 23386 11112
rect 23442 11056 23447 11112
rect 19057 11054 23447 11056
rect 19057 11051 19123 11054
rect 23381 11051 23447 11054
rect 12985 10976 14658 10978
rect 12985 10920 12990 10976
rect 13046 10920 14658 10976
rect 12985 10918 14658 10920
rect 14917 10978 14983 10981
rect 15653 10978 15719 10981
rect 17677 10978 17743 10981
rect 14917 10976 17743 10978
rect 14917 10920 14922 10976
rect 14978 10920 15658 10976
rect 15714 10920 17682 10976
rect 17738 10920 17743 10976
rect 14917 10918 17743 10920
rect 12985 10915 13051 10918
rect 14917 10915 14983 10918
rect 15653 10915 15719 10918
rect 17677 10915 17743 10918
rect 4642 10912 4962 10913
rect 4642 10848 4650 10912
rect 4714 10848 4730 10912
rect 4794 10848 4810 10912
rect 4874 10848 4890 10912
rect 4954 10848 4962 10912
rect 4642 10847 4962 10848
rect 12040 10912 12360 10913
rect 12040 10848 12048 10912
rect 12112 10848 12128 10912
rect 12192 10848 12208 10912
rect 12272 10848 12288 10912
rect 12352 10848 12360 10912
rect 12040 10847 12360 10848
rect 19437 10912 19757 10913
rect 19437 10848 19445 10912
rect 19509 10848 19525 10912
rect 19589 10848 19605 10912
rect 19669 10848 19685 10912
rect 19749 10848 19757 10912
rect 19437 10847 19757 10848
rect 5758 10780 5764 10844
rect 5828 10842 5834 10844
rect 11789 10842 11855 10845
rect 5828 10840 11855 10842
rect 5828 10784 11794 10840
rect 11850 10784 11855 10840
rect 5828 10782 11855 10784
rect 5828 10780 5834 10782
rect 11789 10779 11855 10782
rect 12985 10842 13051 10845
rect 13721 10842 13787 10845
rect 12985 10840 13787 10842
rect 12985 10784 12990 10840
rect 13046 10784 13726 10840
rect 13782 10784 13787 10840
rect 12985 10782 13787 10784
rect 12985 10779 13051 10782
rect 13721 10779 13787 10782
rect 15510 10780 15516 10844
rect 15580 10842 15586 10844
rect 15653 10842 15719 10845
rect 15580 10840 15719 10842
rect 15580 10784 15658 10840
rect 15714 10784 15719 10840
rect 15580 10782 15719 10784
rect 15580 10780 15586 10782
rect 15653 10779 15719 10782
rect 20805 10842 20871 10845
rect 23920 10842 24400 10872
rect 20805 10840 24400 10842
rect 20805 10784 20810 10840
rect 20866 10784 24400 10840
rect 20805 10782 24400 10784
rect 20805 10779 20871 10782
rect 23920 10752 24400 10782
rect 7230 10644 7236 10708
rect 7300 10706 7306 10708
rect 11830 10706 11836 10708
rect 7300 10646 11836 10706
rect 7300 10644 7306 10646
rect 11830 10644 11836 10646
rect 11900 10644 11906 10708
rect 17217 10706 17283 10709
rect 12712 10704 17283 10706
rect 12712 10648 17222 10704
rect 17278 10648 17283 10704
rect 12712 10646 17283 10648
rect 3141 10570 3207 10573
rect 8477 10570 8543 10573
rect 3141 10568 8543 10570
rect 3141 10512 3146 10568
rect 3202 10512 8482 10568
rect 8538 10512 8543 10568
rect 3141 10510 8543 10512
rect 3141 10507 3207 10510
rect 8477 10507 8543 10510
rect 9438 10508 9444 10572
rect 9508 10570 9514 10572
rect 12525 10570 12591 10573
rect 9508 10568 12591 10570
rect 9508 10512 12530 10568
rect 12586 10512 12591 10568
rect 9508 10510 12591 10512
rect 9508 10508 9514 10510
rect 12525 10507 12591 10510
rect 9806 10372 9812 10436
rect 9876 10434 9882 10436
rect 12712 10434 12772 10646
rect 17217 10643 17283 10646
rect 19926 10644 19932 10708
rect 19996 10706 20002 10708
rect 20621 10706 20687 10709
rect 19996 10704 20687 10706
rect 19996 10648 20626 10704
rect 20682 10648 20687 10704
rect 19996 10646 20687 10648
rect 19996 10644 20002 10646
rect 20621 10643 20687 10646
rect 12934 10508 12940 10572
rect 13004 10570 13010 10572
rect 21449 10570 21515 10573
rect 13004 10568 21515 10570
rect 13004 10512 21454 10568
rect 21510 10512 21515 10568
rect 13004 10510 21515 10512
rect 13004 10508 13010 10510
rect 21449 10507 21515 10510
rect 9876 10374 12772 10434
rect 13813 10432 13879 10437
rect 13813 10376 13818 10432
rect 13874 10376 13879 10432
rect 9876 10372 9882 10374
rect 13813 10371 13879 10376
rect 8341 10368 8661 10369
rect 8341 10304 8349 10368
rect 8413 10304 8429 10368
rect 8493 10304 8509 10368
rect 8573 10304 8589 10368
rect 8653 10304 8661 10368
rect 8341 10303 8661 10304
rect 4797 10298 4863 10301
rect 5758 10298 5764 10300
rect 4797 10296 5764 10298
rect 4797 10240 4802 10296
rect 4858 10240 5764 10296
rect 4797 10238 5764 10240
rect 4797 10235 4863 10238
rect 5758 10236 5764 10238
rect 5828 10236 5834 10300
rect 11973 10298 12039 10301
rect 13670 10298 13676 10300
rect 11973 10296 13676 10298
rect 11973 10240 11978 10296
rect 12034 10240 13676 10296
rect 11973 10238 13676 10240
rect 11973 10235 12039 10238
rect 13670 10236 13676 10238
rect 13740 10236 13746 10300
rect 13816 10165 13876 10371
rect 15738 10368 16058 10369
rect 15738 10304 15746 10368
rect 15810 10304 15826 10368
rect 15890 10304 15906 10368
rect 15970 10304 15986 10368
rect 16050 10304 16058 10368
rect 15738 10303 16058 10304
rect 7414 10100 7420 10164
rect 7484 10162 7490 10164
rect 8886 10162 8892 10164
rect 7484 10102 8892 10162
rect 7484 10100 7490 10102
rect 8886 10100 8892 10102
rect 8956 10100 8962 10164
rect 12985 10162 13051 10165
rect 12390 10160 13051 10162
rect 12390 10104 12990 10160
rect 13046 10104 13051 10160
rect 12390 10102 13051 10104
rect 6862 9964 6868 10028
rect 6932 10026 6938 10028
rect 12390 10026 12450 10102
rect 12985 10099 13051 10102
rect 13813 10160 13879 10165
rect 13813 10104 13818 10160
rect 13874 10104 13879 10160
rect 13813 10099 13879 10104
rect 16113 10162 16179 10165
rect 16246 10162 16252 10164
rect 16113 10160 16252 10162
rect 16113 10104 16118 10160
rect 16174 10104 16252 10160
rect 16113 10102 16252 10104
rect 16113 10099 16179 10102
rect 16246 10100 16252 10102
rect 16316 10100 16322 10164
rect 20253 10162 20319 10165
rect 23920 10162 24400 10192
rect 20253 10160 24400 10162
rect 20253 10104 20258 10160
rect 20314 10104 24400 10160
rect 20253 10102 24400 10104
rect 20253 10099 20319 10102
rect 23920 10072 24400 10102
rect 6932 9966 12450 10026
rect 12525 10026 12591 10029
rect 15193 10026 15259 10029
rect 12525 10024 15259 10026
rect 12525 9968 12530 10024
rect 12586 9968 15198 10024
rect 15254 9968 15259 10024
rect 12525 9966 15259 9968
rect 6932 9964 6938 9966
rect 12525 9963 12591 9966
rect 15193 9963 15259 9966
rect 16297 10026 16363 10029
rect 18321 10026 18387 10029
rect 19701 10026 19767 10029
rect 16297 10024 19767 10026
rect 16297 9968 16302 10024
rect 16358 9968 18326 10024
rect 18382 9968 19706 10024
rect 19762 9968 19767 10024
rect 16297 9966 19767 9968
rect 16297 9963 16363 9966
rect 18321 9963 18387 9966
rect 19701 9963 19767 9966
rect 7598 9828 7604 9892
rect 7668 9890 7674 9892
rect 8753 9890 8819 9893
rect 7668 9888 8819 9890
rect 7668 9832 8758 9888
rect 8814 9832 8819 9888
rect 7668 9830 8819 9832
rect 7668 9828 7674 9830
rect 8753 9827 8819 9830
rect 8886 9828 8892 9892
rect 8956 9890 8962 9892
rect 9213 9890 9279 9893
rect 18965 9890 19031 9893
rect 8956 9888 9279 9890
rect 8956 9832 9218 9888
rect 9274 9832 9279 9888
rect 8956 9830 9279 9832
rect 8956 9828 8962 9830
rect 9213 9827 9279 9830
rect 12436 9888 19031 9890
rect 12436 9832 18970 9888
rect 19026 9832 19031 9888
rect 12436 9830 19031 9832
rect 4642 9824 4962 9825
rect 4642 9760 4650 9824
rect 4714 9760 4730 9824
rect 4794 9760 4810 9824
rect 4874 9760 4890 9824
rect 4954 9760 4962 9824
rect 4642 9759 4962 9760
rect 12040 9824 12360 9825
rect 12040 9760 12048 9824
rect 12112 9760 12128 9824
rect 12192 9760 12208 9824
rect 12272 9760 12288 9824
rect 12352 9760 12360 9824
rect 12040 9759 12360 9760
rect 7046 9754 7052 9756
rect 6870 9694 7052 9754
rect 4797 9618 4863 9621
rect 6870 9618 6930 9694
rect 7046 9692 7052 9694
rect 7116 9692 7122 9756
rect 7782 9692 7788 9756
rect 7852 9754 7858 9756
rect 8937 9754 9003 9757
rect 7852 9752 9003 9754
rect 7852 9696 8942 9752
rect 8998 9696 9003 9752
rect 7852 9694 9003 9696
rect 7852 9692 7858 9694
rect 8937 9691 9003 9694
rect 9213 9754 9279 9757
rect 10174 9754 10180 9756
rect 9213 9752 10180 9754
rect 9213 9696 9218 9752
rect 9274 9696 10180 9752
rect 9213 9694 10180 9696
rect 9213 9691 9279 9694
rect 10174 9692 10180 9694
rect 10244 9754 10250 9756
rect 10685 9754 10751 9757
rect 10244 9752 10751 9754
rect 10244 9696 10690 9752
rect 10746 9696 10751 9752
rect 10244 9694 10751 9696
rect 10244 9692 10250 9694
rect 10685 9691 10751 9694
rect 4797 9616 6930 9618
rect 4797 9560 4802 9616
rect 4858 9560 6930 9616
rect 4797 9558 6930 9560
rect 7005 9618 7071 9621
rect 8293 9618 8359 9621
rect 7005 9616 8359 9618
rect 7005 9560 7010 9616
rect 7066 9560 8298 9616
rect 8354 9560 8359 9616
rect 7005 9558 8359 9560
rect 4797 9555 4863 9558
rect 7005 9555 7071 9558
rect 8293 9555 8359 9558
rect 8477 9618 8543 9621
rect 12436 9618 12496 9830
rect 18965 9827 19031 9830
rect 19437 9824 19757 9825
rect 19437 9760 19445 9824
rect 19509 9760 19525 9824
rect 19589 9760 19605 9824
rect 19669 9760 19685 9824
rect 19749 9760 19757 9824
rect 19437 9759 19757 9760
rect 17033 9754 17099 9757
rect 17769 9754 17835 9757
rect 17033 9752 17835 9754
rect 17033 9696 17038 9752
rect 17094 9696 17774 9752
rect 17830 9696 17835 9752
rect 17033 9694 17835 9696
rect 17033 9691 17099 9694
rect 17769 9691 17835 9694
rect 18137 9618 18203 9621
rect 8477 9616 12496 9618
rect 8477 9560 8482 9616
rect 8538 9560 12496 9616
rect 8477 9558 12496 9560
rect 15150 9616 18203 9618
rect 15150 9560 18142 9616
rect 18198 9560 18203 9616
rect 15150 9558 18203 9560
rect 8477 9555 8543 9558
rect 4889 9482 4955 9485
rect 5022 9482 5028 9484
rect 4889 9480 5028 9482
rect 4889 9424 4894 9480
rect 4950 9424 5028 9480
rect 4889 9422 5028 9424
rect 4889 9419 4955 9422
rect 5022 9420 5028 9422
rect 5092 9420 5098 9484
rect 6361 9482 6427 9485
rect 15150 9482 15210 9558
rect 18137 9555 18203 9558
rect 18689 9618 18755 9621
rect 19333 9618 19399 9621
rect 18689 9616 19399 9618
rect 18689 9560 18694 9616
rect 18750 9560 19338 9616
rect 19394 9560 19399 9616
rect 18689 9558 19399 9560
rect 18689 9555 18755 9558
rect 19333 9555 19399 9558
rect 6361 9480 15210 9482
rect 6361 9424 6366 9480
rect 6422 9424 15210 9480
rect 6361 9422 15210 9424
rect 17309 9482 17375 9485
rect 19701 9482 19767 9485
rect 17309 9480 19767 9482
rect 17309 9424 17314 9480
rect 17370 9424 19706 9480
rect 19762 9424 19767 9480
rect 17309 9422 19767 9424
rect 6361 9419 6427 9422
rect 17309 9419 17375 9422
rect 19701 9419 19767 9422
rect 21265 9482 21331 9485
rect 23920 9482 24400 9512
rect 21265 9480 24400 9482
rect 21265 9424 21270 9480
rect 21326 9424 24400 9480
rect 21265 9422 24400 9424
rect 21265 9419 21331 9422
rect 23920 9392 24400 9422
rect 8109 9346 8175 9349
rect 7928 9344 8175 9346
rect 7928 9288 8114 9344
rect 8170 9288 8175 9344
rect 7928 9286 8175 9288
rect 7928 9213 7988 9286
rect 8109 9283 8175 9286
rect 8937 9346 9003 9349
rect 11605 9346 11671 9349
rect 8937 9344 11671 9346
rect 8937 9288 8942 9344
rect 8998 9288 11610 9344
rect 11666 9288 11671 9344
rect 8937 9286 11671 9288
rect 8937 9283 9003 9286
rect 11605 9283 11671 9286
rect 11830 9284 11836 9348
rect 11900 9346 11906 9348
rect 12566 9346 12572 9348
rect 11900 9286 12572 9346
rect 11900 9284 11906 9286
rect 12566 9284 12572 9286
rect 12636 9284 12642 9348
rect 17861 9346 17927 9349
rect 19149 9346 19215 9349
rect 17861 9344 19215 9346
rect 17861 9288 17866 9344
rect 17922 9288 19154 9344
rect 19210 9288 19215 9344
rect 17861 9286 19215 9288
rect 17861 9283 17927 9286
rect 19149 9283 19215 9286
rect 8341 9280 8661 9281
rect 8341 9216 8349 9280
rect 8413 9216 8429 9280
rect 8493 9216 8509 9280
rect 8573 9216 8589 9280
rect 8653 9216 8661 9280
rect 8341 9215 8661 9216
rect 15738 9280 16058 9281
rect 15738 9216 15746 9280
rect 15810 9216 15826 9280
rect 15890 9216 15906 9280
rect 15970 9216 15986 9280
rect 16050 9216 16058 9280
rect 15738 9215 16058 9216
rect 6361 9210 6427 9213
rect 7281 9210 7347 9213
rect 6361 9208 7347 9210
rect 6361 9152 6366 9208
rect 6422 9152 7286 9208
rect 7342 9152 7347 9208
rect 6361 9150 7347 9152
rect 6361 9147 6427 9150
rect 7281 9147 7347 9150
rect 7925 9208 7991 9213
rect 10133 9210 10199 9213
rect 7925 9152 7930 9208
rect 7986 9152 7991 9208
rect 7925 9147 7991 9152
rect 9078 9208 10199 9210
rect 9078 9152 10138 9208
rect 10194 9152 10199 9208
rect 9078 9150 10199 9152
rect 0 9074 480 9104
rect 1485 9074 1551 9077
rect 0 9072 1551 9074
rect 0 9016 1490 9072
rect 1546 9016 1551 9072
rect 0 9014 1551 9016
rect 0 8984 480 9014
rect 1485 9011 1551 9014
rect 5533 9074 5599 9077
rect 9078 9074 9138 9150
rect 10133 9147 10199 9150
rect 18505 9210 18571 9213
rect 19241 9210 19307 9213
rect 18505 9208 19307 9210
rect 18505 9152 18510 9208
rect 18566 9152 19246 9208
rect 19302 9152 19307 9208
rect 18505 9150 19307 9152
rect 18505 9147 18571 9150
rect 19241 9147 19307 9150
rect 5533 9072 9138 9074
rect 5533 9016 5538 9072
rect 5594 9016 9138 9072
rect 5533 9014 9138 9016
rect 9489 9074 9555 9077
rect 9622 9074 9628 9076
rect 9489 9072 9628 9074
rect 9489 9016 9494 9072
rect 9550 9016 9628 9072
rect 9489 9014 9628 9016
rect 5533 9011 5599 9014
rect 9489 9011 9555 9014
rect 9622 9012 9628 9014
rect 9692 9012 9698 9076
rect 10225 9074 10291 9077
rect 10409 9074 10475 9077
rect 10225 9072 10475 9074
rect 10225 9016 10230 9072
rect 10286 9016 10414 9072
rect 10470 9016 10475 9072
rect 10225 9014 10475 9016
rect 10225 9011 10291 9014
rect 10409 9011 10475 9014
rect 14733 9074 14799 9077
rect 18137 9074 18203 9077
rect 18873 9074 18939 9077
rect 14733 9072 14842 9074
rect 14733 9016 14738 9072
rect 14794 9016 14842 9072
rect 14733 9011 14842 9016
rect 18137 9072 18939 9074
rect 18137 9016 18142 9072
rect 18198 9016 18878 9072
rect 18934 9016 18939 9072
rect 18137 9014 18939 9016
rect 18137 9011 18203 9014
rect 18873 9011 18939 9014
rect 19057 9074 19123 9077
rect 19885 9074 19951 9077
rect 20161 9074 20227 9077
rect 19057 9072 20227 9074
rect 19057 9016 19062 9072
rect 19118 9016 19890 9072
rect 19946 9016 20166 9072
rect 20222 9016 20227 9072
rect 19057 9014 20227 9016
rect 19057 9011 19123 9014
rect 19885 9011 19951 9014
rect 20161 9011 20227 9014
rect 6862 8876 6868 8940
rect 6932 8938 6938 8940
rect 7005 8938 7071 8941
rect 6932 8936 7071 8938
rect 6932 8880 7010 8936
rect 7066 8880 7071 8936
rect 6932 8878 7071 8880
rect 6932 8876 6938 8878
rect 7005 8875 7071 8878
rect 7189 8938 7255 8941
rect 12709 8938 12775 8941
rect 7189 8936 12775 8938
rect 7189 8880 7194 8936
rect 7250 8880 12714 8936
rect 12770 8880 12775 8936
rect 7189 8878 12775 8880
rect 14782 8938 14842 9011
rect 14917 8938 14983 8941
rect 14782 8936 14983 8938
rect 14782 8880 14922 8936
rect 14978 8880 14983 8936
rect 14782 8878 14983 8880
rect 7189 8875 7255 8878
rect 12709 8875 12775 8878
rect 14917 8875 14983 8878
rect 19190 8876 19196 8940
rect 19260 8938 19266 8940
rect 19333 8938 19399 8941
rect 19260 8936 19399 8938
rect 19260 8880 19338 8936
rect 19394 8880 19399 8936
rect 19260 8878 19399 8880
rect 19260 8876 19266 8878
rect 19333 8875 19399 8878
rect 5390 8802 5396 8804
rect 5030 8742 5396 8802
rect 4642 8736 4962 8737
rect 4642 8672 4650 8736
rect 4714 8672 4730 8736
rect 4794 8672 4810 8736
rect 4874 8672 4890 8736
rect 4954 8672 4962 8736
rect 4642 8671 4962 8672
rect 4337 8530 4403 8533
rect 5030 8530 5090 8742
rect 5390 8740 5396 8742
rect 5460 8802 5466 8804
rect 5460 8742 11898 8802
rect 5460 8740 5466 8742
rect 7649 8668 7715 8669
rect 7598 8604 7604 8668
rect 7668 8666 7715 8668
rect 8937 8666 9003 8669
rect 11421 8666 11487 8669
rect 7668 8664 7760 8666
rect 7710 8608 7760 8664
rect 7668 8606 7760 8608
rect 8937 8664 11487 8666
rect 8937 8608 8942 8664
rect 8998 8608 11426 8664
rect 11482 8608 11487 8664
rect 8937 8606 11487 8608
rect 7668 8604 7715 8606
rect 7649 8603 7715 8604
rect 8937 8603 9003 8606
rect 11421 8603 11487 8606
rect 4337 8528 5090 8530
rect 4337 8472 4342 8528
rect 4398 8472 5090 8528
rect 4337 8470 5090 8472
rect 6729 8530 6795 8533
rect 8150 8530 8156 8532
rect 6729 8528 8156 8530
rect 6729 8472 6734 8528
rect 6790 8472 8156 8528
rect 6729 8470 8156 8472
rect 4337 8467 4403 8470
rect 6729 8467 6795 8470
rect 8150 8468 8156 8470
rect 8220 8468 8226 8532
rect 8385 8530 8451 8533
rect 9857 8530 9923 8533
rect 10358 8530 10364 8532
rect 8385 8528 10364 8530
rect 8385 8472 8390 8528
rect 8446 8472 9862 8528
rect 9918 8472 10364 8528
rect 8385 8470 10364 8472
rect 8385 8467 8451 8470
rect 9857 8467 9923 8470
rect 10358 8468 10364 8470
rect 10428 8468 10434 8532
rect 11838 8530 11898 8742
rect 18638 8740 18644 8804
rect 18708 8802 18714 8804
rect 19241 8802 19307 8805
rect 18708 8800 19307 8802
rect 18708 8744 19246 8800
rect 19302 8744 19307 8800
rect 18708 8742 19307 8744
rect 18708 8740 18714 8742
rect 19241 8739 19307 8742
rect 22461 8802 22527 8805
rect 23920 8802 24400 8832
rect 22461 8800 24400 8802
rect 22461 8744 22466 8800
rect 22522 8744 24400 8800
rect 22461 8742 24400 8744
rect 22461 8739 22527 8742
rect 12040 8736 12360 8737
rect 12040 8672 12048 8736
rect 12112 8672 12128 8736
rect 12192 8672 12208 8736
rect 12272 8672 12288 8736
rect 12352 8672 12360 8736
rect 12040 8671 12360 8672
rect 19437 8736 19757 8737
rect 19437 8672 19445 8736
rect 19509 8672 19525 8736
rect 19589 8672 19605 8736
rect 19669 8672 19685 8736
rect 19749 8672 19757 8736
rect 23920 8712 24400 8742
rect 19437 8671 19757 8672
rect 18454 8604 18460 8668
rect 18524 8666 18530 8668
rect 18873 8666 18939 8669
rect 18524 8664 18939 8666
rect 18524 8608 18878 8664
rect 18934 8608 18939 8664
rect 18524 8606 18939 8608
rect 18524 8604 18530 8606
rect 18873 8603 18939 8606
rect 12157 8530 12223 8533
rect 11838 8528 12223 8530
rect 11838 8472 12162 8528
rect 12218 8472 12223 8528
rect 11838 8470 12223 8472
rect 12157 8467 12223 8470
rect 8293 8394 8359 8397
rect 9990 8394 9996 8396
rect 8293 8392 9996 8394
rect 8293 8336 8298 8392
rect 8354 8336 9996 8392
rect 8293 8334 9996 8336
rect 8293 8331 8359 8334
rect 9990 8332 9996 8334
rect 10060 8332 10066 8396
rect 11789 8394 11855 8397
rect 13353 8396 13419 8397
rect 12934 8394 12940 8396
rect 11789 8392 12940 8394
rect 11789 8336 11794 8392
rect 11850 8336 12940 8392
rect 11789 8334 12940 8336
rect 11789 8331 11855 8334
rect 12934 8332 12940 8334
rect 13004 8332 13010 8396
rect 13302 8394 13308 8396
rect 13262 8334 13308 8394
rect 13372 8392 13419 8396
rect 13414 8336 13419 8392
rect 13302 8332 13308 8334
rect 13372 8332 13419 8336
rect 13353 8331 13419 8332
rect 13629 8394 13695 8397
rect 13629 8392 13922 8394
rect 13629 8336 13634 8392
rect 13690 8336 13922 8392
rect 13629 8334 13922 8336
rect 13629 8331 13695 8334
rect 8753 8258 8819 8261
rect 9254 8258 9260 8260
rect 8753 8256 9260 8258
rect 8753 8200 8758 8256
rect 8814 8200 9260 8256
rect 8753 8198 9260 8200
rect 8753 8195 8819 8198
rect 9254 8196 9260 8198
rect 9324 8196 9330 8260
rect 13862 8258 13922 8334
rect 15518 8334 16314 8394
rect 15518 8258 15578 8334
rect 13862 8198 15578 8258
rect 16254 8258 16314 8334
rect 20478 8258 20484 8260
rect 16254 8198 20484 8258
rect 20478 8196 20484 8198
rect 20548 8196 20554 8260
rect 21265 8258 21331 8261
rect 23920 8258 24400 8288
rect 21265 8256 24400 8258
rect 21265 8200 21270 8256
rect 21326 8200 24400 8256
rect 21265 8198 24400 8200
rect 21265 8195 21331 8198
rect 8341 8192 8661 8193
rect 8341 8128 8349 8192
rect 8413 8128 8429 8192
rect 8493 8128 8509 8192
rect 8573 8128 8589 8192
rect 8653 8128 8661 8192
rect 8341 8127 8661 8128
rect 15738 8192 16058 8193
rect 15738 8128 15746 8192
rect 15810 8128 15826 8192
rect 15890 8128 15906 8192
rect 15970 8128 15986 8192
rect 16050 8128 16058 8192
rect 23920 8168 24400 8198
rect 15738 8127 16058 8128
rect 7005 8122 7071 8125
rect 8845 8124 8911 8125
rect 7230 8122 7236 8124
rect 7005 8120 7236 8122
rect 7005 8064 7010 8120
rect 7066 8064 7236 8120
rect 7005 8062 7236 8064
rect 7005 8059 7071 8062
rect 7230 8060 7236 8062
rect 7300 8060 7306 8124
rect 8845 8120 8892 8124
rect 8956 8122 8962 8124
rect 9121 8122 9187 8125
rect 9990 8122 9996 8124
rect 8845 8064 8850 8120
rect 8845 8060 8892 8064
rect 8956 8062 9002 8122
rect 9121 8120 9996 8122
rect 9121 8064 9126 8120
rect 9182 8064 9996 8120
rect 9121 8062 9996 8064
rect 8956 8060 8962 8062
rect 8845 8059 8911 8060
rect 9121 8059 9187 8062
rect 9990 8060 9996 8062
rect 10060 8060 10066 8124
rect 15009 8122 15075 8125
rect 10182 8120 15075 8122
rect 10182 8064 15014 8120
rect 15070 8064 15075 8120
rect 10182 8062 15075 8064
rect 5625 7986 5691 7989
rect 5758 7986 5764 7988
rect 5625 7984 5764 7986
rect 5625 7928 5630 7984
rect 5686 7928 5764 7984
rect 5625 7926 5764 7928
rect 5625 7923 5691 7926
rect 5758 7924 5764 7926
rect 5828 7924 5834 7988
rect 7925 7986 7991 7989
rect 10182 7986 10242 8062
rect 15009 8059 15075 8062
rect 7925 7984 10242 7986
rect 7925 7928 7930 7984
rect 7986 7928 10242 7984
rect 7925 7926 10242 7928
rect 11605 7986 11671 7989
rect 16573 7986 16639 7989
rect 11605 7984 16639 7986
rect 11605 7928 11610 7984
rect 11666 7928 16578 7984
rect 16634 7928 16639 7984
rect 11605 7926 16639 7928
rect 7925 7923 7991 7926
rect 11605 7923 11671 7926
rect 16573 7923 16639 7926
rect 17217 7986 17283 7989
rect 20989 7986 21055 7989
rect 17217 7984 21055 7986
rect 17217 7928 17222 7984
rect 17278 7928 20994 7984
rect 21050 7928 21055 7984
rect 17217 7926 21055 7928
rect 17217 7923 17283 7926
rect 20989 7923 21055 7926
rect 7557 7850 7623 7853
rect 20110 7850 20116 7852
rect 7557 7848 20116 7850
rect 7557 7792 7562 7848
rect 7618 7792 20116 7848
rect 7557 7790 20116 7792
rect 7557 7787 7623 7790
rect 20110 7788 20116 7790
rect 20180 7788 20186 7852
rect 7189 7714 7255 7717
rect 7414 7714 7420 7716
rect 7189 7712 7420 7714
rect 7189 7656 7194 7712
rect 7250 7656 7420 7712
rect 7189 7654 7420 7656
rect 7189 7651 7255 7654
rect 7414 7652 7420 7654
rect 7484 7652 7490 7716
rect 7557 7714 7623 7717
rect 7782 7714 7788 7716
rect 7557 7712 7788 7714
rect 7557 7656 7562 7712
rect 7618 7656 7788 7712
rect 7557 7654 7788 7656
rect 7557 7651 7623 7654
rect 7782 7652 7788 7654
rect 7852 7652 7858 7716
rect 7925 7714 7991 7717
rect 11605 7714 11671 7717
rect 7925 7712 11671 7714
rect 7925 7656 7930 7712
rect 7986 7656 11610 7712
rect 11666 7656 11671 7712
rect 7925 7654 11671 7656
rect 7925 7651 7991 7654
rect 11605 7651 11671 7654
rect 14457 7714 14523 7717
rect 15009 7714 15075 7717
rect 18597 7714 18663 7717
rect 14457 7712 18663 7714
rect 14457 7656 14462 7712
rect 14518 7656 15014 7712
rect 15070 7656 18602 7712
rect 18658 7656 18663 7712
rect 14457 7654 18663 7656
rect 14457 7651 14523 7654
rect 15009 7651 15075 7654
rect 18597 7651 18663 7654
rect 4642 7648 4962 7649
rect 4642 7584 4650 7648
rect 4714 7584 4730 7648
rect 4794 7584 4810 7648
rect 4874 7584 4890 7648
rect 4954 7584 4962 7648
rect 4642 7583 4962 7584
rect 12040 7648 12360 7649
rect 12040 7584 12048 7648
rect 12112 7584 12128 7648
rect 12192 7584 12208 7648
rect 12272 7584 12288 7648
rect 12352 7584 12360 7648
rect 12040 7583 12360 7584
rect 19437 7648 19757 7649
rect 19437 7584 19445 7648
rect 19509 7584 19525 7648
rect 19589 7584 19605 7648
rect 19669 7584 19685 7648
rect 19749 7584 19757 7648
rect 19437 7583 19757 7584
rect 7925 7578 7991 7581
rect 10961 7578 11027 7581
rect 7925 7576 11027 7578
rect 7925 7520 7930 7576
rect 7986 7520 10966 7576
rect 11022 7520 11027 7576
rect 7925 7518 11027 7520
rect 7925 7515 7991 7518
rect 10961 7515 11027 7518
rect 13077 7578 13143 7581
rect 15142 7578 15148 7580
rect 13077 7576 15148 7578
rect 13077 7520 13082 7576
rect 13138 7520 15148 7576
rect 13077 7518 15148 7520
rect 13077 7515 13143 7518
rect 15142 7516 15148 7518
rect 15212 7516 15218 7580
rect 19006 7578 19012 7580
rect 15702 7518 19012 7578
rect 7925 7442 7991 7445
rect 15702 7442 15762 7518
rect 19006 7516 19012 7518
rect 19076 7516 19082 7580
rect 20989 7578 21055 7581
rect 21449 7578 21515 7581
rect 23920 7578 24400 7608
rect 20989 7576 24400 7578
rect 20989 7520 20994 7576
rect 21050 7520 21454 7576
rect 21510 7520 24400 7576
rect 20989 7518 24400 7520
rect 20989 7515 21055 7518
rect 21449 7515 21515 7518
rect 23920 7488 24400 7518
rect 7925 7440 15762 7442
rect 7925 7384 7930 7440
rect 7986 7384 15762 7440
rect 7925 7382 15762 7384
rect 15837 7442 15903 7445
rect 18045 7442 18111 7445
rect 18413 7442 18479 7445
rect 20253 7442 20319 7445
rect 20713 7442 20779 7445
rect 15837 7440 18479 7442
rect 15837 7384 15842 7440
rect 15898 7384 18050 7440
rect 18106 7384 18418 7440
rect 18474 7384 18479 7440
rect 15837 7382 18479 7384
rect 7925 7379 7991 7382
rect 15837 7379 15903 7382
rect 18045 7379 18111 7382
rect 18413 7379 18479 7382
rect 20118 7440 20319 7442
rect 20118 7384 20258 7440
rect 20314 7384 20319 7440
rect 20118 7382 20319 7384
rect 8937 7306 9003 7309
rect 19241 7306 19307 7309
rect 8937 7304 19307 7306
rect 8937 7248 8942 7304
rect 8998 7248 19246 7304
rect 19302 7248 19307 7304
rect 8937 7246 19307 7248
rect 8937 7243 9003 7246
rect 19241 7243 19307 7246
rect 9806 7170 9812 7172
rect 8756 7110 9812 7170
rect 8341 7104 8661 7105
rect 8341 7040 8349 7104
rect 8413 7040 8429 7104
rect 8493 7040 8509 7104
rect 8573 7040 8589 7104
rect 8653 7040 8661 7104
rect 8341 7039 8661 7040
rect 8756 7037 8816 7110
rect 9806 7108 9812 7110
rect 9876 7108 9882 7172
rect 9990 7108 9996 7172
rect 10060 7170 10066 7172
rect 15009 7170 15075 7173
rect 10060 7168 15075 7170
rect 10060 7112 15014 7168
rect 15070 7112 15075 7168
rect 10060 7110 15075 7112
rect 10060 7108 10066 7110
rect 15009 7107 15075 7110
rect 15738 7104 16058 7105
rect 15738 7040 15746 7104
rect 15810 7040 15826 7104
rect 15890 7040 15906 7104
rect 15970 7040 15986 7104
rect 16050 7040 16058 7104
rect 15738 7039 16058 7040
rect 8753 7032 8819 7037
rect 10685 7034 10751 7037
rect 8753 6976 8758 7032
rect 8814 6976 8819 7032
rect 8753 6971 8819 6976
rect 9630 7032 10751 7034
rect 9630 6976 10690 7032
rect 10746 6976 10751 7032
rect 9630 6974 10751 6976
rect 9630 6901 9690 6974
rect 10685 6971 10751 6974
rect 11789 7034 11855 7037
rect 13629 7036 13695 7037
rect 13629 7034 13676 7036
rect 11789 7032 13676 7034
rect 11789 6976 11794 7032
rect 11850 6976 13634 7032
rect 11789 6974 13676 6976
rect 11789 6971 11855 6974
rect 13629 6972 13676 6974
rect 13740 6972 13746 7036
rect 13629 6971 13695 6972
rect 5165 6898 5231 6901
rect 7966 6898 7972 6900
rect 5165 6896 7972 6898
rect 5165 6840 5170 6896
rect 5226 6840 7972 6896
rect 5165 6838 7972 6840
rect 5165 6835 5231 6838
rect 7966 6836 7972 6838
rect 8036 6836 8042 6900
rect 9581 6896 9690 6901
rect 9581 6840 9586 6896
rect 9642 6840 9690 6896
rect 9581 6838 9690 6840
rect 10041 6898 10107 6901
rect 10593 6898 10659 6901
rect 10041 6896 10659 6898
rect 10041 6840 10046 6896
rect 10102 6840 10598 6896
rect 10654 6840 10659 6896
rect 10041 6838 10659 6840
rect 9581 6835 9647 6838
rect 10041 6835 10107 6838
rect 10593 6835 10659 6838
rect 12341 6898 12407 6901
rect 17033 6898 17099 6901
rect 12341 6896 17099 6898
rect 12341 6840 12346 6896
rect 12402 6840 17038 6896
rect 17094 6840 17099 6896
rect 12341 6838 17099 6840
rect 12341 6835 12407 6838
rect 16300 6765 16360 6838
rect 17033 6835 17099 6838
rect 20118 6765 20178 7382
rect 20253 7379 20319 7382
rect 20670 7440 20779 7442
rect 20670 7384 20718 7440
rect 20774 7384 20779 7440
rect 20670 7379 20779 7384
rect 20670 7306 20730 7379
rect 20624 7246 20730 7306
rect 20624 7173 20684 7246
rect 20621 7168 20687 7173
rect 20621 7112 20626 7168
rect 20682 7112 20687 7168
rect 20621 7107 20687 7112
rect 22737 6898 22803 6901
rect 23920 6898 24400 6928
rect 22737 6896 24400 6898
rect 22737 6840 22742 6896
rect 22798 6840 24400 6896
rect 22737 6838 24400 6840
rect 22737 6835 22803 6838
rect 23920 6808 24400 6838
rect 8569 6762 8635 6765
rect 9489 6762 9555 6765
rect 8569 6760 9555 6762
rect 8569 6704 8574 6760
rect 8630 6704 9494 6760
rect 9550 6704 9555 6760
rect 8569 6702 9555 6704
rect 8569 6699 8635 6702
rect 9489 6699 9555 6702
rect 10133 6762 10199 6765
rect 10133 6760 12818 6762
rect 10133 6704 10138 6760
rect 10194 6704 12818 6760
rect 10133 6702 12818 6704
rect 10133 6699 10199 6702
rect 9029 6628 9095 6629
rect 9489 6628 9555 6629
rect 9029 6626 9076 6628
rect 8984 6624 9076 6626
rect 8984 6568 9034 6624
rect 8984 6566 9076 6568
rect 9029 6564 9076 6566
rect 9140 6564 9146 6628
rect 9438 6564 9444 6628
rect 9508 6626 9555 6628
rect 12758 6626 12818 6702
rect 16297 6760 16363 6765
rect 16297 6704 16302 6760
rect 16358 6704 16363 6760
rect 16297 6699 16363 6704
rect 20069 6760 20178 6765
rect 20069 6704 20074 6760
rect 20130 6704 20178 6760
rect 20069 6702 20178 6704
rect 20069 6699 20135 6702
rect 18822 6626 18828 6628
rect 9508 6624 9600 6626
rect 9550 6568 9600 6624
rect 9508 6566 9600 6568
rect 12758 6566 18828 6626
rect 9508 6564 9555 6566
rect 18822 6564 18828 6566
rect 18892 6564 18898 6628
rect 9029 6563 9095 6564
rect 9489 6563 9555 6564
rect 4642 6560 4962 6561
rect 4642 6496 4650 6560
rect 4714 6496 4730 6560
rect 4794 6496 4810 6560
rect 4874 6496 4890 6560
rect 4954 6496 4962 6560
rect 4642 6495 4962 6496
rect 12040 6560 12360 6561
rect 12040 6496 12048 6560
rect 12112 6496 12128 6560
rect 12192 6496 12208 6560
rect 12272 6496 12288 6560
rect 12352 6496 12360 6560
rect 12040 6495 12360 6496
rect 19437 6560 19757 6561
rect 19437 6496 19445 6560
rect 19509 6496 19525 6560
rect 19589 6496 19605 6560
rect 19669 6496 19685 6560
rect 19749 6496 19757 6560
rect 19437 6495 19757 6496
rect 8385 6490 8451 6493
rect 10501 6490 10567 6493
rect 8385 6488 10567 6490
rect 8385 6432 8390 6488
rect 8446 6432 10506 6488
rect 10562 6432 10567 6488
rect 8385 6430 10567 6432
rect 8385 6427 8451 6430
rect 10501 6427 10567 6430
rect 12617 6490 12683 6493
rect 16849 6490 16915 6493
rect 12617 6488 16915 6490
rect 12617 6432 12622 6488
rect 12678 6432 16854 6488
rect 16910 6432 16915 6488
rect 12617 6430 16915 6432
rect 12617 6427 12683 6430
rect 8661 6354 8727 6357
rect 13854 6354 13860 6356
rect 8661 6352 13860 6354
rect 8661 6296 8666 6352
rect 8722 6296 13860 6352
rect 8661 6294 13860 6296
rect 8661 6291 8727 6294
rect 13854 6292 13860 6294
rect 13924 6292 13930 6356
rect 6494 6156 6500 6220
rect 6564 6218 6570 6220
rect 7925 6218 7991 6221
rect 6564 6216 7991 6218
rect 6564 6160 7930 6216
rect 7986 6160 7991 6216
rect 6564 6158 7991 6160
rect 6564 6156 6570 6158
rect 7925 6155 7991 6158
rect 10174 6156 10180 6220
rect 10244 6218 10250 6220
rect 10317 6218 10383 6221
rect 10244 6216 10383 6218
rect 10244 6160 10322 6216
rect 10378 6160 10383 6216
rect 10244 6158 10383 6160
rect 10244 6156 10250 6158
rect 10317 6155 10383 6158
rect 13813 6082 13879 6085
rect 14000 6082 14060 6430
rect 16849 6427 16915 6430
rect 15009 6354 15075 6357
rect 20989 6354 21055 6357
rect 15009 6352 21055 6354
rect 15009 6296 15014 6352
rect 15070 6296 20994 6352
rect 21050 6296 21055 6352
rect 15009 6294 21055 6296
rect 15009 6291 15075 6294
rect 20989 6291 21055 6294
rect 22461 6218 22527 6221
rect 23920 6218 24400 6248
rect 22461 6216 24400 6218
rect 22461 6160 22466 6216
rect 22522 6160 24400 6216
rect 22461 6158 24400 6160
rect 22461 6155 22527 6158
rect 23920 6128 24400 6158
rect 14457 6082 14523 6085
rect 13813 6080 14060 6082
rect 13813 6024 13818 6080
rect 13874 6024 14060 6080
rect 13813 6022 14060 6024
rect 14414 6080 14523 6082
rect 14414 6024 14462 6080
rect 14518 6024 14523 6080
rect 13813 6019 13879 6022
rect 14414 6019 14523 6024
rect 8341 6016 8661 6017
rect 8341 5952 8349 6016
rect 8413 5952 8429 6016
rect 8493 5952 8509 6016
rect 8573 5952 8589 6016
rect 8653 5952 8661 6016
rect 8341 5951 8661 5952
rect 6545 5946 6611 5949
rect 9305 5948 9371 5949
rect 6678 5946 6684 5948
rect 6545 5944 6684 5946
rect 6545 5888 6550 5944
rect 6606 5888 6684 5944
rect 6545 5886 6684 5888
rect 6545 5883 6611 5886
rect 6678 5884 6684 5886
rect 6748 5884 6754 5948
rect 9254 5884 9260 5948
rect 9324 5946 9371 5948
rect 9673 5946 9739 5949
rect 14181 5946 14247 5949
rect 9324 5944 9416 5946
rect 9366 5888 9416 5944
rect 9324 5886 9416 5888
rect 9673 5944 14247 5946
rect 9673 5888 9678 5944
rect 9734 5888 14186 5944
rect 14242 5888 14247 5944
rect 9673 5886 14247 5888
rect 9324 5884 9371 5886
rect 9305 5883 9371 5884
rect 9673 5883 9739 5886
rect 14181 5883 14247 5886
rect 14414 5813 14474 6019
rect 15738 6016 16058 6017
rect 15738 5952 15746 6016
rect 15810 5952 15826 6016
rect 15890 5952 15906 6016
rect 15970 5952 15986 6016
rect 16050 5952 16058 6016
rect 15738 5951 16058 5952
rect 13629 5812 13695 5813
rect 13629 5808 13676 5812
rect 13740 5810 13746 5812
rect 13629 5752 13634 5808
rect 13629 5748 13676 5752
rect 13740 5750 13786 5810
rect 14365 5808 14474 5813
rect 14365 5752 14370 5808
rect 14426 5752 14474 5808
rect 14365 5750 14474 5752
rect 13740 5748 13746 5750
rect 13629 5747 13695 5748
rect 14365 5747 14431 5750
rect 9397 5674 9463 5677
rect 11830 5674 11836 5676
rect 9397 5672 11836 5674
rect 9397 5616 9402 5672
rect 9458 5616 11836 5672
rect 9397 5614 11836 5616
rect 9397 5611 9463 5614
rect 11830 5612 11836 5614
rect 11900 5612 11906 5676
rect 19149 5674 19215 5677
rect 20345 5674 20411 5677
rect 19149 5672 20411 5674
rect 19149 5616 19154 5672
rect 19210 5616 20350 5672
rect 20406 5616 20411 5672
rect 19149 5614 20411 5616
rect 19149 5611 19215 5614
rect 20345 5611 20411 5614
rect 22829 5538 22895 5541
rect 23920 5538 24400 5568
rect 22829 5536 24400 5538
rect 22829 5480 22834 5536
rect 22890 5480 24400 5536
rect 22829 5478 24400 5480
rect 22829 5475 22895 5478
rect 4642 5472 4962 5473
rect 4642 5408 4650 5472
rect 4714 5408 4730 5472
rect 4794 5408 4810 5472
rect 4874 5408 4890 5472
rect 4954 5408 4962 5472
rect 4642 5407 4962 5408
rect 12040 5472 12360 5473
rect 12040 5408 12048 5472
rect 12112 5408 12128 5472
rect 12192 5408 12208 5472
rect 12272 5408 12288 5472
rect 12352 5408 12360 5472
rect 12040 5407 12360 5408
rect 19437 5472 19757 5473
rect 19437 5408 19445 5472
rect 19509 5408 19525 5472
rect 19589 5408 19605 5472
rect 19669 5408 19685 5472
rect 19749 5408 19757 5472
rect 23920 5448 24400 5478
rect 19437 5407 19757 5408
rect 13721 5402 13787 5405
rect 17677 5402 17743 5405
rect 13721 5400 17743 5402
rect 13721 5344 13726 5400
rect 13782 5344 17682 5400
rect 17738 5344 17743 5400
rect 13721 5342 17743 5344
rect 13721 5339 13787 5342
rect 17677 5339 17743 5342
rect 9857 5266 9923 5269
rect 15561 5266 15627 5269
rect 9857 5264 15627 5266
rect 9857 5208 9862 5264
rect 9918 5208 15566 5264
rect 15622 5208 15627 5264
rect 9857 5206 15627 5208
rect 9857 5203 9923 5206
rect 15561 5203 15627 5206
rect 20069 5266 20135 5269
rect 21357 5266 21423 5269
rect 22093 5266 22159 5269
rect 20069 5264 22159 5266
rect 20069 5208 20074 5264
rect 20130 5208 21362 5264
rect 21418 5208 22098 5264
rect 22154 5208 22159 5264
rect 20069 5206 22159 5208
rect 20069 5203 20135 5206
rect 21357 5203 21423 5206
rect 22093 5203 22159 5206
rect 11697 5130 11763 5133
rect 12433 5130 12499 5133
rect 11697 5128 12499 5130
rect 11697 5072 11702 5128
rect 11758 5072 12438 5128
rect 12494 5072 12499 5128
rect 11697 5070 12499 5072
rect 11697 5067 11763 5070
rect 12433 5067 12499 5070
rect 13813 5130 13879 5133
rect 15653 5130 15719 5133
rect 13813 5128 15719 5130
rect 13813 5072 13818 5128
rect 13874 5072 15658 5128
rect 15714 5072 15719 5128
rect 13813 5070 15719 5072
rect 13813 5067 13879 5070
rect 15653 5067 15719 5070
rect 19425 5130 19491 5133
rect 20713 5130 20779 5133
rect 19425 5128 20779 5130
rect 19425 5072 19430 5128
rect 19486 5072 20718 5128
rect 20774 5072 20779 5128
rect 19425 5070 20779 5072
rect 19425 5067 19491 5070
rect 20713 5067 20779 5070
rect 12249 4994 12315 4997
rect 13905 4994 13971 4997
rect 12249 4992 13971 4994
rect 12249 4936 12254 4992
rect 12310 4936 13910 4992
rect 13966 4936 13971 4992
rect 12249 4934 13971 4936
rect 12249 4931 12315 4934
rect 13905 4931 13971 4934
rect 8341 4928 8661 4929
rect 8341 4864 8349 4928
rect 8413 4864 8429 4928
rect 8493 4864 8509 4928
rect 8573 4864 8589 4928
rect 8653 4864 8661 4928
rect 8341 4863 8661 4864
rect 15738 4928 16058 4929
rect 15738 4864 15746 4928
rect 15810 4864 15826 4928
rect 15890 4864 15906 4928
rect 15970 4864 15986 4928
rect 16050 4864 16058 4928
rect 15738 4863 16058 4864
rect 11697 4858 11763 4861
rect 12341 4858 12407 4861
rect 11697 4856 12407 4858
rect 11697 4800 11702 4856
rect 11758 4800 12346 4856
rect 12402 4800 12407 4856
rect 11697 4798 12407 4800
rect 11697 4795 11763 4798
rect 12341 4795 12407 4798
rect 13353 4858 13419 4861
rect 13997 4858 14063 4861
rect 13353 4856 14063 4858
rect 13353 4800 13358 4856
rect 13414 4800 14002 4856
rect 14058 4800 14063 4856
rect 13353 4798 14063 4800
rect 13353 4795 13419 4798
rect 13997 4795 14063 4798
rect 19885 4858 19951 4861
rect 23920 4858 24400 4888
rect 19885 4856 24400 4858
rect 19885 4800 19890 4856
rect 19946 4800 24400 4856
rect 19885 4798 24400 4800
rect 19885 4795 19951 4798
rect 23920 4768 24400 4798
rect 10317 4722 10383 4725
rect 14641 4722 14707 4725
rect 10317 4720 14707 4722
rect 10317 4664 10322 4720
rect 10378 4664 14646 4720
rect 14702 4664 14707 4720
rect 10317 4662 14707 4664
rect 10317 4659 10383 4662
rect 14641 4659 14707 4662
rect 13905 4586 13971 4589
rect 17401 4586 17467 4589
rect 13905 4584 17467 4586
rect 13905 4528 13910 4584
rect 13966 4528 17406 4584
rect 17462 4528 17467 4584
rect 13905 4526 17467 4528
rect 13905 4523 13971 4526
rect 17401 4523 17467 4526
rect 4642 4384 4962 4385
rect 4642 4320 4650 4384
rect 4714 4320 4730 4384
rect 4794 4320 4810 4384
rect 4874 4320 4890 4384
rect 4954 4320 4962 4384
rect 4642 4319 4962 4320
rect 12040 4384 12360 4385
rect 12040 4320 12048 4384
rect 12112 4320 12128 4384
rect 12192 4320 12208 4384
rect 12272 4320 12288 4384
rect 12352 4320 12360 4384
rect 12040 4319 12360 4320
rect 19437 4384 19757 4385
rect 19437 4320 19445 4384
rect 19509 4320 19525 4384
rect 19589 4320 19605 4384
rect 19669 4320 19685 4384
rect 19749 4320 19757 4384
rect 19437 4319 19757 4320
rect 12985 4314 13051 4317
rect 19241 4314 19307 4317
rect 12985 4312 19307 4314
rect 12985 4256 12990 4312
rect 13046 4256 19246 4312
rect 19302 4256 19307 4312
rect 12985 4254 19307 4256
rect 12985 4251 13051 4254
rect 19241 4251 19307 4254
rect 20161 4314 20227 4317
rect 23920 4314 24400 4344
rect 20161 4312 24400 4314
rect 20161 4256 20166 4312
rect 20222 4256 24400 4312
rect 20161 4254 24400 4256
rect 20161 4251 20227 4254
rect 23920 4224 24400 4254
rect 11881 4180 11947 4181
rect 11830 4116 11836 4180
rect 11900 4178 11947 4180
rect 14365 4178 14431 4181
rect 18413 4178 18479 4181
rect 11900 4176 11992 4178
rect 11942 4120 11992 4176
rect 11900 4118 11992 4120
rect 14365 4176 18479 4178
rect 14365 4120 14370 4176
rect 14426 4120 18418 4176
rect 18474 4120 18479 4176
rect 14365 4118 18479 4120
rect 11900 4116 11947 4118
rect 11881 4115 11947 4116
rect 14365 4115 14431 4118
rect 18413 4115 18479 4118
rect 22001 4178 22067 4181
rect 22369 4178 22435 4181
rect 22001 4176 22435 4178
rect 22001 4120 22006 4176
rect 22062 4120 22374 4176
rect 22430 4120 22435 4176
rect 22001 4118 22435 4120
rect 22001 4115 22067 4118
rect 22369 4115 22435 4118
rect 13997 4044 14063 4045
rect 13997 4042 14044 4044
rect 13952 4040 14044 4042
rect 13952 3984 14002 4040
rect 13952 3982 14044 3984
rect 13997 3980 14044 3982
rect 14108 3980 14114 4044
rect 14641 4042 14707 4045
rect 17125 4042 17191 4045
rect 14641 4040 17191 4042
rect 14641 3984 14646 4040
rect 14702 3984 17130 4040
rect 17186 3984 17191 4040
rect 14641 3982 17191 3984
rect 13997 3979 14063 3980
rect 14641 3979 14707 3982
rect 17125 3979 17191 3982
rect 13077 3906 13143 3909
rect 14406 3906 14412 3908
rect 13077 3904 14412 3906
rect 13077 3848 13082 3904
rect 13138 3848 14412 3904
rect 13077 3846 14412 3848
rect 13077 3843 13143 3846
rect 14406 3844 14412 3846
rect 14476 3844 14482 3908
rect 8341 3840 8661 3841
rect 8341 3776 8349 3840
rect 8413 3776 8429 3840
rect 8493 3776 8509 3840
rect 8573 3776 8589 3840
rect 8653 3776 8661 3840
rect 8341 3775 8661 3776
rect 15738 3840 16058 3841
rect 15738 3776 15746 3840
rect 15810 3776 15826 3840
rect 15890 3776 15906 3840
rect 15970 3776 15986 3840
rect 16050 3776 16058 3840
rect 15738 3775 16058 3776
rect 15561 3634 15627 3637
rect 17953 3634 18019 3637
rect 15561 3632 18019 3634
rect 15561 3576 15566 3632
rect 15622 3576 17958 3632
rect 18014 3576 18019 3632
rect 15561 3574 18019 3576
rect 15561 3571 15627 3574
rect 17953 3571 18019 3574
rect 20529 3634 20595 3637
rect 23920 3634 24400 3664
rect 20529 3632 24400 3634
rect 20529 3576 20534 3632
rect 20590 3576 24400 3632
rect 20529 3574 24400 3576
rect 20529 3571 20595 3574
rect 23920 3544 24400 3574
rect 12617 3362 12683 3365
rect 17534 3362 17540 3364
rect 12617 3360 17540 3362
rect 12617 3304 12622 3360
rect 12678 3304 17540 3360
rect 12617 3302 17540 3304
rect 12617 3299 12683 3302
rect 17534 3300 17540 3302
rect 17604 3300 17610 3364
rect 4642 3296 4962 3297
rect 4642 3232 4650 3296
rect 4714 3232 4730 3296
rect 4794 3232 4810 3296
rect 4874 3232 4890 3296
rect 4954 3232 4962 3296
rect 4642 3231 4962 3232
rect 12040 3296 12360 3297
rect 12040 3232 12048 3296
rect 12112 3232 12128 3296
rect 12192 3232 12208 3296
rect 12272 3232 12288 3296
rect 12352 3232 12360 3296
rect 12040 3231 12360 3232
rect 19437 3296 19757 3297
rect 19437 3232 19445 3296
rect 19509 3232 19525 3296
rect 19589 3232 19605 3296
rect 19669 3232 19685 3296
rect 19749 3232 19757 3296
rect 19437 3231 19757 3232
rect 14089 3226 14155 3229
rect 14222 3226 14228 3228
rect 14089 3224 14228 3226
rect 14089 3168 14094 3224
rect 14150 3168 14228 3224
rect 14089 3166 14228 3168
rect 14089 3163 14155 3166
rect 14222 3164 14228 3166
rect 14292 3164 14298 3228
rect 0 3090 480 3120
rect 1945 3090 2011 3093
rect 0 3088 2011 3090
rect 0 3032 1950 3088
rect 2006 3032 2011 3088
rect 0 3030 2011 3032
rect 0 3000 480 3030
rect 1945 3027 2011 3030
rect 15101 3090 15167 3093
rect 21817 3090 21883 3093
rect 15101 3088 21883 3090
rect 15101 3032 15106 3088
rect 15162 3032 21822 3088
rect 21878 3032 21883 3088
rect 15101 3030 21883 3032
rect 15101 3027 15167 3030
rect 21817 3027 21883 3030
rect 14365 2954 14431 2957
rect 17309 2954 17375 2957
rect 14365 2952 17375 2954
rect 14365 2896 14370 2952
rect 14426 2896 17314 2952
rect 17370 2896 17375 2952
rect 14365 2894 17375 2896
rect 14365 2891 14431 2894
rect 17309 2891 17375 2894
rect 21725 2954 21791 2957
rect 23920 2954 24400 2984
rect 21725 2952 24400 2954
rect 21725 2896 21730 2952
rect 21786 2896 24400 2952
rect 21725 2894 24400 2896
rect 21725 2891 21791 2894
rect 23920 2864 24400 2894
rect 8341 2752 8661 2753
rect 8341 2688 8349 2752
rect 8413 2688 8429 2752
rect 8493 2688 8509 2752
rect 8573 2688 8589 2752
rect 8653 2688 8661 2752
rect 8341 2687 8661 2688
rect 15738 2752 16058 2753
rect 15738 2688 15746 2752
rect 15810 2688 15826 2752
rect 15890 2688 15906 2752
rect 15970 2688 15986 2752
rect 16050 2688 16058 2752
rect 15738 2687 16058 2688
rect 8569 2546 8635 2549
rect 8886 2546 8892 2548
rect 8569 2544 8892 2546
rect 8569 2488 8574 2544
rect 8630 2488 8892 2544
rect 8569 2486 8892 2488
rect 8569 2483 8635 2486
rect 8886 2484 8892 2486
rect 8956 2484 8962 2548
rect 12525 2546 12591 2549
rect 18321 2546 18387 2549
rect 12525 2544 18387 2546
rect 12525 2488 12530 2544
rect 12586 2488 18326 2544
rect 18382 2488 18387 2544
rect 12525 2486 18387 2488
rect 12525 2483 12591 2486
rect 18321 2483 18387 2486
rect 19885 2274 19951 2277
rect 23920 2274 24400 2304
rect 19885 2272 24400 2274
rect 19885 2216 19890 2272
rect 19946 2216 24400 2272
rect 19885 2214 24400 2216
rect 19885 2211 19951 2214
rect 4642 2208 4962 2209
rect 4642 2144 4650 2208
rect 4714 2144 4730 2208
rect 4794 2144 4810 2208
rect 4874 2144 4890 2208
rect 4954 2144 4962 2208
rect 4642 2143 4962 2144
rect 12040 2208 12360 2209
rect 12040 2144 12048 2208
rect 12112 2144 12128 2208
rect 12192 2144 12208 2208
rect 12272 2144 12288 2208
rect 12352 2144 12360 2208
rect 12040 2143 12360 2144
rect 19437 2208 19757 2209
rect 19437 2144 19445 2208
rect 19509 2144 19525 2208
rect 19589 2144 19605 2208
rect 19669 2144 19685 2208
rect 19749 2144 19757 2208
rect 23920 2184 24400 2214
rect 19437 2143 19757 2144
rect 22093 1594 22159 1597
rect 23920 1594 24400 1624
rect 22093 1592 24400 1594
rect 22093 1536 22098 1592
rect 22154 1536 24400 1592
rect 22093 1534 24400 1536
rect 22093 1531 22159 1534
rect 23920 1504 24400 1534
rect 19333 914 19399 917
rect 23920 914 24400 944
rect 19333 912 24400 914
rect 19333 856 19338 912
rect 19394 856 24400 912
rect 19333 854 24400 856
rect 19333 851 19399 854
rect 23920 824 24400 854
rect 22645 370 22711 373
rect 23920 370 24400 400
rect 22645 368 24400 370
rect 22645 312 22650 368
rect 22706 312 24400 368
rect 22645 310 24400 312
rect 22645 307 22711 310
rect 23920 280 24400 310
<< via3 >>
rect 4650 21788 4714 21792
rect 4650 21732 4654 21788
rect 4654 21732 4710 21788
rect 4710 21732 4714 21788
rect 4650 21728 4714 21732
rect 4730 21788 4794 21792
rect 4730 21732 4734 21788
rect 4734 21732 4790 21788
rect 4790 21732 4794 21788
rect 4730 21728 4794 21732
rect 4810 21788 4874 21792
rect 4810 21732 4814 21788
rect 4814 21732 4870 21788
rect 4870 21732 4874 21788
rect 4810 21728 4874 21732
rect 4890 21788 4954 21792
rect 4890 21732 4894 21788
rect 4894 21732 4950 21788
rect 4950 21732 4954 21788
rect 4890 21728 4954 21732
rect 12048 21788 12112 21792
rect 12048 21732 12052 21788
rect 12052 21732 12108 21788
rect 12108 21732 12112 21788
rect 12048 21728 12112 21732
rect 12128 21788 12192 21792
rect 12128 21732 12132 21788
rect 12132 21732 12188 21788
rect 12188 21732 12192 21788
rect 12128 21728 12192 21732
rect 12208 21788 12272 21792
rect 12208 21732 12212 21788
rect 12212 21732 12268 21788
rect 12268 21732 12272 21788
rect 12208 21728 12272 21732
rect 12288 21788 12352 21792
rect 12288 21732 12292 21788
rect 12292 21732 12348 21788
rect 12348 21732 12352 21788
rect 12288 21728 12352 21732
rect 19445 21788 19509 21792
rect 19445 21732 19449 21788
rect 19449 21732 19505 21788
rect 19505 21732 19509 21788
rect 19445 21728 19509 21732
rect 19525 21788 19589 21792
rect 19525 21732 19529 21788
rect 19529 21732 19585 21788
rect 19585 21732 19589 21788
rect 19525 21728 19589 21732
rect 19605 21788 19669 21792
rect 19605 21732 19609 21788
rect 19609 21732 19665 21788
rect 19665 21732 19669 21788
rect 19605 21728 19669 21732
rect 19685 21788 19749 21792
rect 19685 21732 19689 21788
rect 19689 21732 19745 21788
rect 19745 21732 19749 21788
rect 19685 21728 19749 21732
rect 8349 21244 8413 21248
rect 8349 21188 8353 21244
rect 8353 21188 8409 21244
rect 8409 21188 8413 21244
rect 8349 21184 8413 21188
rect 8429 21244 8493 21248
rect 8429 21188 8433 21244
rect 8433 21188 8489 21244
rect 8489 21188 8493 21244
rect 8429 21184 8493 21188
rect 8509 21244 8573 21248
rect 8509 21188 8513 21244
rect 8513 21188 8569 21244
rect 8569 21188 8573 21244
rect 8509 21184 8573 21188
rect 8589 21244 8653 21248
rect 8589 21188 8593 21244
rect 8593 21188 8649 21244
rect 8649 21188 8653 21244
rect 8589 21184 8653 21188
rect 15746 21244 15810 21248
rect 15746 21188 15750 21244
rect 15750 21188 15806 21244
rect 15806 21188 15810 21244
rect 15746 21184 15810 21188
rect 15826 21244 15890 21248
rect 15826 21188 15830 21244
rect 15830 21188 15886 21244
rect 15886 21188 15890 21244
rect 15826 21184 15890 21188
rect 15906 21244 15970 21248
rect 15906 21188 15910 21244
rect 15910 21188 15966 21244
rect 15966 21188 15970 21244
rect 15906 21184 15970 21188
rect 15986 21244 16050 21248
rect 15986 21188 15990 21244
rect 15990 21188 16046 21244
rect 16046 21188 16050 21244
rect 15986 21184 16050 21188
rect 14228 20844 14292 20908
rect 4650 20700 4714 20704
rect 4650 20644 4654 20700
rect 4654 20644 4710 20700
rect 4710 20644 4714 20700
rect 4650 20640 4714 20644
rect 4730 20700 4794 20704
rect 4730 20644 4734 20700
rect 4734 20644 4790 20700
rect 4790 20644 4794 20700
rect 4730 20640 4794 20644
rect 4810 20700 4874 20704
rect 4810 20644 4814 20700
rect 4814 20644 4870 20700
rect 4870 20644 4874 20700
rect 4810 20640 4874 20644
rect 4890 20700 4954 20704
rect 4890 20644 4894 20700
rect 4894 20644 4950 20700
rect 4950 20644 4954 20700
rect 4890 20640 4954 20644
rect 12048 20700 12112 20704
rect 12048 20644 12052 20700
rect 12052 20644 12108 20700
rect 12108 20644 12112 20700
rect 12048 20640 12112 20644
rect 12128 20700 12192 20704
rect 12128 20644 12132 20700
rect 12132 20644 12188 20700
rect 12188 20644 12192 20700
rect 12128 20640 12192 20644
rect 12208 20700 12272 20704
rect 12208 20644 12212 20700
rect 12212 20644 12268 20700
rect 12268 20644 12272 20700
rect 12208 20640 12272 20644
rect 12288 20700 12352 20704
rect 12288 20644 12292 20700
rect 12292 20644 12348 20700
rect 12348 20644 12352 20700
rect 12288 20640 12352 20644
rect 19445 20700 19509 20704
rect 19445 20644 19449 20700
rect 19449 20644 19505 20700
rect 19505 20644 19509 20700
rect 19445 20640 19509 20644
rect 19525 20700 19589 20704
rect 19525 20644 19529 20700
rect 19529 20644 19585 20700
rect 19585 20644 19589 20700
rect 19525 20640 19589 20644
rect 19605 20700 19669 20704
rect 19605 20644 19609 20700
rect 19609 20644 19665 20700
rect 19665 20644 19669 20700
rect 19605 20640 19669 20644
rect 19685 20700 19749 20704
rect 19685 20644 19689 20700
rect 19689 20644 19745 20700
rect 19745 20644 19749 20700
rect 19685 20640 19749 20644
rect 15332 20300 15396 20364
rect 8349 20156 8413 20160
rect 8349 20100 8353 20156
rect 8353 20100 8409 20156
rect 8409 20100 8413 20156
rect 8349 20096 8413 20100
rect 8429 20156 8493 20160
rect 8429 20100 8433 20156
rect 8433 20100 8489 20156
rect 8489 20100 8493 20156
rect 8429 20096 8493 20100
rect 8509 20156 8573 20160
rect 8509 20100 8513 20156
rect 8513 20100 8569 20156
rect 8569 20100 8573 20156
rect 8509 20096 8573 20100
rect 8589 20156 8653 20160
rect 8589 20100 8593 20156
rect 8593 20100 8649 20156
rect 8649 20100 8653 20156
rect 8589 20096 8653 20100
rect 15746 20156 15810 20160
rect 15746 20100 15750 20156
rect 15750 20100 15806 20156
rect 15806 20100 15810 20156
rect 15746 20096 15810 20100
rect 15826 20156 15890 20160
rect 15826 20100 15830 20156
rect 15830 20100 15886 20156
rect 15886 20100 15890 20156
rect 15826 20096 15890 20100
rect 15906 20156 15970 20160
rect 15906 20100 15910 20156
rect 15910 20100 15966 20156
rect 15966 20100 15970 20156
rect 15906 20096 15970 20100
rect 15986 20156 16050 20160
rect 15986 20100 15990 20156
rect 15990 20100 16046 20156
rect 16046 20100 16050 20156
rect 15986 20096 16050 20100
rect 14412 19620 14476 19684
rect 4650 19612 4714 19616
rect 4650 19556 4654 19612
rect 4654 19556 4710 19612
rect 4710 19556 4714 19612
rect 4650 19552 4714 19556
rect 4730 19612 4794 19616
rect 4730 19556 4734 19612
rect 4734 19556 4790 19612
rect 4790 19556 4794 19612
rect 4730 19552 4794 19556
rect 4810 19612 4874 19616
rect 4810 19556 4814 19612
rect 4814 19556 4870 19612
rect 4870 19556 4874 19612
rect 4810 19552 4874 19556
rect 4890 19612 4954 19616
rect 4890 19556 4894 19612
rect 4894 19556 4950 19612
rect 4950 19556 4954 19612
rect 4890 19552 4954 19556
rect 12048 19612 12112 19616
rect 12048 19556 12052 19612
rect 12052 19556 12108 19612
rect 12108 19556 12112 19612
rect 12048 19552 12112 19556
rect 12128 19612 12192 19616
rect 12128 19556 12132 19612
rect 12132 19556 12188 19612
rect 12188 19556 12192 19612
rect 12128 19552 12192 19556
rect 12208 19612 12272 19616
rect 12208 19556 12212 19612
rect 12212 19556 12268 19612
rect 12268 19556 12272 19612
rect 12208 19552 12272 19556
rect 12288 19612 12352 19616
rect 12288 19556 12292 19612
rect 12292 19556 12348 19612
rect 12348 19556 12352 19612
rect 12288 19552 12352 19556
rect 19445 19612 19509 19616
rect 19445 19556 19449 19612
rect 19449 19556 19505 19612
rect 19505 19556 19509 19612
rect 19445 19552 19509 19556
rect 19525 19612 19589 19616
rect 19525 19556 19529 19612
rect 19529 19556 19585 19612
rect 19585 19556 19589 19612
rect 19525 19552 19589 19556
rect 19605 19612 19669 19616
rect 19605 19556 19609 19612
rect 19609 19556 19665 19612
rect 19665 19556 19669 19612
rect 19605 19552 19669 19556
rect 19685 19612 19749 19616
rect 19685 19556 19689 19612
rect 19689 19556 19745 19612
rect 19745 19556 19749 19612
rect 19685 19552 19749 19556
rect 6684 19484 6748 19548
rect 11652 19076 11716 19140
rect 8349 19068 8413 19072
rect 8349 19012 8353 19068
rect 8353 19012 8409 19068
rect 8409 19012 8413 19068
rect 8349 19008 8413 19012
rect 8429 19068 8493 19072
rect 8429 19012 8433 19068
rect 8433 19012 8489 19068
rect 8489 19012 8493 19068
rect 8429 19008 8493 19012
rect 8509 19068 8573 19072
rect 8509 19012 8513 19068
rect 8513 19012 8569 19068
rect 8569 19012 8573 19068
rect 8509 19008 8573 19012
rect 8589 19068 8653 19072
rect 8589 19012 8593 19068
rect 8593 19012 8649 19068
rect 8649 19012 8653 19068
rect 8589 19008 8653 19012
rect 15746 19068 15810 19072
rect 15746 19012 15750 19068
rect 15750 19012 15806 19068
rect 15806 19012 15810 19068
rect 15746 19008 15810 19012
rect 15826 19068 15890 19072
rect 15826 19012 15830 19068
rect 15830 19012 15886 19068
rect 15886 19012 15890 19068
rect 15826 19008 15890 19012
rect 15906 19068 15970 19072
rect 15906 19012 15910 19068
rect 15910 19012 15966 19068
rect 15966 19012 15970 19068
rect 15906 19008 15970 19012
rect 15986 19068 16050 19072
rect 15986 19012 15990 19068
rect 15990 19012 16046 19068
rect 16046 19012 16050 19068
rect 15986 19008 16050 19012
rect 4650 18524 4714 18528
rect 4650 18468 4654 18524
rect 4654 18468 4710 18524
rect 4710 18468 4714 18524
rect 4650 18464 4714 18468
rect 4730 18524 4794 18528
rect 4730 18468 4734 18524
rect 4734 18468 4790 18524
rect 4790 18468 4794 18524
rect 4730 18464 4794 18468
rect 4810 18524 4874 18528
rect 4810 18468 4814 18524
rect 4814 18468 4870 18524
rect 4870 18468 4874 18524
rect 4810 18464 4874 18468
rect 4890 18524 4954 18528
rect 4890 18468 4894 18524
rect 4894 18468 4950 18524
rect 4950 18468 4954 18524
rect 4890 18464 4954 18468
rect 12048 18524 12112 18528
rect 12048 18468 12052 18524
rect 12052 18468 12108 18524
rect 12108 18468 12112 18524
rect 12048 18464 12112 18468
rect 12128 18524 12192 18528
rect 12128 18468 12132 18524
rect 12132 18468 12188 18524
rect 12188 18468 12192 18524
rect 12128 18464 12192 18468
rect 12208 18524 12272 18528
rect 12208 18468 12212 18524
rect 12212 18468 12268 18524
rect 12268 18468 12272 18524
rect 12208 18464 12272 18468
rect 12288 18524 12352 18528
rect 12288 18468 12292 18524
rect 12292 18468 12348 18524
rect 12348 18468 12352 18524
rect 12288 18464 12352 18468
rect 19445 18524 19509 18528
rect 19445 18468 19449 18524
rect 19449 18468 19505 18524
rect 19505 18468 19509 18524
rect 19445 18464 19509 18468
rect 19525 18524 19589 18528
rect 19525 18468 19529 18524
rect 19529 18468 19585 18524
rect 19585 18468 19589 18524
rect 19525 18464 19589 18468
rect 19605 18524 19669 18528
rect 19605 18468 19609 18524
rect 19609 18468 19665 18524
rect 19665 18468 19669 18524
rect 19605 18464 19669 18468
rect 19685 18524 19749 18528
rect 19685 18468 19689 18524
rect 19689 18468 19745 18524
rect 19745 18468 19749 18524
rect 19685 18464 19749 18468
rect 14044 18124 14108 18188
rect 4476 18048 4540 18052
rect 4476 17992 4490 18048
rect 4490 17992 4540 18048
rect 4476 17988 4540 17992
rect 8349 17980 8413 17984
rect 8349 17924 8353 17980
rect 8353 17924 8409 17980
rect 8409 17924 8413 17980
rect 8349 17920 8413 17924
rect 8429 17980 8493 17984
rect 8429 17924 8433 17980
rect 8433 17924 8489 17980
rect 8489 17924 8493 17980
rect 8429 17920 8493 17924
rect 8509 17980 8573 17984
rect 8509 17924 8513 17980
rect 8513 17924 8569 17980
rect 8569 17924 8573 17980
rect 8509 17920 8573 17924
rect 8589 17980 8653 17984
rect 8589 17924 8593 17980
rect 8593 17924 8649 17980
rect 8649 17924 8653 17980
rect 8589 17920 8653 17924
rect 17540 17988 17604 18052
rect 20300 18048 20364 18052
rect 20300 17992 20350 18048
rect 20350 17992 20364 18048
rect 20300 17988 20364 17992
rect 15746 17980 15810 17984
rect 15746 17924 15750 17980
rect 15750 17924 15806 17980
rect 15806 17924 15810 17980
rect 15746 17920 15810 17924
rect 15826 17980 15890 17984
rect 15826 17924 15830 17980
rect 15830 17924 15886 17980
rect 15886 17924 15890 17980
rect 15826 17920 15890 17924
rect 15906 17980 15970 17984
rect 15906 17924 15910 17980
rect 15910 17924 15966 17980
rect 15966 17924 15970 17980
rect 15906 17920 15970 17924
rect 15986 17980 16050 17984
rect 15986 17924 15990 17980
rect 15990 17924 16046 17980
rect 16046 17924 16050 17980
rect 15986 17920 16050 17924
rect 19196 17580 19260 17644
rect 7972 17444 8036 17508
rect 4650 17436 4714 17440
rect 4650 17380 4654 17436
rect 4654 17380 4710 17436
rect 4710 17380 4714 17436
rect 4650 17376 4714 17380
rect 4730 17436 4794 17440
rect 4730 17380 4734 17436
rect 4734 17380 4790 17436
rect 4790 17380 4794 17436
rect 4730 17376 4794 17380
rect 4810 17436 4874 17440
rect 4810 17380 4814 17436
rect 4814 17380 4870 17436
rect 4870 17380 4874 17436
rect 4810 17376 4874 17380
rect 4890 17436 4954 17440
rect 4890 17380 4894 17436
rect 4894 17380 4950 17436
rect 4950 17380 4954 17436
rect 4890 17376 4954 17380
rect 12048 17436 12112 17440
rect 12048 17380 12052 17436
rect 12052 17380 12108 17436
rect 12108 17380 12112 17436
rect 12048 17376 12112 17380
rect 12128 17436 12192 17440
rect 12128 17380 12132 17436
rect 12132 17380 12188 17436
rect 12188 17380 12192 17436
rect 12128 17376 12192 17380
rect 12208 17436 12272 17440
rect 12208 17380 12212 17436
rect 12212 17380 12268 17436
rect 12268 17380 12272 17436
rect 12208 17376 12272 17380
rect 12288 17436 12352 17440
rect 12288 17380 12292 17436
rect 12292 17380 12348 17436
rect 12348 17380 12352 17436
rect 12288 17376 12352 17380
rect 19445 17436 19509 17440
rect 19445 17380 19449 17436
rect 19449 17380 19505 17436
rect 19505 17380 19509 17436
rect 19445 17376 19509 17380
rect 19525 17436 19589 17440
rect 19525 17380 19529 17436
rect 19529 17380 19585 17436
rect 19585 17380 19589 17436
rect 19525 17376 19589 17380
rect 19605 17436 19669 17440
rect 19605 17380 19609 17436
rect 19609 17380 19665 17436
rect 19665 17380 19669 17436
rect 19605 17376 19669 17380
rect 19685 17436 19749 17440
rect 19685 17380 19689 17436
rect 19689 17380 19745 17436
rect 19745 17380 19749 17436
rect 19685 17376 19749 17380
rect 8892 17172 8956 17236
rect 8349 16892 8413 16896
rect 8349 16836 8353 16892
rect 8353 16836 8409 16892
rect 8409 16836 8413 16892
rect 8349 16832 8413 16836
rect 8429 16892 8493 16896
rect 8429 16836 8433 16892
rect 8433 16836 8489 16892
rect 8489 16836 8493 16892
rect 8429 16832 8493 16836
rect 8509 16892 8573 16896
rect 8509 16836 8513 16892
rect 8513 16836 8569 16892
rect 8569 16836 8573 16892
rect 8509 16832 8573 16836
rect 8589 16892 8653 16896
rect 8589 16836 8593 16892
rect 8593 16836 8649 16892
rect 8649 16836 8653 16892
rect 8589 16832 8653 16836
rect 15746 16892 15810 16896
rect 15746 16836 15750 16892
rect 15750 16836 15806 16892
rect 15806 16836 15810 16892
rect 15746 16832 15810 16836
rect 15826 16892 15890 16896
rect 15826 16836 15830 16892
rect 15830 16836 15886 16892
rect 15886 16836 15890 16892
rect 15826 16832 15890 16836
rect 15906 16892 15970 16896
rect 15906 16836 15910 16892
rect 15910 16836 15966 16892
rect 15966 16836 15970 16892
rect 15906 16832 15970 16836
rect 15986 16892 16050 16896
rect 15986 16836 15990 16892
rect 15990 16836 16046 16892
rect 16046 16836 16050 16892
rect 15986 16832 16050 16836
rect 4650 16348 4714 16352
rect 4650 16292 4654 16348
rect 4654 16292 4710 16348
rect 4710 16292 4714 16348
rect 4650 16288 4714 16292
rect 4730 16348 4794 16352
rect 4730 16292 4734 16348
rect 4734 16292 4790 16348
rect 4790 16292 4794 16348
rect 4730 16288 4794 16292
rect 4810 16348 4874 16352
rect 4810 16292 4814 16348
rect 4814 16292 4870 16348
rect 4870 16292 4874 16348
rect 4810 16288 4874 16292
rect 4890 16348 4954 16352
rect 4890 16292 4894 16348
rect 4894 16292 4950 16348
rect 4950 16292 4954 16348
rect 4890 16288 4954 16292
rect 12048 16348 12112 16352
rect 12048 16292 12052 16348
rect 12052 16292 12108 16348
rect 12108 16292 12112 16348
rect 12048 16288 12112 16292
rect 12128 16348 12192 16352
rect 12128 16292 12132 16348
rect 12132 16292 12188 16348
rect 12188 16292 12192 16348
rect 12128 16288 12192 16292
rect 12208 16348 12272 16352
rect 12208 16292 12212 16348
rect 12212 16292 12268 16348
rect 12268 16292 12272 16348
rect 12208 16288 12272 16292
rect 12288 16348 12352 16352
rect 12288 16292 12292 16348
rect 12292 16292 12348 16348
rect 12348 16292 12352 16348
rect 12288 16288 12352 16292
rect 19445 16348 19509 16352
rect 19445 16292 19449 16348
rect 19449 16292 19505 16348
rect 19505 16292 19509 16348
rect 19445 16288 19509 16292
rect 19525 16348 19589 16352
rect 19525 16292 19529 16348
rect 19529 16292 19585 16348
rect 19585 16292 19589 16348
rect 19525 16288 19589 16292
rect 19605 16348 19669 16352
rect 19605 16292 19609 16348
rect 19609 16292 19665 16348
rect 19665 16292 19669 16348
rect 19605 16288 19669 16292
rect 19685 16348 19749 16352
rect 19685 16292 19689 16348
rect 19689 16292 19745 16348
rect 19745 16292 19749 16348
rect 19685 16288 19749 16292
rect 11836 16084 11900 16148
rect 13676 15812 13740 15876
rect 8349 15804 8413 15808
rect 8349 15748 8353 15804
rect 8353 15748 8409 15804
rect 8409 15748 8413 15804
rect 8349 15744 8413 15748
rect 8429 15804 8493 15808
rect 8429 15748 8433 15804
rect 8433 15748 8489 15804
rect 8489 15748 8493 15804
rect 8429 15744 8493 15748
rect 8509 15804 8573 15808
rect 8509 15748 8513 15804
rect 8513 15748 8569 15804
rect 8569 15748 8573 15804
rect 8509 15744 8573 15748
rect 8589 15804 8653 15808
rect 8589 15748 8593 15804
rect 8593 15748 8649 15804
rect 8649 15748 8653 15804
rect 8589 15744 8653 15748
rect 15746 15804 15810 15808
rect 15746 15748 15750 15804
rect 15750 15748 15806 15804
rect 15806 15748 15810 15804
rect 15746 15744 15810 15748
rect 15826 15804 15890 15808
rect 15826 15748 15830 15804
rect 15830 15748 15886 15804
rect 15886 15748 15890 15804
rect 15826 15744 15890 15748
rect 15906 15804 15970 15808
rect 15906 15748 15910 15804
rect 15910 15748 15966 15804
rect 15966 15748 15970 15804
rect 15906 15744 15970 15748
rect 15986 15804 16050 15808
rect 15986 15748 15990 15804
rect 15990 15748 16046 15804
rect 16046 15748 16050 15804
rect 15986 15744 16050 15748
rect 5396 15736 5460 15740
rect 5396 15680 5410 15736
rect 5410 15680 5460 15736
rect 5396 15676 5460 15680
rect 19932 15540 19996 15604
rect 15516 15404 15580 15468
rect 13860 15328 13924 15332
rect 13860 15272 13874 15328
rect 13874 15272 13924 15328
rect 13860 15268 13924 15272
rect 4650 15260 4714 15264
rect 4650 15204 4654 15260
rect 4654 15204 4710 15260
rect 4710 15204 4714 15260
rect 4650 15200 4714 15204
rect 4730 15260 4794 15264
rect 4730 15204 4734 15260
rect 4734 15204 4790 15260
rect 4790 15204 4794 15260
rect 4730 15200 4794 15204
rect 4810 15260 4874 15264
rect 4810 15204 4814 15260
rect 4814 15204 4870 15260
rect 4870 15204 4874 15260
rect 4810 15200 4874 15204
rect 4890 15260 4954 15264
rect 4890 15204 4894 15260
rect 4894 15204 4950 15260
rect 4950 15204 4954 15260
rect 4890 15200 4954 15204
rect 12048 15260 12112 15264
rect 12048 15204 12052 15260
rect 12052 15204 12108 15260
rect 12108 15204 12112 15260
rect 12048 15200 12112 15204
rect 12128 15260 12192 15264
rect 12128 15204 12132 15260
rect 12132 15204 12188 15260
rect 12188 15204 12192 15260
rect 12128 15200 12192 15204
rect 12208 15260 12272 15264
rect 12208 15204 12212 15260
rect 12212 15204 12268 15260
rect 12268 15204 12272 15260
rect 12208 15200 12272 15204
rect 12288 15260 12352 15264
rect 12288 15204 12292 15260
rect 12292 15204 12348 15260
rect 12348 15204 12352 15260
rect 12288 15200 12352 15204
rect 19445 15260 19509 15264
rect 19445 15204 19449 15260
rect 19449 15204 19505 15260
rect 19505 15204 19509 15260
rect 19445 15200 19509 15204
rect 19525 15260 19589 15264
rect 19525 15204 19529 15260
rect 19529 15204 19585 15260
rect 19585 15204 19589 15260
rect 19525 15200 19589 15204
rect 19605 15260 19669 15264
rect 19605 15204 19609 15260
rect 19609 15204 19665 15260
rect 19665 15204 19669 15260
rect 19605 15200 19669 15204
rect 19685 15260 19749 15264
rect 19685 15204 19689 15260
rect 19689 15204 19745 15260
rect 19745 15204 19749 15260
rect 19685 15200 19749 15204
rect 18460 15132 18524 15196
rect 7052 14860 7116 14924
rect 9996 14724 10060 14788
rect 8349 14716 8413 14720
rect 8349 14660 8353 14716
rect 8353 14660 8409 14716
rect 8409 14660 8413 14716
rect 8349 14656 8413 14660
rect 8429 14716 8493 14720
rect 8429 14660 8433 14716
rect 8433 14660 8489 14716
rect 8489 14660 8493 14716
rect 8429 14656 8493 14660
rect 8509 14716 8573 14720
rect 8509 14660 8513 14716
rect 8513 14660 8569 14716
rect 8569 14660 8573 14716
rect 8509 14656 8573 14660
rect 8589 14716 8653 14720
rect 8589 14660 8593 14716
rect 8593 14660 8649 14716
rect 8649 14660 8653 14716
rect 8589 14656 8653 14660
rect 15746 14716 15810 14720
rect 15746 14660 15750 14716
rect 15750 14660 15806 14716
rect 15806 14660 15810 14716
rect 15746 14656 15810 14660
rect 15826 14716 15890 14720
rect 15826 14660 15830 14716
rect 15830 14660 15886 14716
rect 15886 14660 15890 14716
rect 15826 14656 15890 14660
rect 15906 14716 15970 14720
rect 15906 14660 15910 14716
rect 15910 14660 15966 14716
rect 15966 14660 15970 14716
rect 15906 14656 15970 14660
rect 15986 14716 16050 14720
rect 15986 14660 15990 14716
rect 15990 14660 16046 14716
rect 16046 14660 16050 14716
rect 15986 14656 16050 14660
rect 16252 14648 16316 14652
rect 16252 14592 16266 14648
rect 16266 14592 16316 14648
rect 16252 14588 16316 14592
rect 18644 14452 18708 14516
rect 15148 14180 15212 14244
rect 4650 14172 4714 14176
rect 4650 14116 4654 14172
rect 4654 14116 4710 14172
rect 4710 14116 4714 14172
rect 4650 14112 4714 14116
rect 4730 14172 4794 14176
rect 4730 14116 4734 14172
rect 4734 14116 4790 14172
rect 4790 14116 4794 14172
rect 4730 14112 4794 14116
rect 4810 14172 4874 14176
rect 4810 14116 4814 14172
rect 4814 14116 4870 14172
rect 4870 14116 4874 14172
rect 4810 14112 4874 14116
rect 4890 14172 4954 14176
rect 4890 14116 4894 14172
rect 4894 14116 4950 14172
rect 4950 14116 4954 14172
rect 4890 14112 4954 14116
rect 12048 14172 12112 14176
rect 12048 14116 12052 14172
rect 12052 14116 12108 14172
rect 12108 14116 12112 14172
rect 12048 14112 12112 14116
rect 12128 14172 12192 14176
rect 12128 14116 12132 14172
rect 12132 14116 12188 14172
rect 12188 14116 12192 14172
rect 12128 14112 12192 14116
rect 12208 14172 12272 14176
rect 12208 14116 12212 14172
rect 12212 14116 12268 14172
rect 12268 14116 12272 14172
rect 12208 14112 12272 14116
rect 12288 14172 12352 14176
rect 12288 14116 12292 14172
rect 12292 14116 12348 14172
rect 12348 14116 12352 14172
rect 12288 14112 12352 14116
rect 19445 14172 19509 14176
rect 19445 14116 19449 14172
rect 19449 14116 19505 14172
rect 19505 14116 19509 14172
rect 19445 14112 19509 14116
rect 19525 14172 19589 14176
rect 19525 14116 19529 14172
rect 19529 14116 19585 14172
rect 19585 14116 19589 14172
rect 19525 14112 19589 14116
rect 19605 14172 19669 14176
rect 19605 14116 19609 14172
rect 19609 14116 19665 14172
rect 19665 14116 19669 14172
rect 19605 14112 19669 14116
rect 19685 14172 19749 14176
rect 19685 14116 19689 14172
rect 19689 14116 19745 14172
rect 19745 14116 19749 14172
rect 19685 14112 19749 14116
rect 12572 14044 12636 14108
rect 9628 13908 9692 13972
rect 8349 13628 8413 13632
rect 8349 13572 8353 13628
rect 8353 13572 8409 13628
rect 8409 13572 8413 13628
rect 8349 13568 8413 13572
rect 8429 13628 8493 13632
rect 8429 13572 8433 13628
rect 8433 13572 8489 13628
rect 8489 13572 8493 13628
rect 8429 13568 8493 13572
rect 8509 13628 8573 13632
rect 8509 13572 8513 13628
rect 8513 13572 8569 13628
rect 8569 13572 8573 13628
rect 8509 13568 8573 13572
rect 8589 13628 8653 13632
rect 8589 13572 8593 13628
rect 8593 13572 8649 13628
rect 8649 13572 8653 13628
rect 8589 13568 8653 13572
rect 15746 13628 15810 13632
rect 15746 13572 15750 13628
rect 15750 13572 15806 13628
rect 15806 13572 15810 13628
rect 15746 13568 15810 13572
rect 15826 13628 15890 13632
rect 15826 13572 15830 13628
rect 15830 13572 15886 13628
rect 15886 13572 15890 13628
rect 15826 13568 15890 13572
rect 15906 13628 15970 13632
rect 15906 13572 15910 13628
rect 15910 13572 15966 13628
rect 15966 13572 15970 13628
rect 15906 13568 15970 13572
rect 15986 13628 16050 13632
rect 15986 13572 15990 13628
rect 15990 13572 16046 13628
rect 16046 13572 16050 13628
rect 15986 13568 16050 13572
rect 10364 13364 10428 13428
rect 6500 13092 6564 13156
rect 4650 13084 4714 13088
rect 4650 13028 4654 13084
rect 4654 13028 4710 13084
rect 4710 13028 4714 13084
rect 4650 13024 4714 13028
rect 4730 13084 4794 13088
rect 4730 13028 4734 13084
rect 4734 13028 4790 13084
rect 4790 13028 4794 13084
rect 4730 13024 4794 13028
rect 4810 13084 4874 13088
rect 4810 13028 4814 13084
rect 4814 13028 4870 13084
rect 4870 13028 4874 13084
rect 4810 13024 4874 13028
rect 4890 13084 4954 13088
rect 4890 13028 4894 13084
rect 4894 13028 4950 13084
rect 4950 13028 4954 13084
rect 4890 13024 4954 13028
rect 12048 13084 12112 13088
rect 12048 13028 12052 13084
rect 12052 13028 12108 13084
rect 12108 13028 12112 13084
rect 12048 13024 12112 13028
rect 12128 13084 12192 13088
rect 12128 13028 12132 13084
rect 12132 13028 12188 13084
rect 12188 13028 12192 13084
rect 12128 13024 12192 13028
rect 12208 13084 12272 13088
rect 12208 13028 12212 13084
rect 12212 13028 12268 13084
rect 12268 13028 12272 13084
rect 12208 13024 12272 13028
rect 12288 13084 12352 13088
rect 12288 13028 12292 13084
rect 12292 13028 12348 13084
rect 12348 13028 12352 13084
rect 12288 13024 12352 13028
rect 19445 13084 19509 13088
rect 19445 13028 19449 13084
rect 19449 13028 19505 13084
rect 19505 13028 19509 13084
rect 19445 13024 19509 13028
rect 19525 13084 19589 13088
rect 19525 13028 19529 13084
rect 19529 13028 19585 13084
rect 19585 13028 19589 13084
rect 19525 13024 19589 13028
rect 19605 13084 19669 13088
rect 19605 13028 19609 13084
rect 19609 13028 19665 13084
rect 19665 13028 19669 13084
rect 19605 13024 19669 13028
rect 19685 13084 19749 13088
rect 19685 13028 19689 13084
rect 19689 13028 19745 13084
rect 19745 13028 19749 13084
rect 19685 13024 19749 13028
rect 4476 12744 4540 12748
rect 4476 12688 4526 12744
rect 4526 12688 4540 12744
rect 4476 12684 4540 12688
rect 5764 12684 5828 12748
rect 11652 12548 11716 12612
rect 8349 12540 8413 12544
rect 8349 12484 8353 12540
rect 8353 12484 8409 12540
rect 8409 12484 8413 12540
rect 8349 12480 8413 12484
rect 8429 12540 8493 12544
rect 8429 12484 8433 12540
rect 8433 12484 8489 12540
rect 8489 12484 8493 12540
rect 8429 12480 8493 12484
rect 8509 12540 8573 12544
rect 8509 12484 8513 12540
rect 8513 12484 8569 12540
rect 8569 12484 8573 12540
rect 8509 12480 8573 12484
rect 8589 12540 8653 12544
rect 8589 12484 8593 12540
rect 8593 12484 8649 12540
rect 8649 12484 8653 12540
rect 8589 12480 8653 12484
rect 6316 12412 6380 12476
rect 12756 12548 12820 12612
rect 15746 12540 15810 12544
rect 15746 12484 15750 12540
rect 15750 12484 15806 12540
rect 15806 12484 15810 12540
rect 15746 12480 15810 12484
rect 15826 12540 15890 12544
rect 15826 12484 15830 12540
rect 15830 12484 15886 12540
rect 15886 12484 15890 12540
rect 15826 12480 15890 12484
rect 15906 12540 15970 12544
rect 15906 12484 15910 12540
rect 15910 12484 15966 12540
rect 15966 12484 15970 12540
rect 15906 12480 15970 12484
rect 15986 12540 16050 12544
rect 15986 12484 15990 12540
rect 15990 12484 16046 12540
rect 16046 12484 16050 12540
rect 15986 12480 16050 12484
rect 12940 12412 13004 12476
rect 20116 12608 20180 12612
rect 20116 12552 20130 12608
rect 20130 12552 20180 12608
rect 20116 12548 20180 12552
rect 20484 12472 20548 12476
rect 20484 12416 20534 12472
rect 20534 12416 20548 12472
rect 20484 12412 20548 12416
rect 5764 12140 5828 12204
rect 6316 12004 6380 12068
rect 4650 11996 4714 12000
rect 4650 11940 4654 11996
rect 4654 11940 4710 11996
rect 4710 11940 4714 11996
rect 4650 11936 4714 11940
rect 4730 11996 4794 12000
rect 4730 11940 4734 11996
rect 4734 11940 4790 11996
rect 4790 11940 4794 11996
rect 4730 11936 4794 11940
rect 4810 11996 4874 12000
rect 4810 11940 4814 11996
rect 4814 11940 4870 11996
rect 4870 11940 4874 11996
rect 4810 11936 4874 11940
rect 4890 11996 4954 12000
rect 4890 11940 4894 11996
rect 4894 11940 4950 11996
rect 4950 11940 4954 11996
rect 4890 11936 4954 11940
rect 13308 12276 13372 12340
rect 12756 12200 12820 12204
rect 12756 12144 12770 12200
rect 12770 12144 12820 12200
rect 12756 12140 12820 12144
rect 18828 12004 18892 12068
rect 12048 11996 12112 12000
rect 12048 11940 12052 11996
rect 12052 11940 12108 11996
rect 12108 11940 12112 11996
rect 12048 11936 12112 11940
rect 12128 11996 12192 12000
rect 12128 11940 12132 11996
rect 12132 11940 12188 11996
rect 12188 11940 12192 11996
rect 12128 11936 12192 11940
rect 12208 11996 12272 12000
rect 12208 11940 12212 11996
rect 12212 11940 12268 11996
rect 12268 11940 12272 11996
rect 12208 11936 12272 11940
rect 12288 11996 12352 12000
rect 12288 11940 12292 11996
rect 12292 11940 12348 11996
rect 12348 11940 12352 11996
rect 12288 11936 12352 11940
rect 19445 11996 19509 12000
rect 19445 11940 19449 11996
rect 19449 11940 19505 11996
rect 19505 11940 19509 11996
rect 19445 11936 19509 11940
rect 19525 11996 19589 12000
rect 19525 11940 19529 11996
rect 19529 11940 19585 11996
rect 19585 11940 19589 11996
rect 19525 11936 19589 11940
rect 19605 11996 19669 12000
rect 19605 11940 19609 11996
rect 19609 11940 19665 11996
rect 19665 11940 19669 11996
rect 19605 11936 19669 11940
rect 19685 11996 19749 12000
rect 19685 11940 19689 11996
rect 19689 11940 19745 11996
rect 19745 11940 19749 11996
rect 19685 11936 19749 11940
rect 19012 11928 19076 11932
rect 19012 11872 19026 11928
rect 19026 11872 19076 11928
rect 19012 11868 19076 11872
rect 8349 11452 8413 11456
rect 8349 11396 8353 11452
rect 8353 11396 8409 11452
rect 8409 11396 8413 11452
rect 8349 11392 8413 11396
rect 8429 11452 8493 11456
rect 8429 11396 8433 11452
rect 8433 11396 8489 11452
rect 8489 11396 8493 11452
rect 8429 11392 8493 11396
rect 8509 11452 8573 11456
rect 8509 11396 8513 11452
rect 8513 11396 8569 11452
rect 8569 11396 8573 11452
rect 8509 11392 8573 11396
rect 8589 11452 8653 11456
rect 8589 11396 8593 11452
rect 8593 11396 8649 11452
rect 8649 11396 8653 11452
rect 8589 11392 8653 11396
rect 15746 11452 15810 11456
rect 15746 11396 15750 11452
rect 15750 11396 15806 11452
rect 15806 11396 15810 11452
rect 15746 11392 15810 11396
rect 15826 11452 15890 11456
rect 15826 11396 15830 11452
rect 15830 11396 15886 11452
rect 15886 11396 15890 11452
rect 15826 11392 15890 11396
rect 15906 11452 15970 11456
rect 15906 11396 15910 11452
rect 15910 11396 15966 11452
rect 15966 11396 15970 11452
rect 15906 11392 15970 11396
rect 15986 11452 16050 11456
rect 15986 11396 15990 11452
rect 15990 11396 16046 11452
rect 16046 11396 16050 11452
rect 15986 11392 16050 11396
rect 8156 11188 8220 11252
rect 15332 11324 15396 11388
rect 20300 11324 20364 11388
rect 5028 11052 5092 11116
rect 15148 11052 15212 11116
rect 4650 10908 4714 10912
rect 4650 10852 4654 10908
rect 4654 10852 4710 10908
rect 4710 10852 4714 10908
rect 4650 10848 4714 10852
rect 4730 10908 4794 10912
rect 4730 10852 4734 10908
rect 4734 10852 4790 10908
rect 4790 10852 4794 10908
rect 4730 10848 4794 10852
rect 4810 10908 4874 10912
rect 4810 10852 4814 10908
rect 4814 10852 4870 10908
rect 4870 10852 4874 10908
rect 4810 10848 4874 10852
rect 4890 10908 4954 10912
rect 4890 10852 4894 10908
rect 4894 10852 4950 10908
rect 4950 10852 4954 10908
rect 4890 10848 4954 10852
rect 12048 10908 12112 10912
rect 12048 10852 12052 10908
rect 12052 10852 12108 10908
rect 12108 10852 12112 10908
rect 12048 10848 12112 10852
rect 12128 10908 12192 10912
rect 12128 10852 12132 10908
rect 12132 10852 12188 10908
rect 12188 10852 12192 10908
rect 12128 10848 12192 10852
rect 12208 10908 12272 10912
rect 12208 10852 12212 10908
rect 12212 10852 12268 10908
rect 12268 10852 12272 10908
rect 12208 10848 12272 10852
rect 12288 10908 12352 10912
rect 12288 10852 12292 10908
rect 12292 10852 12348 10908
rect 12348 10852 12352 10908
rect 12288 10848 12352 10852
rect 19445 10908 19509 10912
rect 19445 10852 19449 10908
rect 19449 10852 19505 10908
rect 19505 10852 19509 10908
rect 19445 10848 19509 10852
rect 19525 10908 19589 10912
rect 19525 10852 19529 10908
rect 19529 10852 19585 10908
rect 19585 10852 19589 10908
rect 19525 10848 19589 10852
rect 19605 10908 19669 10912
rect 19605 10852 19609 10908
rect 19609 10852 19665 10908
rect 19665 10852 19669 10908
rect 19605 10848 19669 10852
rect 19685 10908 19749 10912
rect 19685 10852 19689 10908
rect 19689 10852 19745 10908
rect 19745 10852 19749 10908
rect 19685 10848 19749 10852
rect 5764 10780 5828 10844
rect 15516 10780 15580 10844
rect 7236 10644 7300 10708
rect 11836 10644 11900 10708
rect 9444 10508 9508 10572
rect 9812 10372 9876 10436
rect 19932 10644 19996 10708
rect 12940 10508 13004 10572
rect 8349 10364 8413 10368
rect 8349 10308 8353 10364
rect 8353 10308 8409 10364
rect 8409 10308 8413 10364
rect 8349 10304 8413 10308
rect 8429 10364 8493 10368
rect 8429 10308 8433 10364
rect 8433 10308 8489 10364
rect 8489 10308 8493 10364
rect 8429 10304 8493 10308
rect 8509 10364 8573 10368
rect 8509 10308 8513 10364
rect 8513 10308 8569 10364
rect 8569 10308 8573 10364
rect 8509 10304 8573 10308
rect 8589 10364 8653 10368
rect 8589 10308 8593 10364
rect 8593 10308 8649 10364
rect 8649 10308 8653 10364
rect 8589 10304 8653 10308
rect 5764 10236 5828 10300
rect 13676 10236 13740 10300
rect 15746 10364 15810 10368
rect 15746 10308 15750 10364
rect 15750 10308 15806 10364
rect 15806 10308 15810 10364
rect 15746 10304 15810 10308
rect 15826 10364 15890 10368
rect 15826 10308 15830 10364
rect 15830 10308 15886 10364
rect 15886 10308 15890 10364
rect 15826 10304 15890 10308
rect 15906 10364 15970 10368
rect 15906 10308 15910 10364
rect 15910 10308 15966 10364
rect 15966 10308 15970 10364
rect 15906 10304 15970 10308
rect 15986 10364 16050 10368
rect 15986 10308 15990 10364
rect 15990 10308 16046 10364
rect 16046 10308 16050 10364
rect 15986 10304 16050 10308
rect 7420 10100 7484 10164
rect 8892 10100 8956 10164
rect 6868 9964 6932 10028
rect 16252 10100 16316 10164
rect 7604 9828 7668 9892
rect 8892 9828 8956 9892
rect 4650 9820 4714 9824
rect 4650 9764 4654 9820
rect 4654 9764 4710 9820
rect 4710 9764 4714 9820
rect 4650 9760 4714 9764
rect 4730 9820 4794 9824
rect 4730 9764 4734 9820
rect 4734 9764 4790 9820
rect 4790 9764 4794 9820
rect 4730 9760 4794 9764
rect 4810 9820 4874 9824
rect 4810 9764 4814 9820
rect 4814 9764 4870 9820
rect 4870 9764 4874 9820
rect 4810 9760 4874 9764
rect 4890 9820 4954 9824
rect 4890 9764 4894 9820
rect 4894 9764 4950 9820
rect 4950 9764 4954 9820
rect 4890 9760 4954 9764
rect 12048 9820 12112 9824
rect 12048 9764 12052 9820
rect 12052 9764 12108 9820
rect 12108 9764 12112 9820
rect 12048 9760 12112 9764
rect 12128 9820 12192 9824
rect 12128 9764 12132 9820
rect 12132 9764 12188 9820
rect 12188 9764 12192 9820
rect 12128 9760 12192 9764
rect 12208 9820 12272 9824
rect 12208 9764 12212 9820
rect 12212 9764 12268 9820
rect 12268 9764 12272 9820
rect 12208 9760 12272 9764
rect 12288 9820 12352 9824
rect 12288 9764 12292 9820
rect 12292 9764 12348 9820
rect 12348 9764 12352 9820
rect 12288 9760 12352 9764
rect 7052 9692 7116 9756
rect 7788 9692 7852 9756
rect 10180 9692 10244 9756
rect 19445 9820 19509 9824
rect 19445 9764 19449 9820
rect 19449 9764 19505 9820
rect 19505 9764 19509 9820
rect 19445 9760 19509 9764
rect 19525 9820 19589 9824
rect 19525 9764 19529 9820
rect 19529 9764 19585 9820
rect 19585 9764 19589 9820
rect 19525 9760 19589 9764
rect 19605 9820 19669 9824
rect 19605 9764 19609 9820
rect 19609 9764 19665 9820
rect 19665 9764 19669 9820
rect 19605 9760 19669 9764
rect 19685 9820 19749 9824
rect 19685 9764 19689 9820
rect 19689 9764 19745 9820
rect 19745 9764 19749 9820
rect 19685 9760 19749 9764
rect 5028 9420 5092 9484
rect 11836 9284 11900 9348
rect 12572 9284 12636 9348
rect 8349 9276 8413 9280
rect 8349 9220 8353 9276
rect 8353 9220 8409 9276
rect 8409 9220 8413 9276
rect 8349 9216 8413 9220
rect 8429 9276 8493 9280
rect 8429 9220 8433 9276
rect 8433 9220 8489 9276
rect 8489 9220 8493 9276
rect 8429 9216 8493 9220
rect 8509 9276 8573 9280
rect 8509 9220 8513 9276
rect 8513 9220 8569 9276
rect 8569 9220 8573 9276
rect 8509 9216 8573 9220
rect 8589 9276 8653 9280
rect 8589 9220 8593 9276
rect 8593 9220 8649 9276
rect 8649 9220 8653 9276
rect 8589 9216 8653 9220
rect 15746 9276 15810 9280
rect 15746 9220 15750 9276
rect 15750 9220 15806 9276
rect 15806 9220 15810 9276
rect 15746 9216 15810 9220
rect 15826 9276 15890 9280
rect 15826 9220 15830 9276
rect 15830 9220 15886 9276
rect 15886 9220 15890 9276
rect 15826 9216 15890 9220
rect 15906 9276 15970 9280
rect 15906 9220 15910 9276
rect 15910 9220 15966 9276
rect 15966 9220 15970 9276
rect 15906 9216 15970 9220
rect 15986 9276 16050 9280
rect 15986 9220 15990 9276
rect 15990 9220 16046 9276
rect 16046 9220 16050 9276
rect 15986 9216 16050 9220
rect 9628 9012 9692 9076
rect 6868 8876 6932 8940
rect 19196 8876 19260 8940
rect 4650 8732 4714 8736
rect 4650 8676 4654 8732
rect 4654 8676 4710 8732
rect 4710 8676 4714 8732
rect 4650 8672 4714 8676
rect 4730 8732 4794 8736
rect 4730 8676 4734 8732
rect 4734 8676 4790 8732
rect 4790 8676 4794 8732
rect 4730 8672 4794 8676
rect 4810 8732 4874 8736
rect 4810 8676 4814 8732
rect 4814 8676 4870 8732
rect 4870 8676 4874 8732
rect 4810 8672 4874 8676
rect 4890 8732 4954 8736
rect 4890 8676 4894 8732
rect 4894 8676 4950 8732
rect 4950 8676 4954 8732
rect 4890 8672 4954 8676
rect 5396 8740 5460 8804
rect 7604 8664 7668 8668
rect 7604 8608 7654 8664
rect 7654 8608 7668 8664
rect 7604 8604 7668 8608
rect 8156 8468 8220 8532
rect 10364 8468 10428 8532
rect 18644 8740 18708 8804
rect 12048 8732 12112 8736
rect 12048 8676 12052 8732
rect 12052 8676 12108 8732
rect 12108 8676 12112 8732
rect 12048 8672 12112 8676
rect 12128 8732 12192 8736
rect 12128 8676 12132 8732
rect 12132 8676 12188 8732
rect 12188 8676 12192 8732
rect 12128 8672 12192 8676
rect 12208 8732 12272 8736
rect 12208 8676 12212 8732
rect 12212 8676 12268 8732
rect 12268 8676 12272 8732
rect 12208 8672 12272 8676
rect 12288 8732 12352 8736
rect 12288 8676 12292 8732
rect 12292 8676 12348 8732
rect 12348 8676 12352 8732
rect 12288 8672 12352 8676
rect 19445 8732 19509 8736
rect 19445 8676 19449 8732
rect 19449 8676 19505 8732
rect 19505 8676 19509 8732
rect 19445 8672 19509 8676
rect 19525 8732 19589 8736
rect 19525 8676 19529 8732
rect 19529 8676 19585 8732
rect 19585 8676 19589 8732
rect 19525 8672 19589 8676
rect 19605 8732 19669 8736
rect 19605 8676 19609 8732
rect 19609 8676 19665 8732
rect 19665 8676 19669 8732
rect 19605 8672 19669 8676
rect 19685 8732 19749 8736
rect 19685 8676 19689 8732
rect 19689 8676 19745 8732
rect 19745 8676 19749 8732
rect 19685 8672 19749 8676
rect 18460 8604 18524 8668
rect 9996 8332 10060 8396
rect 12940 8332 13004 8396
rect 13308 8392 13372 8396
rect 13308 8336 13358 8392
rect 13358 8336 13372 8392
rect 13308 8332 13372 8336
rect 9260 8196 9324 8260
rect 20484 8196 20548 8260
rect 8349 8188 8413 8192
rect 8349 8132 8353 8188
rect 8353 8132 8409 8188
rect 8409 8132 8413 8188
rect 8349 8128 8413 8132
rect 8429 8188 8493 8192
rect 8429 8132 8433 8188
rect 8433 8132 8489 8188
rect 8489 8132 8493 8188
rect 8429 8128 8493 8132
rect 8509 8188 8573 8192
rect 8509 8132 8513 8188
rect 8513 8132 8569 8188
rect 8569 8132 8573 8188
rect 8509 8128 8573 8132
rect 8589 8188 8653 8192
rect 8589 8132 8593 8188
rect 8593 8132 8649 8188
rect 8649 8132 8653 8188
rect 8589 8128 8653 8132
rect 15746 8188 15810 8192
rect 15746 8132 15750 8188
rect 15750 8132 15806 8188
rect 15806 8132 15810 8188
rect 15746 8128 15810 8132
rect 15826 8188 15890 8192
rect 15826 8132 15830 8188
rect 15830 8132 15886 8188
rect 15886 8132 15890 8188
rect 15826 8128 15890 8132
rect 15906 8188 15970 8192
rect 15906 8132 15910 8188
rect 15910 8132 15966 8188
rect 15966 8132 15970 8188
rect 15906 8128 15970 8132
rect 15986 8188 16050 8192
rect 15986 8132 15990 8188
rect 15990 8132 16046 8188
rect 16046 8132 16050 8188
rect 15986 8128 16050 8132
rect 7236 8060 7300 8124
rect 8892 8120 8956 8124
rect 8892 8064 8906 8120
rect 8906 8064 8956 8120
rect 8892 8060 8956 8064
rect 9996 8060 10060 8124
rect 5764 7924 5828 7988
rect 20116 7788 20180 7852
rect 7420 7652 7484 7716
rect 7788 7652 7852 7716
rect 4650 7644 4714 7648
rect 4650 7588 4654 7644
rect 4654 7588 4710 7644
rect 4710 7588 4714 7644
rect 4650 7584 4714 7588
rect 4730 7644 4794 7648
rect 4730 7588 4734 7644
rect 4734 7588 4790 7644
rect 4790 7588 4794 7644
rect 4730 7584 4794 7588
rect 4810 7644 4874 7648
rect 4810 7588 4814 7644
rect 4814 7588 4870 7644
rect 4870 7588 4874 7644
rect 4810 7584 4874 7588
rect 4890 7644 4954 7648
rect 4890 7588 4894 7644
rect 4894 7588 4950 7644
rect 4950 7588 4954 7644
rect 4890 7584 4954 7588
rect 12048 7644 12112 7648
rect 12048 7588 12052 7644
rect 12052 7588 12108 7644
rect 12108 7588 12112 7644
rect 12048 7584 12112 7588
rect 12128 7644 12192 7648
rect 12128 7588 12132 7644
rect 12132 7588 12188 7644
rect 12188 7588 12192 7644
rect 12128 7584 12192 7588
rect 12208 7644 12272 7648
rect 12208 7588 12212 7644
rect 12212 7588 12268 7644
rect 12268 7588 12272 7644
rect 12208 7584 12272 7588
rect 12288 7644 12352 7648
rect 12288 7588 12292 7644
rect 12292 7588 12348 7644
rect 12348 7588 12352 7644
rect 12288 7584 12352 7588
rect 19445 7644 19509 7648
rect 19445 7588 19449 7644
rect 19449 7588 19505 7644
rect 19505 7588 19509 7644
rect 19445 7584 19509 7588
rect 19525 7644 19589 7648
rect 19525 7588 19529 7644
rect 19529 7588 19585 7644
rect 19585 7588 19589 7644
rect 19525 7584 19589 7588
rect 19605 7644 19669 7648
rect 19605 7588 19609 7644
rect 19609 7588 19665 7644
rect 19665 7588 19669 7644
rect 19605 7584 19669 7588
rect 19685 7644 19749 7648
rect 19685 7588 19689 7644
rect 19689 7588 19745 7644
rect 19745 7588 19749 7644
rect 19685 7584 19749 7588
rect 15148 7516 15212 7580
rect 19012 7516 19076 7580
rect 8349 7100 8413 7104
rect 8349 7044 8353 7100
rect 8353 7044 8409 7100
rect 8409 7044 8413 7100
rect 8349 7040 8413 7044
rect 8429 7100 8493 7104
rect 8429 7044 8433 7100
rect 8433 7044 8489 7100
rect 8489 7044 8493 7100
rect 8429 7040 8493 7044
rect 8509 7100 8573 7104
rect 8509 7044 8513 7100
rect 8513 7044 8569 7100
rect 8569 7044 8573 7100
rect 8509 7040 8573 7044
rect 8589 7100 8653 7104
rect 8589 7044 8593 7100
rect 8593 7044 8649 7100
rect 8649 7044 8653 7100
rect 8589 7040 8653 7044
rect 9812 7108 9876 7172
rect 9996 7108 10060 7172
rect 15746 7100 15810 7104
rect 15746 7044 15750 7100
rect 15750 7044 15806 7100
rect 15806 7044 15810 7100
rect 15746 7040 15810 7044
rect 15826 7100 15890 7104
rect 15826 7044 15830 7100
rect 15830 7044 15886 7100
rect 15886 7044 15890 7100
rect 15826 7040 15890 7044
rect 15906 7100 15970 7104
rect 15906 7044 15910 7100
rect 15910 7044 15966 7100
rect 15966 7044 15970 7100
rect 15906 7040 15970 7044
rect 15986 7100 16050 7104
rect 15986 7044 15990 7100
rect 15990 7044 16046 7100
rect 16046 7044 16050 7100
rect 15986 7040 16050 7044
rect 13676 7032 13740 7036
rect 13676 6976 13690 7032
rect 13690 6976 13740 7032
rect 13676 6972 13740 6976
rect 7972 6836 8036 6900
rect 9076 6624 9140 6628
rect 9076 6568 9090 6624
rect 9090 6568 9140 6624
rect 9076 6564 9140 6568
rect 9444 6624 9508 6628
rect 9444 6568 9494 6624
rect 9494 6568 9508 6624
rect 9444 6564 9508 6568
rect 18828 6564 18892 6628
rect 4650 6556 4714 6560
rect 4650 6500 4654 6556
rect 4654 6500 4710 6556
rect 4710 6500 4714 6556
rect 4650 6496 4714 6500
rect 4730 6556 4794 6560
rect 4730 6500 4734 6556
rect 4734 6500 4790 6556
rect 4790 6500 4794 6556
rect 4730 6496 4794 6500
rect 4810 6556 4874 6560
rect 4810 6500 4814 6556
rect 4814 6500 4870 6556
rect 4870 6500 4874 6556
rect 4810 6496 4874 6500
rect 4890 6556 4954 6560
rect 4890 6500 4894 6556
rect 4894 6500 4950 6556
rect 4950 6500 4954 6556
rect 4890 6496 4954 6500
rect 12048 6556 12112 6560
rect 12048 6500 12052 6556
rect 12052 6500 12108 6556
rect 12108 6500 12112 6556
rect 12048 6496 12112 6500
rect 12128 6556 12192 6560
rect 12128 6500 12132 6556
rect 12132 6500 12188 6556
rect 12188 6500 12192 6556
rect 12128 6496 12192 6500
rect 12208 6556 12272 6560
rect 12208 6500 12212 6556
rect 12212 6500 12268 6556
rect 12268 6500 12272 6556
rect 12208 6496 12272 6500
rect 12288 6556 12352 6560
rect 12288 6500 12292 6556
rect 12292 6500 12348 6556
rect 12348 6500 12352 6556
rect 12288 6496 12352 6500
rect 19445 6556 19509 6560
rect 19445 6500 19449 6556
rect 19449 6500 19505 6556
rect 19505 6500 19509 6556
rect 19445 6496 19509 6500
rect 19525 6556 19589 6560
rect 19525 6500 19529 6556
rect 19529 6500 19585 6556
rect 19585 6500 19589 6556
rect 19525 6496 19589 6500
rect 19605 6556 19669 6560
rect 19605 6500 19609 6556
rect 19609 6500 19665 6556
rect 19665 6500 19669 6556
rect 19605 6496 19669 6500
rect 19685 6556 19749 6560
rect 19685 6500 19689 6556
rect 19689 6500 19745 6556
rect 19745 6500 19749 6556
rect 19685 6496 19749 6500
rect 13860 6292 13924 6356
rect 6500 6156 6564 6220
rect 10180 6156 10244 6220
rect 8349 6012 8413 6016
rect 8349 5956 8353 6012
rect 8353 5956 8409 6012
rect 8409 5956 8413 6012
rect 8349 5952 8413 5956
rect 8429 6012 8493 6016
rect 8429 5956 8433 6012
rect 8433 5956 8489 6012
rect 8489 5956 8493 6012
rect 8429 5952 8493 5956
rect 8509 6012 8573 6016
rect 8509 5956 8513 6012
rect 8513 5956 8569 6012
rect 8569 5956 8573 6012
rect 8509 5952 8573 5956
rect 8589 6012 8653 6016
rect 8589 5956 8593 6012
rect 8593 5956 8649 6012
rect 8649 5956 8653 6012
rect 8589 5952 8653 5956
rect 6684 5884 6748 5948
rect 9260 5944 9324 5948
rect 9260 5888 9310 5944
rect 9310 5888 9324 5944
rect 9260 5884 9324 5888
rect 15746 6012 15810 6016
rect 15746 5956 15750 6012
rect 15750 5956 15806 6012
rect 15806 5956 15810 6012
rect 15746 5952 15810 5956
rect 15826 6012 15890 6016
rect 15826 5956 15830 6012
rect 15830 5956 15886 6012
rect 15886 5956 15890 6012
rect 15826 5952 15890 5956
rect 15906 6012 15970 6016
rect 15906 5956 15910 6012
rect 15910 5956 15966 6012
rect 15966 5956 15970 6012
rect 15906 5952 15970 5956
rect 15986 6012 16050 6016
rect 15986 5956 15990 6012
rect 15990 5956 16046 6012
rect 16046 5956 16050 6012
rect 15986 5952 16050 5956
rect 13676 5808 13740 5812
rect 13676 5752 13690 5808
rect 13690 5752 13740 5808
rect 13676 5748 13740 5752
rect 11836 5612 11900 5676
rect 4650 5468 4714 5472
rect 4650 5412 4654 5468
rect 4654 5412 4710 5468
rect 4710 5412 4714 5468
rect 4650 5408 4714 5412
rect 4730 5468 4794 5472
rect 4730 5412 4734 5468
rect 4734 5412 4790 5468
rect 4790 5412 4794 5468
rect 4730 5408 4794 5412
rect 4810 5468 4874 5472
rect 4810 5412 4814 5468
rect 4814 5412 4870 5468
rect 4870 5412 4874 5468
rect 4810 5408 4874 5412
rect 4890 5468 4954 5472
rect 4890 5412 4894 5468
rect 4894 5412 4950 5468
rect 4950 5412 4954 5468
rect 4890 5408 4954 5412
rect 12048 5468 12112 5472
rect 12048 5412 12052 5468
rect 12052 5412 12108 5468
rect 12108 5412 12112 5468
rect 12048 5408 12112 5412
rect 12128 5468 12192 5472
rect 12128 5412 12132 5468
rect 12132 5412 12188 5468
rect 12188 5412 12192 5468
rect 12128 5408 12192 5412
rect 12208 5468 12272 5472
rect 12208 5412 12212 5468
rect 12212 5412 12268 5468
rect 12268 5412 12272 5468
rect 12208 5408 12272 5412
rect 12288 5468 12352 5472
rect 12288 5412 12292 5468
rect 12292 5412 12348 5468
rect 12348 5412 12352 5468
rect 12288 5408 12352 5412
rect 19445 5468 19509 5472
rect 19445 5412 19449 5468
rect 19449 5412 19505 5468
rect 19505 5412 19509 5468
rect 19445 5408 19509 5412
rect 19525 5468 19589 5472
rect 19525 5412 19529 5468
rect 19529 5412 19585 5468
rect 19585 5412 19589 5468
rect 19525 5408 19589 5412
rect 19605 5468 19669 5472
rect 19605 5412 19609 5468
rect 19609 5412 19665 5468
rect 19665 5412 19669 5468
rect 19605 5408 19669 5412
rect 19685 5468 19749 5472
rect 19685 5412 19689 5468
rect 19689 5412 19745 5468
rect 19745 5412 19749 5468
rect 19685 5408 19749 5412
rect 8349 4924 8413 4928
rect 8349 4868 8353 4924
rect 8353 4868 8409 4924
rect 8409 4868 8413 4924
rect 8349 4864 8413 4868
rect 8429 4924 8493 4928
rect 8429 4868 8433 4924
rect 8433 4868 8489 4924
rect 8489 4868 8493 4924
rect 8429 4864 8493 4868
rect 8509 4924 8573 4928
rect 8509 4868 8513 4924
rect 8513 4868 8569 4924
rect 8569 4868 8573 4924
rect 8509 4864 8573 4868
rect 8589 4924 8653 4928
rect 8589 4868 8593 4924
rect 8593 4868 8649 4924
rect 8649 4868 8653 4924
rect 8589 4864 8653 4868
rect 15746 4924 15810 4928
rect 15746 4868 15750 4924
rect 15750 4868 15806 4924
rect 15806 4868 15810 4924
rect 15746 4864 15810 4868
rect 15826 4924 15890 4928
rect 15826 4868 15830 4924
rect 15830 4868 15886 4924
rect 15886 4868 15890 4924
rect 15826 4864 15890 4868
rect 15906 4924 15970 4928
rect 15906 4868 15910 4924
rect 15910 4868 15966 4924
rect 15966 4868 15970 4924
rect 15906 4864 15970 4868
rect 15986 4924 16050 4928
rect 15986 4868 15990 4924
rect 15990 4868 16046 4924
rect 16046 4868 16050 4924
rect 15986 4864 16050 4868
rect 4650 4380 4714 4384
rect 4650 4324 4654 4380
rect 4654 4324 4710 4380
rect 4710 4324 4714 4380
rect 4650 4320 4714 4324
rect 4730 4380 4794 4384
rect 4730 4324 4734 4380
rect 4734 4324 4790 4380
rect 4790 4324 4794 4380
rect 4730 4320 4794 4324
rect 4810 4380 4874 4384
rect 4810 4324 4814 4380
rect 4814 4324 4870 4380
rect 4870 4324 4874 4380
rect 4810 4320 4874 4324
rect 4890 4380 4954 4384
rect 4890 4324 4894 4380
rect 4894 4324 4950 4380
rect 4950 4324 4954 4380
rect 4890 4320 4954 4324
rect 12048 4380 12112 4384
rect 12048 4324 12052 4380
rect 12052 4324 12108 4380
rect 12108 4324 12112 4380
rect 12048 4320 12112 4324
rect 12128 4380 12192 4384
rect 12128 4324 12132 4380
rect 12132 4324 12188 4380
rect 12188 4324 12192 4380
rect 12128 4320 12192 4324
rect 12208 4380 12272 4384
rect 12208 4324 12212 4380
rect 12212 4324 12268 4380
rect 12268 4324 12272 4380
rect 12208 4320 12272 4324
rect 12288 4380 12352 4384
rect 12288 4324 12292 4380
rect 12292 4324 12348 4380
rect 12348 4324 12352 4380
rect 12288 4320 12352 4324
rect 19445 4380 19509 4384
rect 19445 4324 19449 4380
rect 19449 4324 19505 4380
rect 19505 4324 19509 4380
rect 19445 4320 19509 4324
rect 19525 4380 19589 4384
rect 19525 4324 19529 4380
rect 19529 4324 19585 4380
rect 19585 4324 19589 4380
rect 19525 4320 19589 4324
rect 19605 4380 19669 4384
rect 19605 4324 19609 4380
rect 19609 4324 19665 4380
rect 19665 4324 19669 4380
rect 19605 4320 19669 4324
rect 19685 4380 19749 4384
rect 19685 4324 19689 4380
rect 19689 4324 19745 4380
rect 19745 4324 19749 4380
rect 19685 4320 19749 4324
rect 11836 4176 11900 4180
rect 11836 4120 11886 4176
rect 11886 4120 11900 4176
rect 11836 4116 11900 4120
rect 14044 4040 14108 4044
rect 14044 3984 14058 4040
rect 14058 3984 14108 4040
rect 14044 3980 14108 3984
rect 14412 3844 14476 3908
rect 8349 3836 8413 3840
rect 8349 3780 8353 3836
rect 8353 3780 8409 3836
rect 8409 3780 8413 3836
rect 8349 3776 8413 3780
rect 8429 3836 8493 3840
rect 8429 3780 8433 3836
rect 8433 3780 8489 3836
rect 8489 3780 8493 3836
rect 8429 3776 8493 3780
rect 8509 3836 8573 3840
rect 8509 3780 8513 3836
rect 8513 3780 8569 3836
rect 8569 3780 8573 3836
rect 8509 3776 8573 3780
rect 8589 3836 8653 3840
rect 8589 3780 8593 3836
rect 8593 3780 8649 3836
rect 8649 3780 8653 3836
rect 8589 3776 8653 3780
rect 15746 3836 15810 3840
rect 15746 3780 15750 3836
rect 15750 3780 15806 3836
rect 15806 3780 15810 3836
rect 15746 3776 15810 3780
rect 15826 3836 15890 3840
rect 15826 3780 15830 3836
rect 15830 3780 15886 3836
rect 15886 3780 15890 3836
rect 15826 3776 15890 3780
rect 15906 3836 15970 3840
rect 15906 3780 15910 3836
rect 15910 3780 15966 3836
rect 15966 3780 15970 3836
rect 15906 3776 15970 3780
rect 15986 3836 16050 3840
rect 15986 3780 15990 3836
rect 15990 3780 16046 3836
rect 16046 3780 16050 3836
rect 15986 3776 16050 3780
rect 17540 3300 17604 3364
rect 4650 3292 4714 3296
rect 4650 3236 4654 3292
rect 4654 3236 4710 3292
rect 4710 3236 4714 3292
rect 4650 3232 4714 3236
rect 4730 3292 4794 3296
rect 4730 3236 4734 3292
rect 4734 3236 4790 3292
rect 4790 3236 4794 3292
rect 4730 3232 4794 3236
rect 4810 3292 4874 3296
rect 4810 3236 4814 3292
rect 4814 3236 4870 3292
rect 4870 3236 4874 3292
rect 4810 3232 4874 3236
rect 4890 3292 4954 3296
rect 4890 3236 4894 3292
rect 4894 3236 4950 3292
rect 4950 3236 4954 3292
rect 4890 3232 4954 3236
rect 12048 3292 12112 3296
rect 12048 3236 12052 3292
rect 12052 3236 12108 3292
rect 12108 3236 12112 3292
rect 12048 3232 12112 3236
rect 12128 3292 12192 3296
rect 12128 3236 12132 3292
rect 12132 3236 12188 3292
rect 12188 3236 12192 3292
rect 12128 3232 12192 3236
rect 12208 3292 12272 3296
rect 12208 3236 12212 3292
rect 12212 3236 12268 3292
rect 12268 3236 12272 3292
rect 12208 3232 12272 3236
rect 12288 3292 12352 3296
rect 12288 3236 12292 3292
rect 12292 3236 12348 3292
rect 12348 3236 12352 3292
rect 12288 3232 12352 3236
rect 19445 3292 19509 3296
rect 19445 3236 19449 3292
rect 19449 3236 19505 3292
rect 19505 3236 19509 3292
rect 19445 3232 19509 3236
rect 19525 3292 19589 3296
rect 19525 3236 19529 3292
rect 19529 3236 19585 3292
rect 19585 3236 19589 3292
rect 19525 3232 19589 3236
rect 19605 3292 19669 3296
rect 19605 3236 19609 3292
rect 19609 3236 19665 3292
rect 19665 3236 19669 3292
rect 19605 3232 19669 3236
rect 19685 3292 19749 3296
rect 19685 3236 19689 3292
rect 19689 3236 19745 3292
rect 19745 3236 19749 3292
rect 19685 3232 19749 3236
rect 14228 3164 14292 3228
rect 8349 2748 8413 2752
rect 8349 2692 8353 2748
rect 8353 2692 8409 2748
rect 8409 2692 8413 2748
rect 8349 2688 8413 2692
rect 8429 2748 8493 2752
rect 8429 2692 8433 2748
rect 8433 2692 8489 2748
rect 8489 2692 8493 2748
rect 8429 2688 8493 2692
rect 8509 2748 8573 2752
rect 8509 2692 8513 2748
rect 8513 2692 8569 2748
rect 8569 2692 8573 2748
rect 8509 2688 8573 2692
rect 8589 2748 8653 2752
rect 8589 2692 8593 2748
rect 8593 2692 8649 2748
rect 8649 2692 8653 2748
rect 8589 2688 8653 2692
rect 15746 2748 15810 2752
rect 15746 2692 15750 2748
rect 15750 2692 15806 2748
rect 15806 2692 15810 2748
rect 15746 2688 15810 2692
rect 15826 2748 15890 2752
rect 15826 2692 15830 2748
rect 15830 2692 15886 2748
rect 15886 2692 15890 2748
rect 15826 2688 15890 2692
rect 15906 2748 15970 2752
rect 15906 2692 15910 2748
rect 15910 2692 15966 2748
rect 15966 2692 15970 2748
rect 15906 2688 15970 2692
rect 15986 2748 16050 2752
rect 15986 2692 15990 2748
rect 15990 2692 16046 2748
rect 16046 2692 16050 2748
rect 15986 2688 16050 2692
rect 8892 2484 8956 2548
rect 4650 2204 4714 2208
rect 4650 2148 4654 2204
rect 4654 2148 4710 2204
rect 4710 2148 4714 2204
rect 4650 2144 4714 2148
rect 4730 2204 4794 2208
rect 4730 2148 4734 2204
rect 4734 2148 4790 2204
rect 4790 2148 4794 2204
rect 4730 2144 4794 2148
rect 4810 2204 4874 2208
rect 4810 2148 4814 2204
rect 4814 2148 4870 2204
rect 4870 2148 4874 2204
rect 4810 2144 4874 2148
rect 4890 2204 4954 2208
rect 4890 2148 4894 2204
rect 4894 2148 4950 2204
rect 4950 2148 4954 2204
rect 4890 2144 4954 2148
rect 12048 2204 12112 2208
rect 12048 2148 12052 2204
rect 12052 2148 12108 2204
rect 12108 2148 12112 2204
rect 12048 2144 12112 2148
rect 12128 2204 12192 2208
rect 12128 2148 12132 2204
rect 12132 2148 12188 2204
rect 12188 2148 12192 2204
rect 12128 2144 12192 2148
rect 12208 2204 12272 2208
rect 12208 2148 12212 2204
rect 12212 2148 12268 2204
rect 12268 2148 12272 2204
rect 12208 2144 12272 2148
rect 12288 2204 12352 2208
rect 12288 2148 12292 2204
rect 12292 2148 12348 2204
rect 12348 2148 12352 2204
rect 12288 2144 12352 2148
rect 19445 2204 19509 2208
rect 19445 2148 19449 2204
rect 19449 2148 19505 2204
rect 19505 2148 19509 2204
rect 19445 2144 19509 2148
rect 19525 2204 19589 2208
rect 19525 2148 19529 2204
rect 19529 2148 19585 2204
rect 19585 2148 19589 2204
rect 19525 2144 19589 2148
rect 19605 2204 19669 2208
rect 19605 2148 19609 2204
rect 19609 2148 19665 2204
rect 19665 2148 19669 2204
rect 19605 2144 19669 2148
rect 19685 2204 19749 2208
rect 19685 2148 19689 2204
rect 19689 2148 19745 2204
rect 19745 2148 19749 2204
rect 19685 2144 19749 2148
<< metal4 >>
rect 4642 21792 4963 21808
rect 4642 21728 4650 21792
rect 4714 21728 4730 21792
rect 4794 21728 4810 21792
rect 4874 21728 4890 21792
rect 4954 21728 4963 21792
rect 4642 20704 4963 21728
rect 4642 20640 4650 20704
rect 4714 20640 4730 20704
rect 4794 20640 4810 20704
rect 4874 20640 4890 20704
rect 4954 20640 4963 20704
rect 4642 19616 4963 20640
rect 4642 19552 4650 19616
rect 4714 19552 4730 19616
rect 4794 19552 4810 19616
rect 4874 19552 4890 19616
rect 4954 19552 4963 19616
rect 4642 18528 4963 19552
rect 8341 21248 8661 21808
rect 8341 21184 8349 21248
rect 8413 21184 8429 21248
rect 8493 21184 8509 21248
rect 8573 21184 8589 21248
rect 8653 21184 8661 21248
rect 8341 20160 8661 21184
rect 8341 20096 8349 20160
rect 8413 20096 8429 20160
rect 8493 20096 8509 20160
rect 8573 20096 8589 20160
rect 8653 20096 8661 20160
rect 6683 19548 6749 19549
rect 6683 19484 6684 19548
rect 6748 19484 6749 19548
rect 6683 19483 6749 19484
rect 4642 18464 4650 18528
rect 4714 18464 4730 18528
rect 4794 18464 4810 18528
rect 4874 18464 4890 18528
rect 4954 18464 4963 18528
rect 4475 18052 4541 18053
rect 4475 17988 4476 18052
rect 4540 17988 4541 18052
rect 4475 17987 4541 17988
rect 4478 12749 4538 17987
rect 4642 17440 4963 18464
rect 4642 17376 4650 17440
rect 4714 17376 4730 17440
rect 4794 17376 4810 17440
rect 4874 17376 4890 17440
rect 4954 17376 4963 17440
rect 4642 16352 4963 17376
rect 4642 16288 4650 16352
rect 4714 16288 4730 16352
rect 4794 16288 4810 16352
rect 4874 16288 4890 16352
rect 4954 16288 4963 16352
rect 4642 15264 4963 16288
rect 5395 15740 5461 15741
rect 5395 15676 5396 15740
rect 5460 15676 5461 15740
rect 5395 15675 5461 15676
rect 4642 15200 4650 15264
rect 4714 15200 4730 15264
rect 4794 15200 4810 15264
rect 4874 15200 4890 15264
rect 4954 15200 4963 15264
rect 4642 14176 4963 15200
rect 4642 14112 4650 14176
rect 4714 14112 4730 14176
rect 4794 14112 4810 14176
rect 4874 14112 4890 14176
rect 4954 14112 4963 14176
rect 4642 13088 4963 14112
rect 4642 13024 4650 13088
rect 4714 13024 4730 13088
rect 4794 13024 4810 13088
rect 4874 13024 4890 13088
rect 4954 13024 4963 13088
rect 4475 12748 4541 12749
rect 4475 12684 4476 12748
rect 4540 12684 4541 12748
rect 4475 12683 4541 12684
rect 4642 12000 4963 13024
rect 4642 11936 4650 12000
rect 4714 11936 4730 12000
rect 4794 11936 4810 12000
rect 4874 11936 4890 12000
rect 4954 11936 4963 12000
rect 4642 10912 4963 11936
rect 5027 11116 5093 11117
rect 5027 11052 5028 11116
rect 5092 11052 5093 11116
rect 5027 11051 5093 11052
rect 4642 10848 4650 10912
rect 4714 10848 4730 10912
rect 4794 10848 4810 10912
rect 4874 10848 4890 10912
rect 4954 10848 4963 10912
rect 4642 9824 4963 10848
rect 4642 9760 4650 9824
rect 4714 9760 4730 9824
rect 4794 9760 4810 9824
rect 4874 9760 4890 9824
rect 4954 9760 4963 9824
rect 4642 8736 4963 9760
rect 5030 9485 5090 11051
rect 5027 9484 5093 9485
rect 5027 9420 5028 9484
rect 5092 9420 5093 9484
rect 5027 9419 5093 9420
rect 5398 8805 5458 15675
rect 6499 13156 6565 13157
rect 6499 13092 6500 13156
rect 6564 13092 6565 13156
rect 6499 13091 6565 13092
rect 5763 12748 5829 12749
rect 5763 12684 5764 12748
rect 5828 12684 5829 12748
rect 5763 12683 5829 12684
rect 5766 12205 5826 12683
rect 6315 12476 6381 12477
rect 6315 12412 6316 12476
rect 6380 12412 6381 12476
rect 6315 12411 6381 12412
rect 5763 12204 5829 12205
rect 5763 12140 5764 12204
rect 5828 12140 5829 12204
rect 5763 12139 5829 12140
rect 6318 12069 6378 12411
rect 6315 12068 6381 12069
rect 6315 12004 6316 12068
rect 6380 12004 6381 12068
rect 6315 12003 6381 12004
rect 5763 10844 5829 10845
rect 5763 10780 5764 10844
rect 5828 10780 5829 10844
rect 5763 10779 5829 10780
rect 5766 10301 5826 10779
rect 5763 10300 5829 10301
rect 5763 10236 5764 10300
rect 5828 10236 5829 10300
rect 5763 10235 5829 10236
rect 5395 8804 5461 8805
rect 5395 8740 5396 8804
rect 5460 8740 5461 8804
rect 5395 8739 5461 8740
rect 4642 8672 4650 8736
rect 4714 8672 4730 8736
rect 4794 8672 4810 8736
rect 4874 8672 4890 8736
rect 4954 8672 4963 8736
rect 4642 7648 4963 8672
rect 5766 7989 5826 10235
rect 5763 7988 5829 7989
rect 5763 7924 5764 7988
rect 5828 7924 5829 7988
rect 5763 7923 5829 7924
rect 4642 7584 4650 7648
rect 4714 7584 4730 7648
rect 4794 7584 4810 7648
rect 4874 7584 4890 7648
rect 4954 7584 4963 7648
rect 4642 6560 4963 7584
rect 4642 6496 4650 6560
rect 4714 6496 4730 6560
rect 4794 6496 4810 6560
rect 4874 6496 4890 6560
rect 4954 6496 4963 6560
rect 4642 5472 4963 6496
rect 6502 6221 6562 13091
rect 6499 6220 6565 6221
rect 6499 6156 6500 6220
rect 6564 6156 6565 6220
rect 6499 6155 6565 6156
rect 6686 5949 6746 19483
rect 8341 19072 8661 20096
rect 12040 21792 12360 21808
rect 12040 21728 12048 21792
rect 12112 21728 12128 21792
rect 12192 21728 12208 21792
rect 12272 21728 12288 21792
rect 12352 21728 12360 21792
rect 12040 20704 12360 21728
rect 15738 21248 16058 21808
rect 15738 21184 15746 21248
rect 15810 21184 15826 21248
rect 15890 21184 15906 21248
rect 15970 21184 15986 21248
rect 16050 21184 16058 21248
rect 14227 20908 14293 20909
rect 14227 20844 14228 20908
rect 14292 20844 14293 20908
rect 14227 20843 14293 20844
rect 12040 20640 12048 20704
rect 12112 20640 12128 20704
rect 12192 20640 12208 20704
rect 12272 20640 12288 20704
rect 12352 20640 12360 20704
rect 12040 19616 12360 20640
rect 12040 19552 12048 19616
rect 12112 19552 12128 19616
rect 12192 19552 12208 19616
rect 12272 19552 12288 19616
rect 12352 19552 12360 19616
rect 11651 19140 11717 19141
rect 11651 19076 11652 19140
rect 11716 19076 11717 19140
rect 11651 19075 11717 19076
rect 8341 19008 8349 19072
rect 8413 19008 8429 19072
rect 8493 19008 8509 19072
rect 8573 19008 8589 19072
rect 8653 19008 8661 19072
rect 8341 17984 8661 19008
rect 8341 17920 8349 17984
rect 8413 17920 8429 17984
rect 8493 17920 8509 17984
rect 8573 17920 8589 17984
rect 8653 17920 8661 17984
rect 7971 17508 8037 17509
rect 7971 17444 7972 17508
rect 8036 17444 8037 17508
rect 7971 17443 8037 17444
rect 7051 14924 7117 14925
rect 7051 14860 7052 14924
rect 7116 14860 7117 14924
rect 7051 14859 7117 14860
rect 6867 10028 6933 10029
rect 6867 9964 6868 10028
rect 6932 9964 6933 10028
rect 6867 9963 6933 9964
rect 6870 8941 6930 9963
rect 7054 9757 7114 14859
rect 7235 10708 7301 10709
rect 7235 10644 7236 10708
rect 7300 10644 7301 10708
rect 7235 10643 7301 10644
rect 7051 9756 7117 9757
rect 7051 9692 7052 9756
rect 7116 9692 7117 9756
rect 7051 9691 7117 9692
rect 6867 8940 6933 8941
rect 6867 8876 6868 8940
rect 6932 8876 6933 8940
rect 6867 8875 6933 8876
rect 7238 8125 7298 10643
rect 7419 10164 7485 10165
rect 7419 10100 7420 10164
rect 7484 10100 7485 10164
rect 7419 10099 7485 10100
rect 7235 8124 7301 8125
rect 7235 8060 7236 8124
rect 7300 8060 7301 8124
rect 7235 8059 7301 8060
rect 7422 7717 7482 10099
rect 7603 9892 7669 9893
rect 7603 9828 7604 9892
rect 7668 9828 7669 9892
rect 7603 9827 7669 9828
rect 7606 8669 7666 9827
rect 7787 9756 7853 9757
rect 7787 9692 7788 9756
rect 7852 9692 7853 9756
rect 7787 9691 7853 9692
rect 7603 8668 7669 8669
rect 7603 8604 7604 8668
rect 7668 8604 7669 8668
rect 7603 8603 7669 8604
rect 7790 7717 7850 9691
rect 7419 7716 7485 7717
rect 7419 7652 7420 7716
rect 7484 7652 7485 7716
rect 7419 7651 7485 7652
rect 7787 7716 7853 7717
rect 7787 7652 7788 7716
rect 7852 7652 7853 7716
rect 7787 7651 7853 7652
rect 7974 6901 8034 17443
rect 8341 16896 8661 17920
rect 8891 17236 8957 17237
rect 8891 17172 8892 17236
rect 8956 17172 8957 17236
rect 8891 17171 8957 17172
rect 8341 16832 8349 16896
rect 8413 16832 8429 16896
rect 8493 16832 8509 16896
rect 8573 16832 8589 16896
rect 8653 16832 8661 16896
rect 8341 15808 8661 16832
rect 8341 15744 8349 15808
rect 8413 15744 8429 15808
rect 8493 15744 8509 15808
rect 8573 15744 8589 15808
rect 8653 15744 8661 15808
rect 8341 14720 8661 15744
rect 8341 14656 8349 14720
rect 8413 14656 8429 14720
rect 8493 14656 8509 14720
rect 8573 14656 8589 14720
rect 8653 14656 8661 14720
rect 8341 13632 8661 14656
rect 8341 13568 8349 13632
rect 8413 13568 8429 13632
rect 8493 13568 8509 13632
rect 8573 13568 8589 13632
rect 8653 13568 8661 13632
rect 8341 12544 8661 13568
rect 8341 12480 8349 12544
rect 8413 12480 8429 12544
rect 8493 12480 8509 12544
rect 8573 12480 8589 12544
rect 8653 12480 8661 12544
rect 8341 11456 8661 12480
rect 8341 11392 8349 11456
rect 8413 11392 8429 11456
rect 8493 11392 8509 11456
rect 8573 11392 8589 11456
rect 8653 11392 8661 11456
rect 8155 11252 8221 11253
rect 8155 11188 8156 11252
rect 8220 11188 8221 11252
rect 8155 11187 8221 11188
rect 8158 8533 8218 11187
rect 8341 10368 8661 11392
rect 8341 10304 8349 10368
rect 8413 10304 8429 10368
rect 8493 10304 8509 10368
rect 8573 10304 8589 10368
rect 8653 10304 8661 10368
rect 8341 9280 8661 10304
rect 8894 10165 8954 17171
rect 9995 14788 10061 14789
rect 9995 14724 9996 14788
rect 10060 14724 10061 14788
rect 9995 14723 10061 14724
rect 9627 13972 9693 13973
rect 9627 13908 9628 13972
rect 9692 13908 9693 13972
rect 9627 13907 9693 13908
rect 9443 10572 9509 10573
rect 9443 10508 9444 10572
rect 9508 10508 9509 10572
rect 9443 10507 9509 10508
rect 8891 10164 8957 10165
rect 8891 10100 8892 10164
rect 8956 10100 8957 10164
rect 8891 10099 8957 10100
rect 8891 9892 8957 9893
rect 8891 9828 8892 9892
rect 8956 9828 8957 9892
rect 8891 9827 8957 9828
rect 8341 9216 8349 9280
rect 8413 9216 8429 9280
rect 8493 9216 8509 9280
rect 8573 9216 8589 9280
rect 8653 9216 8661 9280
rect 8155 8532 8221 8533
rect 8155 8468 8156 8532
rect 8220 8468 8221 8532
rect 8155 8467 8221 8468
rect 8341 8192 8661 9216
rect 8894 9210 8954 9827
rect 8756 9150 8954 9210
rect 8756 8530 8816 9150
rect 8756 8470 9138 8530
rect 8341 8128 8349 8192
rect 8413 8128 8429 8192
rect 8493 8128 8509 8192
rect 8573 8128 8589 8192
rect 8653 8128 8661 8192
rect 8341 7104 8661 8128
rect 8891 8124 8957 8125
rect 8891 8060 8892 8124
rect 8956 8060 8957 8124
rect 8891 8059 8957 8060
rect 8341 7040 8349 7104
rect 8413 7040 8429 7104
rect 8493 7040 8509 7104
rect 8573 7040 8589 7104
rect 8653 7040 8661 7104
rect 7971 6900 8037 6901
rect 7971 6836 7972 6900
rect 8036 6836 8037 6900
rect 7971 6835 8037 6836
rect 8341 6016 8661 7040
rect 8341 5952 8349 6016
rect 8413 5952 8429 6016
rect 8493 5952 8509 6016
rect 8573 5952 8589 6016
rect 8653 5952 8661 6016
rect 6683 5948 6749 5949
rect 6683 5884 6684 5948
rect 6748 5884 6749 5948
rect 6683 5883 6749 5884
rect 4642 5408 4650 5472
rect 4714 5408 4730 5472
rect 4794 5408 4810 5472
rect 4874 5408 4890 5472
rect 4954 5408 4963 5472
rect 4642 4384 4963 5408
rect 4642 4320 4650 4384
rect 4714 4320 4730 4384
rect 4794 4320 4810 4384
rect 4874 4320 4890 4384
rect 4954 4320 4963 4384
rect 4642 3296 4963 4320
rect 4642 3232 4650 3296
rect 4714 3232 4730 3296
rect 4794 3232 4810 3296
rect 4874 3232 4890 3296
rect 4954 3232 4963 3296
rect 4642 2208 4963 3232
rect 4642 2144 4650 2208
rect 4714 2144 4730 2208
rect 4794 2144 4810 2208
rect 4874 2144 4890 2208
rect 4954 2144 4963 2208
rect 4642 2128 4963 2144
rect 8341 4928 8661 5952
rect 8341 4864 8349 4928
rect 8413 4864 8429 4928
rect 8493 4864 8509 4928
rect 8573 4864 8589 4928
rect 8653 4864 8661 4928
rect 8341 3840 8661 4864
rect 8341 3776 8349 3840
rect 8413 3776 8429 3840
rect 8493 3776 8509 3840
rect 8573 3776 8589 3840
rect 8653 3776 8661 3840
rect 8341 2752 8661 3776
rect 8341 2688 8349 2752
rect 8413 2688 8429 2752
rect 8493 2688 8509 2752
rect 8573 2688 8589 2752
rect 8653 2688 8661 2752
rect 8341 2128 8661 2688
rect 8894 2549 8954 8059
rect 9078 6629 9138 8470
rect 9259 8260 9325 8261
rect 9259 8196 9260 8260
rect 9324 8196 9325 8260
rect 9259 8195 9325 8196
rect 9075 6628 9141 6629
rect 9075 6564 9076 6628
rect 9140 6564 9141 6628
rect 9075 6563 9141 6564
rect 9262 5949 9322 8195
rect 9446 6629 9506 10507
rect 9630 9077 9690 13907
rect 9811 10436 9877 10437
rect 9811 10372 9812 10436
rect 9876 10372 9877 10436
rect 9811 10371 9877 10372
rect 9627 9076 9693 9077
rect 9627 9012 9628 9076
rect 9692 9012 9693 9076
rect 9627 9011 9693 9012
rect 9814 7173 9874 10371
rect 9998 8397 10058 14723
rect 10363 13428 10429 13429
rect 10363 13364 10364 13428
rect 10428 13364 10429 13428
rect 10363 13363 10429 13364
rect 10179 9756 10245 9757
rect 10179 9692 10180 9756
rect 10244 9692 10245 9756
rect 10179 9691 10245 9692
rect 9995 8396 10061 8397
rect 9995 8332 9996 8396
rect 10060 8332 10061 8396
rect 9995 8331 10061 8332
rect 9995 8124 10061 8125
rect 9995 8060 9996 8124
rect 10060 8060 10061 8124
rect 9995 8059 10061 8060
rect 9998 7173 10058 8059
rect 9811 7172 9877 7173
rect 9811 7108 9812 7172
rect 9876 7108 9877 7172
rect 9811 7107 9877 7108
rect 9995 7172 10061 7173
rect 9995 7108 9996 7172
rect 10060 7108 10061 7172
rect 9995 7107 10061 7108
rect 9443 6628 9509 6629
rect 9443 6564 9444 6628
rect 9508 6564 9509 6628
rect 9443 6563 9509 6564
rect 10182 6221 10242 9691
rect 10366 8533 10426 13363
rect 11654 12613 11714 19075
rect 12040 18528 12360 19552
rect 12040 18464 12048 18528
rect 12112 18464 12128 18528
rect 12192 18464 12208 18528
rect 12272 18464 12288 18528
rect 12352 18464 12360 18528
rect 12040 17440 12360 18464
rect 14043 18188 14109 18189
rect 14043 18124 14044 18188
rect 14108 18124 14109 18188
rect 14043 18123 14109 18124
rect 12040 17376 12048 17440
rect 12112 17376 12128 17440
rect 12192 17376 12208 17440
rect 12272 17376 12288 17440
rect 12352 17376 12360 17440
rect 12040 16352 12360 17376
rect 12040 16288 12048 16352
rect 12112 16288 12128 16352
rect 12192 16288 12208 16352
rect 12272 16288 12288 16352
rect 12352 16288 12360 16352
rect 11835 16148 11901 16149
rect 11835 16084 11836 16148
rect 11900 16084 11901 16148
rect 11835 16083 11901 16084
rect 11651 12612 11717 12613
rect 11651 12548 11652 12612
rect 11716 12548 11717 12612
rect 11651 12547 11717 12548
rect 11838 10709 11898 16083
rect 12040 15264 12360 16288
rect 13675 15876 13741 15877
rect 13675 15812 13676 15876
rect 13740 15812 13741 15876
rect 13675 15811 13741 15812
rect 12040 15200 12048 15264
rect 12112 15200 12128 15264
rect 12192 15200 12208 15264
rect 12272 15200 12288 15264
rect 12352 15200 12360 15264
rect 12040 14176 12360 15200
rect 12040 14112 12048 14176
rect 12112 14112 12128 14176
rect 12192 14112 12208 14176
rect 12272 14112 12288 14176
rect 12352 14112 12360 14176
rect 12040 13088 12360 14112
rect 12571 14108 12637 14109
rect 12571 14044 12572 14108
rect 12636 14044 12637 14108
rect 12571 14043 12637 14044
rect 12040 13024 12048 13088
rect 12112 13024 12128 13088
rect 12192 13024 12208 13088
rect 12272 13024 12288 13088
rect 12352 13024 12360 13088
rect 12040 12000 12360 13024
rect 12040 11936 12048 12000
rect 12112 11936 12128 12000
rect 12192 11936 12208 12000
rect 12272 11936 12288 12000
rect 12352 11936 12360 12000
rect 12040 10912 12360 11936
rect 12040 10848 12048 10912
rect 12112 10848 12128 10912
rect 12192 10848 12208 10912
rect 12272 10848 12288 10912
rect 12352 10848 12360 10912
rect 11835 10708 11901 10709
rect 11835 10644 11836 10708
rect 11900 10644 11901 10708
rect 11835 10643 11901 10644
rect 12040 9824 12360 10848
rect 12040 9760 12048 9824
rect 12112 9760 12128 9824
rect 12192 9760 12208 9824
rect 12272 9760 12288 9824
rect 12352 9760 12360 9824
rect 11835 9348 11901 9349
rect 11835 9284 11836 9348
rect 11900 9284 11901 9348
rect 11835 9283 11901 9284
rect 10363 8532 10429 8533
rect 10363 8468 10364 8532
rect 10428 8468 10429 8532
rect 10363 8467 10429 8468
rect 10179 6220 10245 6221
rect 10179 6156 10180 6220
rect 10244 6156 10245 6220
rect 10179 6155 10245 6156
rect 9259 5948 9325 5949
rect 9259 5884 9260 5948
rect 9324 5884 9325 5948
rect 9259 5883 9325 5884
rect 11838 5677 11898 9283
rect 12040 8736 12360 9760
rect 12574 9349 12634 14043
rect 12755 12612 12821 12613
rect 12755 12548 12756 12612
rect 12820 12548 12821 12612
rect 12755 12547 12821 12548
rect 12758 12205 12818 12547
rect 12939 12476 13005 12477
rect 12939 12412 12940 12476
rect 13004 12412 13005 12476
rect 12939 12411 13005 12412
rect 12755 12204 12821 12205
rect 12755 12140 12756 12204
rect 12820 12140 12821 12204
rect 12755 12139 12821 12140
rect 12942 10573 13002 12411
rect 13307 12340 13373 12341
rect 13307 12276 13308 12340
rect 13372 12276 13373 12340
rect 13307 12275 13373 12276
rect 12939 10572 13005 10573
rect 12939 10508 12940 10572
rect 13004 10508 13005 10572
rect 12939 10507 13005 10508
rect 12571 9348 12637 9349
rect 12571 9284 12572 9348
rect 12636 9284 12637 9348
rect 12571 9283 12637 9284
rect 12040 8672 12048 8736
rect 12112 8672 12128 8736
rect 12192 8672 12208 8736
rect 12272 8672 12288 8736
rect 12352 8672 12360 8736
rect 12040 7648 12360 8672
rect 12942 8397 13002 10507
rect 13310 8397 13370 12275
rect 13678 10301 13738 15811
rect 13859 15332 13925 15333
rect 13859 15268 13860 15332
rect 13924 15268 13925 15332
rect 13859 15267 13925 15268
rect 13675 10300 13741 10301
rect 13675 10236 13676 10300
rect 13740 10236 13741 10300
rect 13675 10235 13741 10236
rect 12939 8396 13005 8397
rect 12939 8332 12940 8396
rect 13004 8332 13005 8396
rect 12939 8331 13005 8332
rect 13307 8396 13373 8397
rect 13307 8332 13308 8396
rect 13372 8332 13373 8396
rect 13307 8331 13373 8332
rect 12040 7584 12048 7648
rect 12112 7584 12128 7648
rect 12192 7584 12208 7648
rect 12272 7584 12288 7648
rect 12352 7584 12360 7648
rect 12040 6560 12360 7584
rect 13675 7036 13741 7037
rect 13675 6972 13676 7036
rect 13740 6972 13741 7036
rect 13675 6971 13741 6972
rect 12040 6496 12048 6560
rect 12112 6496 12128 6560
rect 12192 6496 12208 6560
rect 12272 6496 12288 6560
rect 12352 6496 12360 6560
rect 11835 5676 11901 5677
rect 11835 5612 11836 5676
rect 11900 5612 11901 5676
rect 11835 5611 11901 5612
rect 11838 4181 11898 5611
rect 12040 5472 12360 6496
rect 13678 5813 13738 6971
rect 13862 6357 13922 15267
rect 13859 6356 13925 6357
rect 13859 6292 13860 6356
rect 13924 6292 13925 6356
rect 13859 6291 13925 6292
rect 13675 5812 13741 5813
rect 13675 5748 13676 5812
rect 13740 5748 13741 5812
rect 13675 5747 13741 5748
rect 12040 5408 12048 5472
rect 12112 5408 12128 5472
rect 12192 5408 12208 5472
rect 12272 5408 12288 5472
rect 12352 5408 12360 5472
rect 12040 4384 12360 5408
rect 12040 4320 12048 4384
rect 12112 4320 12128 4384
rect 12192 4320 12208 4384
rect 12272 4320 12288 4384
rect 12352 4320 12360 4384
rect 11835 4180 11901 4181
rect 11835 4116 11836 4180
rect 11900 4116 11901 4180
rect 11835 4115 11901 4116
rect 12040 3296 12360 4320
rect 14046 4045 14106 18123
rect 14043 4044 14109 4045
rect 14043 3980 14044 4044
rect 14108 3980 14109 4044
rect 14043 3979 14109 3980
rect 12040 3232 12048 3296
rect 12112 3232 12128 3296
rect 12192 3232 12208 3296
rect 12272 3232 12288 3296
rect 12352 3232 12360 3296
rect 8891 2548 8957 2549
rect 8891 2484 8892 2548
rect 8956 2484 8957 2548
rect 8891 2483 8957 2484
rect 12040 2208 12360 3232
rect 14230 3229 14290 20843
rect 15331 20364 15397 20365
rect 15331 20300 15332 20364
rect 15396 20300 15397 20364
rect 15331 20299 15397 20300
rect 14411 19684 14477 19685
rect 14411 19620 14412 19684
rect 14476 19620 14477 19684
rect 14411 19619 14477 19620
rect 14414 3909 14474 19619
rect 15147 14244 15213 14245
rect 15147 14180 15148 14244
rect 15212 14180 15213 14244
rect 15147 14179 15213 14180
rect 15150 11117 15210 14179
rect 15334 11389 15394 20299
rect 15738 20160 16058 21184
rect 15738 20096 15746 20160
rect 15810 20096 15826 20160
rect 15890 20096 15906 20160
rect 15970 20096 15986 20160
rect 16050 20096 16058 20160
rect 15738 19072 16058 20096
rect 15738 19008 15746 19072
rect 15810 19008 15826 19072
rect 15890 19008 15906 19072
rect 15970 19008 15986 19072
rect 16050 19008 16058 19072
rect 15738 17984 16058 19008
rect 19437 21792 19757 21808
rect 19437 21728 19445 21792
rect 19509 21728 19525 21792
rect 19589 21728 19605 21792
rect 19669 21728 19685 21792
rect 19749 21728 19757 21792
rect 19437 20704 19757 21728
rect 19437 20640 19445 20704
rect 19509 20640 19525 20704
rect 19589 20640 19605 20704
rect 19669 20640 19685 20704
rect 19749 20640 19757 20704
rect 19437 19616 19757 20640
rect 19437 19552 19445 19616
rect 19509 19552 19525 19616
rect 19589 19552 19605 19616
rect 19669 19552 19685 19616
rect 19749 19552 19757 19616
rect 19437 18528 19757 19552
rect 19437 18464 19445 18528
rect 19509 18464 19525 18528
rect 19589 18464 19605 18528
rect 19669 18464 19685 18528
rect 19749 18464 19757 18528
rect 17539 18052 17605 18053
rect 17539 17988 17540 18052
rect 17604 17988 17605 18052
rect 17539 17987 17605 17988
rect 15738 17920 15746 17984
rect 15810 17920 15826 17984
rect 15890 17920 15906 17984
rect 15970 17920 15986 17984
rect 16050 17920 16058 17984
rect 15738 16896 16058 17920
rect 15738 16832 15746 16896
rect 15810 16832 15826 16896
rect 15890 16832 15906 16896
rect 15970 16832 15986 16896
rect 16050 16832 16058 16896
rect 15738 15808 16058 16832
rect 15738 15744 15746 15808
rect 15810 15744 15826 15808
rect 15890 15744 15906 15808
rect 15970 15744 15986 15808
rect 16050 15744 16058 15808
rect 15515 15468 15581 15469
rect 15515 15404 15516 15468
rect 15580 15404 15581 15468
rect 15515 15403 15581 15404
rect 15331 11388 15397 11389
rect 15331 11324 15332 11388
rect 15396 11324 15397 11388
rect 15331 11323 15397 11324
rect 15147 11116 15213 11117
rect 15147 11052 15148 11116
rect 15212 11052 15213 11116
rect 15147 11051 15213 11052
rect 15150 7581 15210 11051
rect 15518 10845 15578 15403
rect 15738 14720 16058 15744
rect 15738 14656 15746 14720
rect 15810 14656 15826 14720
rect 15890 14656 15906 14720
rect 15970 14656 15986 14720
rect 16050 14656 16058 14720
rect 15738 13632 16058 14656
rect 16251 14652 16317 14653
rect 16251 14588 16252 14652
rect 16316 14588 16317 14652
rect 16251 14587 16317 14588
rect 15738 13568 15746 13632
rect 15810 13568 15826 13632
rect 15890 13568 15906 13632
rect 15970 13568 15986 13632
rect 16050 13568 16058 13632
rect 15738 12544 16058 13568
rect 15738 12480 15746 12544
rect 15810 12480 15826 12544
rect 15890 12480 15906 12544
rect 15970 12480 15986 12544
rect 16050 12480 16058 12544
rect 15738 11456 16058 12480
rect 15738 11392 15746 11456
rect 15810 11392 15826 11456
rect 15890 11392 15906 11456
rect 15970 11392 15986 11456
rect 16050 11392 16058 11456
rect 15515 10844 15581 10845
rect 15515 10780 15516 10844
rect 15580 10780 15581 10844
rect 15515 10779 15581 10780
rect 15738 10368 16058 11392
rect 15738 10304 15746 10368
rect 15810 10304 15826 10368
rect 15890 10304 15906 10368
rect 15970 10304 15986 10368
rect 16050 10304 16058 10368
rect 15738 9280 16058 10304
rect 16254 10165 16314 14587
rect 16251 10164 16317 10165
rect 16251 10100 16252 10164
rect 16316 10100 16317 10164
rect 16251 10099 16317 10100
rect 15738 9216 15746 9280
rect 15810 9216 15826 9280
rect 15890 9216 15906 9280
rect 15970 9216 15986 9280
rect 16050 9216 16058 9280
rect 15738 8192 16058 9216
rect 15738 8128 15746 8192
rect 15810 8128 15826 8192
rect 15890 8128 15906 8192
rect 15970 8128 15986 8192
rect 16050 8128 16058 8192
rect 15147 7580 15213 7581
rect 15147 7516 15148 7580
rect 15212 7516 15213 7580
rect 15147 7515 15213 7516
rect 15738 7104 16058 8128
rect 15738 7040 15746 7104
rect 15810 7040 15826 7104
rect 15890 7040 15906 7104
rect 15970 7040 15986 7104
rect 16050 7040 16058 7104
rect 15738 6016 16058 7040
rect 15738 5952 15746 6016
rect 15810 5952 15826 6016
rect 15890 5952 15906 6016
rect 15970 5952 15986 6016
rect 16050 5952 16058 6016
rect 15738 4928 16058 5952
rect 15738 4864 15746 4928
rect 15810 4864 15826 4928
rect 15890 4864 15906 4928
rect 15970 4864 15986 4928
rect 16050 4864 16058 4928
rect 14411 3908 14477 3909
rect 14411 3844 14412 3908
rect 14476 3844 14477 3908
rect 14411 3843 14477 3844
rect 15738 3840 16058 4864
rect 15738 3776 15746 3840
rect 15810 3776 15826 3840
rect 15890 3776 15906 3840
rect 15970 3776 15986 3840
rect 16050 3776 16058 3840
rect 14227 3228 14293 3229
rect 14227 3164 14228 3228
rect 14292 3164 14293 3228
rect 14227 3163 14293 3164
rect 12040 2144 12048 2208
rect 12112 2144 12128 2208
rect 12192 2144 12208 2208
rect 12272 2144 12288 2208
rect 12352 2144 12360 2208
rect 12040 2128 12360 2144
rect 15738 2752 16058 3776
rect 17542 3365 17602 17987
rect 19195 17644 19261 17645
rect 19195 17580 19196 17644
rect 19260 17580 19261 17644
rect 19195 17579 19261 17580
rect 18459 15196 18525 15197
rect 18459 15132 18460 15196
rect 18524 15132 18525 15196
rect 18459 15131 18525 15132
rect 18462 8669 18522 15131
rect 18643 14516 18709 14517
rect 18643 14452 18644 14516
rect 18708 14452 18709 14516
rect 18643 14451 18709 14452
rect 18646 8805 18706 14451
rect 18827 12068 18893 12069
rect 18827 12004 18828 12068
rect 18892 12004 18893 12068
rect 18827 12003 18893 12004
rect 18643 8804 18709 8805
rect 18643 8740 18644 8804
rect 18708 8740 18709 8804
rect 18643 8739 18709 8740
rect 18459 8668 18525 8669
rect 18459 8604 18460 8668
rect 18524 8604 18525 8668
rect 18459 8603 18525 8604
rect 18830 6629 18890 12003
rect 19011 11932 19077 11933
rect 19011 11868 19012 11932
rect 19076 11868 19077 11932
rect 19011 11867 19077 11868
rect 19014 7581 19074 11867
rect 19198 8941 19258 17579
rect 19437 17440 19757 18464
rect 20299 18052 20365 18053
rect 20299 17988 20300 18052
rect 20364 17988 20365 18052
rect 20299 17987 20365 17988
rect 19437 17376 19445 17440
rect 19509 17376 19525 17440
rect 19589 17376 19605 17440
rect 19669 17376 19685 17440
rect 19749 17376 19757 17440
rect 19437 16352 19757 17376
rect 19437 16288 19445 16352
rect 19509 16288 19525 16352
rect 19589 16288 19605 16352
rect 19669 16288 19685 16352
rect 19749 16288 19757 16352
rect 19437 15264 19757 16288
rect 19931 15604 19997 15605
rect 19931 15540 19932 15604
rect 19996 15540 19997 15604
rect 19931 15539 19997 15540
rect 19437 15200 19445 15264
rect 19509 15200 19525 15264
rect 19589 15200 19605 15264
rect 19669 15200 19685 15264
rect 19749 15200 19757 15264
rect 19437 14176 19757 15200
rect 19437 14112 19445 14176
rect 19509 14112 19525 14176
rect 19589 14112 19605 14176
rect 19669 14112 19685 14176
rect 19749 14112 19757 14176
rect 19437 13088 19757 14112
rect 19437 13024 19445 13088
rect 19509 13024 19525 13088
rect 19589 13024 19605 13088
rect 19669 13024 19685 13088
rect 19749 13024 19757 13088
rect 19437 12000 19757 13024
rect 19437 11936 19445 12000
rect 19509 11936 19525 12000
rect 19589 11936 19605 12000
rect 19669 11936 19685 12000
rect 19749 11936 19757 12000
rect 19437 10912 19757 11936
rect 19437 10848 19445 10912
rect 19509 10848 19525 10912
rect 19589 10848 19605 10912
rect 19669 10848 19685 10912
rect 19749 10848 19757 10912
rect 19437 9824 19757 10848
rect 19934 10709 19994 15539
rect 20115 12612 20181 12613
rect 20115 12548 20116 12612
rect 20180 12548 20181 12612
rect 20115 12547 20181 12548
rect 19931 10708 19997 10709
rect 19931 10644 19932 10708
rect 19996 10644 19997 10708
rect 19931 10643 19997 10644
rect 19437 9760 19445 9824
rect 19509 9760 19525 9824
rect 19589 9760 19605 9824
rect 19669 9760 19685 9824
rect 19749 9760 19757 9824
rect 19195 8940 19261 8941
rect 19195 8876 19196 8940
rect 19260 8876 19261 8940
rect 19195 8875 19261 8876
rect 19437 8736 19757 9760
rect 19437 8672 19445 8736
rect 19509 8672 19525 8736
rect 19589 8672 19605 8736
rect 19669 8672 19685 8736
rect 19749 8672 19757 8736
rect 19437 7648 19757 8672
rect 20118 7853 20178 12547
rect 20302 11389 20362 17987
rect 20483 12476 20549 12477
rect 20483 12412 20484 12476
rect 20548 12412 20549 12476
rect 20483 12411 20549 12412
rect 20299 11388 20365 11389
rect 20299 11324 20300 11388
rect 20364 11324 20365 11388
rect 20299 11323 20365 11324
rect 20486 8261 20546 12411
rect 20483 8260 20549 8261
rect 20483 8196 20484 8260
rect 20548 8196 20549 8260
rect 20483 8195 20549 8196
rect 20115 7852 20181 7853
rect 20115 7788 20116 7852
rect 20180 7788 20181 7852
rect 20115 7787 20181 7788
rect 19437 7584 19445 7648
rect 19509 7584 19525 7648
rect 19589 7584 19605 7648
rect 19669 7584 19685 7648
rect 19749 7584 19757 7648
rect 19011 7580 19077 7581
rect 19011 7516 19012 7580
rect 19076 7516 19077 7580
rect 19011 7515 19077 7516
rect 18827 6628 18893 6629
rect 18827 6564 18828 6628
rect 18892 6564 18893 6628
rect 18827 6563 18893 6564
rect 19437 6560 19757 7584
rect 19437 6496 19445 6560
rect 19509 6496 19525 6560
rect 19589 6496 19605 6560
rect 19669 6496 19685 6560
rect 19749 6496 19757 6560
rect 19437 5472 19757 6496
rect 19437 5408 19445 5472
rect 19509 5408 19525 5472
rect 19589 5408 19605 5472
rect 19669 5408 19685 5472
rect 19749 5408 19757 5472
rect 19437 4384 19757 5408
rect 19437 4320 19445 4384
rect 19509 4320 19525 4384
rect 19589 4320 19605 4384
rect 19669 4320 19685 4384
rect 19749 4320 19757 4384
rect 17539 3364 17605 3365
rect 17539 3300 17540 3364
rect 17604 3300 17605 3364
rect 17539 3299 17605 3300
rect 15738 2688 15746 2752
rect 15810 2688 15826 2752
rect 15890 2688 15906 2752
rect 15970 2688 15986 2752
rect 16050 2688 16058 2752
rect 15738 2128 16058 2688
rect 19437 3296 19757 4320
rect 19437 3232 19445 3296
rect 19509 3232 19525 3296
rect 19589 3232 19605 3296
rect 19669 3232 19685 3296
rect 19749 3232 19757 3296
rect 19437 2208 19757 3232
rect 19437 2144 19445 2208
rect 19509 2144 19525 2208
rect 19589 2144 19605 2208
rect 19669 2144 19685 2208
rect 19749 2144 19757 2208
rect 19437 2128 19757 2144
use sky130_fd_sc_hd__buf_2  _68_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2484 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1748 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606256979
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606256979
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_13 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_19
timestamp 1606256979
transform 1 0 2852 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _64_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 4876 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1606256979
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1606256979
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_31 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3956 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_39
timestamp 1606256979
transform 1 0 4692 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606256979
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606256979
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1606256979
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1606256979
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1606256979
transform 1 0 5152 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_56
timestamp 1606256979
transform 1 0 6256 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1606256979
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1606256979
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1606256979
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1606256979
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1606256979
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606256979
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1606256979
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1606256979
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1606256979
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606256979
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606256979
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1606256979
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125
timestamp 1606256979
transform 1 0 12604 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1606256979
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_123
timestamp 1606256979
transform 1 0 12420 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_131
timestamp 1606256979
transform 1 0 13156 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 14352 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1606256979
transform 1 0 13248 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1606256979
transform 1 0 13340 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1606256979
transform 1 0 14076 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 15088 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_142
timestamp 1606256979
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_150
timestamp 1606256979
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15272 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1606256979
transform 1 0 16192 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 16284 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606256979
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1606256979
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_156
timestamp 1606256979
transform 1 0 15456 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_173
timestamp 1606256979
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_163
timestamp 1606256979
transform 1 0 16100 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1606256979
transform 1 0 17204 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1606256979
transform 1 0 18308 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1606256979
transform 1 0 18216 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606256979
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606256979
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1606256979
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1606256979
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_184
timestamp 1606256979
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1606256979
transform 1 0 21160 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1606256979
transform 1 0 20700 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 20056 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1606256979
transform 1 0 19964 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606256979
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_203
timestamp 1606256979
transform 1 0 19780 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1606256979
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_202
timestamp 1606256979
transform 1 0 19688 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_211
timestamp 1606256979
transform 1 0 20516 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1606256979
transform 1 0 22356 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606256979
transform -1 0 23276 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606256979
transform -1 0 23276 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_234
timestamp 1606256979
transform 1 0 22632 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_229
timestamp 1606256979
transform 1 0 22172 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_235
timestamp 1606256979
transform 1 0 22724 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606256979
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606256979
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1606256979
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606256979
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1606256979
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1606256979
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1606256979
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1606256979
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1606256979
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1606256979
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1606256979
transform 1 0 11132 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606256979
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1606256979
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_105
timestamp 1606256979
transform 1 0 10764 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13156 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1606256979
transform 1 0 12144 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_118
timestamp 1606256979
transform 1 0 11960 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_129
timestamp 1606256979
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1606256979
transform 1 0 14168 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_140
timestamp 1606256979
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1606256979
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1606256979
transform 1 0 15548 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1606256979
transform 1 0 17112 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16100 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606256979
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1606256979
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_161
timestamp 1606256979
transform 1 0 15916 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_172
timestamp 1606256979
transform 1 0 16928 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1606256979
transform 1 0 18952 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_190
timestamp 1606256979
transform 1 0 18584 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1606256979
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606256979
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_210
timestamp 1606256979
transform 1 0 20424 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_218
timestamp 1606256979
transform 1 0 21160 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1606256979
transform 1 0 21344 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606256979
transform -1 0 23276 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_236
timestamp 1606256979
transform 1 0 22816 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606256979
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606256979
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1606256979
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1606256979
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1606256979
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606256979
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1606256979
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606256979
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1606256979
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1606256979
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1606256979
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1606256979
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1606256979
transform 1 0 11316 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12604 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606256979
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_110
timestamp 1606256979
transform 1 0 11224 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1606256979
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_123
timestamp 1606256979
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 14628 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1606256979
transform 1 0 13616 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_134
timestamp 1606256979
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_145
timestamp 1606256979
transform 1 0 14444 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606256979
transform 1 0 16284 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_163
timestamp 1606256979
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1606256979
transform 1 0 19044 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1606256979
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606256979
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1606256979
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp 1606256979
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1606256979
transform 1 0 19504 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_198
timestamp 1606256979
transform 1 0 19320 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_216
timestamp 1606256979
transform 1 0 20976 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1606256979
transform 1 0 21344 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606256979
transform -1 0 23276 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_236
timestamp 1606256979
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606256979
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606256979
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1606256979
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606256979
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1606256979
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1606256979
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1606256979
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1606256979
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1606256979
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1606256979
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10856 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1606256979
transform 1 0 9844 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606256979
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1606256979
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_104
timestamp 1606256979
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11868 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12880 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_115
timestamp 1606256979
transform 1 0 11684 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_126
timestamp 1606256979
transform 1 0 12696 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1606256979
transform 1 0 13892 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_137
timestamp 1606256979
transform 1 0 13708 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1606256979
transform 1 0 14720 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1606256979
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1606256979
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 15824 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606256979
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_158
timestamp 1606256979
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1606256979
transform 1 0 18768 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1606256979
transform 1 0 17756 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_176
timestamp 1606256979
transform 1 0 17296 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_180
timestamp 1606256979
transform 1 0 17664 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_190
timestamp 1606256979
transform 1 0 18584 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1606256979
transform 1 0 19780 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1606256979
transform 1 0 21068 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606256979
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_201
timestamp 1606256979
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1606256979
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_215
timestamp 1606256979
transform 1 0 20884 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606256979
transform -1 0 23276 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_233
timestamp 1606256979
transform 1 0 22540 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_237
timestamp 1606256979
transform 1 0 22908 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606256979
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606256979
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606256979
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1606256979
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1606256979
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606256979
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1606256979
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606256979
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_62
timestamp 1606256979
transform 1 0 6808 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1606256979
transform 1 0 7636 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1606256979
transform 1 0 9108 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_70
timestamp 1606256979
transform 1 0 7544 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_80
timestamp 1606256979
transform 1 0 8464 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_86
timestamp 1606256979
transform 1 0 9016 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1606256979
transform 1 0 11132 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1606256979
transform 1 0 10120 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_96
timestamp 1606256979
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_107
timestamp 1606256979
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1606256979
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606256979
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1606256979
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13524 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_5_132
timestamp 1606256979
transform 1 0 13248 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_151
timestamp 1606256979
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16836 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15180 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1606256979
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1606256979
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1606256979
transform 1 0 18492 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606256979
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_180
timestamp 1606256979
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_187
timestamp 1606256979
transform 1 0 18308 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1606256979
transform 1 0 19596 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606256979
transform 1 0 20608 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1606256979
transform 1 0 21160 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_5_198
timestamp 1606256979
transform 1 0 19320 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_210
timestamp 1606256979
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_216
timestamp 1606256979
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606256979
transform -1 0 23276 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_234
timestamp 1606256979
transform 1 0 22632 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606256979
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606256979
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606256979
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606256979
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606256979
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1606256979
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606256979
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606256979
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1606256979
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1606256979
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_39
timestamp 1606256979
transform 1 0 4692 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5520 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6532 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5612 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606256979
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_44
timestamp 1606256979
transform 1 0 5152 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_57
timestamp 1606256979
transform 1 0 6348 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_47
timestamp 1606256979
transform 1 0 5428 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_58
timestamp 1606256979
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_62
timestamp 1606256979
transform 1 0 6808 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1606256979
transform 1 0 7544 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1606256979
transform 1 0 7636 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8648 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8556 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_68
timestamp 1606256979
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_79
timestamp 1606256979
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_70
timestamp 1606256979
transform 1 0 7544 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_80
timestamp 1606256979
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1606256979
transform 1 0 9660 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1606256979
transform 1 0 10672 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1606256979
transform 1 0 10580 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606256979
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1606256979
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_93
timestamp 1606256979
transform 1 0 9660 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_101
timestamp 1606256979
transform 1 0 10396 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_91
timestamp 1606256979
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_102
timestamp 1606256979
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606256979
transform 1 0 12512 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1606256979
transform 1 0 12236 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1606256979
transform 1 0 13064 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606256979
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_119
timestamp 1606256979
transform 1 0 12052 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1606256979
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_123
timestamp 1606256979
transform 1 0 12420 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_128
timestamp 1606256979
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1606256979
transform 1 0 13892 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1606256979
transform 1 0 14720 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_137
timestamp 1606256979
transform 1 0 13708 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_148
timestamp 1606256979
transform 1 0 14720 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_146
timestamp 1606256979
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_161
timestamp 1606256979
transform 1 0 15916 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1606256979
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606256979
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16100 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1606256979
transform 1 0 15548 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_170
timestamp 1606256979
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_164
timestamp 1606256979
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_172
timestamp 1606256979
transform 1 0 16928 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16928 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606256979
transform 1 0 16376 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 17112 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606256979
transform 1 0 18216 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18768 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 18768 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606256979
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_190
timestamp 1606256979
transform 1 0 18584 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1606256979
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1606256979
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_190
timestamp 1606256979
transform 1 0 18584 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1606256979
transform 1 0 19780 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606256979
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 20700 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606256979
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_201
timestamp 1606256979
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1606256979
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_208
timestamp 1606256979
transform 1 0 20240 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_212
timestamp 1606256979
transform 1 0 20608 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_218
timestamp 1606256979
transform 1 0 21160 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1606256979
transform 1 0 21436 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1606256979
transform 1 0 22448 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 21344 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606256979
transform -1 0 23276 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606256979
transform -1 0 23276 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_219
timestamp 1606256979
transform 1 0 21252 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_230
timestamp 1606256979
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_236
timestamp 1606256979
transform 1 0 22816 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_236
timestamp 1606256979
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606256979
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1606256979
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1606256979
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4508 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606256979
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606256979
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 1606256979
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_36
timestamp 1606256979
transform 1 0 4416 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5520 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1606256979
transform 1 0 6532 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_46
timestamp 1606256979
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_57
timestamp 1606256979
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1606256979
transform 1 0 7544 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1606256979
transform 1 0 8556 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_68
timestamp 1606256979
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_79
timestamp 1606256979
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1606256979
transform 1 0 10396 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606256979
transform 1 0 9844 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606256979
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1606256979
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1606256979
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_99
timestamp 1606256979
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12512 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_117
timestamp 1606256979
transform 1 0 11868 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_123
timestamp 1606256979
transform 1 0 12420 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1606256979
transform 1 0 13524 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_133
timestamp 1606256979
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1606256979
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15640 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606256979
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_154
timestamp 1606256979
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_174
timestamp 1606256979
transform 1 0 17112 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1606256979
transform 1 0 17296 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 17756 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_179
timestamp 1606256979
transform 1 0 17572 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 19412 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 20884 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606256979
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 20424 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1606256979
transform 1 0 19228 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_208
timestamp 1606256979
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1606256979
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1606256979
transform 1 0 22540 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606256979
transform -1 0 23276 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_231
timestamp 1606256979
transform 1 0 22356 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_236
timestamp 1606256979
transform 1 0 22816 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606256979
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606256979
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1606256979
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 3680 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4692 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1606256979
transform 1 0 3588 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_37
timestamp 1606256979
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1606256979
transform 1 0 5704 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606256979
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_48
timestamp 1606256979
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1606256979
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_62
timestamp 1606256979
transform 1 0 6808 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8556 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1606256979
transform 1 0 7544 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_79
timestamp 1606256979
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606256979
transform 1 0 10212 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_97
timestamp 1606256979
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12512 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606256979
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_115
timestamp 1606256979
transform 1 0 11684 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1606256979
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_123
timestamp 1606256979
transform 1 0 12420 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1606256979
transform 1 0 13524 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_133
timestamp 1606256979
transform 1 0 13340 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_151
timestamp 1606256979
transform 1 0 14996 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 15824 0 1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606256979
transform 1 0 15272 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_158
timestamp 1606256979
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606256979
transform 1 0 18400 0 1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606256979
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1606256979
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp 1606256979
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 20516 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_209
timestamp 1606256979
transform 1 0 20332 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  Test_en_E_FTB01
timestamp 1606256979
transform 1 0 22172 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606256979
transform -1 0 23276 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_227
timestamp 1606256979
transform 1 0 21988 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_235
timestamp 1606256979
transform 1 0 22724 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606256979
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1606256979
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_11
timestamp 1606256979
transform 1 0 2116 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  Test_en_FTB00
timestamp 1606256979
transform 1 0 4416 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606256979
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_25
timestamp 1606256979
transform 1 0 3404 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1606256979
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606256979
transform 1 0 5704 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6532 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_48
timestamp 1606256979
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_54
timestamp 1606256979
transform 1 0 6072 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_58
timestamp 1606256979
transform 1 0 6440 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1606256979
transform 1 0 8556 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1606256979
transform 1 0 7544 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_68
timestamp 1606256979
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_79
timestamp 1606256979
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 9752 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606256979
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1606256979
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_93
timestamp 1606256979
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1606256979
transform 1 0 13064 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 11408 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_110
timestamp 1606256979
transform 1 0 11224 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_128
timestamp 1606256979
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1606256979
transform 1 0 14720 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_146
timestamp 1606256979
transform 1 0 14536 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1606256979
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15640 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606256979
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1606256979
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_174
timestamp 1606256979
transform 1 0 17112 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606256979
transform 1 0 17296 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 17940 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_10_180
timestamp 1606256979
transform 1 0 17664 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 19596 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_E_FTB01
timestamp 1606256979
transform 1 0 20976 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606256979
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_199
timestamp 1606256979
transform 1 0 19412 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_210
timestamp 1606256979
transform 1 0 20424 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_215
timestamp 1606256979
transform 1 0 20884 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 21712 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606256979
transform -1 0 23276 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_222
timestamp 1606256979
transform 1 0 21528 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_233
timestamp 1606256979
transform 1 0 22540 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_237
timestamp 1606256979
transform 1 0 22908 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1606256979
transform 1 0 2944 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 1932 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606256979
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1606256979
transform 1 0 1380 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_18
timestamp 1606256979
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1606256979
transform 1 0 3956 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1606256979
transform 1 0 4692 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_29
timestamp 1606256979
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_35
timestamp 1606256979
transform 1 0 4324 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1606256979
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5704 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606256979
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_48
timestamp 1606256979
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1606256979
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8740 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1606256979
transform 1 0 7728 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_11_66
timestamp 1606256979
transform 1 0 7176 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_81
timestamp 1606256979
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 9752 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_92
timestamp 1606256979
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606256979
transform 1 0 11408 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1606256979
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606256979
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 13064 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 11960 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1606256979
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_116
timestamp 1606256979
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1606256979
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_127
timestamp 1606256979
transform 1 0 12788 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606256979
transform 1 0 14996 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1606256979
transform 1 0 13340 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_149
timestamp 1606256979
transform 1 0 14812 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15548 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_155
timestamp 1606256979
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_173
timestamp 1606256979
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 19136 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18124 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1606256979
transform 1 0 17204 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606256979
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1606256979
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_184
timestamp 1606256979
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_194
timestamp 1606256979
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 20792 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_212
timestamp 1606256979
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606256979
transform 1 0 22448 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606256979
transform -1 0 23276 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_230
timestamp 1606256979
transform 1 0 22264 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_236
timestamp 1606256979
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1606256979
transform 1 0 2852 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 1840 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606256979
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1606256979
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1606256979
transform 1 0 1748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_17
timestamp 1606256979
transform 1 0 2668 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1606256979
transform 1 0 5060 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606256979
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_28
timestamp 1606256979
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1606256979
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1606256979
transform 1 0 6532 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_12_52
timestamp 1606256979
transform 1 0 5888 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_58
timestamp 1606256979
transform 1 0 6440 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1606256979
transform 1 0 7544 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1606256979
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_68
timestamp 1606256979
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_79
timestamp 1606256979
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10580 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1606256979
transform 1 0 10028 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606256979
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1606256979
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1606256979
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_101
timestamp 1606256979
transform 1 0 10396 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1606256979
transform 1 0 11592 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1606256979
transform 1 0 12972 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 12696 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_112
timestamp 1606256979
transform 1 0 11408 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_123
timestamp 1606256979
transform 1 0 12420 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1606256979
transform 1 0 13524 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_133
timestamp 1606256979
transform 1 0 13340 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1606256979
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16468 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15456 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606256979
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_154
timestamp 1606256979
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_165
timestamp 1606256979
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606256979
transform 1 0 18308 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_12_183
timestamp 1606256979
transform 1 0 17940 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606256979
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_208
timestamp 1606256979
transform 1 0 20240 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1606256979
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 21252 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606256979
transform -1 0 23276 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_235
timestamp 1606256979
transform 1 0 22724 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1606256979
transform 1 0 1472 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 1380 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 2024 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 3036 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606256979
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606256979
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1606256979
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_19
timestamp 1606256979
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1606256979
transform 1 0 1380 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _51_
timestamp 1606256979
transform 1 0 4692 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606256979
transform 1 0 4140 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606256979
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_37
timestamp 1606256979
transform 1 0 4508 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_42
timestamp 1606256979
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_26
timestamp 1606256979
transform 1 0 3496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1606256979
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_32
timestamp 1606256979
transform 1 0 4048 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1606256979
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1606256979
transform 1 0 5796 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606256979
transform 1 0 6164 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606256979
transform 1 0 7084 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606256979
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_53
timestamp 1606256979
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606256979
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_62
timestamp 1606256979
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_49
timestamp 1606256979
transform 1 0 5612 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1606256979
transform 1 0 7636 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1606256979
transform 1 0 7912 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1606256979
transform 1 0 8648 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_13_69
timestamp 1606256979
transform 1 0 7452 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_80
timestamp 1606256979
transform 1 0 8464 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_67
timestamp 1606256979
transform 1 0 7268 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_73
timestamp 1606256979
transform 1 0 7820 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1606256979
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1606256979
transform 1 0 10304 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606256979
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_98
timestamp 1606256979
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1606256979
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_109
timestamp 1606256979
transform 1 0 11132 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1606256979
transform 1 0 11684 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1606256979
transform 1 0 12696 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1606256979
transform 1 0 12696 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606256979
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_116
timestamp 1606256979
transform 1 0 11776 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_123
timestamp 1606256979
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_124
timestamp 1606256979
transform 1 0 12512 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1606256979
transform 1 0 14352 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1606256979
transform 1 0 14628 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 14352 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_142
timestamp 1606256979
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_152
timestamp 1606256979
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_142
timestamp 1606256979
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_148
timestamp 1606256979
transform 1 0 14720 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16928 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15272 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15456 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606256979
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_170
timestamp 1606256979
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1606256979
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_172
timestamp 1606256979
transform 1 0 16928 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606256979
transform 1 0 19136 0 1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 18216 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 17204 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 18124 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606256979
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1606256979
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_184
timestamp 1606256979
transform 1 0 18032 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_194
timestamp 1606256979
transform 1 0 18952 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_184
timestamp 1606256979
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606256979
transform 1 0 19872 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606256979
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 20424 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_217
timestamp 1606256979
transform 1 0 21068 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_202
timestamp 1606256979
transform 1 0 19688 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_208
timestamp 1606256979
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1606256979
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1606256979
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606256979
transform 1 0 21252 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 21344 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 21804 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606256979
transform -1 0 23276 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606256979
transform -1 0 23276 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_236
timestamp 1606256979
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_223
timestamp 1606256979
transform 1 0 21620 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_234
timestamp 1606256979
transform 1 0 22632 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1606256979
transform 1 0 1748 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606256979
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1606256979
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 3404 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1606256979
transform 1 0 5060 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_23
timestamp 1606256979
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_41
timestamp 1606256979
transform 1 0 4876 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606256979
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606256979
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1606256979
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1606256979
transform 1 0 9108 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1606256979
transform 1 0 7452 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_15_66
timestamp 1606256979
transform 1 0 7176 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_85
timestamp 1606256979
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1606256979
transform 1 0 9936 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 9660 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_91
timestamp 1606256979
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606256979
transform 1 0 11776 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606256979
transform 1 0 12512 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606256979
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_112
timestamp 1606256979
transform 1 0 11408 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1606256979
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_123
timestamp 1606256979
transform 1 0 12420 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1606256979
transform 1 0 14168 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_140
timestamp 1606256979
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 15824 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_158
timestamp 1606256979
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1606256979
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606256979
transform 1 0 17296 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 18216 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606256979
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1606256979
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_195
timestamp 1606256979
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1606256979
transform 1 0 19228 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 19688 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_200
timestamp 1606256979
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_218
timestamp 1606256979
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606256979
transform 1 0 22356 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 21344 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606256979
transform -1 0 23276 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_229
timestamp 1606256979
transform 1 0 22172 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_235
timestamp 1606256979
transform 1 0 22724 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1606256979
transform 1 0 1380 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606256979
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_19
timestamp 1606256979
transform 1 0 2852 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1606256979
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606256979
transform 1 0 3404 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606256979
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 3128 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1606256979
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_41
timestamp 1606256979
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _56_
timestamp 1606256979
transform 1 0 6808 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1606256979
transform 1 0 5152 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_60
timestamp 1606256979
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_65
timestamp 1606256979
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1606256979
transform 1 0 9016 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1606256979
transform 1 0 7268 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_83
timestamp 1606256979
transform 1 0 8740 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1606256979
transform 1 0 9844 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1606256979
transform 1 0 10396 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606256979
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1606256979
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1606256979
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_99
timestamp 1606256979
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1606256979
transform 1 0 12236 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1606256979
transform 1 0 12788 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_117
timestamp 1606256979
transform 1 0 11868 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_125
timestamp 1606256979
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1606256979
transform 1 0 14628 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_143
timestamp 1606256979
transform 1 0 14260 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1606256979
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1606256979
transform 1 0 17112 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 15640 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606256979
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_154
timestamp 1606256979
transform 1 0 15272 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606256979
transform 1 0 17940 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606256979
transform 1 0 20240 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606256979
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_204
timestamp 1606256979
transform 1 0 19872 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1606256979
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1606256979
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 21252 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606256979
transform -1 0 23276 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_235
timestamp 1606256979
transform 1 0 22724 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1606256979
transform 1 0 3036 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1606256979
transform 1 0 1380 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606256979
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_19
timestamp 1606256979
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1606256979
transform 1 0 4048 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1606256979
transform 1 0 5060 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_30
timestamp 1606256979
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_41
timestamp 1606256979
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606256979
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1606256979
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_62
timestamp 1606256979
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1606256979
transform 1 0 7176 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 8832 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_82
timestamp 1606256979
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_87
timestamp 1606256979
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1606256979
transform 1 0 9292 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1606256979
transform 1 0 10304 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_98
timestamp 1606256979
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606256979
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606256979
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ltile_clb_mode__0.clb_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 12604 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_17_116
timestamp 1606256979
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1606256979
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1606256979
transform 1 0 14444 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16928 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15916 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1606256979
transform 1 0 15272 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_158
timestamp 1606256979
transform 1 0 15640 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_170
timestamp 1606256979
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606256979
transform 1 0 19044 0 1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606256979
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1606256979
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1606256979
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_216
timestamp 1606256979
transform 1 0 20976 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 21344 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606256979
transform -1 0 23276 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1606256979
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1606256979
transform 1 0 1564 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606256979
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1606256979
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_21
timestamp 1606256979
transform 1 0 3036 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1606256979
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1606256979
transform 1 0 3404 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606256979
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 5060 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1606256979
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_41
timestamp 1606256979
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1606256979
transform 1 0 5336 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606256979
transform 1 0 6440 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606256979
transform 1 0 6992 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_55
timestamp 1606256979
transform 1 0 6164 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_62
timestamp 1606256979
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606256979
transform 1 0 9016 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 8648 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_80
timestamp 1606256979
transform 1 0 8464 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1606256979
transform 1 0 8924 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606256979
transform 1 0 9752 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606256979
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_ltile_clb_mode__0.clb_clk
timestamp 1606256979
transform 1 0 10488 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 10948 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1606256979
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_93
timestamp 1606256979
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1606256979
transform 1 0 10120 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_105
timestamp 1606256979
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 11408 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_18_110
timestamp 1606256979
transform 1 0 11224 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1606256979
transform 1 0 13248 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_ltile_clb_mode__0.clb_clk
timestamp 1606256979
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_148
timestamp 1606256979
transform 1 0 14720 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1606256979
transform 1 0 17020 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1606256979
transform 1 0 16008 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1606256979
transform 1 0 15456 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606256979
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1606256979
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_160
timestamp 1606256979
transform 1 0 15824 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_171
timestamp 1606256979
transform 1 0 16836 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 17480 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_176
timestamp 1606256979
transform 1 0 17296 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_194
timestamp 1606256979
transform 1 0 18952 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 20884 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 19412 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606256979
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_198
timestamp 1606256979
transform 1 0 19320 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_208
timestamp 1606256979
transform 1 0 20240 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1606256979
transform 1 0 22540 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606256979
transform -1 0 23276 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_231
timestamp 1606256979
transform 1 0 22356 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_236
timestamp 1606256979
transform 1 0 22816 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_10
timestamp 1606256979
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1606256979
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 1606256979
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606256979
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606256979
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606256979
transform 1 0 1656 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1606256979
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_21
timestamp 1606256979
transform 1 0 3036 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 2208 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1606256979
transform 1 0 1932 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606256979
transform 1 0 3404 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1606256979
transform 1 0 3588 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1606256979
transform 1 0 4416 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606256979
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_25
timestamp 1606256979
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_43
timestamp 1606256979
transform 1 0 5060 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1606256979
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_32
timestamp 1606256979
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_52
timestamp 1606256979
transform 1 0 5888 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1606256979
transform 1 0 6072 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1606256979
transform 1 0 6072 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1606256979
transform 1 0 5244 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_59
timestamp 1606256979
transform 1 0 6532 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1606256979
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606256979
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _55_
timestamp 1606256979
transform 1 0 6256 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 6716 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1606256979
transform 1 0 8464 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1606256979
transform 1 0 8372 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_78
timestamp 1606256979
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_77
timestamp 1606256979
transform 1 0 8188 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _59_
timestamp 1606256979
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1606256979
transform 1 0 9476 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1606256979
transform 1 0 9844 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1606256979
transform 1 0 10304 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1606256979
transform 1 0 10672 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606256979
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_89
timestamp 1606256979
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_88
timestamp 1606256979
transform 1 0 9200 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_93
timestamp 1606256979
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1606256979
transform 1 0 11868 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 12144 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1606256979
transform 1 0 12604 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606256979
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_116
timestamp 1606256979
transform 1 0 11776 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1606256979
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1606256979
transform 1 0 14168 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1606256979
transform 1 0 13616 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_19_141
timestamp 1606256979
transform 1 0 14076 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_151
timestamp 1606256979
transform 1 0 14996 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1606256979
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1606256979
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1606256979
transform 1 0 16652 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1606256979
transform 1 0 15180 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1606256979
transform 1 0 15732 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606256979
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_157
timestamp 1606256979
transform 1 0 15548 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_181
timestamp 1606256979
transform 1 0 17756 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_175
timestamp 1606256979
transform 1 0 17204 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_178
timestamp 1606256979
transform 1 0 17480 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606256979
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606256979
transform 1 0 17388 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606256979
transform 1 0 18032 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_188
timestamp 1606256979
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 18584 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 17940 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_199
timestamp 1606256979
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_206
timestamp 1606256979
transform 1 0 20056 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 19596 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_210
timestamp 1606256979
transform 1 0 20424 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_212
timestamp 1606256979
transform 1 0 20608 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606256979
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606256979
transform 1 0 20240 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _50_
timestamp 1606256979
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_218
timestamp 1606256979
transform 1 0 21160 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 21160 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1606256979
transform 1 0 22172 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 21344 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606256979
transform -1 0 23276 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606256979
transform -1 0 23276 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_227
timestamp 1606256979
transform 1 0 21988 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_233
timestamp 1606256979
transform 1 0 22540 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_237
timestamp 1606256979
transform 1 0 22908 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_236
timestamp 1606256979
transform 1 0 22816 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 1472 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606256979
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1606256979
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_20
timestamp 1606256979
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1606256979
transform 1 0 4140 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1606256979
transform 1 0 4876 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 3128 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_31
timestamp 1606256979
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_37
timestamp 1606256979
transform 1 0 4508 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606256979
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1606256979
transform 1 0 6348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _54_
timestamp 1606256979
transform 1 0 7820 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8280 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1606256979
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_76
timestamp 1606256979
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1606256979
transform 1 0 9936 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1606256979
transform 1 0 10948 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_94
timestamp 1606256979
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_105
timestamp 1606256979
transform 1 0 10764 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1606256979
transform 1 0 12788 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606256979
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 11960 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_116
timestamp 1606256979
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1606256979
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_123
timestamp 1606256979
transform 1 0 12420 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1606256979
transform 1 0 14536 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_21_143
timestamp 1606256979
transform 1 0 14260 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1606256979
transform 1 0 16284 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_21_162
timestamp 1606256979
transform 1 0 16008 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18216 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606256979
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1606256979
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_184
timestamp 1606256979
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_195
timestamp 1606256979
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606256979
transform 1 0 19596 0 1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 19228 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_200
timestamp 1606256979
transform 1 0 19504 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 21712 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606256979
transform -1 0 23276 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1606256979
transform 1 0 21528 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_233
timestamp 1606256979
transform 1 0 22540 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_237
timestamp 1606256979
transform 1 0 22908 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 1656 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606256979
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1606256979
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606256979
transform 1 0 3404 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5060 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606256979
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_22
timestamp 1606256979
transform 1 0 3128 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1606256979
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_41
timestamp 1606256979
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606256979
transform 1 0 6072 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6624 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_52
timestamp 1606256979
transform 1 0 5888 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_58
timestamp 1606256979
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8556 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 8280 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_76
timestamp 1606256979
transform 1 0 8096 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9844 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606256979
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1606256979
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1606256979
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1606256979
transform 1 0 11500 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1606256979
transform 1 0 12420 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_111
timestamp 1606256979
transform 1 0 11316 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_122
timestamp 1606256979
transform 1 0 12328 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13892 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606256979
transform 1 0 14720 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1606256979
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1606256979
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1606256979
transform 1 0 15732 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606256979
transform 1 0 16744 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606256979
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_157
timestamp 1606256979
transform 1 0 15548 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_168
timestamp 1606256979
transform 1 0 16560 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_174
timestamp 1606256979
transform 1 0 17112 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1606256979
transform 1 0 19136 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 17480 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1606256979
transform 1 0 18952 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 21160 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 19780 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606256979
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_201
timestamp 1606256979
transform 1 0 19596 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1606256979
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_215
timestamp 1606256979
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606256979
transform -1 0 23276 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_234
timestamp 1606256979
transform 1 0 22632 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _52_
timestamp 1606256979
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 1840 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606256979
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_6
timestamp 1606256979
transform 1 0 1656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606256979
transform 1 0 4140 0 1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606256979
transform 1 0 3588 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_24
timestamp 1606256979
transform 1 0 3312 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_31
timestamp 1606256979
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _58_
timestamp 1606256979
transform 1 0 6256 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606256979
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1606256979
transform 1 0 6072 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1606256979
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _60_
timestamp 1606256979
transform 1 0 8464 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8924 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_78
timestamp 1606256979
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_83
timestamp 1606256979
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10672 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_23_101
timestamp 1606256979
transform 1 0 10396 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1606256979
transform 1 0 12512 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606256979
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1606256979
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_123
timestamp 1606256979
transform 1 0 12420 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13432 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_23_133
timestamp 1606256979
transform 1 0 13340 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_150
timestamp 1606256979
transform 1 0 14904 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1606256979
transform 1 0 15272 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 16284 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_163
timestamp 1606256979
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  clk_0_FTB00
timestamp 1606256979
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606256979
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1606256979
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_196
timestamp 1606256979
transform 1 0 19136 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606256979
transform 1 0 19320 0 1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606256979
transform 1 0 22448 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 21436 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606256979
transform -1 0 23276 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_219
timestamp 1606256979
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_230
timestamp 1606256979
transform 1 0 22264 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_236
timestamp 1606256979
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 1472 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606256979
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1606256979
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_20
timestamp 1606256979
transform 1 0 2944 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  Test_en_W_FTB01
timestamp 1606256979
transform 1 0 3128 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606256979
transform 1 0 4968 0 -1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606256979
transform 1 0 4416 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606256979
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_28
timestamp 1606256979
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_32
timestamp 1606256979
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_40
timestamp 1606256979
transform 1 0 4784 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7084 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_63
timestamp 1606256979
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606256979
transform 1 0 9016 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 8740 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_81
timestamp 1606256979
transform 1 0 8556 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606256979
transform 1 0 11040 0 -1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606256979
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 10764 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1606256979
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_102
timestamp 1606256979
transform 1 0 10488 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13156 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_129
timestamp 1606256979
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_147
timestamp 1606256979
transform 1 0 14628 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606256979
transform 1 0 15272 0 -1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606256979
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606256979
transform 1 0 17388 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 17940 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_175
timestamp 1606256979
transform 1 0 17204 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_181
timestamp 1606256979
transform 1 0 17756 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 20884 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 19780 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606256979
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_199
timestamp 1606256979
transform 1 0 19412 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1606256979
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _49_
timestamp 1606256979
transform 1 0 22540 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606256979
transform -1 0 23276 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_231
timestamp 1606256979
transform 1 0 22356 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_236
timestamp 1606256979
transform 1 0 22816 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1606256979
transform 1 0 1472 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2024 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606256979
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1606256979
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_8
timestamp 1606256979
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606256979
transform 1 0 4048 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 3772 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_26
timestamp 1606256979
transform 1 0 3496 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606256979
transform 1 0 6808 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606256979
transform 1 0 6164 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606256979
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1606256979
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1606256979
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606256979
transform 1 0 8924 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_25_83
timestamp 1606256979
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11040 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_106
timestamp 1606256979
transform 1 0 10856 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606256979
transform 1 0 11960 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606256979
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_117
timestamp 1606256979
transform 1 0 11868 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606256979
transform 1 0 13340 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_25_132
timestamp 1606256979
transform 1 0 13248 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15548 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_25_154
timestamp 1606256979
transform 1 0 15272 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_173
timestamp 1606256979
transform 1 0 17020 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1606256979
transform 1 0 17296 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 18032 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606256979
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1606256979
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 19872 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_200
timestamp 1606256979
transform 1 0 19504 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _48_
timestamp 1606256979
transform 1 0 22540 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 21528 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606256979
transform -1 0 23276 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_220
timestamp 1606256979
transform 1 0 21344 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_231
timestamp 1606256979
transform 1 0 22356 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1606256979
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606256979
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 1932 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2116 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606256979
transform 1 0 1564 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606256979
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606256979
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_7
timestamp 1606256979
transform 1 0 1748 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1606256979
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_9
timestamp 1606256979
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5060 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4784 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 3772 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606256979
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_25
timestamp 1606256979
transform 1 0 3404 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_41
timestamp 1606256979
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_27
timestamp 1606256979
transform 1 0 3588 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_38
timestamp 1606256979
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1606256979
transform 1 0 6164 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6808 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6256 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606256979
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 5888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_52
timestamp 1606256979
transform 1 0 5888 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_49
timestamp 1606256979
transform 1 0 5612 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1606256979
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8464 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7912 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_26_72
timestamp 1606256979
transform 1 0 7728 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_78
timestamp 1606256979
transform 1 0 8280 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9660 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10304 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606256979
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1606256979
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_109
timestamp 1606256979
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_96
timestamp 1606256979
transform 1 0 9936 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 11684 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 12604 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606256979
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 11316 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_114
timestamp 1606256979
transform 1 0 11592 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_131
timestamp 1606256979
transform 1 0 13156 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_116
timestamp 1606256979
transform 1 0 11776 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_123
timestamp 1606256979
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_141
timestamp 1606256979
transform 1 0 14076 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13340 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_147
timestamp 1606256979
transform 1 0 14628 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_151
timestamp 1606256979
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_142
timestamp 1606256979
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 14812 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 14352 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606256979
transform 1 0 14260 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606256979
transform 1 0 14628 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15088 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15272 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16928 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606256979
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 16928 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_170
timestamp 1606256979
transform 1 0 16744 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_168
timestamp 1606256979
transform 1 0 16560 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1606256979
transform 1 0 18584 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606256979
transform 1 0 18032 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606256979
transform 1 0 17204 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 17756 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606256979
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_179
timestamp 1606256979
transform 1 0 17572 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1606256979
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_188
timestamp 1606256979
transform 1 0 18400 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_199
timestamp 1606256979
transform 1 0 19412 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1606256979
transform 1 0 19228 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 19780 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1606256979
transform 1 0 19412 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_212
timestamp 1606256979
transform 1 0 20608 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_218
timestamp 1606256979
transform 1 0 21160 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_208
timestamp 1606256979
transform 1 0 20240 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606256979
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1606256979
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 20792 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606256979
transform 1 0 22448 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 21344 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606256979
transform -1 0 23276 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606256979
transform -1 0 23276 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_236
timestamp 1606256979
transform 1 0 22816 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_230
timestamp 1606256979
transform 1 0 22264 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_236
timestamp 1606256979
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 2208 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1606256979
transform 1 0 1656 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606256979
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1606256979
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_10
timestamp 1606256979
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606256979
transform 1 0 4232 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4784 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606256979
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_28
timestamp 1606256979
transform 1 0 3680 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_32
timestamp 1606256979
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_38
timestamp 1606256979
transform 1 0 4600 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6440 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_56
timestamp 1606256979
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _57_
timestamp 1606256979
transform 1 0 9108 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8096 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_74
timestamp 1606256979
transform 1 0 7912 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1606256979
transform 1 0 8924 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1606256979
transform 1 0 9660 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1606256979
transform 1 0 10304 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606256979
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1606256979
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_97
timestamp 1606256979
transform 1 0 10028 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606256979
transform 1 0 12328 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 12880 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_28_116
timestamp 1606256979
transform 1 0 11776 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_126
timestamp 1606256979
transform 1 0 12696 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606256979
transform 1 0 14628 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_144
timestamp 1606256979
transform 1 0 14352 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1606256979
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1606256979
transform 1 0 16928 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15272 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606256979
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_170
timestamp 1606256979
transform 1 0 16744 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1606256979
transform 1 0 19044 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606256979
transform 1 0 17388 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_175
timestamp 1606256979
transform 1 0 17204 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_193
timestamp 1606256979
transform 1 0 18860 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606256979
transform 1 0 20240 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 20884 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606256979
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_204
timestamp 1606256979
transform 1 0 19872 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1606256979
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1606256979
transform 1 0 22540 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606256979
transform -1 0 23276 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_231
timestamp 1606256979
transform 1 0 22356 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_236
timestamp 1606256979
transform 1 0 22816 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2300 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606256979
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606256979
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1606256979
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1606256979
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1606256979
transform 1 0 3956 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4508 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_29
timestamp 1606256979
transform 1 0 3772 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_35
timestamp 1606256979
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _62_
timestamp 1606256979
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606256979
transform 1 0 6164 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606256979
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1606256979
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1606256979
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_65
timestamp 1606256979
transform 1 0 7084 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8280 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 7268 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_76
timestamp 1606256979
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1606256979
transform 1 0 10212 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 9936 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_94
timestamp 1606256979
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _61_
timestamp 1606256979
transform 1 0 11868 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606256979
transform 1 0 12420 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606256979
transform 1 0 12972 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606256979
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_115
timestamp 1606256979
transform 1 0 11684 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1606256979
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_127
timestamp 1606256979
transform 1 0 12788 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1606256979
transform 1 0 14628 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_145
timestamp 1606256979
transform 1 0 14444 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16652 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1606256979
transform 1 0 15640 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_156
timestamp 1606256979
transform 1 0 15456 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_167
timestamp 1606256979
transform 1 0 16468 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1606256979
transform 1 0 18032 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606256979
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_178
timestamp 1606256979
transform 1 0 17480 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606256979
transform 1 0 19780 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 20332 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_29_200
timestamp 1606256979
transform 1 0 19504 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_207
timestamp 1606256979
transform 1 0 20148 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_218
timestamp 1606256979
transform 1 0 21160 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 21344 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606256979
transform -1 0 23276 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_236
timestamp 1606256979
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606256979
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 2300 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606256979
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1606256979
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1606256979
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1606256979
transform 1 0 5060 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606256979
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1606256979
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_41
timestamp 1606256979
transform 1 0 4876 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1606256979
transform 1 0 6808 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606256979
transform 1 0 6256 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_52
timestamp 1606256979
transform 1 0 5888 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_60
timestamp 1606256979
transform 1 0 6624 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1606256979
transform 1 0 7912 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_30_71
timestamp 1606256979
transform 1 0 7636 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606256979
transform 1 0 9660 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1606256979
transform 1 0 10212 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606256979
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1606256979
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_97
timestamp 1606256979
transform 1 0 10028 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 11868 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_115
timestamp 1606256979
transform 1 0 11684 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1606256979
transform 1 0 14628 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13524 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_133
timestamp 1606256979
transform 1 0 13340 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_144
timestamp 1606256979
transform 1 0 14352 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1606256979
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1606256979
transform 1 0 17020 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15364 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606256979
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_154
timestamp 1606256979
transform 1 0 15272 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_171
timestamp 1606256979
transform 1 0 16836 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1606256979
transform 1 0 19136 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1606256979
transform 1 0 17480 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_176
timestamp 1606256979
transform 1 0 17296 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1606256979
transform 1 0 18952 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1606256979
transform 1 0 20148 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606256979
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_205
timestamp 1606256979
transform 1 0 19964 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_211
timestamp 1606256979
transform 1 0 20516 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606256979
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1606256979
transform 1 0 21252 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606256979
transform -1 0 23276 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_235
timestamp 1606256979
transform 1 0 22724 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 1380 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1606256979
transform 1 0 3036 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606256979
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_19
timestamp 1606256979
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1606256979
transform 1 0 4692 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_37
timestamp 1606256979
transform 1 0 4508 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5704 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606256979
transform 1 0 6992 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606256979
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_48
timestamp 1606256979
transform 1 0 5520 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1606256979
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1606256979
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1606256979
transform 1 0 7544 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1606256979
transform 1 0 8556 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_68
timestamp 1606256979
transform 1 0 7360 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_79
timestamp 1606256979
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1606256979
transform 1 0 10304 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_31_97
timestamp 1606256979
transform 1 0 10028 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_109
timestamp 1606256979
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1606256979
transform 1 0 11316 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606256979
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1606256979
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1606256979
transform 1 0 13708 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1606256979
transform 1 0 14260 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_31_132
timestamp 1606256979
transform 1 0 13248 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_136
timestamp 1606256979
transform 1 0 13616 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_141
timestamp 1606256979
transform 1 0 14076 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_152
timestamp 1606256979
transform 1 0 15088 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1606256979
transform 1 0 15272 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1606256979
transform 1 0 16284 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_163
timestamp 1606256979
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_174
timestamp 1606256979
transform 1 0 17112 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1606256979
transform 1 0 17388 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1606256979
transform 1 0 18032 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606256979
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1606256979
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 19688 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1606256979
transform 1 0 20976 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_200
timestamp 1606256979
transform 1 0 19504 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_211
timestamp 1606256979
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_215
timestamp 1606256979
transform 1 0 20884 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606256979
transform -1 0 23276 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_232
timestamp 1606256979
transform 1 0 22448 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1606256979
transform 1 0 3036 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 1380 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606256979
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_19
timestamp 1606256979
transform 1 0 2852 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1606256979
transform 1 0 4416 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606256979
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_25
timestamp 1606256979
transform 1 0 3404 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_32
timestamp 1606256979
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1606256979
transform 1 0 6164 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_32_52
timestamp 1606256979
transform 1 0 5888 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_64
timestamp 1606256979
transform 1 0 6992 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606256979
transform 1 0 7360 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1606256979
transform 1 0 7912 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_72
timestamp 1606256979
transform 1 0 7728 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1606256979
transform 1 0 9660 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1606256979
transform 1 0 10396 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1606256979
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_90
timestamp 1606256979
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_98
timestamp 1606256979
transform 1 0 10120 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1606256979
transform 1 0 12052 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_117
timestamp 1606256979
transform 1 0 11868 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _63_
timestamp 1606256979
transform 1 0 14720 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1606256979
transform 1 0 13524 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1606256979
transform 1 0 14536 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_144
timestamp 1606256979
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_151
timestamp 1606256979
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1606256979
transform 1 0 17020 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15364 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1606256979
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_154
timestamp 1606256979
transform 1 0 15272 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_171
timestamp 1606256979
transform 1 0 16836 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1606256979
transform 1 0 17756 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_32_178
timestamp 1606256979
transform 1 0 17480 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1606256979
transform 1 0 19412 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1606256979
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1606256979
transform 1 0 19228 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_208
timestamp 1606256979
transform 1 0 20240 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_215
timestamp 1606256979
transform 1 0 20884 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1606256979
transform 1 0 21252 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1606256979
transform 1 0 22264 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606256979
transform -1 0 23276 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_228
timestamp 1606256979
transform 1 0 22080 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_235
timestamp 1606256979
transform 1 0 22724 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1606256979
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606256979
transform 1 0 1656 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1606256979
transform 1 0 1932 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1606256979
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1606256979
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_3
timestamp 1606256979
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_7
timestamp 1606256979
transform 1 0 1748 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1606256979
transform 1 0 5060 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1606256979
transform 1 0 4048 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1606256979
transform 1 0 3404 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1606256979
transform 1 0 5060 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1606256979
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_22
timestamp 1606256979
transform 1 0 3128 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_41
timestamp 1606256979
transform 1 0 4876 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_25
timestamp 1606256979
transform 1 0 3404 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_41
timestamp 1606256979
transform 1 0 4876 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1606256979
transform 1 0 5796 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1606256979
transform 1 0 6808 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1606256979
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1606256979
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1606256979
transform 1 0 5428 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1606256979
transform 1 0 7544 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1606256979
transform 1 0 8464 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_33_78
timestamp 1606256979
transform 1 0 8280 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_67
timestamp 1606256979
transform 1 0 7268 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_86
timestamp 1606256979
transform 1 0 9016 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1606256979
transform 1 0 9660 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1606256979
transform 1 0 11040 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1606256979
transform 1 0 10396 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1606256979
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_96
timestamp 1606256979
transform 1 0 9936 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_100
timestamp 1606256979
transform 1 0 10304 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_102
timestamp 1606256979
transform 1 0 10488 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1606256979
transform 1 0 12696 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1606256979
transform 1 0 13064 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1606256979
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_117
timestamp 1606256979
transform 1 0 11868 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1606256979
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_123
timestamp 1606256979
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_130
timestamp 1606256979
transform 1 0 13064 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_124
timestamp 1606256979
transform 1 0 12512 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1606256979
transform 1 0 13248 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1606256979
transform 1 0 14904 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_33_148
timestamp 1606256979
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_146
timestamp 1606256979
transform 1 0 14536 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_152
timestamp 1606256979
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1606256979
transform 1 0 16928 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1606256979
transform 1 0 16560 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1606256979
transform 1 0 15272 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1606256979
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1606256979
transform 1 0 16376 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_170
timestamp 1606256979
transform 1 0 16744 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1606256979
transform 1 0 17480 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1606256979
transform 1 0 19136 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1606256979
transform 1 0 18032 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1606256979
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_177
timestamp 1606256979
transform 1 0 17388 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_176
timestamp 1606256979
transform 1 0 17296 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1606256979
transform 1 0 18952 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1606256979
transform 1 0 19688 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1606256979
transform 1 0 20884 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1606256979
transform 1 0 20792 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1606256979
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_200
timestamp 1606256979
transform 1 0 19504 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_211
timestamp 1606256979
transform 1 0 20516 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1606256979
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606256979
transform 1 0 22448 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1606256979
transform -1 0 23276 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1606256979
transform -1 0 23276 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_230
timestamp 1606256979
transform 1 0 22264 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_236
timestamp 1606256979
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_231
timestamp 1606256979
transform 1 0 22356 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_237
timestamp 1606256979
transform 1 0 22908 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1606256979
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1606256979
transform 1 0 2944 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 1932 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1606256979
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_7
timestamp 1606256979
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_18
timestamp 1606256979
transform 1 0 2760 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1606256979
transform 1 0 5060 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1606256979
transform 1 0 4048 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1606256979
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_29
timestamp 1606256979
transform 1 0 3772 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_41
timestamp 1606256979
transform 1 0 4876 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1606256979
transform 1 0 5796 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1606256979
transform 1 0 6900 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1606256979
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_47
timestamp 1606256979
transform 1 0 5428 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_60
timestamp 1606256979
transform 1 0 6624 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _53_
timestamp 1606256979
transform 1 0 7912 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1606256979
transform 1 0 8372 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_35_72
timestamp 1606256979
transform 1 0 7728 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_77
timestamp 1606256979
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1606256979
transform 1 0 9752 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1606256979
transform 1 0 10672 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1606256979
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_88
timestamp 1606256979
transform 1 0 9200 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_92
timestamp 1606256979
transform 1 0 9568 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_98
timestamp 1606256979
transform 1 0 10120 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1606256979
transform 1 0 12604 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1606256979
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_120
timestamp 1606256979
transform 1 0 12144 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1606256979
transform 1 0 14812 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1606256979
transform 1 0 13616 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_35_134
timestamp 1606256979
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_145
timestamp 1606256979
transform 1 0 14444 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1606256979
transform 1 0 15456 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16468 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1606256979
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_153
timestamp 1606256979
transform 1 0 15180 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_165
timestamp 1606256979
transform 1 0 16284 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1606256979
transform 1 0 17664 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1606256979
transform 1 0 18308 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1606256979
transform 1 0 18860 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1606256979
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_176
timestamp 1606256979
transform 1 0 17296 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_184
timestamp 1606256979
transform 1 0 18032 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_191
timestamp 1606256979
transform 1 0 18676 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1606256979
transform 1 0 21160 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1606256979
transform 1 0 20516 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1606256979
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_209
timestamp 1606256979
transform 1 0 20332 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_215
timestamp 1606256979
transform 1 0 20884 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606256979
transform 1 0 22172 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1606256979
transform -1 0 23276 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_227
timestamp 1606256979
transform 1 0 21988 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_233
timestamp 1606256979
transform 1 0 22540 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_237
timestamp 1606256979
transform 1 0 22908 0 1 21216
box -38 -48 130 592
<< labels >>
rlabel metal2 s 8574 0 8630 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 16946 23920 17002 24400 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 12070 0 12126 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 17590 23920 17646 24400 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal3 s 23920 6808 24400 6928 6 Test_en_E_in
port 4 nsew default input
rlabel metal3 s 23920 6128 24400 6248 6 Test_en_E_out
port 5 nsew default tristate
rlabel metal3 s 0 21224 480 21344 6 Test_en_W_in
port 6 nsew default input
rlabel metal3 s 0 15104 480 15224 6 Test_en_W_out
port 7 nsew default tristate
rlabel metal2 s 1674 0 1730 480 6 bottom_width_0_height_0__pin_50_
port 8 nsew default tristate
rlabel metal2 s 5078 0 5134 480 6 bottom_width_0_height_0__pin_51_
port 9 nsew default tristate
rlabel metal3 s 0 8984 480 9104 6 ccff_head
port 10 nsew default input
rlabel metal3 s 23920 5448 24400 5568 6 ccff_tail
port 11 nsew default tristate
rlabel metal2 s 18234 23920 18290 24400 6 clk_0_N_in
port 12 nsew default input
rlabel metal2 s 15566 0 15622 480 6 clk_0_S_in
port 13 nsew default input
rlabel metal3 s 23920 8168 24400 8288 6 prog_clk_0_E_out
port 14 nsew default tristate
rlabel metal3 s 23920 7488 24400 7608 6 prog_clk_0_N_in
port 15 nsew default input
rlabel metal2 s 18878 23920 18934 24400 6 prog_clk_0_N_out
port 16 nsew default tristate
rlabel metal2 s 19062 0 19118 480 6 prog_clk_0_S_in
port 17 nsew default input
rlabel metal2 s 22558 0 22614 480 6 prog_clk_0_S_out
port 18 nsew default tristate
rlabel metal3 s 0 3000 480 3120 6 prog_clk_0_W_out
port 19 nsew default tristate
rlabel metal3 s 23920 8712 24400 8832 6 right_width_0_height_0__pin_16_
port 20 nsew default input
rlabel metal3 s 23920 9392 24400 9512 6 right_width_0_height_0__pin_17_
port 21 nsew default input
rlabel metal3 s 23920 10072 24400 10192 6 right_width_0_height_0__pin_18_
port 22 nsew default input
rlabel metal3 s 23920 10752 24400 10872 6 right_width_0_height_0__pin_19_
port 23 nsew default input
rlabel metal3 s 23920 11432 24400 11552 6 right_width_0_height_0__pin_20_
port 24 nsew default input
rlabel metal3 s 23920 12112 24400 12232 6 right_width_0_height_0__pin_21_
port 25 nsew default input
rlabel metal3 s 23920 12656 24400 12776 6 right_width_0_height_0__pin_22_
port 26 nsew default input
rlabel metal3 s 23920 13336 24400 13456 6 right_width_0_height_0__pin_23_
port 27 nsew default input
rlabel metal3 s 23920 14016 24400 14136 6 right_width_0_height_0__pin_24_
port 28 nsew default input
rlabel metal3 s 23920 14696 24400 14816 6 right_width_0_height_0__pin_25_
port 29 nsew default input
rlabel metal3 s 23920 15376 24400 15496 6 right_width_0_height_0__pin_26_
port 30 nsew default input
rlabel metal3 s 23920 16056 24400 16176 6 right_width_0_height_0__pin_27_
port 31 nsew default input
rlabel metal3 s 23920 16600 24400 16720 6 right_width_0_height_0__pin_28_
port 32 nsew default input
rlabel metal3 s 23920 17280 24400 17400 6 right_width_0_height_0__pin_29_
port 33 nsew default input
rlabel metal3 s 23920 17960 24400 18080 6 right_width_0_height_0__pin_30_
port 34 nsew default input
rlabel metal3 s 23920 18640 24400 18760 6 right_width_0_height_0__pin_31_
port 35 nsew default input
rlabel metal3 s 23920 280 24400 400 6 right_width_0_height_0__pin_42_lower
port 36 nsew default tristate
rlabel metal3 s 23920 19320 24400 19440 6 right_width_0_height_0__pin_42_upper
port 37 nsew default tristate
rlabel metal3 s 23920 824 24400 944 6 right_width_0_height_0__pin_43_lower
port 38 nsew default tristate
rlabel metal3 s 23920 20000 24400 20120 6 right_width_0_height_0__pin_43_upper
port 39 nsew default tristate
rlabel metal3 s 23920 1504 24400 1624 6 right_width_0_height_0__pin_44_lower
port 40 nsew default tristate
rlabel metal3 s 23920 20544 24400 20664 6 right_width_0_height_0__pin_44_upper
port 41 nsew default tristate
rlabel metal3 s 23920 2184 24400 2304 6 right_width_0_height_0__pin_45_lower
port 42 nsew default tristate
rlabel metal3 s 23920 21224 24400 21344 6 right_width_0_height_0__pin_45_upper
port 43 nsew default tristate
rlabel metal3 s 23920 2864 24400 2984 6 right_width_0_height_0__pin_46_lower
port 44 nsew default tristate
rlabel metal3 s 23920 21904 24400 22024 6 right_width_0_height_0__pin_46_upper
port 45 nsew default tristate
rlabel metal3 s 23920 3544 24400 3664 6 right_width_0_height_0__pin_47_lower
port 46 nsew default tristate
rlabel metal3 s 23920 22584 24400 22704 6 right_width_0_height_0__pin_47_upper
port 47 nsew default tristate
rlabel metal3 s 23920 4224 24400 4344 6 right_width_0_height_0__pin_48_lower
port 48 nsew default tristate
rlabel metal3 s 23920 23264 24400 23384 6 right_width_0_height_0__pin_48_upper
port 49 nsew default tristate
rlabel metal3 s 23920 4768 24400 4888 6 right_width_0_height_0__pin_49_lower
port 50 nsew default tristate
rlabel metal3 s 23920 23944 24400 24064 6 right_width_0_height_0__pin_49_upper
port 51 nsew default tristate
rlabel metal2 s 5354 23920 5410 24400 6 top_width_0_height_0__pin_0_
port 52 nsew default input
rlabel metal2 s 11794 23920 11850 24400 6 top_width_0_height_0__pin_10_
port 53 nsew default input
rlabel metal2 s 12438 23920 12494 24400 6 top_width_0_height_0__pin_11_
port 54 nsew default input
rlabel metal2 s 13082 23920 13138 24400 6 top_width_0_height_0__pin_12_
port 55 nsew default input
rlabel metal2 s 13726 23920 13782 24400 6 top_width_0_height_0__pin_13_
port 56 nsew default input
rlabel metal2 s 14370 23920 14426 24400 6 top_width_0_height_0__pin_14_
port 57 nsew default input
rlabel metal2 s 15014 23920 15070 24400 6 top_width_0_height_0__pin_15_
port 58 nsew default input
rlabel metal2 s 5998 23920 6054 24400 6 top_width_0_height_0__pin_1_
port 59 nsew default input
rlabel metal2 s 6642 23920 6698 24400 6 top_width_0_height_0__pin_2_
port 60 nsew default input
rlabel metal2 s 15658 23920 15714 24400 6 top_width_0_height_0__pin_32_
port 61 nsew default input
rlabel metal2 s 16302 23920 16358 24400 6 top_width_0_height_0__pin_33_
port 62 nsew default input
rlabel metal2 s 19522 23920 19578 24400 6 top_width_0_height_0__pin_34_lower
port 63 nsew default tristate
rlabel metal2 s 294 23920 350 24400 6 top_width_0_height_0__pin_34_upper
port 64 nsew default tristate
rlabel metal2 s 20166 23920 20222 24400 6 top_width_0_height_0__pin_35_lower
port 65 nsew default tristate
rlabel metal2 s 846 23920 902 24400 6 top_width_0_height_0__pin_35_upper
port 66 nsew default tristate
rlabel metal2 s 20810 23920 20866 24400 6 top_width_0_height_0__pin_36_lower
port 67 nsew default tristate
rlabel metal2 s 1490 23920 1546 24400 6 top_width_0_height_0__pin_36_upper
port 68 nsew default tristate
rlabel metal2 s 21454 23920 21510 24400 6 top_width_0_height_0__pin_37_lower
port 69 nsew default tristate
rlabel metal2 s 2134 23920 2190 24400 6 top_width_0_height_0__pin_37_upper
port 70 nsew default tristate
rlabel metal2 s 22098 23920 22154 24400 6 top_width_0_height_0__pin_38_lower
port 71 nsew default tristate
rlabel metal2 s 2778 23920 2834 24400 6 top_width_0_height_0__pin_38_upper
port 72 nsew default tristate
rlabel metal2 s 22742 23920 22798 24400 6 top_width_0_height_0__pin_39_lower
port 73 nsew default tristate
rlabel metal2 s 3422 23920 3478 24400 6 top_width_0_height_0__pin_39_upper
port 74 nsew default tristate
rlabel metal2 s 7286 23920 7342 24400 6 top_width_0_height_0__pin_3_
port 75 nsew default input
rlabel metal2 s 23386 23920 23442 24400 6 top_width_0_height_0__pin_40_lower
port 76 nsew default tristate
rlabel metal2 s 4066 23920 4122 24400 6 top_width_0_height_0__pin_40_upper
port 77 nsew default tristate
rlabel metal2 s 24030 23920 24086 24400 6 top_width_0_height_0__pin_41_lower
port 78 nsew default tristate
rlabel metal2 s 4710 23920 4766 24400 6 top_width_0_height_0__pin_41_upper
port 79 nsew default tristate
rlabel metal2 s 7930 23920 7986 24400 6 top_width_0_height_0__pin_4_
port 80 nsew default input
rlabel metal2 s 8574 23920 8630 24400 6 top_width_0_height_0__pin_5_
port 81 nsew default input
rlabel metal2 s 9218 23920 9274 24400 6 top_width_0_height_0__pin_6_
port 82 nsew default input
rlabel metal2 s 9862 23920 9918 24400 6 top_width_0_height_0__pin_7_
port 83 nsew default input
rlabel metal2 s 10506 23920 10562 24400 6 top_width_0_height_0__pin_8_
port 84 nsew default input
rlabel metal2 s 11150 23920 11206 24400 6 top_width_0_height_0__pin_9_
port 85 nsew default input
rlabel metal4 s 4643 2128 4963 21808 6 VPWR
port 86 nsew default input
rlabel metal4 s 8341 2128 8661 21808 6 VGND
port 87 nsew default input
<< properties >>
string FIXED_BBOX 0 0 24400 24400
<< end >>
