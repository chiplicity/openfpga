* NGSPICE file created from sb_3__3_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

.subckt sb_3__3_ address[0] address[1] address[2] address[3] address[4] address[5]
+ bottom_left_grid_pin_13_ bottom_right_grid_pin_11_ bottom_right_grid_pin_13_ bottom_right_grid_pin_15_
+ bottom_right_grid_pin_1_ bottom_right_grid_pin_3_ bottom_right_grid_pin_5_ bottom_right_grid_pin_7_
+ bottom_right_grid_pin_9_ chanx_left_in[0] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_out[0] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4]
+ chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chany_bottom_in[0]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_out[0] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] data_in enable left_bottom_grid_pin_12_
+ left_top_grid_pin_11_ left_top_grid_pin_13_ left_top_grid_pin_15_ left_top_grid_pin_1_
+ left_top_grid_pin_3_ left_top_grid_pin_5_ left_top_grid_pin_7_ left_top_grid_pin_9_
+ vpwr vgnd
XFILLER_22_166 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_41 vgnd vpwr scs8hd_decap_12
XFILLER_13_177 vgnd vpwr scs8hd_fill_1
XFILLER_13_144 vgnd vpwr scs8hd_fill_1
XFILLER_3_12 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _35_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_86 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_49_ _49_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _49_/A vgnd vpwr scs8hd_inv_1
XFILLER_29_63 vgnd vpwr scs8hd_fill_1
Xmux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _33_/HI mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_161 vgnd vpwr scs8hd_fill_1
XFILLER_25_175 vgnd vpwr scs8hd_decap_3
XFILLER_25_131 vgnd vpwr scs8hd_decap_4
XFILLER_15_98 vgnd vpwr scs8hd_decap_12
XFILLER_16_175 vgnd vpwr scs8hd_decap_3
XFILLER_13_123 vgnd vpwr scs8hd_decap_12
XFILLER_3_24 vgnd vpwr scs8hd_decap_12
XFILLER_9_149 vgnd vpwr scs8hd_decap_12
Xmux_left_track_13.tap_buf4_0_.scs8hd_inv_1 mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _38_/A vgnd vpwr scs8hd_inv_1
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XFILLER_12_11 vgnd vpwr scs8hd_decap_4
XFILLER_5_130 vgnd vpwr scs8hd_decap_12
XFILLER_23_21 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_23_65 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_48_ _48_/A chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
Xmux_left_track_5.tap_buf4_0_.scs8hd_inv_1 mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _42_/A vgnd vpwr scs8hd_inv_1
XFILLER_20_11 vgnd vpwr scs8hd_decap_4
XFILLER_1_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_173 vgnd vpwr scs8hd_decap_4
XFILLER_19_151 vgnd vpwr scs8hd_decap_3
XFILLER_25_154 vpwr vgnd scs8hd_fill_2
XFILLER_25_121 vgnd vpwr scs8hd_fill_1
XFILLER_25_110 vgnd vpwr scs8hd_decap_3
XFILLER_16_154 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_12_ mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_32 vpwr vgnd scs8hd_fill_2
XFILLER_13_135 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _45_/A vgnd vpwr scs8hd_inv_1
Xmux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_36 vgnd vpwr scs8hd_decap_12
XFILLER_12_56 vgnd vpwr scs8hd_decap_12
XFILLER_10_105 vgnd vpwr scs8hd_decap_12
XFILLER_5_142 vgnd vpwr scs8hd_decap_12
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
X_47_ _47_/A chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_29_10 vgnd vpwr scs8hd_decap_4
XFILLER_29_21 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_3_48 vgnd vpwr scs8hd_decap_12
XFILLER_8_140 vgnd vpwr scs8hd_decap_12
XFILLER_12_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_15_ mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_117 vpwr vgnd scs8hd_fill_2
XFILLER_5_121 vgnd vpwr scs8hd_fill_1
XFILLER_5_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_56 vgnd vpwr scs8hd_decap_4
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XFILLER_2_102 vgnd vpwr scs8hd_decap_8
X_46_ _46_/A chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_18_89 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
X_29_ _29_/HI _29_/LO vgnd vpwr scs8hd_conb_1
XFILLER_29_99 vgnd vpwr scs8hd_decap_8
XFILLER_20_35 vgnd vpwr scs8hd_decap_12
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XFILLER_6_59 vgnd vpwr scs8hd_decap_12
XFILLER_19_164 vgnd vpwr scs8hd_fill_1
XFILLER_20_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_25_167 vgnd vpwr scs8hd_decap_8
XFILLER_25_123 vgnd vpwr scs8hd_fill_1
XFILLER_15_46 vgnd vpwr scs8hd_decap_12
Xmux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _32_/HI mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_16_167 vgnd vpwr scs8hd_decap_8
XFILLER_11_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_148 vgnd vpwr scs8hd_decap_6
XFILLER_12_170 vgnd vpwr scs8hd_decap_8
XFILLER_8_152 vgnd vpwr scs8hd_fill_1
XFILLER_5_166 vgnd vpwr scs8hd_decap_12
Xmux_left_track_13.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_13_ mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_35 vgnd vpwr scs8hd_decap_6
XFILLER_9_15 vpwr vgnd scs8hd_fill_2
X_45_ _45_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[3] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_57 vgnd vpwr scs8hd_decap_12
XFILLER_18_46 vgnd vpwr scs8hd_decap_8
XFILLER_18_35 vgnd vpwr scs8hd_decap_8
XFILLER_18_13 vpwr vgnd scs8hd_fill_2
X_28_ _28_/HI _28_/LO vgnd vpwr scs8hd_conb_1
XFILLER_29_78 vpwr vgnd scs8hd_fill_2
XFILLER_29_67 vgnd vpwr scs8hd_decap_8
XFILLER_28_154 vgnd vpwr scs8hd_fill_1
XFILLER_28_121 vgnd vpwr scs8hd_decap_8
XFILLER_20_47 vgnd vpwr scs8hd_decap_12
XFILLER_19_143 vgnd vpwr scs8hd_decap_8
XFILLER_19_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _28_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_10_80 vgnd vpwr scs8hd_decap_12
XFILLER_15_58 vgnd vpwr scs8hd_decap_3
XFILLER_15_14 vpwr vgnd scs8hd_fill_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_90 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_26_57 vgnd vpwr scs8hd_decap_12
XFILLER_21_171 vgnd vpwr scs8hd_decap_6
XFILLER_5_123 vgnd vpwr scs8hd_decap_4
Xmux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_44_ _44_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_18_69 vgnd vpwr scs8hd_decap_12
XFILLER_1_3 vpwr vgnd scs8hd_fill_2
X_27_ _27_/HI _27_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_94 vpwr vgnd scs8hd_fill_2
XFILLER_1_83 vpwr vgnd scs8hd_fill_2
Xmux_left_track_11.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_11_ mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_46 vpwr vgnd scs8hd_fill_2
XFILLER_29_35 vgnd vpwr scs8hd_decap_8
XFILLER_28_177 vgnd vpwr scs8hd_fill_1
Xmux_left_track_7.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[2] mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_59 vgnd vpwr scs8hd_decap_12
XFILLER_19_177 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_103 vpwr vgnd scs8hd_fill_2
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_117 vgnd vpwr scs8hd_decap_12
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_26_69 vgnd vpwr scs8hd_decap_6
XFILLER_26_36 vgnd vpwr scs8hd_fill_1
XFILLER_16_80 vgnd vpwr scs8hd_decap_12
XFILLER_8_154 vgnd vpwr scs8hd_decap_12
XANTENNA__42__A _42_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_113 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__37__A _37_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_39 vgnd vpwr scs8hd_decap_3
XFILLER_29_6 vpwr vgnd scs8hd_fill_2
X_43_ _43_/A chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_1_171 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_3 vpwr vgnd scs8hd_fill_2
XFILLER_28_101 vgnd vpwr scs8hd_decap_8
X_26_ _26_/HI _26_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_73 vgnd vpwr scs8hd_fill_1
XFILLER_1_62 vgnd vpwr scs8hd_decap_3
XANTENNA__50__A _50_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_93 vgnd vpwr scs8hd_decap_12
XFILLER_25_137 vgnd vpwr scs8hd_decap_12
XFILLER_25_115 vgnd vpwr scs8hd_decap_6
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__45__A _45_/A vgnd vpwr scs8hd_diode_2
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_129 vgnd vpwr scs8hd_decap_12
XPHY_1 vgnd vpwr scs8hd_decap_3
Xmux_left_track_5.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_94 vgnd vpwr scs8hd_decap_12
XFILLER_8_166 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _27_/HI mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _51_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__53__A _53_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_150 vgnd vpwr scs8hd_decap_4
X_42_ _42_/A chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__48__A _48_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_81 vgnd vpwr scs8hd_decap_8
XFILLER_24_70 vpwr vgnd scs8hd_fill_2
X_25_ _25_/HI _25_/LO vgnd vpwr scs8hd_conb_1
XFILLER_28_135 vgnd vpwr scs8hd_decap_12
XFILLER_19_157 vgnd vpwr scs8hd_decap_4
XFILLER_19_135 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_149 vgnd vpwr scs8hd_decap_3
XFILLER_25_127 vpwr vgnd scs8hd_fill_2
XFILLER_16_105 vgnd vpwr scs8hd_decap_12
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XFILLER_16_93 vgnd vpwr scs8hd_decap_12
XFILLER_12_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_18 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_15.INVTX1_1_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _44_/A vgnd vpwr scs8hd_inv_1
XFILLER_27_92 vgnd vpwr scs8hd_decap_4
XFILLER_4_96 vgnd vpwr scs8hd_decap_8
XFILLER_23_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_41_ _41_/A chanx_left_out[3] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_9_ mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_19 vgnd vpwr scs8hd_decap_12
XFILLER_18_17 vgnd vpwr scs8hd_decap_12
XFILLER_24_93 vgnd vpwr scs8hd_decap_8
Xmux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_18 vgnd vpwr scs8hd_decap_12
XFILLER_1_31 vgnd vpwr scs8hd_decap_12
X_24_ _24_/HI _24_/LO vgnd vpwr scs8hd_conb_1
XFILLER_28_169 vgnd vpwr scs8hd_decap_8
XFILLER_28_158 vgnd vpwr scs8hd_decap_8
XFILLER_28_147 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _29_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_169 vpwr vgnd scs8hd_fill_2
XFILLER_15_18 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _47_/A vgnd vpwr scs8hd_inv_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_117 vgnd vpwr scs8hd_decap_12
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_5_105 vpwr vgnd scs8hd_fill_2
XFILLER_5_127 vgnd vpwr scs8hd_fill_1
XFILLER_2_119 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[8] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_40_ _40_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_13_62 vgnd vpwr scs8hd_decap_12
XFILLER_13_51 vgnd vpwr scs8hd_decap_8
XFILLER_18_29 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.INVTX1_1_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_7 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_7_ mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_23_ _23_/HI _23_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_43 vgnd vpwr scs8hd_decap_12
XFILLER_29_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_3 vpwr vgnd scs8hd_fill_2
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_62 vpwr vgnd scs8hd_fill_2
XFILLER_21_51 vpwr vgnd scs8hd_fill_2
XFILLER_21_40 vgnd vpwr scs8hd_decap_4
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_129 vgnd vpwr scs8hd_decap_12
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_151 vpwr vgnd scs8hd_fill_2
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_12_154 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _22_/HI mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XFILLER_4_150 vgnd vpwr scs8hd_decap_3
XFILLER_13_74 vgnd vpwr scs8hd_decap_12
X_22_ _22_/HI _22_/LO vgnd vpwr scs8hd_conb_1
XFILLER_27_7 vpwr vgnd scs8hd_fill_2
XFILLER_24_62 vgnd vpwr scs8hd_decap_8
XFILLER_1_55 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_29 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_11.INVTX1_1_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_19_62 vgnd vpwr scs8hd_decap_12
XFILLER_19_51 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_20 vgnd vpwr scs8hd_decap_8
XFILLER_18_3 vpwr vgnd scs8hd_fill_2
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_152 vgnd vpwr scs8hd_fill_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_5.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_5_ mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_7_10 vpwr vgnd scs8hd_fill_2
XFILLER_21_177 vgnd vpwr scs8hd_fill_1
XFILLER_16_30 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _18_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_86 vgnd vpwr scs8hd_decap_12
X_21_ _21_/HI _21_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_67 vgnd vpwr scs8hd_decap_6
XFILLER_19_139 vpwr vgnd scs8hd_fill_2
XFILLER_19_74 vgnd vpwr scs8hd_decap_12
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_7_77 vgnd vpwr scs8hd_decap_6
XFILLER_21_123 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_3.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_3_ mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_105 vgnd vpwr scs8hd_decap_12
XFILLER_27_41 vgnd vpwr scs8hd_decap_8
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_98 vgnd vpwr scs8hd_decap_12
XFILLER_1_177 vgnd vpwr scs8hd_fill_1
XFILLER_1_133 vgnd vpwr scs8hd_decap_4
XFILLER_8_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_79 vpwr vgnd scs8hd_fill_2
X_20_ _20_/HI _20_/LO vgnd vpwr scs8hd_conb_1
XFILLER_28_129 vpwr vgnd scs8hd_fill_2
XFILLER_19_42 vgnd vpwr scs8hd_fill_1
XFILLER_10_44 vgnd vpwr scs8hd_decap_12
XFILLER_27_173 vgnd vpwr scs8hd_decap_4
XFILLER_27_162 vgnd vpwr scs8hd_fill_1
XFILLER_19_86 vgnd vpwr scs8hd_decap_12
XFILLER_24_110 vgnd vpwr scs8hd_decap_12
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _30_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_176 vpwr vgnd scs8hd_fill_2
XFILLER_24_154 vgnd vpwr scs8hd_decap_4
XFILLER_21_10 vpwr vgnd scs8hd_fill_2
XFILLER_15_176 vpwr vgnd scs8hd_fill_2
XFILLER_15_143 vgnd vpwr scs8hd_fill_1
XFILLER_15_110 vgnd vpwr scs8hd_decap_12
XPHY_7 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_3 vgnd vpwr scs8hd_decap_3
XFILLER_21_135 vgnd vpwr scs8hd_decap_12
XFILLER_21_102 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XFILLER_8_117 vgnd vpwr scs8hd_decap_3
XFILLER_5_109 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_1_ mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_75 vpwr vgnd scs8hd_fill_2
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XFILLER_27_20 vpwr vgnd scs8hd_fill_2
XFILLER_4_68 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _21_/HI mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_1_167 vpwr vgnd scs8hd_fill_2
XFILLER_1_156 vpwr vgnd scs8hd_fill_2
XFILLER_1_123 vgnd vpwr scs8hd_fill_1
XFILLER_1_112 vgnd vpwr scs8hd_decap_8
XFILLER_10_56 vgnd vpwr scs8hd_decap_12
XFILLER_19_98 vgnd vpwr scs8hd_decap_12
XFILLER_19_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_163 vgnd vpwr scs8hd_decap_12
XFILLER_18_141 vgnd vpwr scs8hd_decap_12
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_122 vgnd vpwr scs8hd_decap_12
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_66 vgnd vpwr scs8hd_decap_12
XFILLER_21_55 vgnd vpwr scs8hd_decap_6
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _53_/A vgnd vpwr scs8hd_inv_1
XFILLER_16_3 vpwr vgnd scs8hd_fill_2
XFILLER_15_155 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_46 vgnd vpwr scs8hd_fill_1
XFILLER_21_147 vgnd vpwr scs8hd_decap_12
XFILLER_21_114 vgnd vpwr scs8hd_decap_8
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XFILLER_12_158 vgnd vpwr scs8hd_decap_3
XFILLER_8_129 vgnd vpwr scs8hd_decap_8
XFILLER_7_151 vgnd vpwr scs8hd_decap_12
XFILLER_27_98 vpwr vgnd scs8hd_fill_2
XFILLER_4_154 vgnd vpwr scs8hd_decap_12
Xmux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_23 vpwr vgnd scs8hd_fill_2
XFILLER_13_12 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_109 vgnd vpwr scs8hd_decap_3
XFILLER_10_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_175 vgnd vpwr scs8hd_decap_3
XFILLER_18_7 vpwr vgnd scs8hd_fill_2
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_134 vgnd vpwr scs8hd_decap_12
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_78 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_14 vgnd vpwr scs8hd_decap_12
XFILLER_21_159 vgnd vpwr scs8hd_decap_12
XFILLER_16_56 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[7] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_163 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _23_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_89 vgnd vpwr scs8hd_decap_3
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XFILLER_27_121 vgnd vpwr scs8hd_fill_1
XFILLER_19_34 vpwr vgnd scs8hd_fill_2
XFILLER_19_23 vgnd vpwr scs8hd_decap_8
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_15.tap_buf4_0_.scs8hd_inv_1 mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _37_/A vgnd vpwr scs8hd_inv_1
XFILLER_24_168 vgnd vpwr scs8hd_decap_8
XFILLER_24_146 vgnd vpwr scs8hd_decap_6
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_168 vgnd vpwr scs8hd_decap_8
XFILLER_15_135 vgnd vpwr scs8hd_decap_8
XFILLER_7_26 vgnd vpwr scs8hd_decap_12
XFILLER_16_68 vgnd vpwr scs8hd_decap_12
XFILLER_12_105 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.tap_buf4_0_.scs8hd_inv_1 mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _41_/A vgnd vpwr scs8hd_inv_1
XFILLER_7_175 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _19_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_15.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[6] mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_35 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _20_/HI mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_27_177 vgnd vpwr scs8hd_fill_1
XFILLER_27_111 vpwr vgnd scs8hd_fill_2
XFILLER_24_158 vgnd vpwr scs8hd_fill_1
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _31_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_47 vpwr vgnd scs8hd_fill_2
XFILLER_21_36 vpwr vgnd scs8hd_fill_2
XFILLER_21_25 vgnd vpwr scs8hd_decap_6
XFILLER_21_14 vpwr vgnd scs8hd_fill_2
XFILLER_15_147 vpwr vgnd scs8hd_fill_2
XFILLER_7_38 vgnd vpwr scs8hd_decap_8
XFILLER_7_49 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_14 vgnd vpwr scs8hd_decap_12
XFILLER_12_117 vgnd vpwr scs8hd_decap_12
XFILLER_11_172 vgnd vpwr scs8hd_decap_6
XFILLER_7_132 vgnd vpwr scs8hd_decap_4
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XFILLER_27_24 vgnd vpwr scs8hd_decap_6
XFILLER_27_79 vpwr vgnd scs8hd_fill_2
XFILLER_13_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
Xmux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_47 vgnd vpwr scs8hd_decap_6
Xmux_left_track_13.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[5] mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_80 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_47 vpwr vgnd scs8hd_fill_2
XFILLER_27_156 vgnd vpwr scs8hd_decap_6
XFILLER_27_123 vgnd vpwr scs8hd_decap_4
XANTENNA__40__A _40_/A vgnd vpwr scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_170 vgnd vpwr scs8hd_decap_8
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _31_/HI mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_16_26 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_129 vgnd vpwr scs8hd_decap_12
XFILLER_22_91 vgnd vpwr scs8hd_fill_1
XFILLER_8_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XFILLER_13_16 vgnd vpwr scs8hd_decap_4
XFILLER_1_139 vpwr vgnd scs8hd_fill_2
XFILLER_28_90 vpwr vgnd scs8hd_fill_2
XANTENNA__43__A _43_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_94 vpwr vgnd scs8hd_fill_2
XANTENNA__38__A _38_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_19 vgnd vpwr scs8hd_decap_12
XFILLER_10_28 vgnd vpwr scs8hd_decap_3
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XFILLER_4_3 vpwr vgnd scs8hd_fill_2
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _26_/HI mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_11.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[4] mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__51__A _51_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_141 vgnd vpwr scs8hd_decap_12
XANTENNA__46__A _46_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_163 vpwr vgnd scs8hd_fill_2
XFILLER_21_6 vpwr vgnd scs8hd_fill_2
XFILLER_8_50 vgnd vpwr scs8hd_decap_12
XFILLER_4_19 vgnd vpwr scs8hd_decap_12
XFILLER_4_126 vgnd vpwr scs8hd_decap_12
XFILLER_13_39 vgnd vpwr scs8hd_decap_12
XFILLER_1_107 vgnd vpwr scs8hd_decap_3
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _24_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XFILLER_5_51 vgnd vpwr scs8hd_decap_4
XFILLER_5_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_93 vgnd vpwr scs8hd_decap_12
XFILLER_27_169 vpwr vgnd scs8hd_fill_2
XFILLER_19_38 vgnd vpwr scs8hd_decap_4
XANTENNA__49__A _49_/A vgnd vpwr scs8hd_diode_2
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_70 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _19_/HI mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_2_30 vgnd vpwr scs8hd_fill_1
XFILLER_23_161 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _27_/HI vgnd vpwr
+ scs8hd_diode_2
X_39_ _39_/A chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_22_93 vgnd vpwr scs8hd_decap_12
XFILLER_14_6 vpwr vgnd scs8hd_fill_2
XFILLER_11_131 vgnd vpwr scs8hd_decap_12
XFILLER_27_49 vgnd vpwr scs8hd_fill_1
XFILLER_8_62 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_60 vgnd vpwr scs8hd_fill_1
XFILLER_4_138 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _20_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_115 vgnd vpwr scs8hd_decap_6
XFILLER_25_82 vpwr vgnd scs8hd_fill_2
XFILLER_25_71 vgnd vpwr scs8hd_decap_4
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_60 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_71 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_64 vgnd vpwr scs8hd_fill_1
XFILLER_11_62 vgnd vpwr scs8hd_decap_12
X_38_ _38_/A chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_20_165 vgnd vpwr scs8hd_decap_12
XFILLER_20_154 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _30_/HI mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_11_143 vgnd vpwr scs8hd_decap_12
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
XFILLER_7_136 vgnd vpwr scs8hd_fill_1
XFILLER_11_110 vgnd vpwr scs8hd_decap_12
XFILLER_8_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_93 vgnd vpwr scs8hd_decap_4
XFILLER_28_71 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_75 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_15.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_15_ mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_127 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_18_105 vgnd vpwr scs8hd_decap_12
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_61 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _50_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_14_163 vgnd vpwr scs8hd_decap_12
XFILLER_14_141 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_74 vgnd vpwr scs8hd_decap_12
XFILLER_20_177 vgnd vpwr scs8hd_fill_1
X_37_ _37_/A chanx_left_out[7] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _25_/HI mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_11_155 vgnd vpwr scs8hd_decap_6
Xmux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_86 vgnd vpwr scs8hd_decap_6
XFILLER_17_62 vgnd vpwr scs8hd_decap_12
XFILLER_4_107 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_143 vgnd vpwr scs8hd_fill_1
XFILLER_0_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_87 vgnd vpwr scs8hd_decap_3
XFILLER_5_98 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_11.tap_buf4_0_.scs8hd_inv_1 mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _39_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_27_139 vgnd vpwr scs8hd_decap_6
XFILLER_18_117 vgnd vpwr scs8hd_decap_12
XFILLER_4_7 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_13.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_13_ mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_53_ _53_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_26_150 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XPHY_62 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_3.tap_buf4_0_.scs8hd_inv_1 mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _43_/A vgnd vpwr scs8hd_inv_1
XFILLER_14_175 vgnd vpwr scs8hd_decap_3
XFILLER_11_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_36_ _36_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_22_63 vgnd vpwr scs8hd_decap_12
XFILLER_22_52 vgnd vpwr scs8hd_decap_8
XFILLER_22_41 vgnd vpwr scs8hd_decap_8
XFILLER_22_30 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
X_19_ _19_/HI _19_/LO vgnd vpwr scs8hd_conb_1
XFILLER_4_119 vgnd vpwr scs8hd_decap_4
XFILLER_17_74 vgnd vpwr scs8hd_decap_12
XFILLER_3_130 vgnd vpwr scs8hd_decap_12
XFILLER_3_152 vpwr vgnd scs8hd_fill_2
XFILLER_3_163 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _46_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _25_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_166 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_55 vgnd vpwr scs8hd_fill_1
XFILLER_10_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_41 vpwr vgnd scs8hd_fill_2
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_18_129 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_52_ _52_/A chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_2_56 vgnd vpwr scs8hd_decap_8
XPHY_63 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_110 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_11.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _32_/HI vgnd vpwr
+ scs8hd_diode_2
X_35_ _35_/HI _35_/LO vgnd vpwr scs8hd_conb_1
XFILLER_22_75 vgnd vpwr scs8hd_decap_12
XFILLER_11_168 vpwr vgnd scs8hd_fill_2
XFILLER_7_106 vgnd vpwr scs8hd_decap_8
XFILLER_7_139 vgnd vpwr scs8hd_decap_12
XFILLER_8_44 vgnd vpwr scs8hd_decap_3
X_18_ _18_/HI _18_/LO vgnd vpwr scs8hd_conb_1
XFILLER_17_86 vgnd vpwr scs8hd_decap_12
XFILLER_17_53 vgnd vpwr scs8hd_fill_1
XFILLER_17_42 vgnd vpwr scs8hd_fill_1
XFILLER_3_120 vpwr vgnd scs8hd_fill_2
XFILLER_3_142 vgnd vpwr scs8hd_decap_6
XFILLER_3_175 vgnd vpwr scs8hd_decap_3
XFILLER_12_7 vpwr vgnd scs8hd_fill_2
Xmux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _29_/HI mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_156 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _21_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
XFILLER_14_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_25_86 vpwr vgnd scs8hd_fill_2
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XFILLER_25_20 vgnd vpwr scs8hd_decap_8
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_64 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_20 vgnd vpwr scs8hd_decap_3
X_51_ _51_/A chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_2_68 vgnd vpwr scs8hd_decap_8
XFILLER_2_79 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_166 vpwr vgnd scs8hd_fill_2
XFILLER_2_6 vgnd vpwr scs8hd_decap_12
XFILLER_11_33 vgnd vpwr scs8hd_decap_12
X_34_ _34_/HI _34_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_87 vgnd vpwr scs8hd_decap_4
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_151 vpwr vgnd scs8hd_fill_2
XFILLER_17_98 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _24_/HI mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_135 vgnd vpwr scs8hd_decap_6
Xmux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_113 vgnd vpwr scs8hd_decap_8
XFILLER_28_42 vgnd vpwr scs8hd_decap_8
XFILLER_5_79 vgnd vpwr scs8hd_decap_8
XFILLER_14_44 vgnd vpwr scs8hd_decap_12
XFILLER_26_175 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_65 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
X_50_ _50_/A chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_17_175 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_123 vgnd vpwr scs8hd_decap_12
XFILLER_11_45 vgnd vpwr scs8hd_decap_12
XFILLER_14_145 vgnd vpwr scs8hd_decap_8
X_33_ _33_/HI _33_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_90 vgnd vpwr scs8hd_decap_8
XFILLER_26_3 vgnd vpwr scs8hd_decap_3
XFILLER_10_170 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_32 vgnd vpwr scs8hd_fill_1
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XFILLER_0_125 vgnd vpwr scs8hd_fill_1
XFILLER_5_58 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_56 vgnd vpwr scs8hd_decap_12
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_154 vgnd vpwr scs8hd_decap_4
XFILLER_26_132 vgnd vpwr scs8hd_decap_3
XFILLER_25_99 vpwr vgnd scs8hd_fill_2
XFILLER_25_77 vpwr vgnd scs8hd_fill_2
XPHY_44 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_66 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XFILLER_17_154 vpwr vgnd scs8hd_fill_2
XFILLER_17_110 vgnd vpwr scs8hd_decap_12
XFILLER_23_135 vgnd vpwr scs8hd_decap_12
XFILLER_11_57 vgnd vpwr scs8hd_decap_4
XFILLER_28_7 vgnd vpwr scs8hd_decap_12
X_32_ _32_/HI _32_/LO vgnd vpwr scs8hd_conb_1
XFILLER_20_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_172 vgnd vpwr scs8hd_decap_6
XFILLER_11_127 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_9_ mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_120 vgnd vpwr scs8hd_decap_8
XFILLER_6_131 vgnd vpwr scs8hd_decap_12
XFILLER_10_160 vgnd vpwr scs8hd_fill_1
XFILLER_17_56 vgnd vpwr scs8hd_decap_4
XFILLER_17_45 vgnd vpwr scs8hd_decap_8
XFILLER_17_12 vpwr vgnd scs8hd_fill_2
XFILLER_3_112 vgnd vpwr scs8hd_decap_8
XFILLER_3_156 vgnd vpwr scs8hd_decap_4
XFILLER_3_167 vgnd vpwr scs8hd_decap_8
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _26_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_68 vgnd vpwr scs8hd_decap_12
XFILLER_29_141 vpwr vgnd scs8hd_fill_2
Xmux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _28_/HI mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_122 vgnd vpwr scs8hd_decap_8
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_25_45 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_17_144 vpwr vgnd scs8hd_fill_2
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_147 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_117 vgnd vpwr scs8hd_decap_12
X_31_ _31_/HI _31_/LO vgnd vpwr scs8hd_conb_1
XFILLER_9_140 vgnd vpwr scs8hd_fill_1
XFILLER_22_13 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _33_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_143 vgnd vpwr scs8hd_decap_8
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_24 vgnd vpwr scs8hd_decap_3
Xmux_left_track_7.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_7_ mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_78 vgnd vpwr scs8hd_decap_12
XFILLER_28_23 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _22_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XFILLER_10_8 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _52_/A vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _23_/HI mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_153 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_26_167 vgnd vpwr scs8hd_decap_8
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_13 vgnd vpwr scs8hd_decap_3
XFILLER_9_3 vgnd vpwr scs8hd_decap_3
XFILLER_17_167 vgnd vpwr scs8hd_decap_8
XFILLER_17_123 vgnd vpwr scs8hd_decap_12
XFILLER_20_129 vgnd vpwr scs8hd_decap_12
X_30_ _30_/HI _30_/LO vgnd vpwr scs8hd_conb_1
Xmux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_60 vgnd vpwr scs8hd_fill_1
XFILLER_9_163 vpwr vgnd scs8hd_fill_2
XFILLER_12_80 vgnd vpwr scs8hd_decap_12
XFILLER_6_166 vgnd vpwr scs8hd_decap_12
XFILLER_8_16 vgnd vpwr scs8hd_decap_12
XFILLER_24_3 vgnd vpwr scs8hd_decap_3
XFILLER_0_94 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_176 vpwr vgnd scs8hd_fill_2
XFILLER_29_110 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_5.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_5_ mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_91 vgnd vpwr scs8hd_fill_1
XFILLER_6_71 vgnd vpwr scs8hd_decap_4
XFILLER_6_93 vgnd vpwr scs8hd_decap_6
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_69 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_14 vgnd vpwr scs8hd_decap_3
XFILLER_17_135 vgnd vpwr scs8hd_decap_4
XFILLER_2_18 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__41__A _41_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__36__A _36_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_28 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _48_/A vgnd vpwr scs8hd_inv_1
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _35_/HI mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_19_6 vpwr vgnd scs8hd_fill_2
XFILLER_3_126 vpwr vgnd scs8hd_fill_2
XFILLER_3_148 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _36_/A vgnd vpwr scs8hd_inv_1
XFILLER_29_122 vpwr vgnd scs8hd_fill_2
XANTENNA__44__A _44_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_90 vgnd vpwr scs8hd_decap_3
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _40_/A vgnd vpwr scs8hd_inv_1
XPHY_59 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
Xmux_left_track_3.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_3_ mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__39__A _39_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_106 vpwr vgnd scs8hd_fill_2
XFILLER_14_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_62 vgnd vpwr scs8hd_decap_4
XFILLER_3_73 vpwr vgnd scs8hd_fill_2
XFILLER_9_110 vgnd vpwr scs8hd_decap_8
XFILLER_9_132 vpwr vgnd scs8hd_fill_2
XFILLER_12_93 vgnd vpwr scs8hd_decap_12
XANTENNA__52__A _52_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_38 vgnd vpwr scs8hd_decap_4
XFILLER_17_16 vgnd vpwr scs8hd_decap_8
XANTENNA__47__A _47_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_28_59 vgnd vpwr scs8hd_decap_12
XFILLER_18_81 vgnd vpwr scs8hd_decap_8
XFILLER_29_156 vgnd vpwr scs8hd_decap_12
XFILLER_29_145 vgnd vpwr scs8hd_decap_8
XFILLER_14_17 vgnd vpwr scs8hd_decap_12
XFILLER_20_93 vgnd vpwr scs8hd_decap_12
XFILLER_20_71 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_16 vpwr vgnd scs8hd_fill_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XFILLER_6_84 vgnd vpwr scs8hd_decap_8
XPHY_16 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _18_/HI mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_17_148 vgnd vpwr scs8hd_decap_4
XFILLER_11_18 vgnd vpwr scs8hd_decap_8
XFILLER_11_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _34_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_1_ mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_103 vgnd vpwr scs8hd_decap_8
XFILLER_10_154 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_7.INVTX1_1_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_71 vgnd vpwr scs8hd_fill_1
XFILLER_23_60 vgnd vpwr scs8hd_fill_1
XFILLER_0_75 vgnd vpwr scs8hd_decap_6
XFILLER_9_62 vgnd vpwr scs8hd_decap_12
XFILLER_18_93 vgnd vpwr scs8hd_decap_12
XFILLER_22_3 vgnd vpwr scs8hd_fill_1
XFILLER_14_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_168 vgnd vpwr scs8hd_decap_8
XFILLER_20_83 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_26_138 vgnd vpwr scs8hd_decap_12
XFILLER_26_105 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_17 vgnd vpwr scs8hd_decap_3
XFILLER_25_28 vpwr vgnd scs8hd_fill_2
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_22_141 vgnd vpwr scs8hd_decap_12
XFILLER_26_93 vgnd vpwr scs8hd_decap_3
XFILLER_13_141 vgnd vpwr scs8hd_fill_1
XFILLER_9_145 vpwr vgnd scs8hd_fill_2
Xmux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_10_122 vgnd vpwr scs8hd_decap_8
XFILLER_10_133 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_2_140 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _34_/HI mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_9_74 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.INVTX1_1_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_3 vpwr vgnd scs8hd_fill_2
XFILLER_29_125 vgnd vpwr scs8hd_decap_12
XFILLER_29_114 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_82 vgnd vpwr scs8hd_decap_8
XPHY_29 vgnd vpwr scs8hd_decap_3
XPHY_18 vgnd vpwr scs8hd_decap_3
XFILLER_17_139 vgnd vpwr scs8hd_fill_1
XFILLER_15_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_98 vgnd vpwr scs8hd_decap_3
XFILLER_9_168 vpwr vgnd scs8hd_fill_2
XFILLER_12_30 vgnd vpwr scs8hd_fill_1
XFILLER_10_145 vgnd vpwr scs8hd_decap_8
XFILLER_23_95 vgnd vpwr scs8hd_decap_6
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
XFILLER_2_152 vgnd vpwr scs8hd_fill_1
XFILLER_2_163 vgnd vpwr scs8hd_decap_12
XFILLER_9_31 vgnd vpwr scs8hd_decap_8
XFILLER_9_53 vgnd vpwr scs8hd_decap_8
XFILLER_9_86 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_137 vgnd vpwr scs8hd_fill_1
XFILLER_29_94 vpwr vgnd scs8hd_fill_2
XFILLER_29_50 vgnd vpwr scs8hd_decap_12
XFILLER_20_30 vgnd vpwr scs8hd_fill_1
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_3.INVTX1_1_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_74 vgnd vpwr scs8hd_decap_12
XFILLER_26_84 vgnd vpwr scs8hd_decap_8
XFILLER_22_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_6 vpwr vgnd scs8hd_fill_2
XFILLER_13_165 vgnd vpwr scs8hd_decap_12
XFILLER_13_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_66 vgnd vpwr scs8hd_fill_1
XFILLER_3_77 vpwr vgnd scs8hd_fill_2
XFILLER_9_136 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_23_74 vgnd vpwr scs8hd_decap_12
XFILLER_23_52 vpwr vgnd scs8hd_fill_2
XFILLER_2_131 vgnd vpwr scs8hd_decap_6
XFILLER_2_175 vgnd vpwr scs8hd_decap_3
XFILLER_28_19 vgnd vpwr scs8hd_fill_1
XFILLER_0_89 vgnd vpwr scs8hd_decap_4
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XFILLER_9_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_6_99 vgnd vpwr scs8hd_fill_1
XFILLER_15_86 vgnd vpwr scs8hd_decap_12
XFILLER_15_42 vpwr vgnd scs8hd_fill_2
XFILLER_15_31 vgnd vpwr scs8hd_decap_8
XFILLER_16_141 vgnd vpwr scs8hd_decap_12
.ends

