magic
tech sky130A
magscale 1 2
timestamp 1608763979
<< checkpaint >>
rect -1260 -1260 21260 18260
<< locali >>
rect 6745 14263 6779 14365
rect 12265 10999 12299 11169
rect 6653 10455 6687 10625
rect 7205 8891 7239 9061
rect 13001 8959 13035 9129
rect 11897 8823 11931 8925
rect 9505 7735 9539 7905
rect 12541 6783 12575 6885
rect 2789 6239 2823 6409
rect 6929 5763 6963 5865
rect 7021 5559 7055 5729
rect 13001 5627 13035 5865
rect 15025 5763 15059 5865
rect 7573 5015 7607 5185
rect 5181 3927 5215 4097
rect 10885 2907 10919 3077
rect 12265 2839 12299 3145
rect 15209 2295 15243 2397
<< viali >>
rect 6193 14569 6227 14603
rect 7665 14569 7699 14603
rect 9045 14569 9079 14603
rect 10149 14569 10183 14603
rect 13369 14569 13403 14603
rect 8125 14501 8159 14535
rect 10517 14501 10551 14535
rect 16129 14501 16163 14535
rect 17049 14501 17083 14535
rect 8033 14433 8067 14467
rect 9137 14433 9171 14467
rect 11529 14433 11563 14467
rect 11621 14433 11655 14467
rect 13737 14433 13771 14467
rect 14749 14433 14783 14467
rect 14841 14433 14875 14467
rect 15520 14433 15554 14467
rect 6285 14365 6319 14399
rect 6469 14365 6503 14399
rect 6745 14365 6779 14399
rect 8217 14365 8251 14399
rect 9229 14365 9263 14399
rect 10609 14365 10643 14399
rect 10793 14365 10827 14399
rect 11713 14365 11747 14399
rect 13829 14365 13863 14399
rect 13921 14365 13955 14399
rect 14933 14365 14967 14399
rect 16037 14365 16071 14399
rect 8677 14297 8711 14331
rect 5825 14229 5859 14263
rect 6745 14229 6779 14263
rect 11161 14229 11195 14263
rect 14381 14229 14415 14263
rect 15623 14229 15657 14263
rect 8585 14025 8619 14059
rect 9597 14025 9631 14059
rect 10609 14025 10643 14059
rect 15025 14025 15059 14059
rect 5181 13957 5215 13991
rect 6837 13957 6871 13991
rect 18245 13957 18279 13991
rect 5733 13889 5767 13923
rect 7481 13889 7515 13923
rect 9229 13889 9263 13923
rect 10241 13889 10275 13923
rect 11161 13889 11195 13923
rect 11897 13889 11931 13923
rect 13737 13889 13771 13923
rect 15669 13889 15703 13923
rect 16129 13889 16163 13923
rect 17141 13889 17175 13923
rect 7297 13821 7331 13855
rect 11069 13821 11103 13855
rect 11621 13821 11655 13855
rect 13093 13821 13127 13855
rect 13461 13821 13495 13855
rect 15485 13821 15519 13855
rect 17417 13821 17451 13855
rect 18061 13821 18095 13855
rect 7205 13753 7239 13787
rect 8953 13753 8987 13787
rect 9045 13753 9079 13787
rect 16221 13753 16255 13787
rect 5549 13685 5583 13719
rect 5641 13685 5675 13719
rect 9965 13685 9999 13719
rect 10057 13685 10091 13719
rect 10977 13685 11011 13719
rect 15393 13685 15427 13719
rect 17601 13685 17635 13719
rect 5641 13481 5675 13515
rect 8033 13481 8067 13515
rect 8585 13481 8619 13515
rect 9689 13481 9723 13515
rect 10517 13481 10551 13515
rect 10885 13481 10919 13515
rect 12173 13481 12207 13515
rect 12633 13481 12667 13515
rect 14197 13481 14231 13515
rect 14565 13481 14599 13515
rect 15485 13481 15519 13515
rect 14657 13413 14691 13447
rect 15945 13413 15979 13447
rect 17969 13413 18003 13447
rect 6009 13345 6043 13379
rect 6101 13345 6135 13379
rect 6920 13345 6954 13379
rect 8953 13345 8987 13379
rect 9045 13345 9079 13379
rect 12541 13345 12575 13379
rect 13553 13345 13587 13379
rect 15853 13345 15887 13379
rect 16865 13345 16899 13379
rect 16957 13345 16991 13379
rect 17877 13345 17911 13379
rect 6285 13277 6319 13311
rect 6653 13277 6687 13311
rect 9229 13277 9263 13311
rect 10977 13277 11011 13311
rect 11069 13277 11103 13311
rect 12817 13277 12851 13311
rect 13645 13277 13679 13311
rect 13829 13277 13863 13311
rect 14841 13277 14875 13311
rect 16129 13277 16163 13311
rect 17049 13277 17083 13311
rect 18153 13277 18187 13311
rect 16497 13209 16531 13243
rect 13185 13141 13219 13175
rect 17509 13141 17543 13175
rect 5549 12937 5583 12971
rect 8309 12937 8343 12971
rect 10333 12937 10367 12971
rect 11345 12937 11379 12971
rect 13829 12937 13863 12971
rect 5089 12801 5123 12835
rect 6009 12801 6043 12835
rect 6193 12801 6227 12835
rect 10885 12801 10919 12835
rect 11805 12801 11839 12835
rect 11989 12801 12023 12835
rect 17417 12801 17451 12835
rect 3157 12733 3191 12767
rect 6929 12733 6963 12767
rect 7196 12733 7230 12767
rect 8585 12733 8619 12767
rect 8852 12733 8886 12767
rect 10701 12733 10735 12767
rect 12449 12733 12483 12767
rect 14933 12733 14967 12767
rect 15200 12733 15234 12767
rect 17233 12733 17267 12767
rect 3424 12665 3458 12699
rect 5917 12665 5951 12699
rect 10793 12665 10827 12699
rect 11713 12665 11747 12699
rect 12716 12665 12750 12699
rect 2513 12597 2547 12631
rect 4537 12597 4571 12631
rect 9965 12597 9999 12631
rect 16313 12597 16347 12631
rect 16865 12597 16899 12631
rect 17325 12597 17359 12631
rect 3341 12393 3375 12427
rect 6101 12393 6135 12427
rect 7573 12393 7607 12427
rect 8125 12393 8159 12427
rect 11713 12393 11747 12427
rect 14657 12393 14691 12427
rect 15301 12393 15335 12427
rect 18153 12393 18187 12427
rect 4344 12325 4378 12359
rect 10578 12325 10612 12359
rect 12633 12325 12667 12359
rect 13544 12325 13578 12359
rect 2237 12257 2271 12291
rect 6469 12257 6503 12291
rect 7481 12257 7515 12291
rect 8493 12257 8527 12291
rect 12725 12257 12759 12291
rect 16129 12257 16163 12291
rect 16773 12257 16807 12291
rect 17040 12257 17074 12291
rect 2329 12189 2363 12223
rect 2513 12189 2547 12223
rect 3433 12189 3467 12223
rect 3617 12189 3651 12223
rect 4077 12189 4111 12223
rect 6561 12189 6595 12223
rect 6745 12189 6779 12223
rect 7665 12189 7699 12223
rect 8585 12189 8619 12223
rect 8769 12189 8803 12223
rect 10333 12189 10367 12223
rect 12909 12189 12943 12223
rect 13277 12189 13311 12223
rect 16221 12189 16255 12223
rect 16405 12189 16439 12223
rect 2973 12121 3007 12155
rect 1869 12053 1903 12087
rect 5457 12053 5491 12087
rect 7113 12053 7147 12087
rect 12265 12053 12299 12087
rect 15761 12053 15795 12087
rect 2237 11849 2271 11883
rect 6837 11849 6871 11883
rect 11345 11849 11379 11883
rect 14105 11849 14139 11883
rect 16221 11849 16255 11883
rect 5733 11781 5767 11815
rect 9321 11781 9355 11815
rect 2789 11713 2823 11747
rect 6285 11713 6319 11747
rect 7481 11713 7515 11747
rect 10149 11713 10183 11747
rect 11805 11713 11839 11747
rect 11989 11713 12023 11747
rect 14657 11713 14691 11747
rect 15669 11713 15703 11747
rect 15853 11713 15887 11747
rect 16773 11713 16807 11747
rect 1685 11645 1719 11679
rect 2605 11645 2639 11679
rect 3249 11645 3283 11679
rect 3801 11645 3835 11679
rect 7205 11645 7239 11679
rect 7297 11645 7331 11679
rect 7941 11645 7975 11679
rect 8208 11645 8242 11679
rect 11713 11645 11747 11679
rect 12449 11645 12483 11679
rect 12716 11645 12750 11679
rect 16589 11645 16623 11679
rect 2697 11577 2731 11611
rect 4068 11577 4102 11611
rect 10057 11577 10091 11611
rect 14473 11577 14507 11611
rect 15577 11577 15611 11611
rect 1869 11509 1903 11543
rect 3433 11509 3467 11543
rect 5181 11509 5215 11543
rect 6101 11509 6135 11543
rect 6193 11509 6227 11543
rect 9597 11509 9631 11543
rect 9965 11509 9999 11543
rect 13829 11509 13863 11543
rect 14565 11509 14599 11543
rect 15209 11509 15243 11543
rect 16681 11509 16715 11543
rect 6561 11305 6595 11339
rect 7573 11305 7607 11339
rect 8033 11305 8067 11339
rect 8585 11305 8619 11339
rect 9689 11305 9723 11339
rect 13737 11305 13771 11339
rect 14013 11305 14047 11339
rect 16221 11305 16255 11339
rect 17417 11305 17451 11339
rect 17877 11305 17911 11339
rect 16589 11237 16623 11271
rect 1685 11169 1719 11203
rect 2504 11169 2538 11203
rect 4344 11169 4378 11203
rect 6929 11169 6963 11203
rect 7021 11169 7055 11203
rect 7941 11169 7975 11203
rect 8953 11169 8987 11203
rect 9045 11169 9079 11203
rect 10057 11169 10091 11203
rect 11253 11169 11287 11203
rect 11713 11169 11747 11203
rect 12265 11169 12299 11203
rect 12357 11169 12391 11203
rect 12624 11169 12658 11203
rect 14381 11169 14415 11203
rect 17785 11169 17819 11203
rect 2237 11101 2271 11135
rect 4077 11101 4111 11135
rect 7205 11101 7239 11135
rect 8125 11101 8159 11135
rect 9137 11101 9171 11135
rect 10149 11101 10183 11135
rect 10241 11101 10275 11135
rect 11805 11101 11839 11135
rect 11989 11101 12023 11135
rect 1869 11033 1903 11067
rect 3617 11033 3651 11067
rect 5457 11033 5491 11067
rect 11345 11033 11379 11067
rect 14473 11101 14507 11135
rect 14565 11101 14599 11135
rect 15301 11101 15335 11135
rect 16681 11101 16715 11135
rect 16865 11101 16899 11135
rect 18061 11101 18095 11135
rect 11069 10965 11103 10999
rect 12265 10965 12299 10999
rect 2237 10761 2271 10795
rect 8769 10761 8803 10795
rect 10425 10761 10459 10795
rect 11345 10761 11379 10795
rect 13645 10761 13679 10795
rect 16037 10761 16071 10795
rect 17693 10761 17727 10795
rect 1869 10693 1903 10727
rect 2881 10625 2915 10659
rect 4077 10625 4111 10659
rect 5089 10625 5123 10659
rect 6009 10625 6043 10659
rect 6653 10625 6687 10659
rect 7389 10625 7423 10659
rect 11989 10625 12023 10659
rect 13093 10625 13127 10659
rect 14197 10625 14231 10659
rect 14657 10625 14691 10659
rect 1685 10557 1719 10591
rect 2697 10557 2731 10591
rect 2605 10489 2639 10523
rect 5917 10489 5951 10523
rect 7297 10557 7331 10591
rect 9045 10557 9079 10591
rect 9301 10557 9335 10591
rect 16313 10557 16347 10591
rect 16569 10557 16603 10591
rect 7634 10489 7668 10523
rect 14013 10489 14047 10523
rect 14924 10489 14958 10523
rect 3433 10421 3467 10455
rect 3801 10421 3835 10455
rect 3893 10421 3927 10455
rect 4445 10421 4479 10455
rect 4813 10421 4847 10455
rect 4905 10421 4939 10455
rect 5457 10421 5491 10455
rect 5825 10421 5859 10455
rect 6653 10421 6687 10455
rect 7113 10421 7147 10455
rect 11713 10421 11747 10455
rect 11805 10421 11839 10455
rect 12449 10421 12483 10455
rect 12817 10421 12851 10455
rect 12909 10421 12943 10455
rect 14105 10421 14139 10455
rect 3617 10217 3651 10251
rect 4445 10217 4479 10251
rect 4813 10217 4847 10251
rect 5549 10217 5583 10251
rect 7849 10217 7883 10251
rect 8493 10217 8527 10251
rect 8861 10217 8895 10251
rect 12633 10217 12667 10251
rect 14565 10217 14599 10251
rect 17509 10217 17543 10251
rect 17877 10217 17911 10251
rect 1676 10149 1710 10183
rect 9934 10149 9968 10183
rect 13430 10149 13464 10183
rect 16396 10149 16430 10183
rect 3065 10081 3099 10115
rect 3801 10081 3835 10115
rect 4905 10081 4939 10115
rect 5733 10081 5767 10115
rect 6092 10081 6126 10115
rect 9689 10081 9723 10115
rect 12541 10081 12575 10115
rect 15669 10081 15703 10115
rect 1409 10013 1443 10047
rect 5089 10013 5123 10047
rect 5825 10013 5859 10047
rect 7941 10013 7975 10047
rect 8033 10013 8067 10047
rect 8953 10013 8987 10047
rect 9045 10013 9079 10047
rect 12817 10013 12851 10047
rect 13185 10013 13219 10047
rect 16129 10013 16163 10047
rect 7481 9945 7515 9979
rect 11069 9945 11103 9979
rect 15485 9945 15519 9979
rect 2789 9877 2823 9911
rect 3249 9877 3283 9911
rect 7205 9877 7239 9911
rect 12173 9877 12207 9911
rect 4445 9605 4479 9639
rect 13461 9605 13495 9639
rect 16773 9605 16807 9639
rect 2145 9537 2179 9571
rect 4905 9537 4939 9571
rect 5089 9537 5123 9571
rect 6377 9537 6411 9571
rect 7757 9537 7791 9571
rect 8769 9537 8803 9571
rect 9229 9537 9263 9571
rect 13093 9537 13127 9571
rect 14197 9537 14231 9571
rect 17417 9537 17451 9571
rect 1593 9469 1627 9503
rect 2412 9469 2446 9503
rect 3801 9469 3835 9503
rect 7573 9469 7607 9503
rect 8677 9469 8711 9503
rect 9873 9469 9907 9503
rect 13645 9469 13679 9503
rect 17233 9469 17267 9503
rect 8585 9401 8619 9435
rect 10140 9401 10174 9435
rect 12909 9401 12943 9435
rect 14464 9401 14498 9435
rect 1777 9333 1811 9367
rect 3525 9333 3559 9367
rect 3985 9333 4019 9367
rect 4813 9333 4847 9367
rect 5733 9333 5767 9367
rect 6101 9333 6135 9367
rect 6193 9333 6227 9367
rect 7205 9333 7239 9367
rect 7665 9333 7699 9367
rect 8217 9333 8251 9367
rect 11253 9333 11287 9367
rect 12449 9333 12483 9367
rect 12817 9333 12851 9367
rect 15577 9333 15611 9367
rect 17141 9333 17175 9367
rect 2237 9129 2271 9163
rect 2329 9129 2363 9163
rect 2973 9129 3007 9163
rect 3433 9129 3467 9163
rect 10241 9129 10275 9163
rect 11437 9129 11471 9163
rect 12081 9129 12115 9163
rect 12541 9129 12575 9163
rect 13001 9129 13035 9163
rect 15301 9129 15335 9163
rect 18245 9129 18279 9163
rect 4322 9061 4356 9095
rect 7205 9061 7239 9095
rect 7656 9061 7690 9095
rect 12449 9061 12483 9095
rect 3341 8993 3375 9027
rect 6000 8993 6034 9027
rect 2513 8925 2547 8959
rect 3525 8925 3559 8959
rect 4077 8925 4111 8959
rect 5733 8925 5767 8959
rect 10333 8993 10367 9027
rect 11529 8993 11563 9027
rect 13360 8993 13394 9027
rect 15669 8993 15703 9027
rect 16865 8993 16899 9027
rect 17132 8993 17166 9027
rect 7389 8925 7423 8959
rect 9045 8925 9079 8959
rect 10425 8925 10459 8959
rect 11713 8925 11747 8959
rect 11897 8925 11931 8959
rect 12633 8925 12667 8959
rect 13001 8925 13035 8959
rect 13093 8925 13127 8959
rect 15761 8925 15795 8959
rect 15945 8925 15979 8959
rect 7113 8857 7147 8891
rect 7205 8857 7239 8891
rect 11069 8857 11103 8891
rect 1869 8789 1903 8823
rect 5457 8789 5491 8823
rect 8769 8789 8803 8823
rect 9873 8789 9907 8823
rect 11897 8789 11931 8823
rect 14473 8789 14507 8823
rect 5641 8585 5675 8619
rect 5917 8585 5951 8619
rect 7021 8585 7055 8619
rect 10425 8585 10459 8619
rect 13829 8585 13863 8619
rect 17417 8585 17451 8619
rect 4353 8517 4387 8551
rect 10977 8517 11011 8551
rect 11989 8517 12023 8551
rect 1409 8449 1443 8483
rect 3893 8449 3927 8483
rect 4997 8449 5031 8483
rect 6561 8449 6595 8483
rect 11437 8449 11471 8483
rect 11621 8449 11655 8483
rect 14933 8449 14967 8483
rect 16037 8449 16071 8483
rect 3709 8381 3743 8415
rect 4813 8381 4847 8415
rect 5825 8381 5859 8415
rect 6837 8381 6871 8415
rect 7481 8381 7515 8415
rect 9137 8381 9171 8415
rect 12173 8381 12207 8415
rect 12449 8381 12483 8415
rect 16304 8381 16338 8415
rect 18061 8381 18095 8415
rect 1676 8313 1710 8347
rect 3801 8313 3835 8347
rect 4721 8313 4755 8347
rect 6377 8313 6411 8347
rect 7748 8313 7782 8347
rect 12694 8313 12728 8347
rect 14749 8313 14783 8347
rect 14841 8313 14875 8347
rect 2789 8245 2823 8279
rect 3341 8245 3375 8279
rect 6285 8245 6319 8279
rect 8861 8245 8895 8279
rect 11345 8245 11379 8279
rect 14381 8245 14415 8279
rect 18245 8245 18279 8279
rect 2421 8041 2455 8075
rect 2973 8041 3007 8075
rect 3433 8041 3467 8075
rect 6285 8041 6319 8075
rect 6653 8041 6687 8075
rect 7113 8041 7147 8075
rect 7481 8041 7515 8075
rect 8125 8041 8159 8075
rect 8493 8041 8527 8075
rect 9137 8041 9171 8075
rect 9689 8041 9723 8075
rect 11897 8041 11931 8075
rect 13185 8041 13219 8075
rect 14197 8041 14231 8075
rect 14657 8041 14691 8075
rect 17417 8041 17451 8075
rect 7573 7973 7607 8007
rect 10149 7973 10183 8007
rect 10784 7973 10818 8007
rect 13553 7973 13587 8007
rect 14565 7973 14599 8007
rect 16282 7973 16316 8007
rect 1409 7905 1443 7939
rect 2329 7905 2363 7939
rect 3341 7905 3375 7939
rect 4077 7905 4111 7939
rect 5080 7905 5114 7939
rect 6745 7905 6779 7939
rect 9505 7905 9539 7939
rect 10057 7905 10091 7939
rect 12541 7905 12575 7939
rect 16037 7905 16071 7939
rect 17877 7905 17911 7939
rect 2605 7837 2639 7871
rect 3617 7837 3651 7871
rect 4813 7837 4847 7871
rect 6929 7837 6963 7871
rect 7665 7837 7699 7871
rect 8585 7837 8619 7871
rect 8769 7837 8803 7871
rect 1593 7769 1627 7803
rect 6193 7769 6227 7803
rect 10241 7837 10275 7871
rect 10517 7837 10551 7871
rect 12633 7837 12667 7871
rect 12817 7837 12851 7871
rect 13645 7837 13679 7871
rect 13829 7837 13863 7871
rect 14841 7837 14875 7871
rect 1961 7701 1995 7735
rect 4261 7701 4295 7735
rect 9505 7701 9539 7735
rect 12173 7701 12207 7735
rect 18061 7701 18095 7735
rect 3249 7497 3283 7531
rect 4445 7497 4479 7531
rect 6377 7497 6411 7531
rect 10333 7497 10367 7531
rect 16865 7497 16899 7531
rect 17601 7497 17635 7531
rect 3893 7361 3927 7395
rect 8125 7361 8159 7395
rect 10793 7361 10827 7395
rect 10977 7361 11011 7395
rect 11897 7361 11931 7395
rect 13093 7361 13127 7395
rect 13277 7361 13311 7395
rect 14289 7361 14323 7395
rect 1593 7293 1627 7327
rect 3617 7293 3651 7327
rect 4261 7293 4295 7327
rect 4997 7293 5031 7327
rect 6837 7293 6871 7327
rect 8585 7293 8619 7327
rect 14105 7293 14139 7327
rect 15485 7293 15519 7327
rect 17417 7293 17451 7327
rect 18061 7293 18095 7327
rect 1860 7225 1894 7259
rect 5264 7225 5298 7259
rect 7849 7225 7883 7259
rect 8852 7225 8886 7259
rect 10701 7225 10735 7259
rect 15730 7225 15764 7259
rect 2973 7157 3007 7191
rect 3709 7157 3743 7191
rect 7021 7157 7055 7191
rect 7481 7157 7515 7191
rect 7941 7157 7975 7191
rect 9965 7157 9999 7191
rect 11345 7157 11379 7191
rect 11713 7157 11747 7191
rect 11805 7157 11839 7191
rect 12633 7157 12667 7191
rect 13001 7157 13035 7191
rect 13645 7157 13679 7191
rect 14013 7157 14047 7191
rect 14749 7157 14783 7191
rect 18245 7157 18279 7191
rect 4077 6953 4111 6987
rect 5825 6953 5859 6987
rect 6377 6953 6411 6987
rect 6745 6953 6779 6987
rect 11621 6953 11655 6987
rect 14013 6953 14047 6987
rect 15669 6953 15703 6987
rect 16313 6953 16347 6987
rect 5733 6885 5767 6919
rect 11989 6885 12023 6919
rect 12541 6885 12575 6919
rect 13001 6885 13035 6919
rect 13093 6885 13127 6919
rect 16681 6885 16715 6919
rect 1685 6817 1719 6851
rect 2596 6817 2630 6851
rect 4445 6817 4479 6851
rect 5273 6817 5307 6851
rect 6837 6817 6871 6851
rect 7389 6817 7423 6851
rect 7656 6817 7690 6851
rect 9873 6817 9907 6851
rect 10140 6817 10174 6851
rect 14841 6817 14875 6851
rect 17877 6817 17911 6851
rect 2329 6749 2363 6783
rect 4537 6749 4571 6783
rect 4721 6749 4755 6783
rect 6009 6749 6043 6783
rect 7021 6749 7055 6783
rect 9045 6749 9079 6783
rect 12081 6749 12115 6783
rect 12265 6749 12299 6783
rect 12541 6749 12575 6783
rect 13185 6749 13219 6783
rect 14105 6749 14139 6783
rect 14197 6749 14231 6783
rect 15761 6749 15795 6783
rect 15853 6749 15887 6783
rect 16773 6749 16807 6783
rect 16865 6749 16899 6783
rect 8769 6681 8803 6715
rect 11253 6681 11287 6715
rect 13645 6681 13679 6715
rect 15301 6681 15335 6715
rect 1869 6613 1903 6647
rect 3709 6613 3743 6647
rect 5089 6613 5123 6647
rect 5365 6613 5399 6647
rect 12633 6613 12667 6647
rect 14657 6613 14691 6647
rect 18061 6613 18095 6647
rect 2789 6409 2823 6443
rect 5549 6409 5583 6443
rect 8217 6409 8251 6443
rect 14657 6409 14691 6443
rect 14933 6409 14967 6443
rect 2329 6273 2363 6307
rect 2513 6273 2547 6307
rect 13001 6341 13035 6375
rect 3433 6273 3467 6307
rect 6101 6273 6135 6307
rect 9045 6273 9079 6307
rect 11897 6273 11931 6307
rect 15485 6273 15519 6307
rect 16405 6273 16439 6307
rect 16497 6273 16531 6307
rect 1409 6205 1443 6239
rect 2789 6205 2823 6239
rect 3249 6205 3283 6239
rect 3893 6205 3927 6239
rect 4149 6205 4183 6239
rect 6009 6205 6043 6239
rect 6837 6205 6871 6239
rect 7093 6205 7127 6239
rect 8493 6205 8527 6239
rect 11805 6205 11839 6239
rect 13185 6205 13219 6239
rect 13277 6205 13311 6239
rect 13533 6205 13567 6239
rect 15301 6205 15335 6239
rect 15393 6205 15427 6239
rect 17417 6205 17451 6239
rect 18061 6205 18095 6239
rect 3341 6137 3375 6171
rect 9312 6137 9346 6171
rect 11713 6137 11747 6171
rect 12541 6137 12575 6171
rect 1869 6069 1903 6103
rect 2237 6069 2271 6103
rect 2881 6069 2915 6103
rect 5273 6069 5307 6103
rect 5917 6069 5951 6103
rect 8677 6069 8711 6103
rect 10425 6069 10459 6103
rect 10701 6069 10735 6103
rect 11345 6069 11379 6103
rect 15945 6069 15979 6103
rect 16313 6069 16347 6103
rect 17601 6069 17635 6103
rect 18245 6069 18279 6103
rect 4537 5865 4571 5899
rect 6837 5865 6871 5899
rect 6929 5865 6963 5899
rect 9321 5865 9355 5899
rect 13001 5865 13035 5899
rect 13645 5865 13679 5899
rect 14197 5865 14231 5899
rect 14565 5865 14599 5899
rect 15025 5865 15059 5899
rect 1593 5729 1627 5763
rect 1860 5729 1894 5763
rect 3249 5729 3283 5763
rect 4445 5729 4479 5763
rect 5273 5729 5307 5763
rect 5724 5729 5758 5763
rect 6929 5729 6963 5763
rect 7021 5729 7055 5763
rect 7113 5729 7147 5763
rect 7849 5729 7883 5763
rect 7941 5729 7975 5763
rect 8208 5729 8242 5763
rect 9873 5729 9907 5763
rect 10140 5729 10174 5763
rect 11529 5729 11563 5763
rect 11796 5729 11830 5763
rect 4629 5661 4663 5695
rect 5457 5661 5491 5695
rect 13553 5797 13587 5831
rect 15025 5729 15059 5763
rect 15669 5729 15703 5763
rect 17325 5729 17359 5763
rect 17877 5729 17911 5763
rect 13737 5661 13771 5695
rect 14657 5661 14691 5695
rect 14841 5661 14875 5695
rect 15761 5661 15795 5695
rect 15853 5661 15887 5695
rect 7665 5593 7699 5627
rect 13001 5593 13035 5627
rect 17509 5593 17543 5627
rect 2973 5525 3007 5559
rect 3433 5525 3467 5559
rect 4077 5525 4111 5559
rect 5089 5525 5123 5559
rect 7021 5525 7055 5559
rect 7297 5525 7331 5559
rect 11253 5525 11287 5559
rect 12909 5525 12943 5559
rect 13185 5525 13219 5559
rect 15301 5525 15335 5559
rect 18061 5525 18095 5559
rect 8677 5321 8711 5355
rect 9689 5321 9723 5355
rect 10701 5321 10735 5355
rect 15301 5321 15335 5355
rect 15577 5321 15611 5355
rect 4261 5185 4295 5219
rect 4353 5185 4387 5219
rect 5365 5185 5399 5219
rect 7205 5185 7239 5219
rect 7573 5185 7607 5219
rect 8217 5185 8251 5219
rect 9137 5185 9171 5219
rect 9321 5185 9355 5219
rect 10241 5185 10275 5219
rect 11253 5185 11287 5219
rect 13553 5185 13587 5219
rect 16129 5185 16163 5219
rect 1409 5117 1443 5151
rect 3065 5117 3099 5151
rect 4169 5117 4203 5151
rect 5825 5117 5859 5151
rect 6929 5117 6963 5151
rect 1676 5049 1710 5083
rect 3341 5049 3375 5083
rect 5273 5049 5307 5083
rect 6101 5049 6135 5083
rect 8125 5117 8159 5151
rect 11069 5117 11103 5151
rect 11161 5117 11195 5151
rect 11713 5117 11747 5151
rect 13921 5117 13955 5151
rect 14188 5117 14222 5151
rect 16037 5117 16071 5151
rect 18061 5117 18095 5151
rect 9045 5049 9079 5083
rect 13277 5049 13311 5083
rect 2789 4981 2823 5015
rect 3801 4981 3835 5015
rect 4813 4981 4847 5015
rect 5181 4981 5215 5015
rect 7573 4981 7607 5015
rect 7665 4981 7699 5015
rect 8033 4981 8067 5015
rect 10057 4981 10091 5015
rect 10149 4981 10183 5015
rect 12909 4981 12943 5015
rect 13369 4981 13403 5015
rect 15945 4981 15979 5015
rect 18245 4981 18279 5015
rect 2329 4777 2363 4811
rect 5457 4777 5491 4811
rect 6745 4777 6779 4811
rect 7757 4777 7791 4811
rect 9689 4777 9723 4811
rect 10701 4777 10735 4811
rect 11437 4777 11471 4811
rect 13369 4777 13403 4811
rect 13645 4777 13679 4811
rect 14657 4777 14691 4811
rect 3341 4709 3375 4743
rect 8125 4709 8159 4743
rect 11345 4709 11379 4743
rect 12234 4709 12268 4743
rect 15761 4709 15795 4743
rect 1409 4641 1443 4675
rect 2421 4641 2455 4675
rect 3433 4641 3467 4675
rect 4344 4641 4378 4675
rect 6101 4641 6135 4675
rect 6193 4641 6227 4675
rect 7113 4641 7147 4675
rect 8769 4641 8803 4675
rect 10057 4641 10091 4675
rect 10885 4641 10919 4675
rect 14013 4641 14047 4675
rect 15669 4641 15703 4675
rect 17325 4641 17359 4675
rect 17877 4641 17911 4675
rect 2605 4573 2639 4607
rect 3525 4573 3559 4607
rect 4077 4573 4111 4607
rect 6377 4573 6411 4607
rect 7205 4573 7239 4607
rect 7297 4573 7331 4607
rect 8217 4573 8251 4607
rect 8309 4573 8343 4607
rect 8953 4573 8987 4607
rect 10149 4573 10183 4607
rect 10241 4573 10275 4607
rect 11621 4573 11655 4607
rect 11989 4573 12023 4607
rect 14105 4573 14139 4607
rect 14289 4573 14323 4607
rect 15853 4573 15887 4607
rect 1961 4505 1995 4539
rect 1593 4437 1627 4471
rect 2973 4437 3007 4471
rect 5733 4437 5767 4471
rect 10977 4437 11011 4471
rect 15301 4437 15335 4471
rect 17509 4437 17543 4471
rect 18061 4437 18095 4471
rect 9137 4233 9171 4267
rect 15025 4233 15059 4267
rect 14749 4165 14783 4199
rect 5181 4097 5215 4131
rect 5917 4097 5951 4131
rect 7757 4097 7791 4131
rect 11805 4097 11839 4131
rect 11897 4097 11931 4131
rect 15577 4097 15611 4131
rect 1501 4029 1535 4063
rect 2053 4029 2087 4063
rect 3709 4029 3743 4063
rect 2320 3961 2354 3995
rect 3954 3961 3988 3995
rect 6837 4029 6871 4063
rect 9689 4029 9723 4063
rect 12449 4029 12483 4063
rect 13369 4029 13403 4063
rect 15485 4029 15519 4063
rect 17417 4029 17451 4063
rect 18061 4029 18095 4063
rect 7113 3961 7147 3995
rect 8024 3961 8058 3995
rect 9956 3961 9990 3995
rect 12725 3961 12759 3995
rect 13636 3961 13670 3995
rect 15393 3961 15427 3995
rect 1685 3893 1719 3927
rect 3433 3893 3467 3927
rect 5089 3893 5123 3927
rect 5181 3893 5215 3927
rect 5365 3893 5399 3927
rect 5733 3893 5767 3927
rect 5825 3893 5859 3927
rect 11069 3893 11103 3927
rect 11345 3893 11379 3927
rect 11713 3893 11747 3927
rect 17601 3893 17635 3927
rect 18245 3893 18279 3927
rect 2697 3689 2731 3723
rect 3157 3689 3191 3723
rect 4077 3689 4111 3723
rect 4537 3689 4571 3723
rect 6837 3689 6871 3723
rect 8493 3689 8527 3723
rect 11805 3689 11839 3723
rect 13737 3689 13771 3723
rect 14197 3689 14231 3723
rect 3065 3621 3099 3655
rect 5702 3621 5736 3655
rect 7358 3621 7392 3655
rect 9965 3621 9999 3655
rect 12326 3621 12360 3655
rect 1409 3553 1443 3587
rect 1961 3553 1995 3587
rect 4445 3553 4479 3587
rect 5457 3553 5491 3587
rect 7113 3553 7147 3587
rect 8769 3553 8803 3587
rect 9689 3553 9723 3587
rect 10425 3553 10459 3587
rect 10692 3553 10726 3587
rect 14105 3553 14139 3587
rect 15669 3553 15703 3587
rect 17141 3553 17175 3587
rect 17693 3553 17727 3587
rect 2237 3485 2271 3519
rect 3249 3485 3283 3519
rect 4721 3485 4755 3519
rect 8953 3485 8987 3519
rect 12081 3485 12115 3519
rect 14381 3485 14415 3519
rect 15761 3485 15795 3519
rect 15853 3485 15887 3519
rect 13461 3417 13495 3451
rect 15301 3417 15335 3451
rect 17877 3417 17911 3451
rect 1593 3349 1627 3383
rect 17325 3349 17359 3383
rect 7849 3145 7883 3179
rect 12265 3145 12299 3179
rect 14473 3145 14507 3179
rect 2145 3077 2179 3111
rect 6837 3077 6871 3111
rect 10885 3077 10919 3111
rect 2697 3009 2731 3043
rect 3801 3009 3835 3043
rect 4997 3009 5031 3043
rect 6009 3009 6043 3043
rect 7389 3009 7423 3043
rect 8401 3009 8435 3043
rect 9321 3009 9355 3043
rect 9505 3009 9539 3043
rect 10609 3009 10643 3043
rect 1409 2941 1443 2975
rect 1685 2941 1719 2975
rect 3617 2941 3651 2975
rect 4813 2941 4847 2975
rect 4905 2941 4939 2975
rect 5825 2941 5859 2975
rect 7205 2941 7239 2975
rect 8309 2941 8343 2975
rect 10425 2941 10459 2975
rect 11621 3009 11655 3043
rect 11437 2941 11471 2975
rect 2513 2873 2547 2907
rect 2605 2873 2639 2907
rect 3525 2873 3559 2907
rect 5917 2873 5951 2907
rect 7297 2873 7331 2907
rect 10517 2873 10551 2907
rect 10885 2873 10919 2907
rect 12449 3077 12483 3111
rect 13093 3009 13127 3043
rect 14013 3009 14047 3043
rect 15025 3009 15059 3043
rect 15669 3009 15703 3043
rect 15485 2941 15519 2975
rect 16405 2941 16439 2975
rect 16957 2941 16991 2975
rect 18061 2941 18095 2975
rect 12909 2873 12943 2907
rect 14933 2873 14967 2907
rect 3157 2805 3191 2839
rect 4445 2805 4479 2839
rect 5457 2805 5491 2839
rect 8217 2805 8251 2839
rect 8861 2805 8895 2839
rect 9229 2805 9263 2839
rect 10057 2805 10091 2839
rect 11069 2805 11103 2839
rect 11529 2805 11563 2839
rect 12265 2805 12299 2839
rect 12817 2805 12851 2839
rect 13461 2805 13495 2839
rect 13829 2805 13863 2839
rect 13921 2805 13955 2839
rect 14841 2805 14875 2839
rect 16589 2805 16623 2839
rect 17141 2805 17175 2839
rect 18245 2805 18279 2839
rect 3341 2601 3375 2635
rect 4077 2601 4111 2635
rect 4537 2601 4571 2635
rect 4905 2601 4939 2635
rect 8033 2601 8067 2635
rect 8677 2601 8711 2635
rect 9045 2601 9079 2635
rect 10149 2601 10183 2635
rect 11161 2601 11195 2635
rect 13001 2601 13035 2635
rect 13645 2601 13679 2635
rect 14013 2601 14047 2635
rect 14105 2601 14139 2635
rect 3433 2533 3467 2567
rect 6377 2533 6411 2567
rect 8125 2533 8159 2567
rect 10241 2533 10275 2567
rect 12081 2533 12115 2567
rect 13093 2533 13127 2567
rect 1593 2465 1627 2499
rect 2421 2465 2455 2499
rect 5733 2465 5767 2499
rect 6929 2465 6963 2499
rect 9137 2465 9171 2499
rect 11805 2465 11839 2499
rect 14657 2465 14691 2499
rect 15485 2465 15519 2499
rect 16221 2465 16255 2499
rect 16957 2465 16991 2499
rect 17693 2465 17727 2499
rect 1777 2397 1811 2431
rect 3617 2397 3651 2431
rect 4997 2397 5031 2431
rect 5181 2397 5215 2431
rect 7113 2397 7147 2431
rect 8217 2397 8251 2431
rect 9321 2397 9355 2431
rect 10333 2397 10367 2431
rect 11253 2397 11287 2431
rect 11345 2397 11379 2431
rect 13277 2397 13311 2431
rect 14197 2397 14231 2431
rect 14841 2397 14875 2431
rect 15209 2397 15243 2431
rect 15669 2397 15703 2431
rect 16405 2397 16439 2431
rect 2973 2329 3007 2363
rect 10793 2329 10827 2363
rect 12633 2329 12667 2363
rect 2605 2261 2639 2295
rect 7665 2261 7699 2295
rect 9781 2261 9815 2295
rect 15209 2261 15243 2295
rect 17141 2261 17175 2295
rect 17877 2261 17911 2295
<< metal1 >>
rect 3970 15308 3976 15360
rect 4028 15348 4034 15360
rect 6362 15348 6368 15360
rect 4028 15320 6368 15348
rect 4028 15308 4034 15320
rect 6362 15308 6368 15320
rect 6420 15308 6426 15360
rect 4062 15240 4068 15292
rect 4120 15280 4126 15292
rect 8846 15280 8852 15292
rect 4120 15252 8852 15280
rect 4120 15240 4126 15252
rect 8846 15240 8852 15252
rect 8904 15240 8910 15292
rect 3510 14968 3516 15020
rect 3568 15008 3574 15020
rect 6270 15008 6276 15020
rect 3568 14980 6276 15008
rect 3568 14968 3574 14980
rect 6270 14968 6276 14980
rect 6328 14968 6334 15020
rect 9030 14832 9036 14884
rect 9088 14872 9094 14884
rect 18230 14872 18236 14884
rect 9088 14844 18236 14872
rect 9088 14832 9094 14844
rect 18230 14832 18236 14844
rect 18288 14832 18294 14884
rect 3694 14764 3700 14816
rect 3752 14804 3758 14816
rect 11514 14804 11520 14816
rect 3752 14776 11520 14804
rect 3752 14764 3758 14776
rect 11514 14764 11520 14776
rect 11572 14764 11578 14816
rect 1104 14714 18860 14736
rect 1104 14662 6912 14714
rect 6964 14662 6976 14714
rect 7028 14662 7040 14714
rect 7092 14662 7104 14714
rect 7156 14662 12843 14714
rect 12895 14662 12907 14714
rect 12959 14662 12971 14714
rect 13023 14662 13035 14714
rect 13087 14662 18860 14714
rect 1104 14640 18860 14662
rect 6181 14603 6239 14609
rect 6181 14569 6193 14603
rect 6227 14600 6239 14603
rect 7653 14603 7711 14609
rect 7653 14600 7665 14603
rect 6227 14572 7665 14600
rect 6227 14569 6239 14572
rect 6181 14563 6239 14569
rect 7653 14569 7665 14572
rect 7699 14569 7711 14603
rect 9033 14603 9091 14609
rect 7653 14563 7711 14569
rect 8036 14572 8708 14600
rect 3786 14492 3792 14544
rect 3844 14532 3850 14544
rect 8036 14532 8064 14572
rect 3844 14504 8064 14532
rect 8113 14535 8171 14541
rect 3844 14492 3850 14504
rect 8113 14501 8125 14535
rect 8159 14532 8171 14535
rect 8570 14532 8576 14544
rect 8159 14504 8576 14532
rect 8159 14501 8171 14504
rect 8113 14495 8171 14501
rect 8570 14492 8576 14504
rect 8628 14492 8634 14544
rect 8680 14532 8708 14572
rect 9033 14569 9045 14603
rect 9079 14600 9091 14603
rect 10137 14603 10195 14609
rect 10137 14600 10149 14603
rect 9079 14572 10149 14600
rect 9079 14569 9091 14572
rect 9033 14563 9091 14569
rect 10137 14569 10149 14572
rect 10183 14569 10195 14603
rect 10137 14563 10195 14569
rect 13357 14603 13415 14609
rect 13357 14569 13369 14603
rect 13403 14600 13415 14603
rect 15470 14600 15476 14612
rect 13403 14572 15476 14600
rect 13403 14569 13415 14572
rect 13357 14563 13415 14569
rect 15470 14560 15476 14572
rect 15528 14560 15534 14612
rect 10505 14535 10563 14541
rect 10505 14532 10517 14535
rect 8680 14504 10517 14532
rect 10505 14501 10517 14504
rect 10551 14532 10563 14535
rect 11330 14532 11336 14544
rect 10551 14504 11336 14532
rect 10551 14501 10563 14504
rect 10505 14495 10563 14501
rect 11330 14492 11336 14504
rect 11388 14492 11394 14544
rect 14366 14492 14372 14544
rect 14424 14532 14430 14544
rect 16117 14535 16175 14541
rect 16117 14532 16129 14535
rect 14424 14504 16129 14532
rect 14424 14492 14430 14504
rect 8021 14467 8079 14473
rect 8021 14433 8033 14467
rect 8067 14464 8079 14467
rect 8662 14464 8668 14476
rect 8067 14436 8668 14464
rect 8067 14433 8079 14436
rect 8021 14427 8079 14433
rect 8662 14424 8668 14436
rect 8720 14424 8726 14476
rect 9125 14467 9183 14473
rect 9125 14433 9137 14467
rect 9171 14464 9183 14467
rect 9582 14464 9588 14476
rect 9171 14436 9588 14464
rect 9171 14433 9183 14436
rect 9125 14427 9183 14433
rect 9582 14424 9588 14436
rect 9640 14424 9646 14476
rect 11422 14424 11428 14476
rect 11480 14464 11486 14476
rect 11517 14467 11575 14473
rect 11517 14464 11529 14467
rect 11480 14436 11529 14464
rect 11480 14424 11486 14436
rect 11517 14433 11529 14436
rect 11563 14433 11575 14467
rect 11517 14427 11575 14433
rect 11609 14467 11667 14473
rect 11609 14433 11621 14467
rect 11655 14464 11667 14467
rect 11974 14464 11980 14476
rect 11655 14436 11980 14464
rect 11655 14433 11667 14436
rect 11609 14427 11667 14433
rect 11974 14424 11980 14436
rect 12032 14424 12038 14476
rect 12434 14424 12440 14476
rect 12492 14464 12498 14476
rect 13725 14467 13783 14473
rect 13725 14464 13737 14467
rect 12492 14436 13737 14464
rect 12492 14424 12498 14436
rect 13725 14433 13737 14436
rect 13771 14433 13783 14467
rect 14734 14464 14740 14476
rect 14695 14436 14740 14464
rect 13725 14427 13783 14433
rect 14734 14424 14740 14436
rect 14792 14424 14798 14476
rect 14829 14467 14887 14473
rect 14829 14433 14841 14467
rect 14875 14464 14887 14467
rect 15102 14464 15108 14476
rect 14875 14436 15108 14464
rect 14875 14433 14887 14436
rect 14829 14427 14887 14433
rect 6273 14399 6331 14405
rect 6273 14365 6285 14399
rect 6319 14365 6331 14399
rect 6273 14359 6331 14365
rect 6457 14399 6515 14405
rect 6457 14365 6469 14399
rect 6503 14396 6515 14399
rect 6733 14399 6791 14405
rect 6733 14396 6745 14399
rect 6503 14368 6745 14396
rect 6503 14365 6515 14368
rect 6457 14359 6515 14365
rect 6733 14365 6745 14368
rect 6779 14365 6791 14399
rect 8202 14396 8208 14408
rect 8163 14368 8208 14396
rect 6733 14359 6791 14365
rect 6288 14328 6316 14359
rect 8202 14356 8208 14368
rect 8260 14396 8266 14408
rect 9217 14399 9275 14405
rect 9217 14396 9229 14399
rect 8260 14368 9229 14396
rect 8260 14356 8266 14368
rect 9217 14365 9229 14368
rect 9263 14365 9275 14399
rect 10594 14396 10600 14408
rect 10555 14368 10600 14396
rect 9217 14359 9275 14365
rect 10594 14356 10600 14368
rect 10652 14356 10658 14408
rect 10778 14396 10784 14408
rect 10739 14368 10784 14396
rect 10778 14356 10784 14368
rect 10836 14356 10842 14408
rect 11054 14356 11060 14408
rect 11112 14396 11118 14408
rect 11701 14399 11759 14405
rect 11701 14396 11713 14399
rect 11112 14368 11713 14396
rect 11112 14356 11118 14368
rect 11701 14365 11713 14368
rect 11747 14365 11759 14399
rect 11701 14359 11759 14365
rect 12526 14356 12532 14408
rect 12584 14396 12590 14408
rect 13817 14399 13875 14405
rect 13817 14396 13829 14399
rect 12584 14368 13829 14396
rect 12584 14356 12590 14368
rect 13817 14365 13829 14368
rect 13863 14365 13875 14399
rect 13817 14359 13875 14365
rect 13909 14399 13967 14405
rect 13909 14365 13921 14399
rect 13955 14365 13967 14399
rect 14918 14396 14924 14408
rect 14879 14368 14924 14396
rect 13909 14359 13967 14365
rect 8665 14331 8723 14337
rect 8665 14328 8677 14331
rect 6288 14300 8677 14328
rect 8665 14297 8677 14300
rect 8711 14297 8723 14331
rect 8665 14291 8723 14297
rect 13722 14288 13728 14340
rect 13780 14328 13786 14340
rect 13924 14328 13952 14359
rect 14918 14356 14924 14368
rect 14976 14356 14982 14408
rect 13780 14300 13952 14328
rect 13780 14288 13786 14300
rect 14182 14288 14188 14340
rect 14240 14328 14246 14340
rect 15028 14328 15056 14436
rect 15102 14424 15108 14436
rect 15160 14424 15166 14476
rect 15396 14464 15424 14504
rect 16117 14501 16129 14504
rect 16163 14501 16175 14535
rect 16117 14495 16175 14501
rect 17037 14535 17095 14541
rect 17037 14501 17049 14535
rect 17083 14532 17095 14535
rect 18782 14532 18788 14544
rect 17083 14504 18788 14532
rect 17083 14501 17095 14504
rect 17037 14495 17095 14501
rect 18782 14492 18788 14504
rect 18840 14492 18846 14544
rect 15508 14467 15566 14473
rect 15508 14464 15520 14467
rect 15396 14436 15520 14464
rect 15508 14433 15520 14436
rect 15554 14433 15566 14467
rect 15508 14427 15566 14433
rect 15654 14356 15660 14408
rect 15712 14396 15718 14408
rect 16025 14399 16083 14405
rect 16025 14396 16037 14399
rect 15712 14368 16037 14396
rect 15712 14356 15718 14368
rect 16025 14365 16037 14368
rect 16071 14365 16083 14399
rect 16025 14359 16083 14365
rect 14240 14300 15056 14328
rect 14240 14288 14246 14300
rect 5718 14220 5724 14272
rect 5776 14260 5782 14272
rect 5813 14263 5871 14269
rect 5813 14260 5825 14263
rect 5776 14232 5825 14260
rect 5776 14220 5782 14232
rect 5813 14229 5825 14232
rect 5859 14229 5871 14263
rect 5813 14223 5871 14229
rect 6733 14263 6791 14269
rect 6733 14229 6745 14263
rect 6779 14260 6791 14263
rect 9766 14260 9772 14272
rect 6779 14232 9772 14260
rect 6779 14229 6791 14232
rect 6733 14223 6791 14229
rect 9766 14220 9772 14232
rect 9824 14220 9830 14272
rect 11146 14260 11152 14272
rect 11107 14232 11152 14260
rect 11146 14220 11152 14232
rect 11204 14220 11210 14272
rect 13538 14220 13544 14272
rect 13596 14260 13602 14272
rect 14369 14263 14427 14269
rect 14369 14260 14381 14263
rect 13596 14232 14381 14260
rect 13596 14220 13602 14232
rect 14369 14229 14381 14232
rect 14415 14229 14427 14263
rect 14369 14223 14427 14229
rect 15611 14263 15669 14269
rect 15611 14229 15623 14263
rect 15657 14260 15669 14263
rect 16206 14260 16212 14272
rect 15657 14232 16212 14260
rect 15657 14229 15669 14232
rect 15611 14223 15669 14229
rect 16206 14220 16212 14232
rect 16264 14220 16270 14272
rect 1104 14170 18860 14192
rect 1104 14118 3947 14170
rect 3999 14118 4011 14170
rect 4063 14118 4075 14170
rect 4127 14118 4139 14170
rect 4191 14118 9878 14170
rect 9930 14118 9942 14170
rect 9994 14118 10006 14170
rect 10058 14118 10070 14170
rect 10122 14118 15808 14170
rect 15860 14118 15872 14170
rect 15924 14118 15936 14170
rect 15988 14118 16000 14170
rect 16052 14118 18860 14170
rect 1104 14096 18860 14118
rect 3418 14016 3424 14068
rect 3476 14056 3482 14068
rect 8573 14059 8631 14065
rect 3476 14028 8432 14056
rect 3476 14016 3482 14028
rect 3326 13948 3332 14000
rect 3384 13988 3390 14000
rect 5169 13991 5227 13997
rect 5169 13988 5181 13991
rect 3384 13960 5181 13988
rect 3384 13948 3390 13960
rect 5169 13957 5181 13960
rect 5215 13957 5227 13991
rect 5169 13951 5227 13957
rect 6825 13991 6883 13997
rect 6825 13957 6837 13991
rect 6871 13988 6883 13991
rect 8294 13988 8300 14000
rect 6871 13960 8300 13988
rect 6871 13957 6883 13960
rect 6825 13951 6883 13957
rect 8294 13948 8300 13960
rect 8352 13948 8358 14000
rect 8404 13988 8432 14028
rect 8573 14025 8585 14059
rect 8619 14056 8631 14059
rect 8662 14056 8668 14068
rect 8619 14028 8668 14056
rect 8619 14025 8631 14028
rect 8573 14019 8631 14025
rect 8662 14016 8668 14028
rect 8720 14016 8726 14068
rect 9582 14056 9588 14068
rect 9543 14028 9588 14056
rect 9582 14016 9588 14028
rect 9640 14016 9646 14068
rect 10594 14056 10600 14068
rect 10555 14028 10600 14056
rect 10594 14016 10600 14028
rect 10652 14016 10658 14068
rect 12066 14016 12072 14068
rect 12124 14056 12130 14068
rect 15013 14059 15071 14065
rect 15013 14056 15025 14059
rect 12124 14028 15025 14056
rect 12124 14016 12130 14028
rect 15013 14025 15025 14028
rect 15059 14025 15071 14059
rect 15013 14019 15071 14025
rect 18233 13991 18291 13997
rect 8404 13960 18092 13988
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 5721 13923 5779 13929
rect 5721 13920 5733 13923
rect 5500 13892 5733 13920
rect 5500 13880 5506 13892
rect 5721 13889 5733 13892
rect 5767 13889 5779 13923
rect 5721 13883 5779 13889
rect 7469 13923 7527 13929
rect 7469 13889 7481 13923
rect 7515 13920 7527 13923
rect 8754 13920 8760 13932
rect 7515 13892 8760 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 8938 13880 8944 13932
rect 8996 13880 9002 13932
rect 9217 13923 9275 13929
rect 9217 13889 9229 13923
rect 9263 13920 9275 13923
rect 9674 13920 9680 13932
rect 9263 13892 9680 13920
rect 9263 13889 9275 13892
rect 9217 13883 9275 13889
rect 9674 13880 9680 13892
rect 9732 13920 9738 13932
rect 10229 13923 10287 13929
rect 10229 13920 10241 13923
rect 9732 13892 10241 13920
rect 9732 13880 9738 13892
rect 10229 13889 10241 13892
rect 10275 13920 10287 13923
rect 10778 13920 10784 13932
rect 10275 13892 10784 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 10778 13880 10784 13892
rect 10836 13880 10842 13932
rect 10870 13880 10876 13932
rect 10928 13920 10934 13932
rect 11149 13923 11207 13929
rect 11149 13920 11161 13923
rect 10928 13892 11161 13920
rect 10928 13880 10934 13892
rect 11149 13889 11161 13892
rect 11195 13889 11207 13923
rect 11149 13883 11207 13889
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 12158 13920 12164 13932
rect 11931 13892 12164 13920
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 12158 13880 12164 13892
rect 12216 13880 12222 13932
rect 13725 13923 13783 13929
rect 13725 13889 13737 13923
rect 13771 13920 13783 13923
rect 14366 13920 14372 13932
rect 13771 13892 14372 13920
rect 13771 13889 13783 13892
rect 13725 13883 13783 13889
rect 14366 13880 14372 13892
rect 14424 13880 14430 13932
rect 15657 13923 15715 13929
rect 15657 13889 15669 13923
rect 15703 13920 15715 13923
rect 15930 13920 15936 13932
rect 15703 13892 15936 13920
rect 15703 13889 15715 13892
rect 15657 13883 15715 13889
rect 15930 13880 15936 13892
rect 15988 13880 15994 13932
rect 16117 13923 16175 13929
rect 16117 13889 16129 13923
rect 16163 13920 16175 13923
rect 16574 13920 16580 13932
rect 16163 13892 16580 13920
rect 16163 13889 16175 13892
rect 16117 13883 16175 13889
rect 16574 13880 16580 13892
rect 16632 13880 16638 13932
rect 17126 13920 17132 13932
rect 17087 13892 17132 13920
rect 17126 13880 17132 13892
rect 17184 13880 17190 13932
rect 7285 13855 7343 13861
rect 7285 13821 7297 13855
rect 7331 13852 7343 13855
rect 8110 13852 8116 13864
rect 7331 13824 8116 13852
rect 7331 13821 7343 13824
rect 7285 13815 7343 13821
rect 8110 13812 8116 13824
rect 8168 13812 8174 13864
rect 7193 13787 7251 13793
rect 7193 13753 7205 13787
rect 7239 13784 7251 13787
rect 8662 13784 8668 13796
rect 7239 13756 8668 13784
rect 7239 13753 7251 13756
rect 7193 13747 7251 13753
rect 8662 13744 8668 13756
rect 8720 13744 8726 13796
rect 8956 13793 8984 13880
rect 9306 13852 9312 13864
rect 9048 13824 9312 13852
rect 9048 13793 9076 13824
rect 9306 13812 9312 13824
rect 9364 13812 9370 13864
rect 10502 13812 10508 13864
rect 10560 13852 10566 13864
rect 11057 13855 11115 13861
rect 11057 13852 11069 13855
rect 10560 13824 11069 13852
rect 10560 13812 10566 13824
rect 11057 13821 11069 13824
rect 11103 13821 11115 13855
rect 11606 13852 11612 13864
rect 11567 13824 11612 13852
rect 11057 13815 11115 13821
rect 11606 13812 11612 13824
rect 11664 13812 11670 13864
rect 13081 13855 13139 13861
rect 13081 13821 13093 13855
rect 13127 13852 13139 13855
rect 13170 13852 13176 13864
rect 13127 13824 13176 13852
rect 13127 13821 13139 13824
rect 13081 13815 13139 13821
rect 13170 13812 13176 13824
rect 13228 13812 13234 13864
rect 13446 13852 13452 13864
rect 13407 13824 13452 13852
rect 13446 13812 13452 13824
rect 13504 13812 13510 13864
rect 15473 13855 15531 13861
rect 15473 13821 15485 13855
rect 15519 13852 15531 13855
rect 17402 13852 17408 13864
rect 15519 13824 15608 13852
rect 17363 13824 17408 13852
rect 15519 13821 15531 13824
rect 15473 13815 15531 13821
rect 8941 13787 8999 13793
rect 8941 13753 8953 13787
rect 8987 13753 8999 13787
rect 8941 13747 8999 13753
rect 9033 13787 9091 13793
rect 9033 13753 9045 13787
rect 9079 13753 9091 13787
rect 9033 13747 9091 13753
rect 10226 13744 10232 13796
rect 10284 13784 10290 13796
rect 13464 13784 13492 13812
rect 15580 13796 15608 13824
rect 17402 13812 17408 13824
rect 17460 13812 17466 13864
rect 18064 13861 18092 13960
rect 18233 13957 18245 13991
rect 18279 13988 18291 13991
rect 18506 13988 18512 14000
rect 18279 13960 18512 13988
rect 18279 13957 18291 13960
rect 18233 13951 18291 13957
rect 18506 13948 18512 13960
rect 18564 13948 18570 14000
rect 18049 13855 18107 13861
rect 18049 13821 18061 13855
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 10284 13756 13492 13784
rect 10284 13744 10290 13756
rect 15562 13744 15568 13796
rect 15620 13744 15626 13796
rect 16206 13744 16212 13796
rect 16264 13784 16270 13796
rect 16264 13756 16309 13784
rect 16264 13744 16270 13756
rect 5534 13716 5540 13728
rect 5495 13688 5540 13716
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 5626 13676 5632 13728
rect 5684 13716 5690 13728
rect 5684 13688 5729 13716
rect 5684 13676 5690 13688
rect 6362 13676 6368 13728
rect 6420 13716 6426 13728
rect 9490 13716 9496 13728
rect 6420 13688 9496 13716
rect 6420 13676 6426 13688
rect 9490 13676 9496 13688
rect 9548 13676 9554 13728
rect 9950 13716 9956 13728
rect 9911 13688 9956 13716
rect 9950 13676 9956 13688
rect 10008 13676 10014 13728
rect 10045 13719 10103 13725
rect 10045 13685 10057 13719
rect 10091 13716 10103 13719
rect 10318 13716 10324 13728
rect 10091 13688 10324 13716
rect 10091 13685 10103 13688
rect 10045 13679 10103 13685
rect 10318 13676 10324 13688
rect 10376 13676 10382 13728
rect 10594 13676 10600 13728
rect 10652 13716 10658 13728
rect 10965 13719 11023 13725
rect 10965 13716 10977 13719
rect 10652 13688 10977 13716
rect 10652 13676 10658 13688
rect 10965 13685 10977 13688
rect 11011 13685 11023 13719
rect 10965 13679 11023 13685
rect 11238 13676 11244 13728
rect 11296 13716 11302 13728
rect 11698 13716 11704 13728
rect 11296 13688 11704 13716
rect 11296 13676 11302 13688
rect 11698 13676 11704 13688
rect 11756 13716 11762 13728
rect 13906 13716 13912 13728
rect 11756 13688 13912 13716
rect 11756 13676 11762 13688
rect 13906 13676 13912 13688
rect 13964 13676 13970 13728
rect 15194 13676 15200 13728
rect 15252 13716 15258 13728
rect 15381 13719 15439 13725
rect 15381 13716 15393 13719
rect 15252 13688 15393 13716
rect 15252 13676 15258 13688
rect 15381 13685 15393 13688
rect 15427 13685 15439 13719
rect 17586 13716 17592 13728
rect 17547 13688 17592 13716
rect 15381 13679 15439 13685
rect 17586 13676 17592 13688
rect 17644 13676 17650 13728
rect 1104 13626 18860 13648
rect 1104 13574 6912 13626
rect 6964 13574 6976 13626
rect 7028 13574 7040 13626
rect 7092 13574 7104 13626
rect 7156 13574 12843 13626
rect 12895 13574 12907 13626
rect 12959 13574 12971 13626
rect 13023 13574 13035 13626
rect 13087 13574 18860 13626
rect 1104 13552 18860 13574
rect 5534 13472 5540 13524
rect 5592 13512 5598 13524
rect 5629 13515 5687 13521
rect 5629 13512 5641 13515
rect 5592 13484 5641 13512
rect 5592 13472 5598 13484
rect 5629 13481 5641 13484
rect 5675 13481 5687 13515
rect 8021 13515 8079 13521
rect 8021 13512 8033 13515
rect 5629 13475 5687 13481
rect 6564 13484 8033 13512
rect 5074 13336 5080 13388
rect 5132 13376 5138 13388
rect 5997 13379 6055 13385
rect 5997 13376 6009 13379
rect 5132 13348 6009 13376
rect 5132 13336 5138 13348
rect 5997 13345 6009 13348
rect 6043 13345 6055 13379
rect 5997 13339 6055 13345
rect 6089 13379 6147 13385
rect 6089 13345 6101 13379
rect 6135 13376 6147 13379
rect 6454 13376 6460 13388
rect 6135 13348 6460 13376
rect 6135 13345 6147 13348
rect 6089 13339 6147 13345
rect 6454 13336 6460 13348
rect 6512 13336 6518 13388
rect 4062 13268 4068 13320
rect 4120 13308 4126 13320
rect 5810 13308 5816 13320
rect 4120 13280 5816 13308
rect 4120 13268 4126 13280
rect 5810 13268 5816 13280
rect 5868 13268 5874 13320
rect 6178 13268 6184 13320
rect 6236 13308 6242 13320
rect 6273 13311 6331 13317
rect 6273 13308 6285 13311
rect 6236 13280 6285 13308
rect 6236 13268 6242 13280
rect 6273 13277 6285 13280
rect 6319 13308 6331 13311
rect 6564 13308 6592 13484
rect 8021 13481 8033 13484
rect 8067 13481 8079 13515
rect 8570 13512 8576 13524
rect 8531 13484 8576 13512
rect 8021 13475 8079 13481
rect 8570 13472 8576 13484
rect 8628 13472 8634 13524
rect 8938 13472 8944 13524
rect 8996 13512 9002 13524
rect 9677 13515 9735 13521
rect 9677 13512 9689 13515
rect 8996 13484 9689 13512
rect 8996 13472 9002 13484
rect 9677 13481 9689 13484
rect 9723 13481 9735 13515
rect 9677 13475 9735 13481
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 10505 13515 10563 13521
rect 10505 13512 10517 13515
rect 10008 13484 10517 13512
rect 10008 13472 10014 13484
rect 10505 13481 10517 13484
rect 10551 13481 10563 13515
rect 10505 13475 10563 13481
rect 10873 13515 10931 13521
rect 10873 13481 10885 13515
rect 10919 13512 10931 13515
rect 11238 13512 11244 13524
rect 10919 13484 11244 13512
rect 10919 13481 10931 13484
rect 10873 13475 10931 13481
rect 11238 13472 11244 13484
rect 11296 13472 11302 13524
rect 12161 13515 12219 13521
rect 12161 13481 12173 13515
rect 12207 13512 12219 13515
rect 12526 13512 12532 13524
rect 12207 13484 12532 13512
rect 12207 13481 12219 13484
rect 12161 13475 12219 13481
rect 12526 13472 12532 13484
rect 12584 13472 12590 13524
rect 12621 13515 12679 13521
rect 12621 13481 12633 13515
rect 12667 13512 12679 13515
rect 14185 13515 14243 13521
rect 14185 13512 14197 13515
rect 12667 13484 14197 13512
rect 12667 13481 12679 13484
rect 12621 13475 12679 13481
rect 14185 13481 14197 13484
rect 14231 13481 14243 13515
rect 14185 13475 14243 13481
rect 14553 13515 14611 13521
rect 14553 13481 14565 13515
rect 14599 13512 14611 13515
rect 15473 13515 15531 13521
rect 15473 13512 15485 13515
rect 14599 13484 15485 13512
rect 14599 13481 14611 13484
rect 14553 13475 14611 13481
rect 15473 13481 15485 13484
rect 15519 13481 15531 13515
rect 15473 13475 15531 13481
rect 7834 13404 7840 13456
rect 7892 13444 7898 13456
rect 11882 13444 11888 13456
rect 7892 13416 11888 13444
rect 7892 13404 7898 13416
rect 11882 13404 11888 13416
rect 11940 13404 11946 13456
rect 14642 13444 14648 13456
rect 11992 13416 13308 13444
rect 14603 13416 14648 13444
rect 6908 13379 6966 13385
rect 6908 13345 6920 13379
rect 6954 13376 6966 13379
rect 7466 13376 7472 13388
rect 6954 13348 7472 13376
rect 6954 13345 6966 13348
rect 6908 13339 6966 13345
rect 7466 13336 7472 13348
rect 7524 13336 7530 13388
rect 8846 13336 8852 13388
rect 8904 13376 8910 13388
rect 8941 13379 8999 13385
rect 8941 13376 8953 13379
rect 8904 13348 8953 13376
rect 8904 13336 8910 13348
rect 8941 13345 8953 13348
rect 8987 13345 8999 13379
rect 8941 13339 8999 13345
rect 9033 13379 9091 13385
rect 9033 13345 9045 13379
rect 9079 13376 9091 13379
rect 9398 13376 9404 13388
rect 9079 13348 9404 13376
rect 9079 13345 9091 13348
rect 9033 13339 9091 13345
rect 9398 13336 9404 13348
rect 9456 13336 9462 13388
rect 9490 13336 9496 13388
rect 9548 13376 9554 13388
rect 11992 13376 12020 13416
rect 13280 13388 13308 13416
rect 14642 13404 14648 13416
rect 14700 13404 14706 13456
rect 14826 13404 14832 13456
rect 14884 13444 14890 13456
rect 15933 13447 15991 13453
rect 15933 13444 15945 13447
rect 14884 13416 15945 13444
rect 14884 13404 14890 13416
rect 15933 13413 15945 13416
rect 15979 13413 15991 13447
rect 15933 13407 15991 13413
rect 16298 13404 16304 13456
rect 16356 13444 16362 13456
rect 17957 13447 18015 13453
rect 17957 13444 17969 13447
rect 16356 13416 17969 13444
rect 16356 13404 16362 13416
rect 17957 13413 17969 13416
rect 18003 13444 18015 13447
rect 18322 13444 18328 13456
rect 18003 13416 18328 13444
rect 18003 13413 18015 13416
rect 17957 13407 18015 13413
rect 18322 13404 18328 13416
rect 18380 13404 18386 13456
rect 9548 13348 12020 13376
rect 9548 13336 9554 13348
rect 12434 13336 12440 13388
rect 12492 13376 12498 13388
rect 12529 13379 12587 13385
rect 12529 13376 12541 13379
rect 12492 13348 12541 13376
rect 12492 13336 12498 13348
rect 12529 13345 12541 13348
rect 12575 13345 12587 13379
rect 12529 13339 12587 13345
rect 13262 13336 13268 13388
rect 13320 13376 13326 13388
rect 13541 13379 13599 13385
rect 13541 13376 13553 13379
rect 13320 13348 13553 13376
rect 13320 13336 13326 13348
rect 13541 13345 13553 13348
rect 13587 13345 13599 13379
rect 13541 13339 13599 13345
rect 13906 13336 13912 13388
rect 13964 13376 13970 13388
rect 15841 13379 15899 13385
rect 15841 13376 15853 13379
rect 13964 13348 15853 13376
rect 13964 13336 13970 13348
rect 15841 13345 15853 13348
rect 15887 13345 15899 13379
rect 15841 13339 15899 13345
rect 16574 13336 16580 13388
rect 16632 13376 16638 13388
rect 16853 13379 16911 13385
rect 16853 13376 16865 13379
rect 16632 13348 16865 13376
rect 16632 13336 16638 13348
rect 16853 13345 16865 13348
rect 16899 13345 16911 13379
rect 16853 13339 16911 13345
rect 16945 13379 17003 13385
rect 16945 13345 16957 13379
rect 16991 13376 17003 13379
rect 17862 13376 17868 13388
rect 16991 13348 17264 13376
rect 17823 13348 17868 13376
rect 16991 13345 17003 13348
rect 16945 13339 17003 13345
rect 6319 13280 6592 13308
rect 6641 13311 6699 13317
rect 6319 13277 6331 13280
rect 6273 13271 6331 13277
rect 6641 13277 6653 13311
rect 6687 13277 6699 13311
rect 6641 13271 6699 13277
rect 6656 13172 6684 13271
rect 7650 13268 7656 13320
rect 7708 13308 7714 13320
rect 9217 13311 9275 13317
rect 7708 13280 9168 13308
rect 7708 13268 7714 13280
rect 9140 13240 9168 13280
rect 9217 13277 9229 13311
rect 9263 13308 9275 13311
rect 9674 13308 9680 13320
rect 9263 13280 9680 13308
rect 9263 13277 9275 13280
rect 9217 13271 9275 13277
rect 9674 13268 9680 13280
rect 9732 13268 9738 13320
rect 10962 13308 10968 13320
rect 10923 13280 10968 13308
rect 10962 13268 10968 13280
rect 11020 13268 11026 13320
rect 11057 13311 11115 13317
rect 11057 13277 11069 13311
rect 11103 13277 11115 13311
rect 11057 13271 11115 13277
rect 12805 13311 12863 13317
rect 12805 13277 12817 13311
rect 12851 13308 12863 13311
rect 12894 13308 12900 13320
rect 12851 13280 12900 13308
rect 12851 13277 12863 13280
rect 12805 13271 12863 13277
rect 10686 13240 10692 13252
rect 9140 13212 10692 13240
rect 10686 13200 10692 13212
rect 10744 13200 10750 13252
rect 10870 13200 10876 13252
rect 10928 13240 10934 13252
rect 11072 13240 11100 13271
rect 12894 13268 12900 13280
rect 12952 13268 12958 13320
rect 13630 13308 13636 13320
rect 13591 13280 13636 13308
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 13814 13308 13820 13320
rect 13727 13280 13820 13308
rect 13814 13268 13820 13280
rect 13872 13308 13878 13320
rect 14829 13311 14887 13317
rect 14829 13308 14841 13311
rect 13872 13280 14841 13308
rect 13872 13268 13878 13280
rect 14829 13277 14841 13280
rect 14875 13308 14887 13311
rect 14918 13308 14924 13320
rect 14875 13280 14924 13308
rect 14875 13277 14887 13280
rect 14829 13271 14887 13277
rect 14918 13268 14924 13280
rect 14976 13268 14982 13320
rect 15930 13268 15936 13320
rect 15988 13308 15994 13320
rect 16117 13311 16175 13317
rect 16117 13308 16129 13311
rect 15988 13280 16129 13308
rect 15988 13268 15994 13280
rect 16117 13277 16129 13280
rect 16163 13308 16175 13311
rect 17034 13308 17040 13320
rect 16163 13280 17040 13308
rect 16163 13277 16175 13280
rect 16117 13271 16175 13277
rect 17034 13268 17040 13280
rect 17092 13308 17098 13320
rect 17092 13280 17137 13308
rect 17092 13268 17098 13280
rect 10928 13212 11100 13240
rect 10928 13200 10934 13212
rect 11882 13200 11888 13252
rect 11940 13240 11946 13252
rect 13648 13240 13676 13268
rect 11940 13212 13676 13240
rect 11940 13200 11946 13212
rect 14642 13200 14648 13252
rect 14700 13240 14706 13252
rect 16485 13243 16543 13249
rect 16485 13240 16497 13243
rect 14700 13212 16497 13240
rect 14700 13200 14706 13212
rect 16485 13209 16497 13212
rect 16531 13209 16543 13243
rect 17236 13240 17264 13348
rect 17862 13336 17868 13348
rect 17920 13336 17926 13388
rect 18141 13311 18199 13317
rect 18141 13277 18153 13311
rect 18187 13308 18199 13311
rect 18322 13308 18328 13320
rect 18187 13280 18328 13308
rect 18187 13277 18199 13280
rect 18141 13271 18199 13277
rect 18322 13268 18328 13280
rect 18380 13268 18386 13320
rect 16485 13203 16543 13209
rect 16592 13212 17264 13240
rect 6914 13172 6920 13184
rect 6656 13144 6920 13172
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 9122 13132 9128 13184
rect 9180 13172 9186 13184
rect 10226 13172 10232 13184
rect 9180 13144 10232 13172
rect 9180 13132 9186 13144
rect 10226 13132 10232 13144
rect 10284 13132 10290 13184
rect 11790 13132 11796 13184
rect 11848 13172 11854 13184
rect 13173 13175 13231 13181
rect 13173 13172 13185 13175
rect 11848 13144 13185 13172
rect 11848 13132 11854 13144
rect 13173 13141 13185 13144
rect 13219 13141 13231 13175
rect 13173 13135 13231 13141
rect 14550 13132 14556 13184
rect 14608 13172 14614 13184
rect 16592 13172 16620 13212
rect 14608 13144 16620 13172
rect 14608 13132 14614 13144
rect 17218 13132 17224 13184
rect 17276 13172 17282 13184
rect 17497 13175 17555 13181
rect 17497 13172 17509 13175
rect 17276 13144 17509 13172
rect 17276 13132 17282 13144
rect 17497 13141 17509 13144
rect 17543 13141 17555 13175
rect 17497 13135 17555 13141
rect 1104 13082 18860 13104
rect 1104 13030 3947 13082
rect 3999 13030 4011 13082
rect 4063 13030 4075 13082
rect 4127 13030 4139 13082
rect 4191 13030 9878 13082
rect 9930 13030 9942 13082
rect 9994 13030 10006 13082
rect 10058 13030 10070 13082
rect 10122 13030 15808 13082
rect 15860 13030 15872 13082
rect 15924 13030 15936 13082
rect 15988 13030 16000 13082
rect 16052 13030 18860 13082
rect 1104 13008 18860 13030
rect 3510 12928 3516 12980
rect 3568 12968 3574 12980
rect 5537 12971 5595 12977
rect 3568 12940 5212 12968
rect 3568 12928 3574 12940
rect 5184 12900 5212 12940
rect 5537 12937 5549 12971
rect 5583 12968 5595 12971
rect 5626 12968 5632 12980
rect 5583 12940 5632 12968
rect 5583 12937 5595 12940
rect 5537 12931 5595 12937
rect 5626 12928 5632 12940
rect 5684 12928 5690 12980
rect 6840 12940 7880 12968
rect 6086 12900 6092 12912
rect 5184 12872 6092 12900
rect 6086 12860 6092 12872
rect 6144 12900 6150 12912
rect 6730 12900 6736 12912
rect 6144 12872 6736 12900
rect 6144 12860 6150 12872
rect 6730 12860 6736 12872
rect 6788 12860 6794 12912
rect 5074 12832 5080 12844
rect 5035 12804 5080 12832
rect 5074 12792 5080 12804
rect 5132 12792 5138 12844
rect 5994 12832 6000 12844
rect 5955 12804 6000 12832
rect 5994 12792 6000 12804
rect 6052 12792 6058 12844
rect 6178 12832 6184 12844
rect 6139 12804 6184 12832
rect 6178 12792 6184 12804
rect 6236 12832 6242 12844
rect 6638 12832 6644 12844
rect 6236 12804 6644 12832
rect 6236 12792 6242 12804
rect 6638 12792 6644 12804
rect 6696 12792 6702 12844
rect 3145 12767 3203 12773
rect 3145 12733 3157 12767
rect 3191 12764 3203 12767
rect 3694 12764 3700 12776
rect 3191 12736 3700 12764
rect 3191 12733 3203 12736
rect 3145 12727 3203 12733
rect 3694 12724 3700 12736
rect 3752 12724 3758 12776
rect 3970 12724 3976 12776
rect 4028 12764 4034 12776
rect 6840 12764 6868 12940
rect 7852 12900 7880 12940
rect 8018 12928 8024 12980
rect 8076 12968 8082 12980
rect 8297 12971 8355 12977
rect 8297 12968 8309 12971
rect 8076 12940 8309 12968
rect 8076 12928 8082 12940
rect 8297 12937 8309 12940
rect 8343 12937 8355 12971
rect 10318 12968 10324 12980
rect 8297 12931 8355 12937
rect 8404 12940 9536 12968
rect 10279 12940 10324 12968
rect 8404 12900 8432 12940
rect 7852 12872 8432 12900
rect 9508 12900 9536 12940
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 11333 12971 11391 12977
rect 11333 12937 11345 12971
rect 11379 12968 11391 12971
rect 12342 12968 12348 12980
rect 11379 12940 12348 12968
rect 11379 12937 11391 12940
rect 11333 12931 11391 12937
rect 12342 12928 12348 12940
rect 12400 12928 12406 12980
rect 12452 12940 13400 12968
rect 10686 12900 10692 12912
rect 9508 12872 10692 12900
rect 10686 12860 10692 12872
rect 10744 12860 10750 12912
rect 12452 12900 12480 12940
rect 10980 12872 12480 12900
rect 13372 12900 13400 12940
rect 13446 12928 13452 12980
rect 13504 12968 13510 12980
rect 13817 12971 13875 12977
rect 13817 12968 13829 12971
rect 13504 12940 13829 12968
rect 13504 12928 13510 12940
rect 13817 12937 13829 12940
rect 13863 12937 13875 12971
rect 13817 12931 13875 12937
rect 14550 12900 14556 12912
rect 13372 12872 14556 12900
rect 10410 12792 10416 12844
rect 10468 12832 10474 12844
rect 10870 12832 10876 12844
rect 10468 12804 10876 12832
rect 10468 12792 10474 12804
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 4028 12736 6868 12764
rect 4028 12724 4034 12736
rect 6914 12724 6920 12776
rect 6972 12764 6978 12776
rect 7184 12767 7242 12773
rect 6972 12736 7065 12764
rect 6972 12724 6978 12736
rect 7184 12733 7196 12767
rect 7230 12764 7242 12767
rect 7742 12764 7748 12776
rect 7230 12736 7748 12764
rect 7230 12733 7242 12736
rect 7184 12727 7242 12733
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 8573 12767 8631 12773
rect 8573 12764 8585 12767
rect 7944 12736 8585 12764
rect 3412 12699 3470 12705
rect 3412 12665 3424 12699
rect 3458 12696 3470 12699
rect 5442 12696 5448 12708
rect 3458 12668 5448 12696
rect 3458 12665 3470 12668
rect 3412 12659 3470 12665
rect 5442 12656 5448 12668
rect 5500 12656 5506 12708
rect 5905 12699 5963 12705
rect 5905 12665 5917 12699
rect 5951 12696 5963 12699
rect 6362 12696 6368 12708
rect 5951 12668 6368 12696
rect 5951 12665 5963 12668
rect 5905 12659 5963 12665
rect 6362 12656 6368 12668
rect 6420 12656 6426 12708
rect 6932 12696 6960 12724
rect 7944 12708 7972 12736
rect 8573 12733 8585 12736
rect 8619 12733 8631 12767
rect 8573 12727 8631 12733
rect 8840 12767 8898 12773
rect 8840 12733 8852 12767
rect 8886 12764 8898 12767
rect 9674 12764 9680 12776
rect 8886 12736 9680 12764
rect 8886 12733 8898 12736
rect 8840 12727 8898 12733
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 10226 12724 10232 12776
rect 10284 12764 10290 12776
rect 10689 12767 10747 12773
rect 10689 12764 10701 12767
rect 10284 12736 10701 12764
rect 10284 12724 10290 12736
rect 10689 12733 10701 12736
rect 10735 12733 10747 12767
rect 10980 12764 11008 12872
rect 14550 12860 14556 12872
rect 14608 12860 14614 12912
rect 11790 12832 11796 12844
rect 11751 12804 11796 12832
rect 11790 12792 11796 12804
rect 11848 12792 11854 12844
rect 11977 12835 12035 12841
rect 11977 12801 11989 12835
rect 12023 12832 12035 12835
rect 12023 12804 12572 12832
rect 12023 12801 12035 12804
rect 11977 12795 12035 12801
rect 10689 12727 10747 12733
rect 10796 12736 11008 12764
rect 12437 12767 12495 12773
rect 7926 12696 7932 12708
rect 6932 12668 7932 12696
rect 7926 12656 7932 12668
rect 7984 12656 7990 12708
rect 10796 12705 10824 12736
rect 12437 12733 12449 12767
rect 12483 12733 12495 12767
rect 12544 12764 12572 12804
rect 16666 12792 16672 12844
rect 16724 12832 16730 12844
rect 17405 12835 17463 12841
rect 17405 12832 17417 12835
rect 16724 12804 17417 12832
rect 16724 12792 16730 12804
rect 17405 12801 17417 12804
rect 17451 12801 17463 12835
rect 17405 12795 17463 12801
rect 14918 12764 14924 12776
rect 12544 12736 12940 12764
rect 14879 12736 14924 12764
rect 12437 12727 12495 12733
rect 10781 12699 10839 12705
rect 10781 12696 10793 12699
rect 8128 12668 10793 12696
rect 2498 12628 2504 12640
rect 2459 12600 2504 12628
rect 2498 12588 2504 12600
rect 2556 12588 2562 12640
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 4525 12631 4583 12637
rect 4525 12628 4537 12631
rect 4212 12600 4537 12628
rect 4212 12588 4218 12600
rect 4525 12597 4537 12600
rect 4571 12597 4583 12631
rect 4525 12591 4583 12597
rect 7742 12588 7748 12640
rect 7800 12628 7806 12640
rect 8128 12628 8156 12668
rect 10781 12665 10793 12668
rect 10827 12665 10839 12699
rect 10781 12659 10839 12665
rect 10870 12656 10876 12708
rect 10928 12696 10934 12708
rect 11422 12696 11428 12708
rect 10928 12668 11428 12696
rect 10928 12656 10934 12668
rect 11422 12656 11428 12668
rect 11480 12656 11486 12708
rect 11701 12699 11759 12705
rect 11701 12665 11713 12699
rect 11747 12696 11759 12699
rect 12452 12696 12480 12727
rect 12912 12708 12940 12736
rect 14918 12724 14924 12736
rect 14976 12724 14982 12776
rect 15010 12724 15016 12776
rect 15068 12764 15074 12776
rect 15188 12767 15246 12773
rect 15188 12764 15200 12767
rect 15068 12736 15200 12764
rect 15068 12724 15074 12736
rect 15188 12733 15200 12736
rect 15234 12764 15246 12767
rect 16942 12764 16948 12776
rect 15234 12736 16948 12764
rect 15234 12733 15246 12736
rect 15188 12727 15246 12733
rect 16942 12724 16948 12736
rect 17000 12724 17006 12776
rect 17218 12764 17224 12776
rect 17179 12736 17224 12764
rect 17218 12724 17224 12736
rect 17276 12724 17282 12776
rect 12526 12696 12532 12708
rect 11747 12668 12112 12696
rect 12452 12668 12532 12696
rect 11747 12665 11759 12668
rect 11701 12659 11759 12665
rect 7800 12600 8156 12628
rect 7800 12588 7806 12600
rect 8202 12588 8208 12640
rect 8260 12628 8266 12640
rect 9953 12631 10011 12637
rect 9953 12628 9965 12631
rect 8260 12600 9965 12628
rect 8260 12588 8266 12600
rect 9953 12597 9965 12600
rect 9999 12597 10011 12631
rect 12084 12628 12112 12668
rect 12526 12656 12532 12668
rect 12584 12656 12590 12708
rect 12704 12699 12762 12705
rect 12704 12665 12716 12699
rect 12750 12696 12762 12699
rect 12802 12696 12808 12708
rect 12750 12668 12808 12696
rect 12750 12665 12762 12668
rect 12704 12659 12762 12665
rect 12802 12656 12808 12668
rect 12860 12656 12866 12708
rect 12894 12656 12900 12708
rect 12952 12696 12958 12708
rect 12952 12668 13676 12696
rect 12952 12656 12958 12668
rect 13648 12640 13676 12668
rect 16574 12656 16580 12708
rect 16632 12696 16638 12708
rect 17586 12696 17592 12708
rect 16632 12668 17592 12696
rect 16632 12656 16638 12668
rect 17586 12656 17592 12668
rect 17644 12656 17650 12708
rect 13538 12628 13544 12640
rect 12084 12600 13544 12628
rect 9953 12591 10011 12597
rect 13538 12588 13544 12600
rect 13596 12588 13602 12640
rect 13630 12588 13636 12640
rect 13688 12628 13694 12640
rect 16301 12631 16359 12637
rect 16301 12628 16313 12631
rect 13688 12600 16313 12628
rect 13688 12588 13694 12600
rect 16301 12597 16313 12600
rect 16347 12597 16359 12631
rect 16850 12628 16856 12640
rect 16811 12600 16856 12628
rect 16301 12591 16359 12597
rect 16850 12588 16856 12600
rect 16908 12588 16914 12640
rect 17310 12628 17316 12640
rect 17271 12600 17316 12628
rect 17310 12588 17316 12600
rect 17368 12588 17374 12640
rect 1104 12538 18860 12560
rect 1104 12486 6912 12538
rect 6964 12486 6976 12538
rect 7028 12486 7040 12538
rect 7092 12486 7104 12538
rect 7156 12486 12843 12538
rect 12895 12486 12907 12538
rect 12959 12486 12971 12538
rect 13023 12486 13035 12538
rect 13087 12486 18860 12538
rect 1104 12464 18860 12486
rect 3326 12424 3332 12436
rect 3287 12396 3332 12424
rect 3326 12384 3332 12396
rect 3384 12384 3390 12436
rect 6089 12427 6147 12433
rect 6089 12393 6101 12427
rect 6135 12424 6147 12427
rect 7561 12427 7619 12433
rect 7561 12424 7573 12427
rect 6135 12396 7573 12424
rect 6135 12393 6147 12396
rect 6089 12387 6147 12393
rect 7561 12393 7573 12396
rect 7607 12393 7619 12427
rect 8110 12424 8116 12436
rect 8071 12396 8116 12424
rect 7561 12387 7619 12393
rect 8110 12384 8116 12396
rect 8168 12384 8174 12436
rect 9214 12384 9220 12436
rect 9272 12424 9278 12436
rect 10318 12424 10324 12436
rect 9272 12396 10324 12424
rect 9272 12384 9278 12396
rect 10318 12384 10324 12396
rect 10376 12384 10382 12436
rect 10778 12384 10784 12436
rect 10836 12424 10842 12436
rect 11701 12427 11759 12433
rect 11701 12424 11713 12427
rect 10836 12396 11713 12424
rect 10836 12384 10842 12396
rect 11701 12393 11713 12396
rect 11747 12393 11759 12427
rect 11701 12387 11759 12393
rect 12158 12384 12164 12436
rect 12216 12424 12222 12436
rect 13814 12424 13820 12436
rect 12216 12396 13820 12424
rect 12216 12384 12222 12396
rect 13814 12384 13820 12396
rect 13872 12384 13878 12436
rect 14645 12427 14703 12433
rect 14645 12393 14657 12427
rect 14691 12393 14703 12427
rect 14645 12387 14703 12393
rect 4332 12359 4390 12365
rect 4332 12325 4344 12359
rect 4378 12356 4390 12359
rect 6178 12356 6184 12368
rect 4378 12328 6184 12356
rect 4378 12325 4390 12328
rect 4332 12319 4390 12325
rect 6178 12316 6184 12328
rect 6236 12316 6242 12368
rect 7834 12316 7840 12368
rect 7892 12356 7898 12368
rect 7892 12328 10364 12356
rect 7892 12316 7898 12328
rect 2222 12288 2228 12300
rect 2183 12260 2228 12288
rect 2222 12248 2228 12260
rect 2280 12248 2286 12300
rect 4154 12288 4160 12300
rect 3620 12260 4160 12288
rect 2314 12220 2320 12232
rect 2275 12192 2320 12220
rect 2314 12180 2320 12192
rect 2372 12180 2378 12232
rect 2501 12223 2559 12229
rect 2501 12189 2513 12223
rect 2547 12220 2559 12223
rect 2590 12220 2596 12232
rect 2547 12192 2596 12220
rect 2547 12189 2559 12192
rect 2501 12183 2559 12189
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 3620 12229 3648 12260
rect 4154 12248 4160 12260
rect 4212 12248 4218 12300
rect 6457 12291 6515 12297
rect 6457 12257 6469 12291
rect 6503 12288 6515 12291
rect 6822 12288 6828 12300
rect 6503 12260 6828 12288
rect 6503 12257 6515 12260
rect 6457 12251 6515 12257
rect 6822 12248 6828 12260
rect 6880 12248 6886 12300
rect 6914 12248 6920 12300
rect 6972 12288 6978 12300
rect 7469 12291 7527 12297
rect 7469 12288 7481 12291
rect 6972 12260 7481 12288
rect 6972 12248 6978 12260
rect 7469 12257 7481 12260
rect 7515 12257 7527 12291
rect 7469 12251 7527 12257
rect 8481 12291 8539 12297
rect 8481 12257 8493 12291
rect 8527 12288 8539 12291
rect 10226 12288 10232 12300
rect 8527 12260 10232 12288
rect 8527 12257 8539 12260
rect 8481 12251 8539 12257
rect 10226 12248 10232 12260
rect 10284 12248 10290 12300
rect 10336 12288 10364 12328
rect 10410 12316 10416 12368
rect 10468 12356 10474 12368
rect 10566 12359 10624 12365
rect 10566 12356 10578 12359
rect 10468 12328 10578 12356
rect 10468 12316 10474 12328
rect 10566 12325 10578 12328
rect 10612 12325 10624 12359
rect 10566 12319 10624 12325
rect 12621 12359 12679 12365
rect 12621 12325 12633 12359
rect 12667 12356 12679 12359
rect 13354 12356 13360 12368
rect 12667 12328 13360 12356
rect 12667 12325 12679 12328
rect 12621 12319 12679 12325
rect 13354 12316 13360 12328
rect 13412 12316 13418 12368
rect 13532 12359 13590 12365
rect 13532 12325 13544 12359
rect 13578 12356 13590 12359
rect 13630 12356 13636 12368
rect 13578 12328 13636 12356
rect 13578 12325 13590 12328
rect 13532 12319 13590 12325
rect 13630 12316 13636 12328
rect 13688 12316 13694 12368
rect 13722 12316 13728 12368
rect 13780 12356 13786 12368
rect 14660 12356 14688 12387
rect 14734 12384 14740 12436
rect 14792 12424 14798 12436
rect 15289 12427 15347 12433
rect 15289 12424 15301 12427
rect 14792 12396 15301 12424
rect 14792 12384 14798 12396
rect 15289 12393 15301 12396
rect 15335 12393 15347 12427
rect 15289 12387 15347 12393
rect 15562 12384 15568 12436
rect 15620 12424 15626 12436
rect 18046 12424 18052 12436
rect 15620 12396 18052 12424
rect 15620 12384 15626 12396
rect 18046 12384 18052 12396
rect 18104 12384 18110 12436
rect 18141 12427 18199 12433
rect 18141 12393 18153 12427
rect 18187 12393 18199 12427
rect 18141 12387 18199 12393
rect 13780 12328 14688 12356
rect 13780 12316 13786 12328
rect 16942 12316 16948 12368
rect 17000 12356 17006 12368
rect 18156 12356 18184 12387
rect 17000 12328 18184 12356
rect 17000 12316 17006 12328
rect 11606 12288 11612 12300
rect 10336 12260 11612 12288
rect 11606 12248 11612 12260
rect 11664 12248 11670 12300
rect 12713 12291 12771 12297
rect 12713 12257 12725 12291
rect 12759 12288 12771 12291
rect 12759 12260 12848 12288
rect 12759 12257 12771 12260
rect 12713 12251 12771 12257
rect 12820 12232 12848 12260
rect 15562 12248 15568 12300
rect 15620 12248 15626 12300
rect 16114 12288 16120 12300
rect 16075 12260 16120 12288
rect 16114 12248 16120 12260
rect 16172 12248 16178 12300
rect 16758 12288 16764 12300
rect 16719 12260 16764 12288
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 17034 12297 17040 12300
rect 17028 12288 17040 12297
rect 16995 12260 17040 12288
rect 17028 12251 17040 12260
rect 17034 12248 17040 12251
rect 17092 12248 17098 12300
rect 3421 12223 3479 12229
rect 3421 12189 3433 12223
rect 3467 12189 3479 12223
rect 3421 12183 3479 12189
rect 3605 12223 3663 12229
rect 3605 12189 3617 12223
rect 3651 12189 3663 12223
rect 3605 12183 3663 12189
rect 2958 12152 2964 12164
rect 2919 12124 2964 12152
rect 2958 12112 2964 12124
rect 3016 12112 3022 12164
rect 1854 12084 1860 12096
rect 1815 12056 1860 12084
rect 1854 12044 1860 12056
rect 1912 12044 1918 12096
rect 3436 12084 3464 12183
rect 3694 12180 3700 12232
rect 3752 12220 3758 12232
rect 4065 12223 4123 12229
rect 4065 12220 4077 12223
rect 3752 12192 4077 12220
rect 3752 12180 3758 12192
rect 4065 12189 4077 12192
rect 4111 12189 4123 12223
rect 6546 12220 6552 12232
rect 6507 12192 6552 12220
rect 4065 12183 4123 12189
rect 6546 12180 6552 12192
rect 6604 12180 6610 12232
rect 6733 12223 6791 12229
rect 6733 12220 6745 12223
rect 6656 12192 6745 12220
rect 6656 12164 6684 12192
rect 6733 12189 6745 12192
rect 6779 12189 6791 12223
rect 6733 12183 6791 12189
rect 7006 12180 7012 12232
rect 7064 12220 7070 12232
rect 7653 12223 7711 12229
rect 7653 12220 7665 12223
rect 7064 12192 7665 12220
rect 7064 12180 7070 12192
rect 7653 12189 7665 12192
rect 7699 12189 7711 12223
rect 8570 12220 8576 12232
rect 8531 12192 8576 12220
rect 7653 12183 7711 12189
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 8757 12223 8815 12229
rect 8757 12189 8769 12223
rect 8803 12220 8815 12223
rect 8938 12220 8944 12232
rect 8803 12192 8944 12220
rect 8803 12189 8815 12192
rect 8757 12183 8815 12189
rect 8938 12180 8944 12192
rect 8996 12180 9002 12232
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12189 10379 12223
rect 10321 12183 10379 12189
rect 5276 12124 5580 12152
rect 5276 12084 5304 12124
rect 5442 12084 5448 12096
rect 3436 12056 5304 12084
rect 5403 12056 5448 12084
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 5552 12084 5580 12124
rect 6638 12112 6644 12164
rect 6696 12112 6702 12164
rect 8478 12112 8484 12164
rect 8536 12152 8542 12164
rect 8846 12152 8852 12164
rect 8536 12124 8852 12152
rect 8536 12112 8542 12124
rect 8846 12112 8852 12124
rect 8904 12112 8910 12164
rect 7101 12087 7159 12093
rect 7101 12084 7113 12087
rect 5552 12056 7113 12084
rect 7101 12053 7113 12056
rect 7147 12053 7159 12087
rect 7101 12047 7159 12053
rect 7190 12044 7196 12096
rect 7248 12084 7254 12096
rect 9306 12084 9312 12096
rect 7248 12056 9312 12084
rect 7248 12044 7254 12056
rect 9306 12044 9312 12056
rect 9364 12044 9370 12096
rect 10336 12084 10364 12183
rect 12802 12180 12808 12232
rect 12860 12180 12866 12232
rect 12897 12223 12955 12229
rect 12897 12189 12909 12223
rect 12943 12220 12955 12223
rect 13170 12220 13176 12232
rect 12943 12192 13176 12220
rect 12943 12189 12955 12192
rect 12897 12183 12955 12189
rect 13170 12180 13176 12192
rect 13228 12180 13234 12232
rect 13265 12223 13323 12229
rect 13265 12189 13277 12223
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 12526 12112 12532 12164
rect 12584 12152 12590 12164
rect 13280 12152 13308 12183
rect 14550 12180 14556 12232
rect 14608 12220 14614 12232
rect 15010 12220 15016 12232
rect 14608 12192 15016 12220
rect 14608 12180 14614 12192
rect 15010 12180 15016 12192
rect 15068 12180 15074 12232
rect 12584 12124 13308 12152
rect 12584 12112 12590 12124
rect 14274 12112 14280 12164
rect 14332 12152 14338 12164
rect 15102 12152 15108 12164
rect 14332 12124 15108 12152
rect 14332 12112 14338 12124
rect 15102 12112 15108 12124
rect 15160 12112 15166 12164
rect 10502 12084 10508 12096
rect 10336 12056 10508 12084
rect 10502 12044 10508 12056
rect 10560 12044 10566 12096
rect 12066 12044 12072 12096
rect 12124 12084 12130 12096
rect 12253 12087 12311 12093
rect 12253 12084 12265 12087
rect 12124 12056 12265 12084
rect 12124 12044 12130 12056
rect 12253 12053 12265 12056
rect 12299 12053 12311 12087
rect 12253 12047 12311 12053
rect 12710 12044 12716 12096
rect 12768 12084 12774 12096
rect 13630 12084 13636 12096
rect 12768 12056 13636 12084
rect 12768 12044 12774 12056
rect 13630 12044 13636 12056
rect 13688 12044 13694 12096
rect 13998 12044 14004 12096
rect 14056 12084 14062 12096
rect 15580 12084 15608 12248
rect 16206 12220 16212 12232
rect 16167 12192 16212 12220
rect 16206 12180 16212 12192
rect 16264 12180 16270 12232
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12220 16451 12223
rect 16574 12220 16580 12232
rect 16439 12192 16580 12220
rect 16439 12189 16451 12192
rect 16393 12183 16451 12189
rect 16574 12180 16580 12192
rect 16632 12180 16638 12232
rect 14056 12056 15608 12084
rect 14056 12044 14062 12056
rect 15654 12044 15660 12096
rect 15712 12084 15718 12096
rect 15749 12087 15807 12093
rect 15749 12084 15761 12087
rect 15712 12056 15761 12084
rect 15712 12044 15718 12056
rect 15749 12053 15761 12056
rect 15795 12053 15807 12087
rect 15749 12047 15807 12053
rect 1104 11994 18860 12016
rect 1104 11942 3947 11994
rect 3999 11942 4011 11994
rect 4063 11942 4075 11994
rect 4127 11942 4139 11994
rect 4191 11942 9878 11994
rect 9930 11942 9942 11994
rect 9994 11942 10006 11994
rect 10058 11942 10070 11994
rect 10122 11942 15808 11994
rect 15860 11942 15872 11994
rect 15924 11942 15936 11994
rect 15988 11942 16000 11994
rect 16052 11942 18860 11994
rect 1104 11920 18860 11942
rect 2222 11880 2228 11892
rect 2183 11852 2228 11880
rect 2222 11840 2228 11852
rect 2280 11840 2286 11892
rect 6822 11880 6828 11892
rect 6783 11852 6828 11880
rect 6822 11840 6828 11852
rect 6880 11840 6886 11892
rect 11333 11883 11391 11889
rect 7300 11852 11284 11880
rect 5721 11815 5779 11821
rect 5721 11781 5733 11815
rect 5767 11812 5779 11815
rect 6914 11812 6920 11824
rect 5767 11784 6920 11812
rect 5767 11781 5779 11784
rect 5721 11775 5779 11781
rect 6914 11772 6920 11784
rect 6972 11772 6978 11824
rect 2406 11704 2412 11756
rect 2464 11744 2470 11756
rect 2777 11747 2835 11753
rect 2777 11744 2789 11747
rect 2464 11716 2789 11744
rect 2464 11704 2470 11716
rect 2777 11713 2789 11716
rect 2823 11713 2835 11747
rect 2777 11707 2835 11713
rect 6178 11704 6184 11756
rect 6236 11744 6242 11756
rect 6273 11747 6331 11753
rect 6273 11744 6285 11747
rect 6236 11716 6285 11744
rect 6236 11704 6242 11716
rect 6273 11713 6285 11716
rect 6319 11713 6331 11747
rect 6273 11707 6331 11713
rect 6638 11704 6644 11756
rect 6696 11744 6702 11756
rect 7300 11744 7328 11852
rect 9309 11815 9367 11821
rect 9309 11781 9321 11815
rect 9355 11812 9367 11815
rect 9766 11812 9772 11824
rect 9355 11784 9772 11812
rect 9355 11781 9367 11784
rect 9309 11775 9367 11781
rect 9766 11772 9772 11784
rect 9824 11772 9830 11824
rect 11256 11812 11284 11852
rect 11333 11849 11345 11883
rect 11379 11880 11391 11883
rect 12250 11880 12256 11892
rect 11379 11852 12256 11880
rect 11379 11849 11391 11852
rect 11333 11843 11391 11849
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 14093 11883 14151 11889
rect 14093 11880 14105 11883
rect 13412 11852 14105 11880
rect 13412 11840 13418 11852
rect 14093 11849 14105 11852
rect 14139 11849 14151 11883
rect 14093 11843 14151 11849
rect 14734 11840 14740 11892
rect 14792 11880 14798 11892
rect 15286 11880 15292 11892
rect 14792 11852 15292 11880
rect 14792 11840 14798 11852
rect 15286 11840 15292 11852
rect 15344 11840 15350 11892
rect 16114 11840 16120 11892
rect 16172 11880 16178 11892
rect 16209 11883 16267 11889
rect 16209 11880 16221 11883
rect 16172 11852 16221 11880
rect 16172 11840 16178 11852
rect 16209 11849 16221 11852
rect 16255 11849 16267 11883
rect 16209 11843 16267 11849
rect 11698 11812 11704 11824
rect 11256 11784 11704 11812
rect 11698 11772 11704 11784
rect 11756 11772 11762 11824
rect 15562 11772 15568 11824
rect 15620 11812 15626 11824
rect 18230 11812 18236 11824
rect 15620 11784 18236 11812
rect 15620 11772 15626 11784
rect 18230 11772 18236 11784
rect 18288 11772 18294 11824
rect 7466 11744 7472 11756
rect 6696 11716 7328 11744
rect 7427 11716 7472 11744
rect 6696 11704 6702 11716
rect 1670 11676 1676 11688
rect 1631 11648 1676 11676
rect 1670 11636 1676 11648
rect 1728 11636 1734 11688
rect 2498 11636 2504 11688
rect 2556 11676 2562 11688
rect 2593 11679 2651 11685
rect 2593 11676 2605 11679
rect 2556 11648 2605 11676
rect 2556 11636 2562 11648
rect 2593 11645 2605 11648
rect 2639 11645 2651 11679
rect 2593 11639 2651 11645
rect 3237 11679 3295 11685
rect 3237 11645 3249 11679
rect 3283 11645 3295 11679
rect 3237 11639 3295 11645
rect 2682 11608 2688 11620
rect 2643 11580 2688 11608
rect 2682 11568 2688 11580
rect 2740 11568 2746 11620
rect 3252 11608 3280 11639
rect 3694 11636 3700 11688
rect 3752 11676 3758 11688
rect 3789 11679 3847 11685
rect 3789 11676 3801 11679
rect 3752 11648 3801 11676
rect 3752 11636 3758 11648
rect 3789 11645 3801 11648
rect 3835 11645 3847 11679
rect 3789 11639 3847 11645
rect 3878 11636 3884 11688
rect 3936 11676 3942 11688
rect 5074 11676 5080 11688
rect 3936 11648 5080 11676
rect 3936 11636 3942 11648
rect 5074 11636 5080 11648
rect 5132 11636 5138 11688
rect 7098 11676 7104 11688
rect 6656 11648 7104 11676
rect 4056 11611 4114 11617
rect 3252 11580 4016 11608
rect 1486 11500 1492 11552
rect 1544 11540 1550 11552
rect 1857 11543 1915 11549
rect 1857 11540 1869 11543
rect 1544 11512 1869 11540
rect 1544 11500 1550 11512
rect 1857 11509 1869 11512
rect 1903 11509 1915 11543
rect 1857 11503 1915 11509
rect 2958 11500 2964 11552
rect 3016 11540 3022 11552
rect 3421 11543 3479 11549
rect 3421 11540 3433 11543
rect 3016 11512 3433 11540
rect 3016 11500 3022 11512
rect 3421 11509 3433 11512
rect 3467 11509 3479 11543
rect 3988 11540 4016 11580
rect 4056 11577 4068 11611
rect 4102 11608 4114 11611
rect 4246 11608 4252 11620
rect 4102 11580 4252 11608
rect 4102 11577 4114 11580
rect 4056 11571 4114 11577
rect 4246 11568 4252 11580
rect 4304 11568 4310 11620
rect 6656 11608 6684 11648
rect 7098 11636 7104 11648
rect 7156 11636 7162 11688
rect 7208 11685 7236 11716
rect 7466 11704 7472 11716
rect 7524 11704 7530 11756
rect 8938 11704 8944 11756
rect 8996 11744 9002 11756
rect 10137 11747 10195 11753
rect 10137 11744 10149 11747
rect 8996 11716 10149 11744
rect 8996 11704 9002 11716
rect 10137 11713 10149 11716
rect 10183 11713 10195 11747
rect 10137 11707 10195 11713
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11744 11851 11747
rect 11882 11744 11888 11756
rect 11839 11716 11888 11744
rect 11839 11713 11851 11716
rect 11793 11707 11851 11713
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 11977 11747 12035 11753
rect 11977 11713 11989 11747
rect 12023 11744 12035 11747
rect 12158 11744 12164 11756
rect 12023 11716 12164 11744
rect 12023 11713 12035 11716
rect 11977 11707 12035 11713
rect 12158 11704 12164 11716
rect 12216 11704 12222 11756
rect 14090 11744 14096 11756
rect 13464 11716 14096 11744
rect 7193 11679 7251 11685
rect 7193 11645 7205 11679
rect 7239 11645 7251 11679
rect 7193 11639 7251 11645
rect 7285 11679 7343 11685
rect 7285 11645 7297 11679
rect 7331 11676 7343 11679
rect 7650 11676 7656 11688
rect 7331 11648 7656 11676
rect 7331 11645 7343 11648
rect 7285 11639 7343 11645
rect 7650 11636 7656 11648
rect 7708 11636 7714 11688
rect 7929 11679 7987 11685
rect 7929 11645 7941 11679
rect 7975 11676 7987 11679
rect 8018 11676 8024 11688
rect 7975 11648 8024 11676
rect 7975 11645 7987 11648
rect 7929 11639 7987 11645
rect 8018 11636 8024 11648
rect 8076 11636 8082 11688
rect 8202 11685 8208 11688
rect 8196 11639 8208 11685
rect 8260 11676 8266 11688
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 8260 11648 8296 11676
rect 9232 11648 11713 11676
rect 8202 11636 8208 11639
rect 8260 11636 8266 11648
rect 5000 11580 6684 11608
rect 5000 11540 5028 11580
rect 6822 11568 6828 11620
rect 6880 11608 6886 11620
rect 9232 11608 9260 11648
rect 11701 11645 11713 11648
rect 11747 11645 11759 11679
rect 11701 11639 11759 11645
rect 12342 11636 12348 11688
rect 12400 11676 12406 11688
rect 12437 11679 12495 11685
rect 12437 11676 12449 11679
rect 12400 11648 12449 11676
rect 12400 11636 12406 11648
rect 12437 11645 12449 11648
rect 12483 11645 12495 11679
rect 12437 11639 12495 11645
rect 12704 11679 12762 11685
rect 12704 11645 12716 11679
rect 12750 11676 12762 11679
rect 13464 11676 13492 11716
rect 14090 11704 14096 11716
rect 14148 11744 14154 11756
rect 14645 11747 14703 11753
rect 14645 11744 14657 11747
rect 14148 11716 14657 11744
rect 14148 11704 14154 11716
rect 14645 11713 14657 11716
rect 14691 11713 14703 11747
rect 15654 11744 15660 11756
rect 15615 11716 15660 11744
rect 14645 11707 14703 11713
rect 15654 11704 15660 11716
rect 15712 11704 15718 11756
rect 15841 11747 15899 11753
rect 15841 11713 15853 11747
rect 15887 11744 15899 11747
rect 16114 11744 16120 11756
rect 15887 11716 16120 11744
rect 15887 11713 15899 11716
rect 15841 11707 15899 11713
rect 16114 11704 16120 11716
rect 16172 11704 16178 11756
rect 16758 11744 16764 11756
rect 16719 11716 16764 11744
rect 16758 11704 16764 11716
rect 16816 11704 16822 11756
rect 16298 11676 16304 11688
rect 12750 11648 13492 11676
rect 14016 11648 16304 11676
rect 12750 11645 12762 11648
rect 12704 11639 12762 11645
rect 6880 11580 9260 11608
rect 6880 11568 6886 11580
rect 9490 11568 9496 11620
rect 9548 11608 9554 11620
rect 10045 11611 10103 11617
rect 10045 11608 10057 11611
rect 9548 11580 10057 11608
rect 9548 11568 9554 11580
rect 10045 11577 10057 11580
rect 10091 11577 10103 11611
rect 10045 11571 10103 11577
rect 11974 11568 11980 11620
rect 12032 11608 12038 11620
rect 12719 11608 12747 11639
rect 14016 11608 14044 11648
rect 16298 11636 16304 11648
rect 16356 11636 16362 11688
rect 16577 11679 16635 11685
rect 16577 11645 16589 11679
rect 16623 11676 16635 11679
rect 17218 11676 17224 11688
rect 16623 11648 17224 11676
rect 16623 11645 16635 11648
rect 16577 11639 16635 11645
rect 17218 11636 17224 11648
rect 17276 11636 17282 11688
rect 14458 11608 14464 11620
rect 12032 11580 12747 11608
rect 13096 11580 14044 11608
rect 14419 11580 14464 11608
rect 12032 11568 12038 11580
rect 5166 11540 5172 11552
rect 3988 11512 5028 11540
rect 5127 11512 5172 11540
rect 3421 11503 3479 11509
rect 5166 11500 5172 11512
rect 5224 11500 5230 11552
rect 5994 11500 6000 11552
rect 6052 11540 6058 11552
rect 6089 11543 6147 11549
rect 6089 11540 6101 11543
rect 6052 11512 6101 11540
rect 6052 11500 6058 11512
rect 6089 11509 6101 11512
rect 6135 11509 6147 11543
rect 6089 11503 6147 11509
rect 6181 11543 6239 11549
rect 6181 11509 6193 11543
rect 6227 11540 6239 11543
rect 6730 11540 6736 11552
rect 6227 11512 6736 11540
rect 6227 11509 6239 11512
rect 6181 11503 6239 11509
rect 6730 11500 6736 11512
rect 6788 11500 6794 11552
rect 8662 11500 8668 11552
rect 8720 11540 8726 11552
rect 9585 11543 9643 11549
rect 9585 11540 9597 11543
rect 8720 11512 9597 11540
rect 8720 11500 8726 11512
rect 9585 11509 9597 11512
rect 9631 11509 9643 11543
rect 9585 11503 9643 11509
rect 9674 11500 9680 11552
rect 9732 11540 9738 11552
rect 9953 11543 10011 11549
rect 9953 11540 9965 11543
rect 9732 11512 9965 11540
rect 9732 11500 9738 11512
rect 9953 11509 9965 11512
rect 9999 11509 10011 11543
rect 9953 11503 10011 11509
rect 10594 11500 10600 11552
rect 10652 11540 10658 11552
rect 13096 11540 13124 11580
rect 14458 11568 14464 11580
rect 14516 11568 14522 11620
rect 15565 11611 15623 11617
rect 15565 11577 15577 11611
rect 15611 11608 15623 11611
rect 16850 11608 16856 11620
rect 15611 11580 16856 11608
rect 15611 11577 15623 11580
rect 15565 11571 15623 11577
rect 16850 11568 16856 11580
rect 16908 11568 16914 11620
rect 10652 11512 13124 11540
rect 10652 11500 10658 11512
rect 13170 11500 13176 11552
rect 13228 11540 13234 11552
rect 13722 11540 13728 11552
rect 13228 11512 13728 11540
rect 13228 11500 13234 11512
rect 13722 11500 13728 11512
rect 13780 11540 13786 11552
rect 13817 11543 13875 11549
rect 13817 11540 13829 11543
rect 13780 11512 13829 11540
rect 13780 11500 13786 11512
rect 13817 11509 13829 11512
rect 13863 11509 13875 11543
rect 13817 11503 13875 11509
rect 14366 11500 14372 11552
rect 14424 11540 14430 11552
rect 14553 11543 14611 11549
rect 14553 11540 14565 11543
rect 14424 11512 14565 11540
rect 14424 11500 14430 11512
rect 14553 11509 14565 11512
rect 14599 11509 14611 11543
rect 15194 11540 15200 11552
rect 15155 11512 15200 11540
rect 14553 11503 14611 11509
rect 15194 11500 15200 11512
rect 15252 11500 15258 11552
rect 16669 11543 16727 11549
rect 16669 11509 16681 11543
rect 16715 11540 16727 11543
rect 16942 11540 16948 11552
rect 16715 11512 16948 11540
rect 16715 11509 16727 11512
rect 16669 11503 16727 11509
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 1104 11450 18860 11472
rect 1104 11398 6912 11450
rect 6964 11398 6976 11450
rect 7028 11398 7040 11450
rect 7092 11398 7104 11450
rect 7156 11398 12843 11450
rect 12895 11398 12907 11450
rect 12959 11398 12971 11450
rect 13023 11398 13035 11450
rect 13087 11398 18860 11450
rect 1104 11376 18860 11398
rect 2130 11296 2136 11348
rect 2188 11336 2194 11348
rect 6362 11336 6368 11348
rect 2188 11308 6368 11336
rect 2188 11296 2194 11308
rect 6362 11296 6368 11308
rect 6420 11296 6426 11348
rect 6546 11336 6552 11348
rect 6507 11308 6552 11336
rect 6546 11296 6552 11308
rect 6604 11296 6610 11348
rect 6730 11296 6736 11348
rect 6788 11336 6794 11348
rect 7561 11339 7619 11345
rect 7561 11336 7573 11339
rect 6788 11308 7573 11336
rect 6788 11296 6794 11308
rect 7561 11305 7573 11308
rect 7607 11305 7619 11339
rect 7561 11299 7619 11305
rect 8021 11339 8079 11345
rect 8021 11305 8033 11339
rect 8067 11336 8079 11339
rect 8110 11336 8116 11348
rect 8067 11308 8116 11336
rect 8067 11305 8079 11308
rect 8021 11299 8079 11305
rect 8110 11296 8116 11308
rect 8168 11296 8174 11348
rect 8573 11339 8631 11345
rect 8573 11305 8585 11339
rect 8619 11336 8631 11339
rect 9490 11336 9496 11348
rect 8619 11308 9496 11336
rect 8619 11305 8631 11308
rect 8573 11299 8631 11305
rect 9490 11296 9496 11308
rect 9548 11296 9554 11348
rect 9674 11336 9680 11348
rect 9635 11308 9680 11336
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 9858 11296 9864 11348
rect 9916 11336 9922 11348
rect 13630 11336 13636 11348
rect 9916 11308 13636 11336
rect 9916 11296 9922 11308
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 13725 11339 13783 11345
rect 13725 11305 13737 11339
rect 13771 11336 13783 11339
rect 13906 11336 13912 11348
rect 13771 11308 13912 11336
rect 13771 11305 13783 11308
rect 13725 11299 13783 11305
rect 13906 11296 13912 11308
rect 13964 11296 13970 11348
rect 14001 11339 14059 11345
rect 14001 11305 14013 11339
rect 14047 11336 14059 11339
rect 14366 11336 14372 11348
rect 14047 11308 14372 11336
rect 14047 11305 14059 11308
rect 14001 11299 14059 11305
rect 14366 11296 14372 11308
rect 14424 11296 14430 11348
rect 16206 11336 16212 11348
rect 16167 11308 16212 11336
rect 16206 11296 16212 11308
rect 16264 11296 16270 11348
rect 17310 11296 17316 11348
rect 17368 11336 17374 11348
rect 17405 11339 17463 11345
rect 17405 11336 17417 11339
rect 17368 11308 17417 11336
rect 17368 11296 17374 11308
rect 17405 11305 17417 11308
rect 17451 11305 17463 11339
rect 17405 11299 17463 11305
rect 17494 11296 17500 11348
rect 17552 11336 17558 11348
rect 17865 11339 17923 11345
rect 17865 11336 17877 11339
rect 17552 11308 17877 11336
rect 17552 11296 17558 11308
rect 17865 11305 17877 11308
rect 17911 11336 17923 11339
rect 18782 11336 18788 11348
rect 17911 11308 18788 11336
rect 17911 11305 17923 11308
rect 17865 11299 17923 11305
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 2682 11268 2688 11280
rect 1688 11240 2688 11268
rect 1688 11209 1716 11240
rect 2682 11228 2688 11240
rect 2740 11228 2746 11280
rect 2498 11209 2504 11212
rect 1673 11203 1731 11209
rect 1673 11169 1685 11203
rect 1719 11169 1731 11203
rect 2492 11200 2504 11209
rect 2459 11172 2504 11200
rect 1673 11163 1731 11169
rect 2492 11163 2504 11172
rect 2498 11160 2504 11163
rect 2556 11160 2562 11212
rect 4332 11203 4390 11209
rect 4332 11169 4344 11203
rect 4378 11200 4390 11203
rect 5166 11200 5172 11212
rect 4378 11172 5172 11200
rect 4378 11169 4390 11172
rect 4332 11163 4390 11169
rect 5166 11160 5172 11172
rect 5224 11160 5230 11212
rect 6380 11200 6408 11296
rect 7834 11228 7840 11280
rect 7892 11268 7898 11280
rect 10962 11268 10968 11280
rect 7892 11240 10968 11268
rect 7892 11228 7898 11240
rect 10962 11228 10968 11240
rect 11020 11228 11026 11280
rect 11882 11228 11888 11280
rect 11940 11268 11946 11280
rect 16577 11271 16635 11277
rect 16577 11268 16589 11271
rect 11940 11240 16589 11268
rect 11940 11228 11946 11240
rect 16577 11237 16589 11240
rect 16623 11237 16635 11271
rect 17954 11268 17960 11280
rect 16577 11231 16635 11237
rect 16776 11240 17960 11268
rect 6546 11200 6552 11212
rect 6380 11172 6552 11200
rect 6546 11160 6552 11172
rect 6604 11160 6610 11212
rect 6914 11200 6920 11212
rect 6875 11172 6920 11200
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 7009 11203 7067 11209
rect 7009 11169 7021 11203
rect 7055 11200 7067 11203
rect 7742 11200 7748 11212
rect 7055 11172 7748 11200
rect 7055 11169 7067 11172
rect 7009 11163 7067 11169
rect 7742 11160 7748 11172
rect 7800 11160 7806 11212
rect 7926 11200 7932 11212
rect 7887 11172 7932 11200
rect 7926 11160 7932 11172
rect 7984 11160 7990 11212
rect 8386 11160 8392 11212
rect 8444 11200 8450 11212
rect 8941 11203 8999 11209
rect 8941 11200 8953 11203
rect 8444 11172 8953 11200
rect 8444 11160 8450 11172
rect 8941 11169 8953 11172
rect 8987 11169 8999 11203
rect 8941 11163 8999 11169
rect 9033 11203 9091 11209
rect 9033 11169 9045 11203
rect 9079 11200 9091 11203
rect 9214 11200 9220 11212
rect 9079 11172 9220 11200
rect 9079 11169 9091 11172
rect 9033 11163 9091 11169
rect 1302 11092 1308 11144
rect 1360 11132 1366 11144
rect 2225 11135 2283 11141
rect 2225 11132 2237 11135
rect 1360 11104 2237 11132
rect 1360 11092 1366 11104
rect 2225 11101 2237 11104
rect 2271 11101 2283 11135
rect 2225 11095 2283 11101
rect 3694 11092 3700 11144
rect 3752 11132 3758 11144
rect 4065 11135 4123 11141
rect 4065 11132 4077 11135
rect 3752 11104 4077 11132
rect 3752 11092 3758 11104
rect 4065 11101 4077 11104
rect 4111 11101 4123 11135
rect 4065 11095 4123 11101
rect 7193 11135 7251 11141
rect 7193 11101 7205 11135
rect 7239 11101 7251 11135
rect 7193 11095 7251 11101
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11101 8171 11135
rect 9048 11132 9076 11163
rect 9214 11160 9220 11172
rect 9272 11160 9278 11212
rect 9674 11160 9680 11212
rect 9732 11200 9738 11212
rect 10045 11203 10103 11209
rect 10045 11200 10057 11203
rect 9732 11172 10057 11200
rect 9732 11160 9738 11172
rect 10045 11169 10057 11172
rect 10091 11169 10103 11203
rect 10045 11163 10103 11169
rect 11241 11203 11299 11209
rect 11241 11169 11253 11203
rect 11287 11169 11299 11203
rect 11698 11200 11704 11212
rect 11659 11172 11704 11200
rect 11241 11163 11299 11169
rect 8113 11095 8171 11101
rect 8211 11104 9076 11132
rect 9125 11135 9183 11141
rect 1394 11024 1400 11076
rect 1452 11064 1458 11076
rect 1857 11067 1915 11073
rect 1857 11064 1869 11067
rect 1452 11036 1869 11064
rect 1452 11024 1458 11036
rect 1857 11033 1869 11036
rect 1903 11033 1915 11067
rect 1857 11027 1915 11033
rect 3234 11024 3240 11076
rect 3292 11064 3298 11076
rect 3605 11067 3663 11073
rect 3605 11064 3617 11067
rect 3292 11036 3617 11064
rect 3292 11024 3298 11036
rect 3605 11033 3617 11036
rect 3651 11033 3663 11067
rect 5442 11064 5448 11076
rect 5403 11036 5448 11064
rect 3605 11027 3663 11033
rect 5442 11024 5448 11036
rect 5500 11024 5506 11076
rect 7208 11064 7236 11095
rect 7466 11064 7472 11076
rect 7208 11036 7472 11064
rect 7466 11024 7472 11036
rect 7524 11064 7530 11076
rect 8128 11064 8156 11095
rect 7524 11036 8156 11064
rect 7524 11024 7530 11036
rect 3510 10956 3516 11008
rect 3568 10996 3574 11008
rect 5258 10996 5264 11008
rect 3568 10968 5264 10996
rect 3568 10956 3574 10968
rect 5258 10956 5264 10968
rect 5316 10956 5322 11008
rect 5350 10956 5356 11008
rect 5408 10996 5414 11008
rect 8211 10996 8239 11104
rect 9125 11101 9137 11135
rect 9171 11101 9183 11135
rect 9125 11095 9183 11101
rect 8846 11024 8852 11076
rect 8904 11064 8910 11076
rect 9140 11064 9168 11095
rect 9306 11092 9312 11144
rect 9364 11132 9370 11144
rect 10137 11135 10195 11141
rect 10137 11132 10149 11135
rect 9364 11104 10149 11132
rect 9364 11092 9370 11104
rect 10137 11101 10149 11104
rect 10183 11101 10195 11135
rect 10137 11095 10195 11101
rect 10229 11135 10287 11141
rect 10229 11101 10241 11135
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 10244 11064 10272 11095
rect 10318 11092 10324 11144
rect 10376 11132 10382 11144
rect 10594 11132 10600 11144
rect 10376 11104 10600 11132
rect 10376 11092 10382 11104
rect 10594 11092 10600 11104
rect 10652 11092 10658 11144
rect 11256 11132 11284 11163
rect 11698 11160 11704 11172
rect 11756 11160 11762 11212
rect 12253 11203 12311 11209
rect 12253 11169 12265 11203
rect 12299 11200 12311 11203
rect 12342 11200 12348 11212
rect 12299 11172 12348 11200
rect 12299 11169 12311 11172
rect 12253 11163 12311 11169
rect 12342 11160 12348 11172
rect 12400 11160 12406 11212
rect 12618 11209 12624 11212
rect 12612 11200 12624 11209
rect 12579 11172 12624 11200
rect 12612 11163 12624 11172
rect 12618 11160 12624 11163
rect 12676 11160 12682 11212
rect 14366 11200 14372 11212
rect 14327 11172 14372 11200
rect 14366 11160 14372 11172
rect 14424 11160 14430 11212
rect 15654 11160 15660 11212
rect 15712 11200 15718 11212
rect 16776 11200 16804 11240
rect 17954 11228 17960 11240
rect 18012 11228 18018 11280
rect 15712 11172 16804 11200
rect 15712 11160 15718 11172
rect 17586 11160 17592 11212
rect 17644 11200 17650 11212
rect 17773 11203 17831 11209
rect 17773 11200 17785 11203
rect 17644 11172 17785 11200
rect 17644 11160 17650 11172
rect 17773 11169 17785 11172
rect 17819 11169 17831 11203
rect 17773 11163 17831 11169
rect 11790 11132 11796 11144
rect 11256 11104 11652 11132
rect 11751 11104 11796 11132
rect 8904 11036 10272 11064
rect 11333 11067 11391 11073
rect 8904 11024 8910 11036
rect 11333 11033 11345 11067
rect 11379 11064 11391 11067
rect 11422 11064 11428 11076
rect 11379 11036 11428 11064
rect 11379 11033 11391 11036
rect 11333 11027 11391 11033
rect 11422 11024 11428 11036
rect 11480 11024 11486 11076
rect 11624 11064 11652 11104
rect 11790 11092 11796 11104
rect 11848 11092 11854 11144
rect 11974 11092 11980 11144
rect 12032 11132 12038 11144
rect 12032 11104 12077 11132
rect 12032 11092 12038 11104
rect 13998 11092 14004 11144
rect 14056 11132 14062 11144
rect 14274 11132 14280 11144
rect 14056 11104 14280 11132
rect 14056 11092 14062 11104
rect 14274 11092 14280 11104
rect 14332 11132 14338 11144
rect 14461 11135 14519 11141
rect 14461 11132 14473 11135
rect 14332 11104 14473 11132
rect 14332 11092 14338 11104
rect 14461 11101 14473 11104
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 14553 11135 14611 11141
rect 14553 11101 14565 11135
rect 14599 11101 14611 11135
rect 15286 11132 15292 11144
rect 15247 11104 15292 11132
rect 14553 11095 14611 11101
rect 11624 11036 12388 11064
rect 5408 10968 8239 10996
rect 5408 10956 5414 10968
rect 8386 10956 8392 11008
rect 8444 10996 8450 11008
rect 9582 10996 9588 11008
rect 8444 10968 9588 10996
rect 8444 10956 8450 10968
rect 9582 10956 9588 10968
rect 9640 10956 9646 11008
rect 10502 10956 10508 11008
rect 10560 10996 10566 11008
rect 11057 10999 11115 11005
rect 11057 10996 11069 10999
rect 10560 10968 11069 10996
rect 10560 10956 10566 10968
rect 11057 10965 11069 10968
rect 11103 10996 11115 10999
rect 12253 10999 12311 11005
rect 12253 10996 12265 10999
rect 11103 10968 12265 10996
rect 11103 10965 11115 10968
rect 11057 10959 11115 10965
rect 12253 10965 12265 10968
rect 12299 10965 12311 10999
rect 12360 10996 12388 11036
rect 14090 11024 14096 11076
rect 14148 11064 14154 11076
rect 14568 11064 14596 11095
rect 15286 11092 15292 11104
rect 15344 11092 15350 11144
rect 16666 11132 16672 11144
rect 16627 11104 16672 11132
rect 16666 11092 16672 11104
rect 16724 11092 16730 11144
rect 16758 11092 16764 11144
rect 16816 11132 16822 11144
rect 16853 11135 16911 11141
rect 16853 11132 16865 11135
rect 16816 11104 16865 11132
rect 16816 11092 16822 11104
rect 16853 11101 16865 11104
rect 16899 11132 16911 11135
rect 18049 11135 18107 11141
rect 18049 11132 18061 11135
rect 16899 11104 18061 11132
rect 16899 11101 16911 11104
rect 16853 11095 16911 11101
rect 18049 11101 18061 11104
rect 18095 11132 18107 11135
rect 18322 11132 18328 11144
rect 18095 11104 18328 11132
rect 18095 11101 18107 11104
rect 18049 11095 18107 11101
rect 18322 11092 18328 11104
rect 18380 11092 18386 11144
rect 14148 11036 14596 11064
rect 14148 11024 14154 11036
rect 13446 10996 13452 11008
rect 12360 10968 13452 10996
rect 12253 10959 12311 10965
rect 13446 10956 13452 10968
rect 13504 10956 13510 11008
rect 13538 10956 13544 11008
rect 13596 10996 13602 11008
rect 17586 10996 17592 11008
rect 13596 10968 17592 10996
rect 13596 10956 13602 10968
rect 17586 10956 17592 10968
rect 17644 10996 17650 11008
rect 18046 10996 18052 11008
rect 17644 10968 18052 10996
rect 17644 10956 17650 10968
rect 18046 10956 18052 10968
rect 18104 10956 18110 11008
rect 1104 10906 18860 10928
rect 1104 10854 3947 10906
rect 3999 10854 4011 10906
rect 4063 10854 4075 10906
rect 4127 10854 4139 10906
rect 4191 10854 9878 10906
rect 9930 10854 9942 10906
rect 9994 10854 10006 10906
rect 10058 10854 10070 10906
rect 10122 10854 15808 10906
rect 15860 10854 15872 10906
rect 15924 10854 15936 10906
rect 15988 10854 16000 10906
rect 16052 10854 18860 10906
rect 1104 10832 18860 10854
rect 2225 10795 2283 10801
rect 2225 10761 2237 10795
rect 2271 10792 2283 10795
rect 2314 10792 2320 10804
rect 2271 10764 2320 10792
rect 2271 10761 2283 10764
rect 2225 10755 2283 10761
rect 2314 10752 2320 10764
rect 2372 10752 2378 10804
rect 4798 10752 4804 10804
rect 4856 10792 4862 10804
rect 6822 10792 6828 10804
rect 4856 10764 6828 10792
rect 4856 10752 4862 10764
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 8018 10792 8024 10804
rect 7392 10764 8024 10792
rect 1857 10727 1915 10733
rect 1857 10693 1869 10727
rect 1903 10724 1915 10727
rect 3326 10724 3332 10736
rect 1903 10696 3332 10724
rect 1903 10693 1915 10696
rect 1857 10687 1915 10693
rect 3326 10684 3332 10696
rect 3384 10684 3390 10736
rect 4080 10696 5488 10724
rect 2498 10616 2504 10668
rect 2556 10656 2562 10668
rect 4080 10665 4108 10696
rect 5460 10668 5488 10696
rect 2869 10659 2927 10665
rect 2869 10656 2881 10659
rect 2556 10628 2881 10656
rect 2556 10616 2562 10628
rect 2869 10625 2881 10628
rect 2915 10656 2927 10659
rect 4065 10659 4123 10665
rect 4065 10656 4077 10659
rect 2915 10628 4077 10656
rect 2915 10625 2927 10628
rect 2869 10619 2927 10625
rect 4065 10625 4077 10628
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10656 5135 10659
rect 5166 10656 5172 10668
rect 5123 10628 5172 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 5166 10616 5172 10628
rect 5224 10616 5230 10668
rect 5350 10616 5356 10668
rect 5408 10616 5414 10668
rect 5442 10616 5448 10668
rect 5500 10656 5506 10668
rect 7392 10665 7420 10764
rect 8018 10752 8024 10764
rect 8076 10752 8082 10804
rect 8754 10792 8760 10804
rect 8715 10764 8760 10792
rect 8754 10752 8760 10764
rect 8812 10752 8818 10804
rect 10410 10792 10416 10804
rect 10371 10764 10416 10792
rect 10410 10752 10416 10764
rect 10468 10752 10474 10804
rect 11333 10795 11391 10801
rect 11333 10761 11345 10795
rect 11379 10792 11391 10795
rect 11698 10792 11704 10804
rect 11379 10764 11704 10792
rect 11379 10761 11391 10764
rect 11333 10755 11391 10761
rect 11698 10752 11704 10764
rect 11756 10752 11762 10804
rect 13633 10795 13691 10801
rect 13633 10761 13645 10795
rect 13679 10792 13691 10795
rect 14458 10792 14464 10804
rect 13679 10764 14464 10792
rect 13679 10761 13691 10764
rect 13633 10755 13691 10761
rect 14458 10752 14464 10764
rect 14516 10752 14522 10804
rect 14550 10752 14556 10804
rect 14608 10752 14614 10804
rect 14918 10792 14924 10804
rect 14660 10764 14924 10792
rect 5997 10659 6055 10665
rect 5997 10656 6009 10659
rect 5500 10628 6009 10656
rect 5500 10616 5506 10628
rect 5997 10625 6009 10628
rect 6043 10625 6055 10659
rect 5997 10619 6055 10625
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 7377 10659 7435 10665
rect 7377 10656 7389 10659
rect 6687 10628 7389 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 7377 10625 7389 10628
rect 7423 10625 7435 10659
rect 8772 10656 8800 10752
rect 12710 10684 12716 10736
rect 12768 10724 12774 10736
rect 14274 10724 14280 10736
rect 12768 10696 14280 10724
rect 12768 10684 12774 10696
rect 14274 10684 14280 10696
rect 14332 10724 14338 10736
rect 14568 10724 14596 10752
rect 14332 10696 14596 10724
rect 14332 10684 14338 10696
rect 11977 10659 12035 10665
rect 8772 10628 9168 10656
rect 7377 10619 7435 10625
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10588 1731 10591
rect 2685 10591 2743 10597
rect 2685 10588 2697 10591
rect 1719 10560 2697 10588
rect 1719 10557 1731 10560
rect 1673 10551 1731 10557
rect 2685 10557 2697 10560
rect 2731 10588 2743 10591
rect 5368 10588 5396 10616
rect 2731 10560 5396 10588
rect 2731 10557 2743 10560
rect 2685 10551 2743 10557
rect 5534 10548 5540 10600
rect 5592 10588 5598 10600
rect 7285 10591 7343 10597
rect 7285 10588 7297 10591
rect 5592 10560 7297 10588
rect 5592 10548 5598 10560
rect 7285 10557 7297 10560
rect 7331 10557 7343 10591
rect 8938 10588 8944 10600
rect 7285 10551 7343 10557
rect 7944 10560 8944 10588
rect 2593 10523 2651 10529
rect 2593 10489 2605 10523
rect 2639 10520 2651 10523
rect 2774 10520 2780 10532
rect 2639 10492 2780 10520
rect 2639 10489 2651 10492
rect 2593 10483 2651 10489
rect 2774 10480 2780 10492
rect 2832 10520 2838 10532
rect 4062 10520 4068 10532
rect 2832 10492 4068 10520
rect 2832 10480 2838 10492
rect 4062 10480 4068 10492
rect 4120 10480 4126 10532
rect 5905 10523 5963 10529
rect 5905 10520 5917 10523
rect 4448 10492 5917 10520
rect 3418 10452 3424 10464
rect 3379 10424 3424 10452
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 3786 10452 3792 10464
rect 3747 10424 3792 10452
rect 3786 10412 3792 10424
rect 3844 10412 3850 10464
rect 3881 10455 3939 10461
rect 3881 10421 3893 10455
rect 3927 10452 3939 10455
rect 4338 10452 4344 10464
rect 3927 10424 4344 10452
rect 3927 10421 3939 10424
rect 3881 10415 3939 10421
rect 4338 10412 4344 10424
rect 4396 10412 4402 10464
rect 4448 10461 4476 10492
rect 5905 10489 5917 10492
rect 5951 10489 5963 10523
rect 5905 10483 5963 10489
rect 6730 10480 6736 10532
rect 6788 10520 6794 10532
rect 7622 10523 7680 10529
rect 7622 10520 7634 10523
rect 6788 10492 7634 10520
rect 6788 10480 6794 10492
rect 7622 10489 7634 10492
rect 7668 10520 7680 10523
rect 7944 10520 7972 10560
rect 8938 10548 8944 10560
rect 8996 10548 9002 10600
rect 9033 10591 9091 10597
rect 9033 10557 9045 10591
rect 9079 10557 9091 10591
rect 9140 10588 9168 10628
rect 11977 10625 11989 10659
rect 12023 10656 12035 10659
rect 12618 10656 12624 10668
rect 12023 10628 12624 10656
rect 12023 10625 12035 10628
rect 11977 10619 12035 10625
rect 12618 10616 12624 10628
rect 12676 10616 12682 10668
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10656 13139 10659
rect 13170 10656 13176 10668
rect 13127 10628 13176 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 14185 10659 14243 10665
rect 14185 10625 14197 10659
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 9289 10591 9347 10597
rect 9289 10588 9301 10591
rect 9140 10560 9301 10588
rect 9033 10551 9091 10557
rect 9289 10557 9301 10560
rect 9335 10557 9347 10591
rect 9289 10551 9347 10557
rect 7668 10492 7972 10520
rect 7668 10489 7680 10492
rect 7622 10483 7680 10489
rect 8018 10480 8024 10532
rect 8076 10520 8082 10532
rect 9048 10520 9076 10551
rect 9582 10548 9588 10600
rect 9640 10588 9646 10600
rect 12342 10588 12348 10600
rect 9640 10560 12348 10588
rect 9640 10548 9646 10560
rect 12342 10548 12348 10560
rect 12400 10548 12406 10600
rect 12636 10588 12664 10616
rect 14090 10588 14096 10600
rect 12636 10560 14096 10588
rect 14090 10548 14096 10560
rect 14148 10588 14154 10600
rect 14200 10588 14228 10619
rect 14550 10616 14556 10668
rect 14608 10656 14614 10668
rect 14660 10665 14688 10764
rect 14918 10752 14924 10764
rect 14976 10792 14982 10804
rect 16025 10795 16083 10801
rect 14976 10764 15700 10792
rect 14976 10752 14982 10764
rect 14645 10659 14703 10665
rect 14645 10656 14657 10659
rect 14608 10628 14657 10656
rect 14608 10616 14614 10628
rect 14645 10625 14657 10628
rect 14691 10625 14703 10659
rect 14645 10619 14703 10625
rect 14458 10588 14464 10600
rect 14148 10560 14464 10588
rect 14148 10548 14154 10560
rect 14458 10548 14464 10560
rect 14516 10548 14522 10600
rect 15286 10588 15292 10600
rect 14752 10560 15292 10588
rect 13906 10520 13912 10532
rect 8076 10492 9076 10520
rect 9140 10492 13912 10520
rect 8076 10480 8082 10492
rect 4433 10455 4491 10461
rect 4433 10421 4445 10455
rect 4479 10421 4491 10455
rect 4798 10452 4804 10464
rect 4759 10424 4804 10452
rect 4433 10415 4491 10421
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 4893 10455 4951 10461
rect 4893 10421 4905 10455
rect 4939 10452 4951 10455
rect 5258 10452 5264 10464
rect 4939 10424 5264 10452
rect 4939 10421 4951 10424
rect 4893 10415 4951 10421
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 5442 10452 5448 10464
rect 5403 10424 5448 10452
rect 5442 10412 5448 10424
rect 5500 10412 5506 10464
rect 5810 10452 5816 10464
rect 5771 10424 5816 10452
rect 5810 10412 5816 10424
rect 5868 10412 5874 10464
rect 6178 10412 6184 10464
rect 6236 10452 6242 10464
rect 6641 10455 6699 10461
rect 6641 10452 6653 10455
rect 6236 10424 6653 10452
rect 6236 10412 6242 10424
rect 6641 10421 6653 10424
rect 6687 10452 6699 10455
rect 7101 10455 7159 10461
rect 7101 10452 7113 10455
rect 6687 10424 7113 10452
rect 6687 10421 6699 10424
rect 6641 10415 6699 10421
rect 7101 10421 7113 10424
rect 7147 10452 7159 10455
rect 7282 10452 7288 10464
rect 7147 10424 7288 10452
rect 7147 10421 7159 10424
rect 7101 10415 7159 10421
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 7926 10412 7932 10464
rect 7984 10452 7990 10464
rect 9140 10452 9168 10492
rect 13906 10480 13912 10492
rect 13964 10480 13970 10532
rect 14001 10523 14059 10529
rect 14001 10489 14013 10523
rect 14047 10520 14059 10523
rect 14752 10520 14780 10560
rect 15286 10548 15292 10560
rect 15344 10548 15350 10600
rect 15672 10588 15700 10764
rect 16025 10761 16037 10795
rect 16071 10792 16083 10795
rect 16114 10792 16120 10804
rect 16071 10764 16120 10792
rect 16071 10761 16083 10764
rect 16025 10755 16083 10761
rect 16114 10752 16120 10764
rect 16172 10752 16178 10804
rect 17034 10752 17040 10804
rect 17092 10792 17098 10804
rect 17681 10795 17739 10801
rect 17681 10792 17693 10795
rect 17092 10764 17693 10792
rect 17092 10752 17098 10764
rect 17681 10761 17693 10764
rect 17727 10761 17739 10795
rect 17681 10755 17739 10761
rect 16132 10656 16160 10752
rect 16132 10628 16436 10656
rect 15746 10588 15752 10600
rect 15659 10560 15752 10588
rect 15746 10548 15752 10560
rect 15804 10588 15810 10600
rect 16301 10591 16359 10597
rect 16301 10588 16313 10591
rect 15804 10560 16313 10588
rect 15804 10548 15810 10560
rect 16301 10557 16313 10560
rect 16347 10557 16359 10591
rect 16408 10588 16436 10628
rect 16557 10591 16615 10597
rect 16557 10588 16569 10591
rect 16408 10560 16569 10588
rect 16301 10551 16359 10557
rect 16557 10557 16569 10560
rect 16603 10557 16615 10591
rect 16557 10551 16615 10557
rect 14047 10492 14780 10520
rect 14912 10523 14970 10529
rect 14047 10489 14059 10492
rect 14001 10483 14059 10489
rect 14912 10489 14924 10523
rect 14958 10520 14970 10523
rect 17494 10520 17500 10532
rect 14958 10492 17500 10520
rect 14958 10489 14970 10492
rect 14912 10483 14970 10489
rect 16592 10464 16620 10492
rect 17494 10480 17500 10492
rect 17552 10480 17558 10532
rect 7984 10424 9168 10452
rect 7984 10412 7990 10424
rect 9214 10412 9220 10464
rect 9272 10452 9278 10464
rect 10962 10452 10968 10464
rect 9272 10424 10968 10452
rect 9272 10412 9278 10424
rect 10962 10412 10968 10424
rect 11020 10412 11026 10464
rect 11698 10452 11704 10464
rect 11659 10424 11704 10452
rect 11698 10412 11704 10424
rect 11756 10412 11762 10464
rect 11793 10455 11851 10461
rect 11793 10421 11805 10455
rect 11839 10452 11851 10455
rect 12437 10455 12495 10461
rect 12437 10452 12449 10455
rect 11839 10424 12449 10452
rect 11839 10421 11851 10424
rect 11793 10415 11851 10421
rect 12437 10421 12449 10424
rect 12483 10421 12495 10455
rect 12437 10415 12495 10421
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 12805 10455 12863 10461
rect 12805 10452 12817 10455
rect 12768 10424 12817 10452
rect 12768 10412 12774 10424
rect 12805 10421 12817 10424
rect 12851 10421 12863 10455
rect 12805 10415 12863 10421
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10452 12955 10455
rect 13354 10452 13360 10464
rect 12943 10424 13360 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 13354 10412 13360 10424
rect 13412 10412 13418 10464
rect 13814 10412 13820 10464
rect 13872 10452 13878 10464
rect 14093 10455 14151 10461
rect 14093 10452 14105 10455
rect 13872 10424 14105 10452
rect 13872 10412 13878 10424
rect 14093 10421 14105 10424
rect 14139 10452 14151 10455
rect 14734 10452 14740 10464
rect 14139 10424 14740 10452
rect 14139 10421 14151 10424
rect 14093 10415 14151 10421
rect 14734 10412 14740 10424
rect 14792 10412 14798 10464
rect 16574 10412 16580 10464
rect 16632 10412 16638 10464
rect 1104 10362 18860 10384
rect 1104 10310 6912 10362
rect 6964 10310 6976 10362
rect 7028 10310 7040 10362
rect 7092 10310 7104 10362
rect 7156 10310 12843 10362
rect 12895 10310 12907 10362
rect 12959 10310 12971 10362
rect 13023 10310 13035 10362
rect 13087 10310 18860 10362
rect 1104 10288 18860 10310
rect 1302 10208 1308 10260
rect 1360 10248 1366 10260
rect 3605 10251 3663 10257
rect 3605 10248 3617 10251
rect 1360 10220 3617 10248
rect 1360 10208 1366 10220
rect 3605 10217 3617 10220
rect 3651 10248 3663 10251
rect 3694 10248 3700 10260
rect 3651 10220 3700 10248
rect 3651 10217 3663 10220
rect 3605 10211 3663 10217
rect 3694 10208 3700 10220
rect 3752 10208 3758 10260
rect 3786 10208 3792 10260
rect 3844 10248 3850 10260
rect 4433 10251 4491 10257
rect 4433 10248 4445 10251
rect 3844 10220 4445 10248
rect 3844 10208 3850 10220
rect 4433 10217 4445 10220
rect 4479 10217 4491 10251
rect 4433 10211 4491 10217
rect 4801 10251 4859 10257
rect 4801 10217 4813 10251
rect 4847 10248 4859 10251
rect 4982 10248 4988 10260
rect 4847 10220 4988 10248
rect 4847 10217 4859 10220
rect 4801 10211 4859 10217
rect 4982 10208 4988 10220
rect 5040 10208 5046 10260
rect 5534 10248 5540 10260
rect 5092 10220 5540 10248
rect 1664 10183 1722 10189
rect 1664 10149 1676 10183
rect 1710 10180 1722 10183
rect 2590 10180 2596 10192
rect 1710 10152 2596 10180
rect 1710 10149 1722 10152
rect 1664 10143 1722 10149
rect 2590 10140 2596 10152
rect 2648 10180 2654 10192
rect 3234 10180 3240 10192
rect 2648 10152 3240 10180
rect 2648 10140 2654 10152
rect 3234 10140 3240 10152
rect 3292 10140 3298 10192
rect 5092 10180 5120 10220
rect 5534 10208 5540 10220
rect 5592 10208 5598 10260
rect 6086 10208 6092 10260
rect 6144 10248 6150 10260
rect 7837 10251 7895 10257
rect 7837 10248 7849 10251
rect 6144 10220 7849 10248
rect 6144 10208 6150 10220
rect 7837 10217 7849 10220
rect 7883 10217 7895 10251
rect 7837 10211 7895 10217
rect 8481 10251 8539 10257
rect 8481 10217 8493 10251
rect 8527 10248 8539 10251
rect 8570 10248 8576 10260
rect 8527 10220 8576 10248
rect 8527 10217 8539 10220
rect 8481 10211 8539 10217
rect 8570 10208 8576 10220
rect 8628 10208 8634 10260
rect 8849 10251 8907 10257
rect 8849 10217 8861 10251
rect 8895 10248 8907 10251
rect 11882 10248 11888 10260
rect 8895 10220 11888 10248
rect 8895 10217 8907 10220
rect 8849 10211 8907 10217
rect 8864 10180 8892 10211
rect 11882 10208 11888 10220
rect 11940 10248 11946 10260
rect 12621 10251 12679 10257
rect 12621 10248 12633 10251
rect 11940 10220 12633 10248
rect 11940 10208 11946 10220
rect 12621 10217 12633 10220
rect 12667 10248 12679 10251
rect 12667 10220 13032 10248
rect 12667 10217 12679 10220
rect 12621 10211 12679 10217
rect 13004 10192 13032 10220
rect 14458 10208 14464 10260
rect 14516 10248 14522 10260
rect 14553 10251 14611 10257
rect 14553 10248 14565 10251
rect 14516 10220 14565 10248
rect 14516 10208 14522 10220
rect 14553 10217 14565 10220
rect 14599 10217 14611 10251
rect 17494 10248 17500 10260
rect 17455 10220 17500 10248
rect 14553 10211 14611 10217
rect 17494 10208 17500 10220
rect 17552 10208 17558 10260
rect 17862 10248 17868 10260
rect 17823 10220 17868 10248
rect 17862 10208 17868 10220
rect 17920 10208 17926 10260
rect 3804 10152 5120 10180
rect 5460 10152 8892 10180
rect 3804 10121 3832 10152
rect 3053 10115 3111 10121
rect 3053 10081 3065 10115
rect 3099 10112 3111 10115
rect 3789 10115 3847 10121
rect 3099 10084 3740 10112
rect 3099 10081 3111 10084
rect 3053 10075 3111 10081
rect 1302 10004 1308 10056
rect 1360 10044 1366 10056
rect 1397 10047 1455 10053
rect 1397 10044 1409 10047
rect 1360 10016 1409 10044
rect 1360 10004 1366 10016
rect 1397 10013 1409 10016
rect 1443 10013 1455 10047
rect 3712 10044 3740 10084
rect 3789 10081 3801 10115
rect 3835 10081 3847 10115
rect 4890 10112 4896 10124
rect 4851 10084 4896 10112
rect 3789 10075 3847 10081
rect 4890 10072 4896 10084
rect 4948 10112 4954 10124
rect 5460 10112 5488 10152
rect 9766 10140 9772 10192
rect 9824 10180 9830 10192
rect 9922 10183 9980 10189
rect 9922 10180 9934 10183
rect 9824 10152 9934 10180
rect 9824 10140 9830 10152
rect 9922 10149 9934 10152
rect 9968 10149 9980 10183
rect 9922 10143 9980 10149
rect 12986 10140 12992 10192
rect 13044 10140 13050 10192
rect 13170 10140 13176 10192
rect 13228 10180 13234 10192
rect 13418 10183 13476 10189
rect 13418 10180 13430 10183
rect 13228 10152 13430 10180
rect 13228 10140 13234 10152
rect 13418 10149 13430 10152
rect 13464 10149 13476 10183
rect 16384 10183 16442 10189
rect 13418 10143 13476 10149
rect 15764 10152 16344 10180
rect 5718 10112 5724 10124
rect 4948 10084 5488 10112
rect 5679 10084 5724 10112
rect 4948 10072 4954 10084
rect 5718 10072 5724 10084
rect 5776 10072 5782 10124
rect 6080 10115 6138 10121
rect 6080 10081 6092 10115
rect 6126 10112 6138 10115
rect 8846 10112 8852 10124
rect 6126 10084 8852 10112
rect 6126 10081 6138 10084
rect 6080 10075 6138 10081
rect 8846 10072 8852 10084
rect 8904 10112 8910 10124
rect 9677 10115 9735 10121
rect 8904 10084 9076 10112
rect 8904 10072 8910 10084
rect 4614 10044 4620 10056
rect 3712 10016 4620 10044
rect 1397 10007 1455 10013
rect 4614 10004 4620 10016
rect 4672 10004 4678 10056
rect 5077 10047 5135 10053
rect 5077 10013 5089 10047
rect 5123 10044 5135 10047
rect 5166 10044 5172 10056
rect 5123 10016 5172 10044
rect 5123 10013 5135 10016
rect 5077 10007 5135 10013
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10013 5871 10047
rect 5813 10007 5871 10013
rect 4798 9936 4804 9988
rect 4856 9976 4862 9988
rect 5534 9976 5540 9988
rect 4856 9948 5540 9976
rect 4856 9936 4862 9948
rect 5534 9936 5540 9948
rect 5592 9936 5598 9988
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 2832 9880 2877 9908
rect 2832 9868 2838 9880
rect 3050 9868 3056 9920
rect 3108 9908 3114 9920
rect 3237 9911 3295 9917
rect 3237 9908 3249 9911
rect 3108 9880 3249 9908
rect 3108 9868 3114 9880
rect 3237 9877 3249 9880
rect 3283 9877 3295 9911
rect 5828 9908 5856 10007
rect 7190 10004 7196 10056
rect 7248 10044 7254 10056
rect 7926 10044 7932 10056
rect 7248 10016 7932 10044
rect 7248 10004 7254 10016
rect 7926 10004 7932 10016
rect 7984 10004 7990 10056
rect 8018 10004 8024 10056
rect 8076 10044 8082 10056
rect 9048 10053 9076 10084
rect 9677 10081 9689 10115
rect 9723 10112 9735 10115
rect 10410 10112 10416 10124
rect 9723 10084 10416 10112
rect 9723 10081 9735 10084
rect 9677 10075 9735 10081
rect 10410 10072 10416 10084
rect 10468 10072 10474 10124
rect 10502 10072 10508 10124
rect 10560 10112 10566 10124
rect 10870 10112 10876 10124
rect 10560 10084 10876 10112
rect 10560 10072 10566 10084
rect 10870 10072 10876 10084
rect 10928 10112 10934 10124
rect 12342 10112 12348 10124
rect 10928 10084 12348 10112
rect 10928 10072 10934 10084
rect 12342 10072 12348 10084
rect 12400 10112 12406 10124
rect 12529 10115 12587 10121
rect 12529 10112 12541 10115
rect 12400 10084 12541 10112
rect 12400 10072 12406 10084
rect 12529 10081 12541 10084
rect 12575 10081 12587 10115
rect 13188 10112 13216 10140
rect 12529 10075 12587 10081
rect 12820 10084 13216 10112
rect 8941 10047 8999 10053
rect 8076 10016 8121 10044
rect 8076 10004 8082 10016
rect 8941 10013 8953 10047
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 9033 10047 9091 10053
rect 9033 10013 9045 10047
rect 9079 10013 9091 10047
rect 9033 10007 9091 10013
rect 7469 9979 7527 9985
rect 7469 9945 7481 9979
rect 7515 9976 7527 9979
rect 8956 9976 8984 10007
rect 10778 10004 10784 10056
rect 10836 10044 10842 10056
rect 12820 10053 12848 10084
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 15657 10115 15715 10121
rect 15657 10112 15669 10115
rect 13872 10084 15669 10112
rect 13872 10072 13878 10084
rect 15657 10081 15669 10084
rect 15703 10081 15715 10115
rect 15657 10075 15715 10081
rect 12805 10047 12863 10053
rect 10836 10016 12572 10044
rect 10836 10004 10842 10016
rect 11054 9976 11060 9988
rect 7515 9948 8984 9976
rect 10967 9948 11060 9976
rect 7515 9945 7527 9948
rect 7469 9939 7527 9945
rect 11054 9936 11060 9948
rect 11112 9976 11118 9988
rect 12250 9976 12256 9988
rect 11112 9948 12256 9976
rect 11112 9936 11118 9948
rect 12250 9936 12256 9948
rect 12308 9936 12314 9988
rect 6178 9908 6184 9920
rect 5828 9880 6184 9908
rect 3237 9871 3295 9877
rect 6178 9868 6184 9880
rect 6236 9868 6242 9920
rect 6730 9868 6736 9920
rect 6788 9908 6794 9920
rect 7193 9911 7251 9917
rect 7193 9908 7205 9911
rect 6788 9880 7205 9908
rect 6788 9868 6794 9880
rect 7193 9877 7205 9880
rect 7239 9877 7251 9911
rect 7193 9871 7251 9877
rect 7926 9868 7932 9920
rect 7984 9908 7990 9920
rect 10870 9908 10876 9920
rect 7984 9880 10876 9908
rect 7984 9868 7990 9880
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 12161 9911 12219 9917
rect 12161 9877 12173 9911
rect 12207 9908 12219 9911
rect 12434 9908 12440 9920
rect 12207 9880 12440 9908
rect 12207 9877 12219 9880
rect 12161 9871 12219 9877
rect 12434 9868 12440 9880
rect 12492 9868 12498 9920
rect 12544 9908 12572 10016
rect 12805 10013 12817 10047
rect 12851 10013 12863 10047
rect 12805 10007 12863 10013
rect 13173 10047 13231 10053
rect 13173 10013 13185 10047
rect 13219 10013 13231 10047
rect 15764 10044 15792 10152
rect 16206 10072 16212 10124
rect 16264 10072 16270 10124
rect 16316 10112 16344 10152
rect 16384 10149 16396 10183
rect 16430 10180 16442 10183
rect 16758 10180 16764 10192
rect 16430 10152 16764 10180
rect 16430 10149 16442 10152
rect 16384 10143 16442 10149
rect 16758 10140 16764 10152
rect 16816 10180 16822 10192
rect 17770 10180 17776 10192
rect 16816 10152 17776 10180
rect 16816 10140 16822 10152
rect 17770 10140 17776 10152
rect 17828 10140 17834 10192
rect 17218 10112 17224 10124
rect 16316 10084 17224 10112
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 13173 10007 13231 10013
rect 14200 10016 15792 10044
rect 16117 10047 16175 10053
rect 12710 9936 12716 9988
rect 12768 9976 12774 9988
rect 13188 9976 13216 10007
rect 12768 9948 13216 9976
rect 12768 9936 12774 9948
rect 14200 9908 14228 10016
rect 16117 10013 16129 10047
rect 16163 10044 16175 10047
rect 16224 10044 16252 10072
rect 16163 10016 16252 10044
rect 16163 10013 16175 10016
rect 16117 10007 16175 10013
rect 15473 9979 15531 9985
rect 15473 9945 15485 9979
rect 15519 9976 15531 9979
rect 15746 9976 15752 9988
rect 15519 9948 15752 9976
rect 15519 9945 15531 9948
rect 15473 9939 15531 9945
rect 15746 9936 15752 9948
rect 15804 9976 15810 9988
rect 16132 9976 16160 10007
rect 15804 9948 16160 9976
rect 15804 9936 15810 9948
rect 12544 9880 14228 9908
rect 14366 9868 14372 9920
rect 14424 9908 14430 9920
rect 17862 9908 17868 9920
rect 14424 9880 17868 9908
rect 14424 9868 14430 9880
rect 17862 9868 17868 9880
rect 17920 9868 17926 9920
rect 1104 9818 18860 9840
rect 1104 9766 3947 9818
rect 3999 9766 4011 9818
rect 4063 9766 4075 9818
rect 4127 9766 4139 9818
rect 4191 9766 9878 9818
rect 9930 9766 9942 9818
rect 9994 9766 10006 9818
rect 10058 9766 10070 9818
rect 10122 9766 15808 9818
rect 15860 9766 15872 9818
rect 15924 9766 15936 9818
rect 15988 9766 16000 9818
rect 16052 9766 18860 9818
rect 1104 9744 18860 9766
rect 3602 9664 3608 9716
rect 3660 9704 3666 9716
rect 5350 9704 5356 9716
rect 3660 9676 5356 9704
rect 3660 9664 3666 9676
rect 5350 9664 5356 9676
rect 5408 9664 5414 9716
rect 5810 9664 5816 9716
rect 5868 9704 5874 9716
rect 9766 9704 9772 9716
rect 5868 9676 9772 9704
rect 5868 9664 5874 9676
rect 9766 9664 9772 9676
rect 9824 9704 9830 9716
rect 10778 9704 10784 9716
rect 9824 9676 10784 9704
rect 9824 9664 9830 9676
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 10962 9664 10968 9716
rect 11020 9704 11026 9716
rect 16482 9704 16488 9716
rect 11020 9676 16488 9704
rect 11020 9664 11026 9676
rect 16482 9664 16488 9676
rect 16540 9664 16546 9716
rect 4338 9596 4344 9648
rect 4396 9636 4402 9648
rect 4433 9639 4491 9645
rect 4433 9636 4445 9639
rect 4396 9608 4445 9636
rect 4396 9596 4402 9608
rect 4433 9605 4445 9608
rect 4479 9605 4491 9639
rect 4433 9599 4491 9605
rect 6380 9608 8800 9636
rect 6380 9580 6408 9608
rect 1302 9528 1308 9580
rect 1360 9568 1366 9580
rect 2133 9571 2191 9577
rect 2133 9568 2145 9571
rect 1360 9540 2145 9568
rect 1360 9528 1366 9540
rect 2133 9537 2145 9540
rect 2179 9537 2191 9571
rect 2133 9531 2191 9537
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 4893 9571 4951 9577
rect 4893 9568 4905 9571
rect 4120 9540 4905 9568
rect 4120 9528 4126 9540
rect 4893 9537 4905 9540
rect 4939 9537 4951 9571
rect 4893 9531 4951 9537
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9568 5135 9571
rect 5166 9568 5172 9580
rect 5123 9540 5172 9568
rect 5123 9537 5135 9540
rect 5077 9531 5135 9537
rect 1581 9503 1639 9509
rect 1581 9469 1593 9503
rect 1627 9469 1639 9503
rect 1581 9463 1639 9469
rect 2400 9503 2458 9509
rect 2400 9469 2412 9503
rect 2446 9500 2458 9503
rect 2774 9500 2780 9512
rect 2446 9472 2780 9500
rect 2446 9469 2458 9472
rect 2400 9463 2458 9469
rect 1596 9432 1624 9463
rect 2774 9460 2780 9472
rect 2832 9460 2838 9512
rect 3789 9503 3847 9509
rect 3789 9469 3801 9503
rect 3835 9500 3847 9503
rect 4522 9500 4528 9512
rect 3835 9472 4528 9500
rect 3835 9469 3847 9472
rect 3789 9463 3847 9469
rect 4522 9460 4528 9472
rect 4580 9460 4586 9512
rect 4908 9500 4936 9531
rect 5166 9528 5172 9540
rect 5224 9528 5230 9580
rect 6362 9568 6368 9580
rect 6275 9540 6368 9568
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 7745 9571 7803 9577
rect 7745 9568 7757 9571
rect 6788 9540 7757 9568
rect 6788 9528 6794 9540
rect 7745 9537 7757 9540
rect 7791 9537 7803 9571
rect 8570 9568 8576 9580
rect 7745 9531 7803 9537
rect 8036 9540 8576 9568
rect 7190 9500 7196 9512
rect 4908 9472 7196 9500
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 7561 9503 7619 9509
rect 7561 9469 7573 9503
rect 7607 9500 7619 9503
rect 8036 9500 8064 9540
rect 8570 9528 8576 9540
rect 8628 9528 8634 9580
rect 8772 9577 8800 9608
rect 12710 9596 12716 9648
rect 12768 9636 12774 9648
rect 13446 9636 13452 9648
rect 12768 9608 13032 9636
rect 13407 9608 13452 9636
rect 12768 9596 12774 9608
rect 8757 9571 8815 9577
rect 8757 9537 8769 9571
rect 8803 9537 8815 9571
rect 8757 9531 8815 9537
rect 9217 9571 9275 9577
rect 9217 9537 9229 9571
rect 9263 9568 9275 9571
rect 9674 9568 9680 9580
rect 9263 9540 9680 9568
rect 9263 9537 9275 9540
rect 9217 9531 9275 9537
rect 9674 9528 9680 9540
rect 9732 9528 9738 9580
rect 10870 9528 10876 9580
rect 10928 9568 10934 9580
rect 10928 9540 12940 9568
rect 10928 9528 10934 9540
rect 7607 9472 8064 9500
rect 7607 9469 7619 9472
rect 7561 9463 7619 9469
rect 8110 9460 8116 9512
rect 8168 9500 8174 9512
rect 8665 9503 8723 9509
rect 8665 9500 8677 9503
rect 8168 9472 8677 9500
rect 8168 9460 8174 9472
rect 8665 9469 8677 9472
rect 8711 9469 8723 9503
rect 8665 9463 8723 9469
rect 9861 9503 9919 9509
rect 9861 9469 9873 9503
rect 9907 9500 9919 9503
rect 10410 9500 10416 9512
rect 9907 9472 10416 9500
rect 9907 9469 9919 9472
rect 9861 9463 9919 9469
rect 10410 9460 10416 9472
rect 10468 9460 10474 9512
rect 11054 9500 11060 9512
rect 10888 9472 11060 9500
rect 5902 9432 5908 9444
rect 1596 9404 5908 9432
rect 5902 9392 5908 9404
rect 5960 9392 5966 9444
rect 8573 9435 8631 9441
rect 8573 9432 8585 9435
rect 7208 9404 8585 9432
rect 1765 9367 1823 9373
rect 1765 9333 1777 9367
rect 1811 9364 1823 9367
rect 3142 9364 3148 9376
rect 1811 9336 3148 9364
rect 1811 9333 1823 9336
rect 1765 9327 1823 9333
rect 3142 9324 3148 9336
rect 3200 9324 3206 9376
rect 3510 9364 3516 9376
rect 3471 9336 3516 9364
rect 3510 9324 3516 9336
rect 3568 9324 3574 9376
rect 3602 9324 3608 9376
rect 3660 9364 3666 9376
rect 3973 9367 4031 9373
rect 3973 9364 3985 9367
rect 3660 9336 3985 9364
rect 3660 9324 3666 9336
rect 3973 9333 3985 9336
rect 4019 9333 4031 9367
rect 3973 9327 4031 9333
rect 4706 9324 4712 9376
rect 4764 9364 4770 9376
rect 4801 9367 4859 9373
rect 4801 9364 4813 9367
rect 4764 9336 4813 9364
rect 4764 9324 4770 9336
rect 4801 9333 4813 9336
rect 4847 9333 4859 9367
rect 4801 9327 4859 9333
rect 5721 9367 5779 9373
rect 5721 9333 5733 9367
rect 5767 9364 5779 9367
rect 5810 9364 5816 9376
rect 5767 9336 5816 9364
rect 5767 9333 5779 9336
rect 5721 9327 5779 9333
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 6086 9364 6092 9376
rect 6047 9336 6092 9364
rect 6086 9324 6092 9336
rect 6144 9324 6150 9376
rect 6178 9324 6184 9376
rect 6236 9364 6242 9376
rect 7208 9373 7236 9404
rect 8573 9401 8585 9404
rect 8619 9401 8631 9435
rect 8573 9395 8631 9401
rect 10128 9435 10186 9441
rect 10128 9401 10140 9435
rect 10174 9432 10186 9435
rect 10888 9432 10916 9472
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 12912 9441 12940 9540
rect 13004 9500 13032 9608
rect 13446 9596 13452 9608
rect 13504 9636 13510 9648
rect 13814 9636 13820 9648
rect 13504 9608 13820 9636
rect 13504 9596 13510 9608
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 16666 9596 16672 9648
rect 16724 9636 16730 9648
rect 16761 9639 16819 9645
rect 16761 9636 16773 9639
rect 16724 9608 16773 9636
rect 16724 9596 16730 9608
rect 16761 9605 16773 9608
rect 16807 9605 16819 9639
rect 16761 9599 16819 9605
rect 13081 9571 13139 9577
rect 13081 9537 13093 9571
rect 13127 9568 13139 9571
rect 13170 9568 13176 9580
rect 13127 9540 13176 9568
rect 13127 9537 13139 9540
rect 13081 9531 13139 9537
rect 13170 9528 13176 9540
rect 13228 9568 13234 9580
rect 13906 9568 13912 9580
rect 13228 9540 13912 9568
rect 13228 9528 13234 9540
rect 13906 9528 13912 9540
rect 13964 9528 13970 9580
rect 14182 9568 14188 9580
rect 14143 9540 14188 9568
rect 14182 9528 14188 9540
rect 14240 9528 14246 9580
rect 17402 9568 17408 9580
rect 17363 9540 17408 9568
rect 17402 9528 17408 9540
rect 17460 9528 17466 9580
rect 13633 9503 13691 9509
rect 13633 9500 13645 9503
rect 13004 9472 13645 9500
rect 13633 9469 13645 9472
rect 13679 9469 13691 9503
rect 17221 9503 17279 9509
rect 17221 9500 17233 9503
rect 13633 9463 13691 9469
rect 14200 9472 17233 9500
rect 10174 9404 10916 9432
rect 12897 9435 12955 9441
rect 10174 9401 10186 9404
rect 10128 9395 10186 9401
rect 12897 9401 12909 9435
rect 12943 9432 12955 9435
rect 14200 9432 14228 9472
rect 17221 9469 17233 9472
rect 17267 9469 17279 9503
rect 17221 9463 17279 9469
rect 14458 9441 14464 9444
rect 14452 9432 14464 9441
rect 12943 9404 14228 9432
rect 14419 9404 14464 9432
rect 12943 9401 12955 9404
rect 12897 9395 12955 9401
rect 14452 9395 14464 9404
rect 14458 9392 14464 9395
rect 14516 9392 14522 9444
rect 15286 9432 15292 9444
rect 14568 9404 15292 9432
rect 7193 9367 7251 9373
rect 6236 9336 6281 9364
rect 6236 9324 6242 9336
rect 7193 9333 7205 9367
rect 7239 9333 7251 9367
rect 7650 9364 7656 9376
rect 7611 9336 7656 9364
rect 7193 9327 7251 9333
rect 7650 9324 7656 9336
rect 7708 9324 7714 9376
rect 8202 9364 8208 9376
rect 8163 9336 8208 9364
rect 8202 9324 8208 9336
rect 8260 9324 8266 9376
rect 8386 9324 8392 9376
rect 8444 9364 8450 9376
rect 9490 9364 9496 9376
rect 8444 9336 9496 9364
rect 8444 9324 8450 9336
rect 9490 9324 9496 9336
rect 9548 9364 9554 9376
rect 11241 9367 11299 9373
rect 11241 9364 11253 9367
rect 9548 9336 11253 9364
rect 9548 9324 9554 9336
rect 11241 9333 11253 9336
rect 11287 9333 11299 9367
rect 11241 9327 11299 9333
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 12526 9364 12532 9376
rect 12483 9336 12532 9364
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 12526 9324 12532 9336
rect 12584 9324 12590 9376
rect 12805 9367 12863 9373
rect 12805 9333 12817 9367
rect 12851 9364 12863 9367
rect 14568 9364 14596 9404
rect 15286 9392 15292 9404
rect 15344 9432 15350 9444
rect 15344 9404 17172 9432
rect 15344 9392 15350 9404
rect 12851 9336 14596 9364
rect 12851 9333 12863 9336
rect 12805 9327 12863 9333
rect 15378 9324 15384 9376
rect 15436 9364 15442 9376
rect 17144 9373 17172 9404
rect 15565 9367 15623 9373
rect 15565 9364 15577 9367
rect 15436 9336 15577 9364
rect 15436 9324 15442 9336
rect 15565 9333 15577 9336
rect 15611 9333 15623 9367
rect 15565 9327 15623 9333
rect 17129 9367 17187 9373
rect 17129 9333 17141 9367
rect 17175 9364 17187 9367
rect 17310 9364 17316 9376
rect 17175 9336 17316 9364
rect 17175 9333 17187 9336
rect 17129 9327 17187 9333
rect 17310 9324 17316 9336
rect 17368 9324 17374 9376
rect 1104 9274 18860 9296
rect 1104 9222 6912 9274
rect 6964 9222 6976 9274
rect 7028 9222 7040 9274
rect 7092 9222 7104 9274
rect 7156 9222 12843 9274
rect 12895 9222 12907 9274
rect 12959 9222 12971 9274
rect 13023 9222 13035 9274
rect 13087 9222 18860 9274
rect 1104 9200 18860 9222
rect 1854 9120 1860 9172
rect 1912 9160 1918 9172
rect 2225 9163 2283 9169
rect 2225 9160 2237 9163
rect 1912 9132 2237 9160
rect 1912 9120 1918 9132
rect 2225 9129 2237 9132
rect 2271 9129 2283 9163
rect 2225 9123 2283 9129
rect 2317 9163 2375 9169
rect 2317 9129 2329 9163
rect 2363 9160 2375 9163
rect 2961 9163 3019 9169
rect 2961 9160 2973 9163
rect 2363 9132 2973 9160
rect 2363 9129 2375 9132
rect 2317 9123 2375 9129
rect 2961 9129 2973 9132
rect 3007 9129 3019 9163
rect 3418 9160 3424 9172
rect 3379 9132 3424 9160
rect 2961 9123 3019 9129
rect 3418 9120 3424 9132
rect 3476 9120 3482 9172
rect 5902 9120 5908 9172
rect 5960 9160 5966 9172
rect 6270 9160 6276 9172
rect 5960 9132 6276 9160
rect 5960 9120 5966 9132
rect 6270 9120 6276 9132
rect 6328 9120 6334 9172
rect 6454 9120 6460 9172
rect 6512 9160 6518 9172
rect 6512 9132 8156 9160
rect 6512 9120 6518 9132
rect 3510 9052 3516 9104
rect 3568 9092 3574 9104
rect 4310 9095 4368 9101
rect 4310 9092 4322 9095
rect 3568 9064 4322 9092
rect 3568 9052 3574 9064
rect 4310 9061 4322 9064
rect 4356 9061 4368 9095
rect 4310 9055 4368 9061
rect 5810 9052 5816 9104
rect 5868 9092 5874 9104
rect 7193 9095 7251 9101
rect 5868 9064 7052 9092
rect 5868 9052 5874 9064
rect 3329 9027 3387 9033
rect 3329 8993 3341 9027
rect 3375 9024 3387 9027
rect 5442 9024 5448 9036
rect 3375 8996 5448 9024
rect 3375 8993 3387 8996
rect 3329 8987 3387 8993
rect 5442 8984 5448 8996
rect 5500 8984 5506 9036
rect 5988 9027 6046 9033
rect 5988 8993 6000 9027
rect 6034 9024 6046 9027
rect 6270 9024 6276 9036
rect 6034 8996 6276 9024
rect 6034 8993 6046 8996
rect 5988 8987 6046 8993
rect 6270 8984 6276 8996
rect 6328 9024 6334 9036
rect 6822 9024 6828 9036
rect 6328 8996 6828 9024
rect 6328 8984 6334 8996
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 7024 9024 7052 9064
rect 7193 9061 7205 9095
rect 7239 9092 7251 9095
rect 7644 9095 7702 9101
rect 7644 9092 7656 9095
rect 7239 9064 7656 9092
rect 7239 9061 7251 9064
rect 7193 9055 7251 9061
rect 7644 9061 7656 9064
rect 7690 9092 7702 9095
rect 8018 9092 8024 9104
rect 7690 9064 8024 9092
rect 7690 9061 7702 9064
rect 7644 9055 7702 9061
rect 8018 9052 8024 9064
rect 8076 9052 8082 9104
rect 8128 9092 8156 9132
rect 8202 9120 8208 9172
rect 8260 9160 8266 9172
rect 10229 9163 10287 9169
rect 10229 9160 10241 9163
rect 8260 9132 10241 9160
rect 8260 9120 8266 9132
rect 10229 9129 10241 9132
rect 10275 9129 10287 9163
rect 10229 9123 10287 9129
rect 11425 9163 11483 9169
rect 11425 9129 11437 9163
rect 11471 9160 11483 9163
rect 11514 9160 11520 9172
rect 11471 9132 11520 9160
rect 11471 9129 11483 9132
rect 11425 9123 11483 9129
rect 11514 9120 11520 9132
rect 11572 9120 11578 9172
rect 11790 9120 11796 9172
rect 11848 9160 11854 9172
rect 12069 9163 12127 9169
rect 12069 9160 12081 9163
rect 11848 9132 12081 9160
rect 11848 9120 11854 9132
rect 12069 9129 12081 9132
rect 12115 9129 12127 9163
rect 12526 9160 12532 9172
rect 12487 9132 12532 9160
rect 12069 9123 12127 9129
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 12989 9163 13047 9169
rect 12989 9129 13001 9163
rect 13035 9160 13047 9163
rect 14182 9160 14188 9172
rect 13035 9132 14188 9160
rect 13035 9129 13047 9132
rect 12989 9123 13047 9129
rect 14182 9120 14188 9132
rect 14240 9160 14246 9172
rect 14550 9160 14556 9172
rect 14240 9132 14556 9160
rect 14240 9120 14246 9132
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 15289 9163 15347 9169
rect 15289 9129 15301 9163
rect 15335 9129 15347 9163
rect 15289 9123 15347 9129
rect 12342 9092 12348 9104
rect 8128 9064 12348 9092
rect 12342 9052 12348 9064
rect 12400 9052 12406 9104
rect 12434 9052 12440 9104
rect 12492 9092 12498 9104
rect 15304 9092 15332 9123
rect 17770 9120 17776 9172
rect 17828 9160 17834 9172
rect 18233 9163 18291 9169
rect 18233 9160 18245 9163
rect 17828 9132 18245 9160
rect 17828 9120 17834 9132
rect 18233 9129 18245 9132
rect 18279 9129 18291 9163
rect 18233 9123 18291 9129
rect 12492 9064 12537 9092
rect 13280 9064 15332 9092
rect 12492 9052 12498 9064
rect 10321 9027 10379 9033
rect 10321 9024 10333 9027
rect 7024 8996 10333 9024
rect 10321 8993 10333 8996
rect 10367 8993 10379 9027
rect 10321 8987 10379 8993
rect 11517 9027 11575 9033
rect 11517 8993 11529 9027
rect 11563 9024 11575 9027
rect 13280 9024 13308 9064
rect 16206 9052 16212 9104
rect 16264 9052 16270 9104
rect 11563 8996 13308 9024
rect 13348 9027 13406 9033
rect 11563 8993 11575 8996
rect 11517 8987 11575 8993
rect 13348 8993 13360 9027
rect 13394 9024 13406 9027
rect 13722 9024 13728 9036
rect 13394 8996 13728 9024
rect 13394 8993 13406 8996
rect 13348 8987 13406 8993
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 13814 8984 13820 9036
rect 13872 9024 13878 9036
rect 15657 9027 15715 9033
rect 15657 9024 15669 9027
rect 13872 8996 15669 9024
rect 13872 8984 13878 8996
rect 15657 8993 15669 8996
rect 15703 8993 15715 9027
rect 16224 9024 16252 9052
rect 16390 9024 16396 9036
rect 16224 8996 16396 9024
rect 15657 8987 15715 8993
rect 16390 8984 16396 8996
rect 16448 9024 16454 9036
rect 16853 9027 16911 9033
rect 16853 9024 16865 9027
rect 16448 8996 16865 9024
rect 16448 8984 16454 8996
rect 16853 8993 16865 8996
rect 16899 8993 16911 9027
rect 16853 8987 16911 8993
rect 17120 9027 17178 9033
rect 17120 8993 17132 9027
rect 17166 9024 17178 9027
rect 17402 9024 17408 9036
rect 17166 8996 17408 9024
rect 17166 8993 17178 8996
rect 17120 8987 17178 8993
rect 17402 8984 17408 8996
rect 17460 8984 17466 9036
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8956 2559 8959
rect 2774 8956 2780 8968
rect 2547 8928 2780 8956
rect 2547 8925 2559 8928
rect 2501 8919 2559 8925
rect 2774 8916 2780 8928
rect 2832 8916 2838 8968
rect 3234 8916 3240 8968
rect 3292 8956 3298 8968
rect 3513 8959 3571 8965
rect 3513 8956 3525 8959
rect 3292 8928 3525 8956
rect 3292 8916 3298 8928
rect 3513 8925 3525 8928
rect 3559 8925 3571 8959
rect 3513 8919 3571 8925
rect 3694 8916 3700 8968
rect 3752 8956 3758 8968
rect 4065 8959 4123 8965
rect 4065 8956 4077 8959
rect 3752 8928 4077 8956
rect 3752 8916 3758 8928
rect 4065 8925 4077 8928
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 5721 8959 5779 8965
rect 5721 8925 5733 8959
rect 5767 8925 5779 8959
rect 7282 8956 7288 8968
rect 5721 8919 5779 8925
rect 7024 8928 7288 8956
rect 1762 8780 1768 8832
rect 1820 8820 1826 8832
rect 1857 8823 1915 8829
rect 1857 8820 1869 8823
rect 1820 8792 1869 8820
rect 1820 8780 1826 8792
rect 1857 8789 1869 8792
rect 1903 8789 1915 8823
rect 1857 8783 1915 8789
rect 4982 8780 4988 8832
rect 5040 8820 5046 8832
rect 5445 8823 5503 8829
rect 5445 8820 5457 8823
rect 5040 8792 5457 8820
rect 5040 8780 5046 8792
rect 5445 8789 5457 8792
rect 5491 8789 5503 8823
rect 5736 8820 5764 8919
rect 7024 8888 7052 8928
rect 7282 8916 7288 8928
rect 7340 8956 7346 8968
rect 7377 8959 7435 8965
rect 7377 8956 7389 8959
rect 7340 8928 7389 8956
rect 7340 8916 7346 8928
rect 7377 8925 7389 8928
rect 7423 8925 7435 8959
rect 9030 8956 9036 8968
rect 8991 8928 9036 8956
rect 7377 8919 7435 8925
rect 9030 8916 9036 8928
rect 9088 8916 9094 8968
rect 10413 8959 10471 8965
rect 10413 8925 10425 8959
rect 10459 8925 10471 8959
rect 10413 8919 10471 8925
rect 11701 8959 11759 8965
rect 11701 8925 11713 8959
rect 11747 8956 11759 8959
rect 11885 8959 11943 8965
rect 11885 8956 11897 8959
rect 11747 8928 11897 8956
rect 11747 8925 11759 8928
rect 11701 8919 11759 8925
rect 11885 8925 11897 8928
rect 11931 8925 11943 8959
rect 12618 8956 12624 8968
rect 12579 8928 12624 8956
rect 11885 8919 11943 8925
rect 6656 8860 7052 8888
rect 7101 8891 7159 8897
rect 6656 8820 6684 8860
rect 7101 8857 7113 8891
rect 7147 8888 7159 8891
rect 7193 8891 7251 8897
rect 7193 8888 7205 8891
rect 7147 8860 7205 8888
rect 7147 8857 7159 8860
rect 7101 8851 7159 8857
rect 7193 8857 7205 8860
rect 7239 8857 7251 8891
rect 10428 8888 10456 8919
rect 12618 8916 12624 8928
rect 12676 8916 12682 8968
rect 12989 8959 13047 8965
rect 12989 8925 13001 8959
rect 13035 8956 13047 8959
rect 13081 8959 13139 8965
rect 13081 8956 13093 8959
rect 13035 8928 13093 8956
rect 13035 8925 13047 8928
rect 12989 8919 13047 8925
rect 13081 8925 13093 8928
rect 13127 8925 13139 8959
rect 13081 8919 13139 8925
rect 14182 8916 14188 8968
rect 14240 8956 14246 8968
rect 15749 8959 15807 8965
rect 15749 8956 15761 8959
rect 14240 8928 15761 8956
rect 14240 8916 14246 8928
rect 15749 8925 15761 8928
rect 15795 8925 15807 8959
rect 15749 8919 15807 8925
rect 15933 8959 15991 8965
rect 15933 8925 15945 8959
rect 15979 8956 15991 8959
rect 16206 8956 16212 8968
rect 15979 8928 16212 8956
rect 15979 8925 15991 8928
rect 15933 8919 15991 8925
rect 16206 8916 16212 8928
rect 16264 8916 16270 8968
rect 7193 8851 7251 8857
rect 8312 8860 10456 8888
rect 11057 8891 11115 8897
rect 5736 8792 6684 8820
rect 5445 8783 5503 8789
rect 6822 8780 6828 8832
rect 6880 8820 6886 8832
rect 8312 8820 8340 8860
rect 11057 8857 11069 8891
rect 11103 8888 11115 8891
rect 12802 8888 12808 8900
rect 11103 8860 12808 8888
rect 11103 8857 11115 8860
rect 11057 8851 11115 8857
rect 12802 8848 12808 8860
rect 12860 8848 12866 8900
rect 16298 8888 16304 8900
rect 14292 8860 16304 8888
rect 6880 8792 8340 8820
rect 8757 8823 8815 8829
rect 6880 8780 6886 8792
rect 8757 8789 8769 8823
rect 8803 8820 8815 8823
rect 8846 8820 8852 8832
rect 8803 8792 8852 8820
rect 8803 8789 8815 8792
rect 8757 8783 8815 8789
rect 8846 8780 8852 8792
rect 8904 8780 8910 8832
rect 9861 8823 9919 8829
rect 9861 8789 9873 8823
rect 9907 8820 9919 8823
rect 10318 8820 10324 8832
rect 9907 8792 10324 8820
rect 9907 8789 9919 8792
rect 9861 8783 9919 8789
rect 10318 8780 10324 8792
rect 10376 8780 10382 8832
rect 11885 8823 11943 8829
rect 11885 8789 11897 8823
rect 11931 8820 11943 8823
rect 14292 8820 14320 8860
rect 16298 8848 16304 8860
rect 16356 8848 16362 8900
rect 14458 8820 14464 8832
rect 11931 8792 14320 8820
rect 14419 8792 14464 8820
rect 11931 8789 11943 8792
rect 11885 8783 11943 8789
rect 14458 8780 14464 8792
rect 14516 8780 14522 8832
rect 1104 8730 18860 8752
rect 1104 8678 3947 8730
rect 3999 8678 4011 8730
rect 4063 8678 4075 8730
rect 4127 8678 4139 8730
rect 4191 8678 9878 8730
rect 9930 8678 9942 8730
rect 9994 8678 10006 8730
rect 10058 8678 10070 8730
rect 10122 8678 15808 8730
rect 15860 8678 15872 8730
rect 15924 8678 15936 8730
rect 15988 8678 16000 8730
rect 16052 8678 18860 8730
rect 1104 8656 18860 8678
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8616 5687 8619
rect 5718 8616 5724 8628
rect 5675 8588 5724 8616
rect 5675 8585 5687 8588
rect 5629 8579 5687 8585
rect 5718 8576 5724 8588
rect 5776 8576 5782 8628
rect 5905 8619 5963 8625
rect 5905 8585 5917 8619
rect 5951 8616 5963 8619
rect 6178 8616 6184 8628
rect 5951 8588 6184 8616
rect 5951 8585 5963 8588
rect 5905 8579 5963 8585
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 7009 8619 7067 8625
rect 7009 8616 7021 8619
rect 6288 8588 7021 8616
rect 3418 8508 3424 8560
rect 3476 8548 3482 8560
rect 4341 8551 4399 8557
rect 4341 8548 4353 8551
rect 3476 8520 4353 8548
rect 3476 8508 3482 8520
rect 4341 8517 4353 8520
rect 4387 8517 4399 8551
rect 4341 8511 4399 8517
rect 5350 8508 5356 8560
rect 5408 8548 5414 8560
rect 6288 8548 6316 8588
rect 7009 8585 7021 8588
rect 7055 8585 7067 8619
rect 10413 8619 10471 8625
rect 10413 8616 10425 8619
rect 7009 8579 7067 8585
rect 7484 8588 10425 8616
rect 7484 8548 7512 8588
rect 10413 8585 10425 8588
rect 10459 8585 10471 8619
rect 12710 8616 12716 8628
rect 10413 8579 10471 8585
rect 11440 8588 12716 8616
rect 5408 8520 6316 8548
rect 6380 8520 7512 8548
rect 5408 8508 5414 8520
rect 1302 8440 1308 8492
rect 1360 8480 1366 8492
rect 1397 8483 1455 8489
rect 1397 8480 1409 8483
rect 1360 8452 1409 8480
rect 1360 8440 1366 8452
rect 1397 8449 1409 8452
rect 1443 8449 1455 8483
rect 1397 8443 1455 8449
rect 3510 8440 3516 8492
rect 3568 8480 3574 8492
rect 3881 8483 3939 8489
rect 3881 8480 3893 8483
rect 3568 8452 3893 8480
rect 3568 8440 3574 8452
rect 3881 8449 3893 8452
rect 3927 8449 3939 8483
rect 4982 8480 4988 8492
rect 4943 8452 4988 8480
rect 3881 8443 3939 8449
rect 4982 8440 4988 8452
rect 5040 8440 5046 8492
rect 2498 8372 2504 8424
rect 2556 8412 2562 8424
rect 3697 8415 3755 8421
rect 2556 8384 3648 8412
rect 2556 8372 2562 8384
rect 1664 8347 1722 8353
rect 1664 8313 1676 8347
rect 1710 8344 1722 8347
rect 2682 8344 2688 8356
rect 1710 8316 2688 8344
rect 1710 8313 1722 8316
rect 1664 8307 1722 8313
rect 2682 8304 2688 8316
rect 2740 8304 2746 8356
rect 3620 8344 3648 8384
rect 3697 8381 3709 8415
rect 3743 8412 3755 8415
rect 4246 8412 4252 8424
rect 3743 8384 4252 8412
rect 3743 8381 3755 8384
rect 3697 8375 3755 8381
rect 4246 8372 4252 8384
rect 4304 8372 4310 8424
rect 4798 8412 4804 8424
rect 4759 8384 4804 8412
rect 4798 8372 4804 8384
rect 4856 8372 4862 8424
rect 5813 8415 5871 8421
rect 5813 8381 5825 8415
rect 5859 8412 5871 8415
rect 6380 8412 6408 8520
rect 6454 8440 6460 8492
rect 6512 8440 6518 8492
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8480 6607 8483
rect 6730 8480 6736 8492
rect 6595 8452 6736 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 5859 8384 6408 8412
rect 6472 8412 6500 8440
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 6472 8384 6837 8412
rect 5859 8381 5871 8384
rect 5813 8375 5871 8381
rect 6825 8381 6837 8384
rect 6871 8381 6883 8415
rect 6825 8375 6883 8381
rect 7190 8372 7196 8424
rect 7248 8412 7254 8424
rect 7469 8415 7527 8421
rect 7469 8412 7481 8415
rect 7248 8384 7481 8412
rect 7248 8372 7254 8384
rect 7469 8381 7481 8384
rect 7515 8381 7527 8415
rect 9125 8415 9183 8421
rect 9125 8412 9137 8415
rect 7469 8375 7527 8381
rect 7576 8384 9137 8412
rect 3789 8347 3847 8353
rect 3789 8344 3801 8347
rect 3620 8316 3801 8344
rect 3789 8313 3801 8316
rect 3835 8344 3847 8347
rect 4062 8344 4068 8356
rect 3835 8316 4068 8344
rect 3835 8313 3847 8316
rect 3789 8307 3847 8313
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 4430 8304 4436 8356
rect 4488 8344 4494 8356
rect 4709 8347 4767 8353
rect 4709 8344 4721 8347
rect 4488 8316 4721 8344
rect 4488 8304 4494 8316
rect 4709 8313 4721 8316
rect 4755 8344 4767 8347
rect 5718 8344 5724 8356
rect 4755 8316 5724 8344
rect 4755 8313 4767 8316
rect 4709 8307 4767 8313
rect 5718 8304 5724 8316
rect 5776 8304 5782 8356
rect 6365 8347 6423 8353
rect 6365 8313 6377 8347
rect 6411 8344 6423 8347
rect 7282 8344 7288 8356
rect 6411 8316 7288 8344
rect 6411 8313 6423 8316
rect 6365 8307 6423 8313
rect 7282 8304 7288 8316
rect 7340 8304 7346 8356
rect 2777 8279 2835 8285
rect 2777 8245 2789 8279
rect 2823 8276 2835 8279
rect 2866 8276 2872 8288
rect 2823 8248 2872 8276
rect 2823 8245 2835 8248
rect 2777 8239 2835 8245
rect 2866 8236 2872 8248
rect 2924 8236 2930 8288
rect 3326 8276 3332 8288
rect 3287 8248 3332 8276
rect 3326 8236 3332 8248
rect 3384 8236 3390 8288
rect 3970 8236 3976 8288
rect 4028 8276 4034 8288
rect 6273 8279 6331 8285
rect 6273 8276 6285 8279
rect 4028 8248 6285 8276
rect 4028 8236 4034 8248
rect 6273 8245 6285 8248
rect 6319 8276 6331 8279
rect 6454 8276 6460 8288
rect 6319 8248 6460 8276
rect 6319 8245 6331 8248
rect 6273 8239 6331 8245
rect 6454 8236 6460 8248
rect 6512 8236 6518 8288
rect 6546 8236 6552 8288
rect 6604 8276 6610 8288
rect 7576 8276 7604 8384
rect 9125 8381 9137 8384
rect 9171 8381 9183 8415
rect 10428 8412 10456 8579
rect 10962 8548 10968 8560
rect 10923 8520 10968 8548
rect 10962 8508 10968 8520
rect 11020 8508 11026 8560
rect 11440 8489 11468 8588
rect 12710 8576 12716 8588
rect 12768 8576 12774 8628
rect 12802 8576 12808 8628
rect 12860 8616 12866 8628
rect 13817 8619 13875 8625
rect 12860 8588 13400 8616
rect 12860 8576 12866 8588
rect 11977 8551 12035 8557
rect 11977 8517 11989 8551
rect 12023 8548 12035 8551
rect 12342 8548 12348 8560
rect 12023 8520 12348 8548
rect 12023 8517 12035 8520
rect 11977 8511 12035 8517
rect 12342 8508 12348 8520
rect 12400 8508 12406 8560
rect 13372 8548 13400 8588
rect 13817 8585 13829 8619
rect 13863 8616 13875 8619
rect 13906 8616 13912 8628
rect 13863 8588 13912 8616
rect 13863 8585 13875 8588
rect 13817 8579 13875 8585
rect 13906 8576 13912 8588
rect 13964 8576 13970 8628
rect 16390 8616 16396 8628
rect 16040 8588 16396 8616
rect 13372 8520 15056 8548
rect 11425 8483 11483 8489
rect 11425 8449 11437 8483
rect 11471 8449 11483 8483
rect 11606 8480 11612 8492
rect 11567 8452 11612 8480
rect 11425 8443 11483 8449
rect 11606 8440 11612 8452
rect 11664 8440 11670 8492
rect 14458 8440 14464 8492
rect 14516 8480 14522 8492
rect 14921 8483 14979 8489
rect 14921 8480 14933 8483
rect 14516 8452 14933 8480
rect 14516 8440 14522 8452
rect 14921 8449 14933 8452
rect 14967 8449 14979 8483
rect 14921 8443 14979 8449
rect 12161 8415 12219 8421
rect 12161 8412 12173 8415
rect 10428 8384 12173 8412
rect 9125 8375 9183 8381
rect 12161 8381 12173 8384
rect 12207 8381 12219 8415
rect 12161 8375 12219 8381
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8412 12495 8415
rect 13906 8412 13912 8424
rect 12483 8384 13912 8412
rect 12483 8381 12495 8384
rect 12437 8375 12495 8381
rect 13906 8372 13912 8384
rect 13964 8372 13970 8424
rect 7736 8347 7794 8353
rect 7736 8313 7748 8347
rect 7782 8344 7794 8347
rect 8386 8344 8392 8356
rect 7782 8316 8392 8344
rect 7782 8313 7794 8316
rect 7736 8307 7794 8313
rect 8386 8304 8392 8316
rect 8444 8304 8450 8356
rect 12526 8304 12532 8356
rect 12584 8344 12590 8356
rect 12682 8347 12740 8353
rect 12682 8344 12694 8347
rect 12584 8316 12694 8344
rect 12584 8304 12590 8316
rect 12682 8313 12694 8316
rect 12728 8313 12740 8347
rect 14734 8344 14740 8356
rect 14695 8316 14740 8344
rect 12682 8307 12740 8313
rect 14734 8304 14740 8316
rect 14792 8304 14798 8356
rect 14829 8347 14887 8353
rect 14829 8313 14841 8347
rect 14875 8344 14887 8347
rect 14918 8344 14924 8356
rect 14875 8316 14924 8344
rect 14875 8313 14887 8316
rect 14829 8307 14887 8313
rect 14918 8304 14924 8316
rect 14976 8304 14982 8356
rect 15028 8344 15056 8520
rect 16040 8492 16068 8588
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 17402 8616 17408 8628
rect 17363 8588 17408 8616
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 16022 8480 16028 8492
rect 15935 8452 16028 8480
rect 16022 8440 16028 8452
rect 16080 8440 16086 8492
rect 15930 8372 15936 8424
rect 15988 8412 15994 8424
rect 16298 8421 16304 8424
rect 16292 8412 16304 8421
rect 15988 8384 16304 8412
rect 15988 8372 15994 8384
rect 16292 8375 16304 8384
rect 16298 8372 16304 8375
rect 16356 8372 16362 8424
rect 18046 8412 18052 8424
rect 18007 8384 18052 8412
rect 18046 8372 18052 8384
rect 18104 8372 18110 8424
rect 16482 8344 16488 8356
rect 15028 8316 16488 8344
rect 16482 8304 16488 8316
rect 16540 8304 16546 8356
rect 6604 8248 7604 8276
rect 6604 8236 6610 8248
rect 7650 8236 7656 8288
rect 7708 8276 7714 8288
rect 8202 8276 8208 8288
rect 7708 8248 8208 8276
rect 7708 8236 7714 8248
rect 8202 8236 8208 8248
rect 8260 8236 8266 8288
rect 8754 8236 8760 8288
rect 8812 8276 8818 8288
rect 8849 8279 8907 8285
rect 8849 8276 8861 8279
rect 8812 8248 8861 8276
rect 8812 8236 8818 8248
rect 8849 8245 8861 8248
rect 8895 8245 8907 8279
rect 8849 8239 8907 8245
rect 8938 8236 8944 8288
rect 8996 8276 9002 8288
rect 11054 8276 11060 8288
rect 8996 8248 11060 8276
rect 8996 8236 9002 8248
rect 11054 8236 11060 8248
rect 11112 8236 11118 8288
rect 11330 8276 11336 8288
rect 11291 8248 11336 8276
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 12434 8236 12440 8288
rect 12492 8276 12498 8288
rect 13170 8276 13176 8288
rect 12492 8248 13176 8276
rect 12492 8236 12498 8248
rect 13170 8236 13176 8248
rect 13228 8236 13234 8288
rect 14366 8276 14372 8288
rect 14327 8248 14372 8276
rect 14366 8236 14372 8248
rect 14424 8236 14430 8288
rect 15654 8236 15660 8288
rect 15712 8276 15718 8288
rect 16574 8276 16580 8288
rect 15712 8248 16580 8276
rect 15712 8236 15718 8248
rect 16574 8236 16580 8248
rect 16632 8236 16638 8288
rect 18230 8276 18236 8288
rect 18191 8248 18236 8276
rect 18230 8236 18236 8248
rect 18288 8236 18294 8288
rect 1104 8186 18860 8208
rect 1104 8134 6912 8186
rect 6964 8134 6976 8186
rect 7028 8134 7040 8186
rect 7092 8134 7104 8186
rect 7156 8134 12843 8186
rect 12895 8134 12907 8186
rect 12959 8134 12971 8186
rect 13023 8134 13035 8186
rect 13087 8134 18860 8186
rect 1104 8112 18860 8134
rect 2409 8075 2467 8081
rect 2409 8041 2421 8075
rect 2455 8072 2467 8075
rect 2961 8075 3019 8081
rect 2961 8072 2973 8075
rect 2455 8044 2973 8072
rect 2455 8041 2467 8044
rect 2409 8035 2467 8041
rect 2961 8041 2973 8044
rect 3007 8041 3019 8075
rect 2961 8035 3019 8041
rect 3326 8032 3332 8084
rect 3384 8072 3390 8084
rect 3421 8075 3479 8081
rect 3421 8072 3433 8075
rect 3384 8044 3433 8072
rect 3384 8032 3390 8044
rect 3421 8041 3433 8044
rect 3467 8041 3479 8075
rect 3421 8035 3479 8041
rect 6086 8032 6092 8084
rect 6144 8072 6150 8084
rect 6273 8075 6331 8081
rect 6273 8072 6285 8075
rect 6144 8044 6285 8072
rect 6144 8032 6150 8044
rect 6273 8041 6285 8044
rect 6319 8041 6331 8075
rect 6273 8035 6331 8041
rect 6454 8032 6460 8084
rect 6512 8072 6518 8084
rect 6641 8075 6699 8081
rect 6641 8072 6653 8075
rect 6512 8044 6653 8072
rect 6512 8032 6518 8044
rect 6641 8041 6653 8044
rect 6687 8072 6699 8075
rect 7101 8075 7159 8081
rect 6687 8044 6960 8072
rect 6687 8041 6699 8044
rect 6641 8035 6699 8041
rect 4798 8004 4804 8016
rect 1412 7976 4804 8004
rect 1412 7945 1440 7976
rect 4798 7964 4804 7976
rect 4856 7964 4862 8016
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7905 1455 7939
rect 2314 7936 2320 7948
rect 2275 7908 2320 7936
rect 1397 7899 1455 7905
rect 2314 7896 2320 7908
rect 2372 7896 2378 7948
rect 2682 7896 2688 7948
rect 2740 7936 2746 7948
rect 2740 7908 3280 7936
rect 2740 7896 2746 7908
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7868 2651 7871
rect 2866 7868 2872 7880
rect 2639 7840 2872 7868
rect 2639 7837 2651 7840
rect 2593 7831 2651 7837
rect 2866 7828 2872 7840
rect 2924 7828 2930 7880
rect 3252 7868 3280 7908
rect 3326 7896 3332 7948
rect 3384 7936 3390 7948
rect 3970 7936 3976 7948
rect 3384 7908 3976 7936
rect 3384 7896 3390 7908
rect 3970 7896 3976 7908
rect 4028 7896 4034 7948
rect 4065 7939 4123 7945
rect 4065 7905 4077 7939
rect 4111 7936 4123 7939
rect 4111 7908 4752 7936
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 3605 7871 3663 7877
rect 3605 7868 3617 7871
rect 3252 7840 3617 7868
rect 3605 7837 3617 7840
rect 3651 7868 3663 7871
rect 4246 7868 4252 7880
rect 3651 7840 4252 7868
rect 3651 7837 3663 7840
rect 3605 7831 3663 7837
rect 4246 7828 4252 7840
rect 4304 7828 4310 7880
rect 1581 7803 1639 7809
rect 1581 7769 1593 7803
rect 1627 7800 1639 7803
rect 2774 7800 2780 7812
rect 1627 7772 2780 7800
rect 1627 7769 1639 7772
rect 1581 7763 1639 7769
rect 2774 7760 2780 7772
rect 2832 7760 2838 7812
rect 1946 7732 1952 7744
rect 1907 7704 1952 7732
rect 1946 7692 1952 7704
rect 2004 7692 2010 7744
rect 2682 7692 2688 7744
rect 2740 7732 2746 7744
rect 3326 7732 3332 7744
rect 2740 7704 3332 7732
rect 2740 7692 2746 7704
rect 3326 7692 3332 7704
rect 3384 7692 3390 7744
rect 3694 7692 3700 7744
rect 3752 7732 3758 7744
rect 4249 7735 4307 7741
rect 4249 7732 4261 7735
rect 3752 7704 4261 7732
rect 3752 7692 3758 7704
rect 4249 7701 4261 7704
rect 4295 7701 4307 7735
rect 4724 7732 4752 7908
rect 4890 7896 4896 7948
rect 4948 7896 4954 7948
rect 5068 7939 5126 7945
rect 5068 7905 5080 7939
rect 5114 7936 5126 7939
rect 6362 7936 6368 7948
rect 5114 7908 6368 7936
rect 5114 7905 5126 7908
rect 5068 7899 5126 7905
rect 6362 7896 6368 7908
rect 6420 7896 6426 7948
rect 6638 7896 6644 7948
rect 6696 7936 6702 7948
rect 6733 7939 6791 7945
rect 6733 7936 6745 7939
rect 6696 7908 6745 7936
rect 6696 7896 6702 7908
rect 6733 7905 6745 7908
rect 6779 7905 6791 7939
rect 6932 7936 6960 8044
rect 7101 8041 7113 8075
rect 7147 8072 7159 8075
rect 7282 8072 7288 8084
rect 7147 8044 7288 8072
rect 7147 8041 7159 8044
rect 7101 8035 7159 8041
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 7466 8072 7472 8084
rect 7427 8044 7472 8072
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 8110 8072 8116 8084
rect 8071 8044 8116 8072
rect 8110 8032 8116 8044
rect 8168 8032 8174 8084
rect 8478 8072 8484 8084
rect 8439 8044 8484 8072
rect 8478 8032 8484 8044
rect 8536 8032 8542 8084
rect 8570 8032 8576 8084
rect 8628 8072 8634 8084
rect 9125 8075 9183 8081
rect 9125 8072 9137 8075
rect 8628 8044 9137 8072
rect 8628 8032 8634 8044
rect 9125 8041 9137 8044
rect 9171 8041 9183 8075
rect 9125 8035 9183 8041
rect 9677 8075 9735 8081
rect 9677 8041 9689 8075
rect 9723 8072 9735 8075
rect 10226 8072 10232 8084
rect 9723 8044 10232 8072
rect 9723 8041 9735 8044
rect 9677 8035 9735 8041
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 10870 8072 10876 8084
rect 10520 8044 10876 8072
rect 10520 8016 10548 8044
rect 10870 8032 10876 8044
rect 10928 8032 10934 8084
rect 11606 8032 11612 8084
rect 11664 8072 11670 8084
rect 11885 8075 11943 8081
rect 11885 8072 11897 8075
rect 11664 8044 11897 8072
rect 11664 8032 11670 8044
rect 11885 8041 11897 8044
rect 11931 8072 11943 8075
rect 12526 8072 12532 8084
rect 11931 8044 12532 8072
rect 11931 8041 11943 8044
rect 11885 8035 11943 8041
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 13173 8075 13231 8081
rect 13173 8041 13185 8075
rect 13219 8072 13231 8075
rect 13814 8072 13820 8084
rect 13219 8044 13820 8072
rect 13219 8041 13231 8044
rect 13173 8035 13231 8041
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 14182 8072 14188 8084
rect 14143 8044 14188 8072
rect 14182 8032 14188 8044
rect 14240 8032 14246 8084
rect 14366 8032 14372 8084
rect 14424 8072 14430 8084
rect 14645 8075 14703 8081
rect 14645 8072 14657 8075
rect 14424 8044 14657 8072
rect 14424 8032 14430 8044
rect 14645 8041 14657 8044
rect 14691 8041 14703 8075
rect 14645 8035 14703 8041
rect 15930 8032 15936 8084
rect 15988 8072 15994 8084
rect 17405 8075 17463 8081
rect 17405 8072 17417 8075
rect 15988 8044 17417 8072
rect 15988 8032 15994 8044
rect 17405 8041 17417 8044
rect 17451 8041 17463 8075
rect 17405 8035 17463 8041
rect 7558 8004 7564 8016
rect 7519 7976 7564 8004
rect 7558 7964 7564 7976
rect 7616 8004 7622 8016
rect 7742 8004 7748 8016
rect 7616 7976 7748 8004
rect 7616 7964 7622 7976
rect 7742 7964 7748 7976
rect 7800 7964 7806 8016
rect 7834 7964 7840 8016
rect 7892 8004 7898 8016
rect 8018 8004 8024 8016
rect 7892 7976 8024 8004
rect 7892 7964 7898 7976
rect 8018 7964 8024 7976
rect 8076 7964 8082 8016
rect 8938 8004 8944 8016
rect 8404 7976 8944 8004
rect 8404 7936 8432 7976
rect 8938 7964 8944 7976
rect 8996 7964 9002 8016
rect 10137 8007 10195 8013
rect 10137 7973 10149 8007
rect 10183 8004 10195 8007
rect 10502 8004 10508 8016
rect 10183 7976 10508 8004
rect 10183 7973 10195 7976
rect 10137 7967 10195 7973
rect 10502 7964 10508 7976
rect 10560 7964 10566 8016
rect 10772 8007 10830 8013
rect 10772 7973 10784 8007
rect 10818 8004 10830 8007
rect 10962 8004 10968 8016
rect 10818 7976 10968 8004
rect 10818 7973 10830 7976
rect 10772 7967 10830 7973
rect 10962 7964 10968 7976
rect 11020 7964 11026 8016
rect 11054 7964 11060 8016
rect 11112 8004 11118 8016
rect 13541 8007 13599 8013
rect 13541 8004 13553 8007
rect 11112 7976 13553 8004
rect 11112 7964 11118 7976
rect 13541 7973 13553 7976
rect 13587 8004 13599 8007
rect 13630 8004 13636 8016
rect 13587 7976 13636 8004
rect 13587 7973 13599 7976
rect 13541 7967 13599 7973
rect 13630 7964 13636 7976
rect 13688 7964 13694 8016
rect 14550 8004 14556 8016
rect 14511 7976 14556 8004
rect 14550 7964 14556 7976
rect 14608 8004 14614 8016
rect 14826 8004 14832 8016
rect 14608 7976 14832 8004
rect 14608 7964 14614 7976
rect 14826 7964 14832 7976
rect 14884 7964 14890 8016
rect 16206 7964 16212 8016
rect 16264 8013 16270 8016
rect 16264 8007 16328 8013
rect 16264 7973 16282 8007
rect 16316 7973 16328 8007
rect 16264 7967 16328 7973
rect 16264 7964 16270 7967
rect 6932 7908 8432 7936
rect 6733 7899 6791 7905
rect 8478 7896 8484 7948
rect 8536 7936 8542 7948
rect 9493 7939 9551 7945
rect 9493 7936 9505 7939
rect 8536 7908 9505 7936
rect 8536 7896 8542 7908
rect 9493 7905 9505 7908
rect 9539 7905 9551 7939
rect 9493 7899 9551 7905
rect 9858 7896 9864 7948
rect 9916 7936 9922 7948
rect 10045 7939 10103 7945
rect 10045 7936 10057 7939
rect 9916 7908 10057 7936
rect 9916 7896 9922 7908
rect 10045 7905 10057 7908
rect 10091 7905 10103 7939
rect 11514 7936 11520 7948
rect 10045 7899 10103 7905
rect 10336 7908 11520 7936
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7868 4859 7871
rect 4908 7868 4936 7896
rect 4847 7840 4936 7868
rect 4847 7837 4859 7840
rect 4801 7831 4859 7837
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 6917 7871 6975 7877
rect 6917 7868 6929 7871
rect 6880 7840 6929 7868
rect 6880 7828 6886 7840
rect 6917 7837 6929 7840
rect 6963 7868 6975 7871
rect 7650 7868 7656 7880
rect 6963 7840 7328 7868
rect 7611 7840 7656 7868
rect 6963 7837 6975 7840
rect 6917 7831 6975 7837
rect 5994 7800 6000 7812
rect 5736 7772 6000 7800
rect 5736 7732 5764 7772
rect 5994 7760 6000 7772
rect 6052 7760 6058 7812
rect 6181 7803 6239 7809
rect 6181 7769 6193 7803
rect 6227 7800 6239 7803
rect 6270 7800 6276 7812
rect 6227 7772 6276 7800
rect 6227 7769 6239 7772
rect 6181 7763 6239 7769
rect 6270 7760 6276 7772
rect 6328 7760 6334 7812
rect 7300 7800 7328 7840
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 8570 7868 8576 7880
rect 8531 7840 8576 7868
rect 8570 7828 8576 7840
rect 8628 7828 8634 7880
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7837 8815 7871
rect 8757 7831 8815 7837
rect 8662 7800 8668 7812
rect 7300 7772 8668 7800
rect 8662 7760 8668 7772
rect 8720 7800 8726 7812
rect 8772 7800 8800 7831
rect 8846 7828 8852 7880
rect 8904 7868 8910 7880
rect 10229 7871 10287 7877
rect 10229 7868 10241 7871
rect 8904 7840 10241 7868
rect 8904 7828 8910 7840
rect 10229 7837 10241 7840
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 8720 7772 8800 7800
rect 8720 7760 8726 7772
rect 8938 7760 8944 7812
rect 8996 7800 9002 7812
rect 10336 7800 10364 7908
rect 11514 7896 11520 7908
rect 11572 7896 11578 7948
rect 12529 7939 12587 7945
rect 12529 7905 12541 7939
rect 12575 7936 12587 7939
rect 13262 7936 13268 7948
rect 12575 7908 13268 7936
rect 12575 7905 12587 7908
rect 12529 7899 12587 7905
rect 13262 7896 13268 7908
rect 13320 7936 13326 7948
rect 16022 7936 16028 7948
rect 13320 7908 15792 7936
rect 15983 7908 16028 7936
rect 13320 7896 13326 7908
rect 10502 7868 10508 7880
rect 10463 7840 10508 7868
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 11606 7828 11612 7880
rect 11664 7868 11670 7880
rect 12621 7871 12679 7877
rect 12621 7868 12633 7871
rect 11664 7840 12633 7868
rect 11664 7828 11670 7840
rect 12621 7837 12633 7840
rect 12667 7837 12679 7871
rect 12621 7831 12679 7837
rect 12805 7871 12863 7877
rect 12805 7837 12817 7871
rect 12851 7837 12863 7871
rect 12805 7831 12863 7837
rect 8996 7772 10364 7800
rect 11992 7772 12296 7800
rect 8996 7760 9002 7772
rect 4724 7704 5764 7732
rect 9493 7735 9551 7741
rect 4249 7695 4307 7701
rect 9493 7701 9505 7735
rect 9539 7732 9551 7735
rect 11992 7732 12020 7772
rect 12158 7732 12164 7744
rect 9539 7704 12020 7732
rect 12119 7704 12164 7732
rect 9539 7701 9551 7704
rect 9493 7695 9551 7701
rect 12158 7692 12164 7704
rect 12216 7692 12222 7744
rect 12268 7732 12296 7772
rect 12342 7760 12348 7812
rect 12400 7800 12406 7812
rect 12820 7800 12848 7831
rect 13446 7828 13452 7880
rect 13504 7868 13510 7880
rect 13633 7871 13691 7877
rect 13633 7868 13645 7871
rect 13504 7840 13645 7868
rect 13504 7828 13510 7840
rect 13633 7837 13645 7840
rect 13679 7868 13691 7871
rect 13722 7868 13728 7880
rect 13679 7840 13728 7868
rect 13679 7837 13691 7840
rect 13633 7831 13691 7837
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 13817 7871 13875 7877
rect 13817 7837 13829 7871
rect 13863 7868 13875 7871
rect 14829 7871 14887 7877
rect 14829 7868 14841 7871
rect 13863 7840 14841 7868
rect 13863 7837 13875 7840
rect 13817 7831 13875 7837
rect 14829 7837 14841 7840
rect 14875 7868 14887 7871
rect 15378 7868 15384 7880
rect 14875 7840 15384 7868
rect 14875 7837 14887 7840
rect 14829 7831 14887 7837
rect 15378 7828 15384 7840
rect 15436 7828 15442 7880
rect 13906 7800 13912 7812
rect 12400 7772 13912 7800
rect 12400 7760 12406 7772
rect 13906 7760 13912 7772
rect 13964 7760 13970 7812
rect 15654 7732 15660 7744
rect 12268 7704 15660 7732
rect 15654 7692 15660 7704
rect 15712 7692 15718 7744
rect 15764 7732 15792 7908
rect 16022 7896 16028 7908
rect 16080 7896 16086 7948
rect 17862 7936 17868 7948
rect 17823 7908 17868 7936
rect 17862 7896 17868 7908
rect 17920 7896 17926 7948
rect 17494 7732 17500 7744
rect 15764 7704 17500 7732
rect 17494 7692 17500 7704
rect 17552 7692 17558 7744
rect 18046 7732 18052 7744
rect 18007 7704 18052 7732
rect 18046 7692 18052 7704
rect 18104 7692 18110 7744
rect 1104 7642 18860 7664
rect 1104 7590 3947 7642
rect 3999 7590 4011 7642
rect 4063 7590 4075 7642
rect 4127 7590 4139 7642
rect 4191 7590 9878 7642
rect 9930 7590 9942 7642
rect 9994 7590 10006 7642
rect 10058 7590 10070 7642
rect 10122 7590 15808 7642
rect 15860 7590 15872 7642
rect 15924 7590 15936 7642
rect 15988 7590 16000 7642
rect 16052 7590 18860 7642
rect 1104 7568 18860 7590
rect 2314 7488 2320 7540
rect 2372 7528 2378 7540
rect 3237 7531 3295 7537
rect 3237 7528 3249 7531
rect 2372 7500 3249 7528
rect 2372 7488 2378 7500
rect 3237 7497 3249 7500
rect 3283 7497 3295 7531
rect 4433 7531 4491 7537
rect 4433 7528 4445 7531
rect 3237 7491 3295 7497
rect 3344 7500 4445 7528
rect 2590 7420 2596 7472
rect 2648 7460 2654 7472
rect 3344 7460 3372 7500
rect 4433 7497 4445 7500
rect 4479 7497 4491 7531
rect 4433 7491 4491 7497
rect 4798 7488 4804 7540
rect 4856 7528 4862 7540
rect 6362 7528 6368 7540
rect 4856 7500 6224 7528
rect 6323 7500 6368 7528
rect 4856 7488 4862 7500
rect 4246 7460 4252 7472
rect 2648 7432 3372 7460
rect 3896 7432 4252 7460
rect 2648 7420 2654 7432
rect 3896 7401 3924 7432
rect 4246 7420 4252 7432
rect 4304 7460 4310 7472
rect 4982 7460 4988 7472
rect 4304 7432 4988 7460
rect 4304 7420 4310 7432
rect 4982 7420 4988 7432
rect 5040 7420 5046 7472
rect 6196 7460 6224 7500
rect 6362 7488 6368 7500
rect 6420 7488 6426 7540
rect 10321 7531 10379 7537
rect 8588 7500 9628 7528
rect 8588 7460 8616 7500
rect 6196 7432 8616 7460
rect 3881 7395 3939 7401
rect 3881 7361 3893 7395
rect 3927 7361 3939 7395
rect 3881 7355 3939 7361
rect 5994 7352 6000 7404
rect 6052 7392 6058 7404
rect 7558 7392 7564 7404
rect 6052 7364 7564 7392
rect 6052 7352 6058 7364
rect 7558 7352 7564 7364
rect 7616 7352 7622 7404
rect 8110 7392 8116 7404
rect 8071 7364 8116 7392
rect 8110 7352 8116 7364
rect 8168 7352 8174 7404
rect 9600 7392 9628 7500
rect 10321 7497 10333 7531
rect 10367 7528 10379 7531
rect 11330 7528 11336 7540
rect 10367 7500 11336 7528
rect 10367 7497 10379 7500
rect 10321 7491 10379 7497
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 11514 7488 11520 7540
rect 11572 7528 11578 7540
rect 14274 7528 14280 7540
rect 11572 7500 14280 7528
rect 11572 7488 11578 7500
rect 14274 7488 14280 7500
rect 14332 7488 14338 7540
rect 14642 7488 14648 7540
rect 14700 7528 14706 7540
rect 15010 7528 15016 7540
rect 14700 7500 15016 7528
rect 14700 7488 14706 7500
rect 15010 7488 15016 7500
rect 15068 7488 15074 7540
rect 15654 7528 15660 7540
rect 15488 7500 15660 7528
rect 12158 7460 12164 7472
rect 10796 7432 12164 7460
rect 10134 7392 10140 7404
rect 9600 7364 10140 7392
rect 10134 7352 10140 7364
rect 10192 7352 10198 7404
rect 10796 7401 10824 7432
rect 12158 7420 12164 7432
rect 12216 7420 12222 7472
rect 12342 7460 12348 7472
rect 12268 7432 12348 7460
rect 10781 7395 10839 7401
rect 10781 7361 10793 7395
rect 10827 7361 10839 7395
rect 10962 7392 10968 7404
rect 10923 7364 10968 7392
rect 10781 7355 10839 7361
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 11238 7352 11244 7404
rect 11296 7392 11302 7404
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 11296 7364 11897 7392
rect 11296 7352 11302 7364
rect 11885 7361 11897 7364
rect 11931 7392 11943 7395
rect 12268 7392 12296 7432
rect 12342 7420 12348 7432
rect 12400 7420 12406 7472
rect 12526 7420 12532 7472
rect 12584 7460 12590 7472
rect 14734 7460 14740 7472
rect 12584 7432 14740 7460
rect 12584 7420 12590 7432
rect 14734 7420 14740 7432
rect 14792 7420 14798 7472
rect 13078 7392 13084 7404
rect 11931 7364 12296 7392
rect 13039 7364 13084 7392
rect 11931 7361 11943 7364
rect 11885 7355 11943 7361
rect 13078 7352 13084 7364
rect 13136 7352 13142 7404
rect 13265 7395 13323 7401
rect 13265 7361 13277 7395
rect 13311 7361 13323 7395
rect 13265 7355 13323 7361
rect 1581 7327 1639 7333
rect 1581 7293 1593 7327
rect 1627 7293 1639 7327
rect 1581 7287 1639 7293
rect 1596 7188 1624 7287
rect 1670 7284 1676 7336
rect 1728 7324 1734 7336
rect 3605 7327 3663 7333
rect 1728 7296 3464 7324
rect 1728 7284 1734 7296
rect 1848 7259 1906 7265
rect 1848 7225 1860 7259
rect 1894 7256 1906 7259
rect 2866 7256 2872 7268
rect 1894 7228 2872 7256
rect 1894 7225 1906 7228
rect 1848 7219 1906 7225
rect 2866 7216 2872 7228
rect 2924 7256 2930 7268
rect 3326 7256 3332 7268
rect 2924 7228 3332 7256
rect 2924 7216 2930 7228
rect 3326 7216 3332 7228
rect 3384 7216 3390 7268
rect 2314 7188 2320 7200
rect 1596 7160 2320 7188
rect 2314 7148 2320 7160
rect 2372 7148 2378 7200
rect 2958 7188 2964 7200
rect 2919 7160 2964 7188
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 3436 7188 3464 7296
rect 3605 7293 3617 7327
rect 3651 7324 3663 7327
rect 3786 7324 3792 7336
rect 3651 7296 3792 7324
rect 3651 7293 3663 7296
rect 3605 7287 3663 7293
rect 3786 7284 3792 7296
rect 3844 7284 3850 7336
rect 4249 7327 4307 7333
rect 4249 7293 4261 7327
rect 4295 7324 4307 7327
rect 4430 7324 4436 7336
rect 4295 7296 4436 7324
rect 4295 7293 4307 7296
rect 4249 7287 4307 7293
rect 4430 7284 4436 7296
rect 4488 7284 4494 7336
rect 4890 7284 4896 7336
rect 4948 7324 4954 7336
rect 4985 7327 5043 7333
rect 4985 7324 4997 7327
rect 4948 7296 4997 7324
rect 4948 7284 4954 7296
rect 4985 7293 4997 7296
rect 5031 7293 5043 7327
rect 4985 7287 5043 7293
rect 5534 7284 5540 7336
rect 5592 7324 5598 7336
rect 6362 7324 6368 7336
rect 5592 7296 6368 7324
rect 5592 7284 5598 7296
rect 6362 7284 6368 7296
rect 6420 7284 6426 7336
rect 6825 7327 6883 7333
rect 6825 7293 6837 7327
rect 6871 7324 6883 7327
rect 8386 7324 8392 7336
rect 6871 7296 8392 7324
rect 6871 7293 6883 7296
rect 6825 7287 6883 7293
rect 8386 7284 8392 7296
rect 8444 7284 8450 7336
rect 8570 7324 8576 7336
rect 8531 7296 8576 7324
rect 8570 7284 8576 7296
rect 8628 7284 8634 7336
rect 10594 7324 10600 7336
rect 8680 7296 10600 7324
rect 5252 7259 5310 7265
rect 5252 7225 5264 7259
rect 5298 7256 5310 7259
rect 6730 7256 6736 7268
rect 5298 7228 6736 7256
rect 5298 7225 5310 7228
rect 5252 7219 5310 7225
rect 6730 7216 6736 7228
rect 6788 7216 6794 7268
rect 7837 7259 7895 7265
rect 7837 7225 7849 7259
rect 7883 7256 7895 7259
rect 8680 7256 8708 7296
rect 10594 7284 10600 7296
rect 10652 7284 10658 7336
rect 13170 7284 13176 7336
rect 13228 7324 13234 7336
rect 13280 7324 13308 7355
rect 13906 7352 13912 7404
rect 13964 7392 13970 7404
rect 14277 7395 14335 7401
rect 14277 7392 14289 7395
rect 13964 7364 14289 7392
rect 13964 7352 13970 7364
rect 14277 7361 14289 7364
rect 14323 7392 14335 7395
rect 14642 7392 14648 7404
rect 14323 7364 14648 7392
rect 14323 7361 14335 7364
rect 14277 7355 14335 7361
rect 14642 7352 14648 7364
rect 14700 7352 14706 7404
rect 15488 7392 15516 7500
rect 15654 7488 15660 7500
rect 15712 7488 15718 7540
rect 16206 7488 16212 7540
rect 16264 7528 16270 7540
rect 16850 7528 16856 7540
rect 16264 7500 16856 7528
rect 16264 7488 16270 7500
rect 16850 7488 16856 7500
rect 16908 7488 16914 7540
rect 17586 7528 17592 7540
rect 17547 7500 17592 7528
rect 17586 7488 17592 7500
rect 17644 7488 17650 7540
rect 15488 7364 15608 7392
rect 14090 7324 14096 7336
rect 13228 7296 13308 7324
rect 14051 7296 14096 7324
rect 13228 7284 13234 7296
rect 14090 7284 14096 7296
rect 14148 7284 14154 7336
rect 14550 7284 14556 7336
rect 14608 7324 14614 7336
rect 15473 7327 15531 7333
rect 15473 7324 15485 7327
rect 14608 7296 15485 7324
rect 14608 7284 14614 7296
rect 15473 7293 15485 7296
rect 15519 7293 15531 7327
rect 15580 7324 15608 7364
rect 17405 7327 17463 7333
rect 17405 7324 17417 7327
rect 15580 7296 17417 7324
rect 15473 7287 15531 7293
rect 17405 7293 17417 7296
rect 17451 7293 17463 7327
rect 17405 7287 17463 7293
rect 17494 7284 17500 7336
rect 17552 7324 17558 7336
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 17552 7296 18061 7324
rect 17552 7284 17558 7296
rect 18049 7293 18061 7296
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 8846 7265 8852 7268
rect 8840 7256 8852 7265
rect 7883 7228 8708 7256
rect 8807 7228 8852 7256
rect 7883 7225 7895 7228
rect 7837 7219 7895 7225
rect 8840 7219 8852 7228
rect 8846 7216 8852 7219
rect 8904 7216 8910 7268
rect 8938 7216 8944 7268
rect 8996 7256 9002 7268
rect 10689 7259 10747 7265
rect 8996 7228 10640 7256
rect 8996 7216 9002 7228
rect 3697 7191 3755 7197
rect 3697 7188 3709 7191
rect 3436 7160 3709 7188
rect 3697 7157 3709 7160
rect 3743 7188 3755 7191
rect 6638 7188 6644 7200
rect 3743 7160 6644 7188
rect 3743 7157 3755 7160
rect 3697 7151 3755 7157
rect 6638 7148 6644 7160
rect 6696 7148 6702 7200
rect 7009 7191 7067 7197
rect 7009 7157 7021 7191
rect 7055 7188 7067 7191
rect 7282 7188 7288 7200
rect 7055 7160 7288 7188
rect 7055 7157 7067 7160
rect 7009 7151 7067 7157
rect 7282 7148 7288 7160
rect 7340 7148 7346 7200
rect 7466 7188 7472 7200
rect 7427 7160 7472 7188
rect 7466 7148 7472 7160
rect 7524 7148 7530 7200
rect 7929 7191 7987 7197
rect 7929 7157 7941 7191
rect 7975 7188 7987 7191
rect 9674 7188 9680 7200
rect 7975 7160 9680 7188
rect 7975 7157 7987 7160
rect 7929 7151 7987 7157
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 9766 7148 9772 7200
rect 9824 7188 9830 7200
rect 9953 7191 10011 7197
rect 9953 7188 9965 7191
rect 9824 7160 9965 7188
rect 9824 7148 9830 7160
rect 9953 7157 9965 7160
rect 9999 7157 10011 7191
rect 10612 7188 10640 7228
rect 10689 7225 10701 7259
rect 10735 7256 10747 7259
rect 10735 7228 13676 7256
rect 10735 7225 10747 7228
rect 10689 7219 10747 7225
rect 10778 7188 10784 7200
rect 10612 7160 10784 7188
rect 9953 7151 10011 7157
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 11330 7188 11336 7200
rect 11291 7160 11336 7188
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 11422 7148 11428 7200
rect 11480 7188 11486 7200
rect 11701 7191 11759 7197
rect 11701 7188 11713 7191
rect 11480 7160 11713 7188
rect 11480 7148 11486 7160
rect 11701 7157 11713 7160
rect 11747 7157 11759 7191
rect 11701 7151 11759 7157
rect 11790 7148 11796 7200
rect 11848 7188 11854 7200
rect 11848 7160 11893 7188
rect 11848 7148 11854 7160
rect 11974 7148 11980 7200
rect 12032 7188 12038 7200
rect 12621 7191 12679 7197
rect 12621 7188 12633 7191
rect 12032 7160 12633 7188
rect 12032 7148 12038 7160
rect 12621 7157 12633 7160
rect 12667 7157 12679 7191
rect 12621 7151 12679 7157
rect 12989 7191 13047 7197
rect 12989 7157 13001 7191
rect 13035 7188 13047 7191
rect 13262 7188 13268 7200
rect 13035 7160 13268 7188
rect 13035 7157 13047 7160
rect 12989 7151 13047 7157
rect 13262 7148 13268 7160
rect 13320 7188 13326 7200
rect 13446 7188 13452 7200
rect 13320 7160 13452 7188
rect 13320 7148 13326 7160
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 13648 7197 13676 7228
rect 15378 7216 15384 7268
rect 15436 7256 15442 7268
rect 15718 7259 15776 7265
rect 15718 7256 15730 7259
rect 15436 7228 15730 7256
rect 15436 7216 15442 7228
rect 15718 7225 15730 7228
rect 15764 7225 15776 7259
rect 15718 7219 15776 7225
rect 13633 7191 13691 7197
rect 13633 7157 13645 7191
rect 13679 7157 13691 7191
rect 13633 7151 13691 7157
rect 13814 7148 13820 7200
rect 13872 7188 13878 7200
rect 14001 7191 14059 7197
rect 14001 7188 14013 7191
rect 13872 7160 14013 7188
rect 13872 7148 13878 7160
rect 14001 7157 14013 7160
rect 14047 7157 14059 7191
rect 14734 7188 14740 7200
rect 14695 7160 14740 7188
rect 14001 7151 14059 7157
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 15194 7148 15200 7200
rect 15252 7188 15258 7200
rect 16206 7188 16212 7200
rect 15252 7160 16212 7188
rect 15252 7148 15258 7160
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 18230 7188 18236 7200
rect 18191 7160 18236 7188
rect 18230 7148 18236 7160
rect 18288 7148 18294 7200
rect 1104 7098 18860 7120
rect 1104 7046 6912 7098
rect 6964 7046 6976 7098
rect 7028 7046 7040 7098
rect 7092 7046 7104 7098
rect 7156 7046 12843 7098
rect 12895 7046 12907 7098
rect 12959 7046 12971 7098
rect 13023 7046 13035 7098
rect 13087 7046 18860 7098
rect 1104 7024 18860 7046
rect 2866 6944 2872 6996
rect 2924 6984 2930 6996
rect 4065 6987 4123 6993
rect 4065 6984 4077 6987
rect 2924 6956 4077 6984
rect 2924 6944 2930 6956
rect 4065 6953 4077 6956
rect 4111 6953 4123 6987
rect 4065 6947 4123 6953
rect 5813 6987 5871 6993
rect 5813 6953 5825 6987
rect 5859 6984 5871 6987
rect 6365 6987 6423 6993
rect 6365 6984 6377 6987
rect 5859 6956 6377 6984
rect 5859 6953 5871 6956
rect 5813 6947 5871 6953
rect 6365 6953 6377 6956
rect 6411 6953 6423 6987
rect 6365 6947 6423 6953
rect 6733 6987 6791 6993
rect 6733 6953 6745 6987
rect 6779 6984 6791 6987
rect 10226 6984 10232 6996
rect 6779 6956 10232 6984
rect 6779 6953 6791 6956
rect 6733 6947 6791 6953
rect 10226 6944 10232 6956
rect 10284 6944 10290 6996
rect 11609 6987 11667 6993
rect 11609 6953 11621 6987
rect 11655 6984 11667 6987
rect 11790 6984 11796 6996
rect 11655 6956 11796 6984
rect 11655 6953 11667 6956
rect 11609 6947 11667 6953
rect 11790 6944 11796 6956
rect 11848 6944 11854 6996
rect 14001 6987 14059 6993
rect 14001 6984 14013 6987
rect 11900 6956 14013 6984
rect 5721 6919 5779 6925
rect 5721 6885 5733 6919
rect 5767 6916 5779 6919
rect 7466 6916 7472 6928
rect 5767 6888 7472 6916
rect 5767 6885 5779 6888
rect 5721 6879 5779 6885
rect 7466 6876 7472 6888
rect 7524 6876 7530 6928
rect 8570 6916 8576 6928
rect 7576 6888 8576 6916
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6848 1731 6851
rect 1854 6848 1860 6860
rect 1719 6820 1860 6848
rect 1719 6817 1731 6820
rect 1673 6811 1731 6817
rect 1854 6808 1860 6820
rect 1912 6808 1918 6860
rect 2584 6851 2642 6857
rect 2584 6817 2596 6851
rect 2630 6848 2642 6851
rect 2958 6848 2964 6860
rect 2630 6820 2964 6848
rect 2630 6817 2642 6820
rect 2584 6811 2642 6817
rect 2958 6808 2964 6820
rect 3016 6808 3022 6860
rect 3786 6808 3792 6860
rect 3844 6808 3850 6860
rect 4246 6808 4252 6860
rect 4304 6848 4310 6860
rect 4433 6851 4491 6857
rect 4433 6848 4445 6851
rect 4304 6820 4445 6848
rect 4304 6808 4310 6820
rect 4433 6817 4445 6820
rect 4479 6817 4491 6851
rect 4433 6811 4491 6817
rect 5261 6851 5319 6857
rect 5261 6817 5273 6851
rect 5307 6848 5319 6851
rect 5626 6848 5632 6860
rect 5307 6820 5632 6848
rect 5307 6817 5319 6820
rect 5261 6811 5319 6817
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 6825 6851 6883 6857
rect 6825 6817 6837 6851
rect 6871 6848 6883 6851
rect 7282 6848 7288 6860
rect 6871 6820 7288 6848
rect 6871 6817 6883 6820
rect 6825 6811 6883 6817
rect 7282 6808 7288 6820
rect 7340 6808 7346 6860
rect 7377 6851 7435 6857
rect 7377 6817 7389 6851
rect 7423 6848 7435 6851
rect 7576 6848 7604 6888
rect 8570 6876 8576 6888
rect 8628 6876 8634 6928
rect 8846 6876 8852 6928
rect 8904 6916 8910 6928
rect 9306 6916 9312 6928
rect 8904 6888 9312 6916
rect 8904 6876 8910 6888
rect 9306 6876 9312 6888
rect 9364 6876 9370 6928
rect 10502 6916 10508 6928
rect 9876 6888 10508 6916
rect 7423 6820 7604 6848
rect 7644 6851 7702 6857
rect 7423 6817 7435 6820
rect 7377 6811 7435 6817
rect 7644 6817 7656 6851
rect 7690 6848 7702 6851
rect 8202 6848 8208 6860
rect 7690 6820 8208 6848
rect 7690 6817 7702 6820
rect 7644 6811 7702 6817
rect 2314 6780 2320 6792
rect 2275 6752 2320 6780
rect 2314 6740 2320 6752
rect 2372 6740 2378 6792
rect 3804 6712 3832 6808
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6780 4583 6783
rect 4614 6780 4620 6792
rect 4571 6752 4620 6780
rect 4571 6749 4583 6752
rect 4525 6743 4583 6749
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6780 4767 6783
rect 4982 6780 4988 6792
rect 4755 6752 4988 6780
rect 4755 6749 4767 6752
rect 4709 6743 4767 6749
rect 4982 6740 4988 6752
rect 5040 6740 5046 6792
rect 5997 6783 6055 6789
rect 5997 6749 6009 6783
rect 6043 6780 6055 6783
rect 6638 6780 6644 6792
rect 6043 6752 6644 6780
rect 6043 6749 6055 6752
rect 5997 6743 6055 6749
rect 6638 6740 6644 6752
rect 6696 6740 6702 6792
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6749 7067 6783
rect 7009 6743 7067 6749
rect 3804 6684 6960 6712
rect 6932 6656 6960 6684
rect 1857 6647 1915 6653
rect 1857 6613 1869 6647
rect 1903 6644 1915 6647
rect 3510 6644 3516 6656
rect 1903 6616 3516 6644
rect 1903 6613 1915 6616
rect 1857 6607 1915 6613
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 3694 6644 3700 6656
rect 3655 6616 3700 6644
rect 3694 6604 3700 6616
rect 3752 6604 3758 6656
rect 5074 6644 5080 6656
rect 5035 6616 5080 6644
rect 5074 6604 5080 6616
rect 5132 6604 5138 6656
rect 5353 6647 5411 6653
rect 5353 6613 5365 6647
rect 5399 6644 5411 6647
rect 6730 6644 6736 6656
rect 5399 6616 6736 6644
rect 5399 6613 5411 6616
rect 5353 6607 5411 6613
rect 6730 6604 6736 6616
rect 6788 6604 6794 6656
rect 6914 6604 6920 6656
rect 6972 6604 6978 6656
rect 7024 6644 7052 6743
rect 7190 6740 7196 6792
rect 7248 6780 7254 6792
rect 7392 6780 7420 6811
rect 8202 6808 8208 6820
rect 8260 6808 8266 6860
rect 9876 6857 9904 6888
rect 10502 6876 10508 6888
rect 10560 6876 10566 6928
rect 11238 6916 11244 6928
rect 10888 6888 11244 6916
rect 9861 6851 9919 6857
rect 9861 6817 9873 6851
rect 9907 6817 9919 6851
rect 9861 6811 9919 6817
rect 10128 6851 10186 6857
rect 10128 6817 10140 6851
rect 10174 6848 10186 6851
rect 10888 6848 10916 6888
rect 11238 6876 11244 6888
rect 11296 6876 11302 6928
rect 11330 6876 11336 6928
rect 11388 6916 11394 6928
rect 11900 6916 11928 6956
rect 14001 6953 14013 6956
rect 14047 6953 14059 6987
rect 14826 6984 14832 6996
rect 14001 6947 14059 6953
rect 14752 6956 14832 6984
rect 11388 6888 11928 6916
rect 11977 6919 12035 6925
rect 11388 6876 11394 6888
rect 11977 6885 11989 6919
rect 12023 6916 12035 6919
rect 12250 6916 12256 6928
rect 12023 6888 12256 6916
rect 12023 6885 12035 6888
rect 11977 6879 12035 6885
rect 12250 6876 12256 6888
rect 12308 6876 12314 6928
rect 12529 6919 12587 6925
rect 12529 6885 12541 6919
rect 12575 6916 12587 6919
rect 12989 6919 13047 6925
rect 12989 6916 13001 6919
rect 12575 6888 13001 6916
rect 12575 6885 12587 6888
rect 12529 6879 12587 6885
rect 12989 6885 13001 6888
rect 13035 6885 13047 6919
rect 12989 6879 13047 6885
rect 13081 6919 13139 6925
rect 13081 6885 13093 6919
rect 13127 6916 13139 6919
rect 13127 6888 14320 6916
rect 13127 6885 13139 6888
rect 13081 6879 13139 6885
rect 10174 6820 10916 6848
rect 10174 6817 10186 6820
rect 10128 6811 10186 6817
rect 10962 6808 10968 6860
rect 11020 6848 11026 6860
rect 14292 6848 14320 6888
rect 14366 6848 14372 6860
rect 11020 6820 14228 6848
rect 14292 6820 14372 6848
rect 11020 6808 11026 6820
rect 7248 6752 7420 6780
rect 7248 6740 7254 6752
rect 8386 6740 8392 6792
rect 8444 6780 8450 6792
rect 9033 6783 9091 6789
rect 9033 6780 9045 6783
rect 8444 6752 9045 6780
rect 8444 6740 8450 6752
rect 9033 6749 9045 6752
rect 9079 6749 9091 6783
rect 9033 6743 9091 6749
rect 8662 6672 8668 6724
rect 8720 6712 8726 6724
rect 8757 6715 8815 6721
rect 8757 6712 8769 6715
rect 8720 6684 8769 6712
rect 8720 6672 8726 6684
rect 8757 6681 8769 6684
rect 8803 6681 8815 6715
rect 8757 6675 8815 6681
rect 11241 6715 11299 6721
rect 11241 6681 11253 6715
rect 11287 6712 11299 6715
rect 11348 6712 11376 6820
rect 11882 6740 11888 6792
rect 11940 6780 11946 6792
rect 12069 6783 12127 6789
rect 12069 6780 12081 6783
rect 11940 6752 12081 6780
rect 11940 6740 11946 6752
rect 12069 6749 12081 6752
rect 12115 6749 12127 6783
rect 12069 6743 12127 6749
rect 12253 6783 12311 6789
rect 12253 6749 12265 6783
rect 12299 6749 12311 6783
rect 12253 6743 12311 6749
rect 11287 6684 11376 6712
rect 12268 6712 12296 6743
rect 12342 6740 12348 6792
rect 12400 6780 12406 6792
rect 12529 6783 12587 6789
rect 12529 6780 12541 6783
rect 12400 6752 12541 6780
rect 12400 6740 12406 6752
rect 12529 6749 12541 6752
rect 12575 6749 12587 6783
rect 13170 6780 13176 6792
rect 12529 6743 12587 6749
rect 12636 6752 13176 6780
rect 12636 6712 12664 6752
rect 13170 6740 13176 6752
rect 13228 6740 13234 6792
rect 14090 6780 14096 6792
rect 14051 6752 14096 6780
rect 14090 6740 14096 6752
rect 14148 6740 14154 6792
rect 14200 6789 14228 6820
rect 14366 6808 14372 6820
rect 14424 6848 14430 6860
rect 14752 6848 14780 6956
rect 14826 6944 14832 6956
rect 14884 6944 14890 6996
rect 15654 6984 15660 6996
rect 15615 6956 15660 6984
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 16298 6984 16304 6996
rect 16259 6956 16304 6984
rect 16298 6944 16304 6956
rect 16356 6944 16362 6996
rect 14918 6876 14924 6928
rect 14976 6916 14982 6928
rect 16669 6919 16727 6925
rect 16669 6916 16681 6919
rect 14976 6888 16681 6916
rect 14976 6876 14982 6888
rect 16669 6885 16681 6888
rect 16715 6885 16727 6919
rect 16669 6879 16727 6885
rect 14424 6820 14780 6848
rect 14424 6808 14430 6820
rect 14826 6808 14832 6860
rect 14884 6848 14890 6860
rect 14884 6820 14929 6848
rect 14884 6808 14890 6820
rect 15378 6808 15384 6860
rect 15436 6848 15442 6860
rect 15436 6820 15884 6848
rect 15436 6808 15442 6820
rect 14185 6783 14243 6789
rect 14185 6749 14197 6783
rect 14231 6749 14243 6783
rect 14185 6743 14243 6749
rect 15010 6740 15016 6792
rect 15068 6780 15074 6792
rect 15856 6789 15884 6820
rect 16298 6808 16304 6860
rect 16356 6848 16362 6860
rect 17865 6851 17923 6857
rect 17865 6848 17877 6851
rect 16356 6820 17877 6848
rect 16356 6808 16362 6820
rect 17865 6817 17877 6820
rect 17911 6817 17923 6851
rect 17865 6811 17923 6817
rect 15749 6783 15807 6789
rect 15749 6780 15761 6783
rect 15068 6752 15761 6780
rect 15068 6740 15074 6752
rect 15749 6749 15761 6752
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 16761 6783 16819 6789
rect 16761 6749 16773 6783
rect 16807 6749 16819 6783
rect 16761 6743 16819 6749
rect 12268 6684 12664 6712
rect 11287 6681 11299 6684
rect 11241 6675 11299 6681
rect 13446 6672 13452 6724
rect 13504 6712 13510 6724
rect 13633 6715 13691 6721
rect 13633 6712 13645 6715
rect 13504 6684 13645 6712
rect 13504 6672 13510 6684
rect 13633 6681 13645 6684
rect 13679 6681 13691 6715
rect 13633 6675 13691 6681
rect 15289 6715 15347 6721
rect 15289 6681 15301 6715
rect 15335 6712 15347 6715
rect 16776 6712 16804 6743
rect 16850 6740 16856 6792
rect 16908 6780 16914 6792
rect 16908 6752 16953 6780
rect 16908 6740 16914 6752
rect 15335 6684 16804 6712
rect 15335 6681 15347 6684
rect 15289 6675 15347 6681
rect 8110 6644 8116 6656
rect 7024 6616 8116 6644
rect 8110 6604 8116 6616
rect 8168 6604 8174 6656
rect 8478 6604 8484 6656
rect 8536 6644 8542 6656
rect 9306 6644 9312 6656
rect 8536 6616 9312 6644
rect 8536 6604 8542 6616
rect 9306 6604 9312 6616
rect 9364 6644 9370 6656
rect 12250 6644 12256 6656
rect 9364 6616 12256 6644
rect 9364 6604 9370 6616
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 12621 6647 12679 6653
rect 12621 6613 12633 6647
rect 12667 6644 12679 6647
rect 12710 6644 12716 6656
rect 12667 6616 12716 6644
rect 12667 6613 12679 6616
rect 12621 6607 12679 6613
rect 12710 6604 12716 6616
rect 12768 6604 12774 6656
rect 13906 6604 13912 6656
rect 13964 6644 13970 6656
rect 14550 6644 14556 6656
rect 13964 6616 14556 6644
rect 13964 6604 13970 6616
rect 14550 6604 14556 6616
rect 14608 6644 14614 6656
rect 14645 6647 14703 6653
rect 14645 6644 14657 6647
rect 14608 6616 14657 6644
rect 14608 6604 14614 6616
rect 14645 6613 14657 6616
rect 14691 6613 14703 6647
rect 18046 6644 18052 6656
rect 18007 6616 18052 6644
rect 14645 6607 14703 6613
rect 18046 6604 18052 6616
rect 18104 6604 18110 6656
rect 1104 6554 18860 6576
rect 1104 6502 3947 6554
rect 3999 6502 4011 6554
rect 4063 6502 4075 6554
rect 4127 6502 4139 6554
rect 4191 6502 9878 6554
rect 9930 6502 9942 6554
rect 9994 6502 10006 6554
rect 10058 6502 10070 6554
rect 10122 6502 15808 6554
rect 15860 6502 15872 6554
rect 15924 6502 15936 6554
rect 15988 6502 16000 6554
rect 16052 6502 18860 6554
rect 1104 6480 18860 6502
rect 2777 6443 2835 6449
rect 2777 6409 2789 6443
rect 2823 6440 2835 6443
rect 4246 6440 4252 6452
rect 2823 6412 4252 6440
rect 2823 6409 2835 6412
rect 2777 6403 2835 6409
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 5537 6443 5595 6449
rect 5537 6409 5549 6443
rect 5583 6440 5595 6443
rect 7466 6440 7472 6452
rect 5583 6412 7472 6440
rect 5583 6409 5595 6412
rect 5537 6403 5595 6409
rect 7466 6400 7472 6412
rect 7524 6400 7530 6452
rect 7558 6400 7564 6452
rect 7616 6440 7622 6452
rect 8202 6440 8208 6452
rect 7616 6412 8064 6440
rect 8163 6412 8208 6440
rect 7616 6400 7622 6412
rect 4890 6332 4896 6384
rect 4948 6372 4954 6384
rect 6822 6372 6828 6384
rect 4948 6344 6828 6372
rect 4948 6332 4954 6344
rect 6822 6332 6828 6344
rect 6880 6332 6886 6384
rect 8036 6372 8064 6412
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 11882 6440 11888 6452
rect 9048 6412 11284 6440
rect 9048 6372 9076 6412
rect 8036 6344 9076 6372
rect 11256 6372 11284 6412
rect 11440 6412 11888 6440
rect 11440 6372 11468 6412
rect 11882 6400 11888 6412
rect 11940 6440 11946 6452
rect 12434 6440 12440 6452
rect 11940 6412 12440 6440
rect 11940 6400 11946 6412
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 13446 6400 13452 6452
rect 13504 6440 13510 6452
rect 14642 6440 14648 6452
rect 13504 6412 14504 6440
rect 14603 6412 14648 6440
rect 13504 6400 13510 6412
rect 11256 6344 11468 6372
rect 11514 6332 11520 6384
rect 11572 6372 11578 6384
rect 12986 6372 12992 6384
rect 11572 6344 12992 6372
rect 11572 6332 11578 6344
rect 12986 6332 12992 6344
rect 13044 6332 13050 6384
rect 13170 6332 13176 6384
rect 13228 6372 13234 6384
rect 14476 6372 14504 6412
rect 14642 6400 14648 6412
rect 14700 6400 14706 6452
rect 14918 6440 14924 6452
rect 14879 6412 14924 6440
rect 14918 6400 14924 6412
rect 14976 6400 14982 6452
rect 15304 6412 16436 6440
rect 15304 6372 15332 6412
rect 13228 6344 13308 6372
rect 14476 6344 15332 6372
rect 13228 6332 13234 6344
rect 1946 6264 1952 6316
rect 2004 6304 2010 6316
rect 2317 6307 2375 6313
rect 2317 6304 2329 6307
rect 2004 6276 2329 6304
rect 2004 6264 2010 6276
rect 2317 6273 2329 6276
rect 2363 6273 2375 6307
rect 2317 6267 2375 6273
rect 2501 6307 2559 6313
rect 2501 6273 2513 6307
rect 2547 6304 2559 6307
rect 2958 6304 2964 6316
rect 2547 6276 2964 6304
rect 2547 6273 2559 6276
rect 2501 6267 2559 6273
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 3326 6264 3332 6316
rect 3384 6304 3390 6316
rect 3421 6307 3479 6313
rect 3421 6304 3433 6307
rect 3384 6276 3433 6304
rect 3384 6264 3390 6276
rect 3421 6273 3433 6276
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 3694 6264 3700 6316
rect 3752 6304 3758 6316
rect 3752 6276 4016 6304
rect 3752 6264 3758 6276
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 2777 6239 2835 6245
rect 2777 6236 2789 6239
rect 1443 6208 2789 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 2777 6205 2789 6208
rect 2823 6205 2835 6239
rect 2777 6199 2835 6205
rect 2866 6196 2872 6248
rect 2924 6236 2930 6248
rect 3237 6239 3295 6245
rect 3237 6236 3249 6239
rect 2924 6208 3249 6236
rect 2924 6196 2930 6208
rect 3237 6205 3249 6208
rect 3283 6205 3295 6239
rect 3237 6199 3295 6205
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6205 3939 6239
rect 3988 6236 4016 6276
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 6089 6307 6147 6313
rect 6089 6304 6101 6307
rect 5592 6276 6101 6304
rect 5592 6264 5598 6276
rect 6089 6273 6101 6276
rect 6135 6273 6147 6307
rect 6089 6267 6147 6273
rect 6638 6264 6644 6316
rect 6696 6304 6702 6316
rect 6696 6276 6960 6304
rect 6696 6264 6702 6276
rect 4154 6245 4160 6248
rect 4137 6239 4160 6245
rect 4137 6236 4149 6239
rect 3988 6208 4149 6236
rect 3881 6199 3939 6205
rect 4137 6205 4149 6208
rect 4212 6236 4218 6248
rect 4212 6208 4285 6236
rect 4137 6199 4160 6205
rect 2314 6128 2320 6180
rect 2372 6168 2378 6180
rect 3329 6171 3387 6177
rect 2372 6140 3004 6168
rect 2372 6128 2378 6140
rect 1394 6060 1400 6112
rect 1452 6100 1458 6112
rect 1857 6103 1915 6109
rect 1857 6100 1869 6103
rect 1452 6072 1869 6100
rect 1452 6060 1458 6072
rect 1857 6069 1869 6072
rect 1903 6069 1915 6103
rect 1857 6063 1915 6069
rect 2225 6103 2283 6109
rect 2225 6069 2237 6103
rect 2271 6100 2283 6103
rect 2869 6103 2927 6109
rect 2869 6100 2881 6103
rect 2271 6072 2881 6100
rect 2271 6069 2283 6072
rect 2225 6063 2283 6069
rect 2869 6069 2881 6072
rect 2915 6069 2927 6103
rect 2976 6100 3004 6140
rect 3329 6137 3341 6171
rect 3375 6168 3387 6171
rect 3418 6168 3424 6180
rect 3375 6140 3424 6168
rect 3375 6137 3387 6140
rect 3329 6131 3387 6137
rect 3418 6128 3424 6140
rect 3476 6128 3482 6180
rect 3896 6100 3924 6199
rect 4154 6196 4160 6199
rect 4212 6196 4218 6208
rect 5350 6196 5356 6248
rect 5408 6236 5414 6248
rect 5997 6239 6055 6245
rect 5997 6236 6009 6239
rect 5408 6208 6009 6236
rect 5408 6196 5414 6208
rect 5997 6205 6009 6208
rect 6043 6205 6055 6239
rect 5997 6199 6055 6205
rect 6825 6239 6883 6245
rect 6825 6205 6837 6239
rect 6871 6205 6883 6239
rect 6932 6236 6960 6276
rect 8312 6276 8616 6304
rect 7081 6239 7139 6245
rect 7081 6236 7093 6239
rect 6932 6208 7093 6236
rect 6825 6199 6883 6205
rect 7081 6205 7093 6208
rect 7127 6205 7139 6239
rect 7081 6199 7139 6205
rect 3970 6128 3976 6180
rect 4028 6168 4034 6180
rect 6840 6168 6868 6199
rect 7650 6196 7656 6248
rect 7708 6236 7714 6248
rect 8312 6236 8340 6276
rect 8478 6236 8484 6248
rect 7708 6208 8340 6236
rect 8439 6208 8484 6236
rect 7708 6196 7714 6208
rect 8478 6196 8484 6208
rect 8536 6196 8542 6248
rect 8588 6236 8616 6276
rect 8662 6264 8668 6316
rect 8720 6304 8726 6316
rect 9033 6307 9091 6313
rect 9033 6304 9045 6307
rect 8720 6276 9045 6304
rect 8720 6264 8726 6276
rect 9033 6273 9045 6276
rect 9079 6273 9091 6307
rect 9033 6267 9091 6273
rect 11238 6264 11244 6316
rect 11296 6304 11302 6316
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 11296 6276 11897 6304
rect 11296 6264 11302 6276
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 12710 6304 12716 6316
rect 11885 6267 11943 6273
rect 12084 6276 12716 6304
rect 10410 6236 10416 6248
rect 8588 6208 10416 6236
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 11793 6239 11851 6245
rect 11793 6205 11805 6239
rect 11839 6236 11851 6239
rect 12084 6236 12112 6276
rect 12710 6264 12716 6276
rect 12768 6264 12774 6316
rect 13280 6304 13308 6344
rect 15378 6332 15384 6384
rect 15436 6372 15442 6384
rect 16408 6372 16436 6412
rect 17218 6372 17224 6384
rect 15436 6344 15516 6372
rect 15436 6332 15442 6344
rect 15488 6313 15516 6344
rect 16408 6344 17224 6372
rect 16408 6313 16436 6344
rect 17218 6332 17224 6344
rect 17276 6332 17282 6384
rect 15473 6307 15531 6313
rect 13280 6276 13400 6304
rect 13372 6248 13400 6276
rect 15473 6273 15485 6307
rect 15519 6273 15531 6307
rect 15473 6267 15531 6273
rect 16393 6307 16451 6313
rect 16393 6273 16405 6307
rect 16439 6273 16451 6307
rect 16393 6267 16451 6273
rect 16485 6307 16543 6313
rect 16485 6273 16497 6307
rect 16531 6273 16543 6307
rect 16485 6267 16543 6273
rect 11839 6208 12112 6236
rect 11839 6205 11851 6208
rect 11793 6199 11851 6205
rect 12618 6196 12624 6248
rect 12676 6236 12682 6248
rect 13173 6239 13231 6245
rect 13173 6236 13185 6239
rect 12676 6208 13185 6236
rect 12676 6196 12682 6208
rect 13173 6205 13185 6208
rect 13219 6205 13231 6239
rect 13173 6199 13231 6205
rect 13265 6239 13323 6245
rect 13265 6205 13277 6239
rect 13311 6205 13323 6239
rect 13265 6199 13323 6205
rect 7190 6168 7196 6180
rect 4028 6140 6132 6168
rect 6840 6140 7196 6168
rect 4028 6128 4034 6140
rect 4982 6100 4988 6112
rect 2976 6072 4988 6100
rect 2869 6063 2927 6069
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 5258 6100 5264 6112
rect 5219 6072 5264 6100
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 5902 6100 5908 6112
rect 5863 6072 5908 6100
rect 5902 6060 5908 6072
rect 5960 6060 5966 6112
rect 6104 6100 6132 6140
rect 7190 6128 7196 6140
rect 7248 6128 7254 6180
rect 9300 6171 9358 6177
rect 9300 6137 9312 6171
rect 9346 6168 9358 6171
rect 9766 6168 9772 6180
rect 9346 6140 9772 6168
rect 9346 6137 9358 6140
rect 9300 6131 9358 6137
rect 9766 6128 9772 6140
rect 9824 6168 9830 6180
rect 11606 6168 11612 6180
rect 9824 6140 11612 6168
rect 9824 6128 9830 6140
rect 11606 6128 11612 6140
rect 11664 6128 11670 6180
rect 11701 6171 11759 6177
rect 11701 6137 11713 6171
rect 11747 6168 11759 6171
rect 11974 6168 11980 6180
rect 11747 6140 11980 6168
rect 11747 6137 11759 6140
rect 11701 6131 11759 6137
rect 11974 6128 11980 6140
rect 12032 6128 12038 6180
rect 12529 6171 12587 6177
rect 12529 6137 12541 6171
rect 12575 6168 12587 6171
rect 12894 6168 12900 6180
rect 12575 6140 12900 6168
rect 12575 6137 12587 6140
rect 12529 6131 12587 6137
rect 12894 6128 12900 6140
rect 12952 6128 12958 6180
rect 13280 6168 13308 6199
rect 13354 6196 13360 6248
rect 13412 6236 13418 6248
rect 13521 6239 13579 6245
rect 13521 6236 13533 6239
rect 13412 6208 13533 6236
rect 13412 6196 13418 6208
rect 13521 6205 13533 6208
rect 13567 6205 13579 6239
rect 13521 6199 13579 6205
rect 14734 6196 14740 6248
rect 14792 6236 14798 6248
rect 15289 6239 15347 6245
rect 15289 6236 15301 6239
rect 14792 6208 15301 6236
rect 14792 6196 14798 6208
rect 15289 6205 15301 6208
rect 15335 6205 15347 6239
rect 15289 6199 15347 6205
rect 15381 6239 15439 6245
rect 15381 6205 15393 6239
rect 15427 6236 15439 6239
rect 15562 6236 15568 6248
rect 15427 6208 15568 6236
rect 15427 6205 15439 6208
rect 15381 6199 15439 6205
rect 15562 6196 15568 6208
rect 15620 6196 15626 6248
rect 13906 6168 13912 6180
rect 13280 6140 13912 6168
rect 13906 6128 13912 6140
rect 13964 6128 13970 6180
rect 16500 6168 16528 6267
rect 17034 6196 17040 6248
rect 17092 6236 17098 6248
rect 17405 6239 17463 6245
rect 17405 6236 17417 6239
rect 17092 6208 17417 6236
rect 17092 6196 17098 6208
rect 17405 6205 17417 6208
rect 17451 6205 17463 6239
rect 17405 6199 17463 6205
rect 17954 6196 17960 6248
rect 18012 6236 18018 6248
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 18012 6208 18061 6236
rect 18012 6196 18018 6208
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 14476 6140 16528 6168
rect 8665 6103 8723 6109
rect 8665 6100 8677 6103
rect 6104 6072 8677 6100
rect 8665 6069 8677 6072
rect 8711 6069 8723 6103
rect 10410 6100 10416 6112
rect 10371 6072 10416 6100
rect 8665 6063 8723 6069
rect 10410 6060 10416 6072
rect 10468 6060 10474 6112
rect 10689 6103 10747 6109
rect 10689 6069 10701 6103
rect 10735 6100 10747 6103
rect 11054 6100 11060 6112
rect 10735 6072 11060 6100
rect 10735 6069 10747 6072
rect 10689 6063 10747 6069
rect 11054 6060 11060 6072
rect 11112 6060 11118 6112
rect 11330 6100 11336 6112
rect 11291 6072 11336 6100
rect 11330 6060 11336 6072
rect 11388 6060 11394 6112
rect 12158 6060 12164 6112
rect 12216 6100 12222 6112
rect 14476 6100 14504 6140
rect 12216 6072 14504 6100
rect 12216 6060 12222 6072
rect 14826 6060 14832 6112
rect 14884 6100 14890 6112
rect 15933 6103 15991 6109
rect 15933 6100 15945 6103
rect 14884 6072 15945 6100
rect 14884 6060 14890 6072
rect 15933 6069 15945 6072
rect 15979 6069 15991 6103
rect 15933 6063 15991 6069
rect 16301 6103 16359 6109
rect 16301 6069 16313 6103
rect 16347 6100 16359 6103
rect 16390 6100 16396 6112
rect 16347 6072 16396 6100
rect 16347 6069 16359 6072
rect 16301 6063 16359 6069
rect 16390 6060 16396 6072
rect 16448 6060 16454 6112
rect 17586 6100 17592 6112
rect 17547 6072 17592 6100
rect 17586 6060 17592 6072
rect 17644 6060 17650 6112
rect 17862 6060 17868 6112
rect 17920 6100 17926 6112
rect 18233 6103 18291 6109
rect 18233 6100 18245 6103
rect 17920 6072 18245 6100
rect 17920 6060 17926 6072
rect 18233 6069 18245 6072
rect 18279 6069 18291 6103
rect 18233 6063 18291 6069
rect 1104 6010 18860 6032
rect 1104 5958 6912 6010
rect 6964 5958 6976 6010
rect 7028 5958 7040 6010
rect 7092 5958 7104 6010
rect 7156 5958 12843 6010
rect 12895 5958 12907 6010
rect 12959 5958 12971 6010
rect 13023 5958 13035 6010
rect 13087 5958 18860 6010
rect 1104 5936 18860 5958
rect 4338 5856 4344 5908
rect 4396 5896 4402 5908
rect 4525 5899 4583 5905
rect 4525 5896 4537 5899
rect 4396 5868 4537 5896
rect 4396 5856 4402 5868
rect 4525 5865 4537 5868
rect 4571 5865 4583 5899
rect 4525 5859 4583 5865
rect 6638 5856 6644 5908
rect 6696 5896 6702 5908
rect 6825 5899 6883 5905
rect 6825 5896 6837 5899
rect 6696 5868 6837 5896
rect 6696 5856 6702 5868
rect 6825 5865 6837 5868
rect 6871 5865 6883 5899
rect 6825 5859 6883 5865
rect 6917 5899 6975 5905
rect 6917 5865 6929 5899
rect 6963 5896 6975 5899
rect 8110 5896 8116 5908
rect 6963 5868 8116 5896
rect 6963 5865 6975 5868
rect 6917 5859 6975 5865
rect 8110 5856 8116 5868
rect 8168 5896 8174 5908
rect 9309 5899 9367 5905
rect 9309 5896 9321 5899
rect 8168 5868 9321 5896
rect 8168 5856 8174 5868
rect 9309 5865 9321 5868
rect 9355 5865 9367 5899
rect 9309 5859 9367 5865
rect 11606 5856 11612 5908
rect 11664 5896 11670 5908
rect 12989 5899 13047 5905
rect 12989 5896 13001 5899
rect 11664 5868 13001 5896
rect 11664 5856 11670 5868
rect 12989 5865 13001 5868
rect 13035 5865 13047 5899
rect 12989 5859 13047 5865
rect 13633 5899 13691 5905
rect 13633 5865 13645 5899
rect 13679 5896 13691 5899
rect 14185 5899 14243 5905
rect 14185 5896 14197 5899
rect 13679 5868 14197 5896
rect 13679 5865 13691 5868
rect 13633 5859 13691 5865
rect 14185 5865 14197 5868
rect 14231 5865 14243 5899
rect 14185 5859 14243 5865
rect 14553 5899 14611 5905
rect 14553 5865 14565 5899
rect 14599 5896 14611 5899
rect 15013 5899 15071 5905
rect 15013 5896 15025 5899
rect 14599 5868 15025 5896
rect 14599 5865 14611 5868
rect 14553 5859 14611 5865
rect 15013 5865 15025 5868
rect 15059 5896 15071 5899
rect 16298 5896 16304 5908
rect 15059 5868 16304 5896
rect 15059 5865 15071 5868
rect 15013 5859 15071 5865
rect 16298 5856 16304 5868
rect 16356 5856 16362 5908
rect 2314 5828 2320 5840
rect 1596 5800 2320 5828
rect 1486 5720 1492 5772
rect 1544 5760 1550 5772
rect 1596 5769 1624 5800
rect 2314 5788 2320 5800
rect 2372 5788 2378 5840
rect 5074 5788 5080 5840
rect 5132 5828 5138 5840
rect 8570 5828 8576 5840
rect 5132 5800 7880 5828
rect 5132 5788 5138 5800
rect 1581 5763 1639 5769
rect 1581 5760 1593 5763
rect 1544 5732 1593 5760
rect 1544 5720 1550 5732
rect 1581 5729 1593 5732
rect 1627 5729 1639 5763
rect 1581 5723 1639 5729
rect 1848 5763 1906 5769
rect 1848 5729 1860 5763
rect 1894 5760 1906 5763
rect 3050 5760 3056 5772
rect 1894 5732 3056 5760
rect 1894 5729 1906 5732
rect 1848 5723 1906 5729
rect 3050 5720 3056 5732
rect 3108 5720 3114 5772
rect 3237 5763 3295 5769
rect 3237 5729 3249 5763
rect 3283 5729 3295 5763
rect 3237 5723 3295 5729
rect 3252 5624 3280 5723
rect 4430 5720 4436 5772
rect 4488 5760 4494 5772
rect 4706 5760 4712 5772
rect 4488 5732 4712 5760
rect 4488 5720 4494 5732
rect 4706 5720 4712 5732
rect 4764 5720 4770 5772
rect 5276 5769 5304 5800
rect 5261 5763 5319 5769
rect 5261 5729 5273 5763
rect 5307 5729 5319 5763
rect 5261 5723 5319 5729
rect 5712 5763 5770 5769
rect 5712 5729 5724 5763
rect 5758 5760 5770 5763
rect 6917 5763 6975 5769
rect 6917 5760 6929 5763
rect 5758 5732 6929 5760
rect 5758 5729 5770 5732
rect 5712 5723 5770 5729
rect 6917 5729 6929 5732
rect 6963 5729 6975 5763
rect 6917 5723 6975 5729
rect 7009 5763 7067 5769
rect 7009 5729 7021 5763
rect 7055 5760 7067 5763
rect 7101 5763 7159 5769
rect 7101 5760 7113 5763
rect 7055 5732 7113 5760
rect 7055 5729 7067 5732
rect 7009 5723 7067 5729
rect 7101 5729 7113 5732
rect 7147 5760 7159 5763
rect 7650 5760 7656 5772
rect 7147 5732 7656 5760
rect 7147 5729 7159 5732
rect 7101 5723 7159 5729
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 7852 5769 7880 5800
rect 7944 5800 8576 5828
rect 7944 5769 7972 5800
rect 8570 5788 8576 5800
rect 8628 5788 8634 5840
rect 10502 5828 10508 5840
rect 9876 5800 10508 5828
rect 7837 5763 7895 5769
rect 7837 5729 7849 5763
rect 7883 5729 7895 5763
rect 7837 5723 7895 5729
rect 7929 5763 7987 5769
rect 7929 5729 7941 5763
rect 7975 5729 7987 5763
rect 7929 5723 7987 5729
rect 8196 5763 8254 5769
rect 8196 5729 8208 5763
rect 8242 5760 8254 5763
rect 9214 5760 9220 5772
rect 8242 5732 9220 5760
rect 8242 5729 8254 5732
rect 8196 5723 8254 5729
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 4617 5695 4675 5701
rect 4617 5692 4629 5695
rect 4212 5664 4629 5692
rect 4212 5652 4218 5664
rect 4617 5661 4629 5664
rect 4663 5661 4675 5695
rect 4617 5655 4675 5661
rect 5445 5695 5503 5701
rect 5445 5661 5457 5695
rect 5491 5661 5503 5695
rect 5445 5655 5503 5661
rect 4890 5624 4896 5636
rect 3252 5596 4896 5624
rect 4890 5584 4896 5596
rect 4948 5584 4954 5636
rect 2958 5556 2964 5568
rect 2919 5528 2964 5556
rect 2958 5516 2964 5528
rect 3016 5516 3022 5568
rect 3421 5559 3479 5565
rect 3421 5525 3433 5559
rect 3467 5556 3479 5559
rect 3786 5556 3792 5568
rect 3467 5528 3792 5556
rect 3467 5525 3479 5528
rect 3421 5519 3479 5525
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 4065 5559 4123 5565
rect 4065 5525 4077 5559
rect 4111 5556 4123 5559
rect 4246 5556 4252 5568
rect 4111 5528 4252 5556
rect 4111 5525 4123 5528
rect 4065 5519 4123 5525
rect 4246 5516 4252 5528
rect 4304 5516 4310 5568
rect 5074 5556 5080 5568
rect 5035 5528 5080 5556
rect 5074 5516 5080 5528
rect 5132 5516 5138 5568
rect 5460 5556 5488 5655
rect 7650 5624 7656 5636
rect 6380 5596 7656 5624
rect 6380 5556 6408 5596
rect 7650 5584 7656 5596
rect 7708 5624 7714 5636
rect 7944 5624 7972 5723
rect 9214 5720 9220 5732
rect 9272 5720 9278 5772
rect 9876 5769 9904 5800
rect 10502 5788 10508 5800
rect 10560 5828 10566 5840
rect 13541 5831 13599 5837
rect 10560 5800 11560 5828
rect 10560 5788 10566 5800
rect 9861 5763 9919 5769
rect 9861 5729 9873 5763
rect 9907 5729 9919 5763
rect 9861 5723 9919 5729
rect 10128 5763 10186 5769
rect 10128 5729 10140 5763
rect 10174 5760 10186 5763
rect 10410 5760 10416 5772
rect 10174 5732 10416 5760
rect 10174 5729 10186 5732
rect 10128 5723 10186 5729
rect 10410 5720 10416 5732
rect 10468 5760 10474 5772
rect 10962 5760 10968 5772
rect 10468 5732 10968 5760
rect 10468 5720 10474 5732
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 11532 5769 11560 5800
rect 11624 5800 13492 5828
rect 11517 5763 11575 5769
rect 11517 5729 11529 5763
rect 11563 5729 11575 5763
rect 11517 5723 11575 5729
rect 11624 5692 11652 5800
rect 11784 5763 11842 5769
rect 11784 5729 11796 5763
rect 11830 5760 11842 5763
rect 13464 5760 13492 5800
rect 13541 5797 13553 5831
rect 13587 5828 13599 5831
rect 15378 5828 15384 5840
rect 13587 5800 15384 5828
rect 13587 5797 13599 5800
rect 13541 5791 13599 5797
rect 15378 5788 15384 5800
rect 15436 5788 15442 5840
rect 15013 5763 15071 5769
rect 15013 5760 15025 5763
rect 11830 5732 13400 5760
rect 13464 5732 15025 5760
rect 11830 5729 11842 5732
rect 11784 5723 11842 5729
rect 7708 5596 7972 5624
rect 11164 5664 11652 5692
rect 13372 5692 13400 5732
rect 15013 5729 15025 5732
rect 15059 5729 15071 5763
rect 15013 5723 15071 5729
rect 15657 5763 15715 5769
rect 15657 5729 15669 5763
rect 15703 5760 15715 5763
rect 16298 5760 16304 5772
rect 15703 5732 16304 5760
rect 15703 5729 15715 5732
rect 15657 5723 15715 5729
rect 16298 5720 16304 5732
rect 16356 5720 16362 5772
rect 17310 5760 17316 5772
rect 17271 5732 17316 5760
rect 17310 5720 17316 5732
rect 17368 5720 17374 5772
rect 17402 5720 17408 5772
rect 17460 5760 17466 5772
rect 17865 5763 17923 5769
rect 17865 5760 17877 5763
rect 17460 5732 17877 5760
rect 17460 5720 17466 5732
rect 17865 5729 17877 5732
rect 17911 5729 17923 5763
rect 17865 5723 17923 5729
rect 13538 5692 13544 5704
rect 13372 5664 13544 5692
rect 7708 5584 7714 5596
rect 5460 5528 6408 5556
rect 6638 5516 6644 5568
rect 6696 5556 6702 5568
rect 7009 5559 7067 5565
rect 7009 5556 7021 5559
rect 6696 5528 7021 5556
rect 6696 5516 6702 5528
rect 7009 5525 7021 5528
rect 7055 5525 7067 5559
rect 7009 5519 7067 5525
rect 7285 5559 7343 5565
rect 7285 5525 7297 5559
rect 7331 5556 7343 5559
rect 7374 5556 7380 5568
rect 7331 5528 7380 5556
rect 7331 5525 7343 5528
rect 7285 5519 7343 5525
rect 7374 5516 7380 5528
rect 7432 5516 7438 5568
rect 7742 5516 7748 5568
rect 7800 5556 7806 5568
rect 9766 5556 9772 5568
rect 7800 5528 9772 5556
rect 7800 5516 7806 5528
rect 9766 5516 9772 5528
rect 9824 5556 9830 5568
rect 11164 5556 11192 5664
rect 13538 5652 13544 5664
rect 13596 5692 13602 5704
rect 13725 5695 13783 5701
rect 13725 5692 13737 5695
rect 13596 5664 13737 5692
rect 13596 5652 13602 5664
rect 13725 5661 13737 5664
rect 13771 5661 13783 5695
rect 13725 5655 13783 5661
rect 14274 5652 14280 5704
rect 14332 5692 14338 5704
rect 14645 5695 14703 5701
rect 14645 5692 14657 5695
rect 14332 5664 14657 5692
rect 14332 5652 14338 5664
rect 14645 5661 14657 5664
rect 14691 5661 14703 5695
rect 14645 5655 14703 5661
rect 14829 5695 14887 5701
rect 14829 5661 14841 5695
rect 14875 5692 14887 5695
rect 15102 5692 15108 5704
rect 14875 5664 15108 5692
rect 14875 5661 14887 5664
rect 14829 5655 14887 5661
rect 15102 5652 15108 5664
rect 15160 5652 15166 5704
rect 15746 5692 15752 5704
rect 15707 5664 15752 5692
rect 15746 5652 15752 5664
rect 15804 5652 15810 5704
rect 15841 5695 15899 5701
rect 15841 5661 15853 5695
rect 15887 5661 15899 5695
rect 15841 5655 15899 5661
rect 12989 5627 13047 5633
rect 12989 5593 13001 5627
rect 13035 5624 13047 5627
rect 15856 5624 15884 5655
rect 17494 5624 17500 5636
rect 13035 5596 15884 5624
rect 17455 5596 17500 5624
rect 13035 5593 13047 5596
rect 12989 5587 13047 5593
rect 17494 5584 17500 5596
rect 17552 5584 17558 5636
rect 9824 5528 11192 5556
rect 11241 5559 11299 5565
rect 9824 5516 9830 5528
rect 11241 5525 11253 5559
rect 11287 5556 11299 5559
rect 11698 5556 11704 5568
rect 11287 5528 11704 5556
rect 11287 5525 11299 5528
rect 11241 5519 11299 5525
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 12618 5516 12624 5568
rect 12676 5556 12682 5568
rect 12897 5559 12955 5565
rect 12897 5556 12909 5559
rect 12676 5528 12909 5556
rect 12676 5516 12682 5528
rect 12897 5525 12909 5528
rect 12943 5525 12955 5559
rect 13170 5556 13176 5568
rect 13131 5528 13176 5556
rect 12897 5519 12955 5525
rect 13170 5516 13176 5528
rect 13228 5516 13234 5568
rect 13814 5516 13820 5568
rect 13872 5556 13878 5568
rect 15289 5559 15347 5565
rect 15289 5556 15301 5559
rect 13872 5528 15301 5556
rect 13872 5516 13878 5528
rect 15289 5525 15301 5528
rect 15335 5525 15347 5559
rect 15289 5519 15347 5525
rect 17770 5516 17776 5568
rect 17828 5556 17834 5568
rect 18049 5559 18107 5565
rect 18049 5556 18061 5559
rect 17828 5528 18061 5556
rect 17828 5516 17834 5528
rect 18049 5525 18061 5528
rect 18095 5525 18107 5559
rect 18049 5519 18107 5525
rect 1104 5466 18860 5488
rect 1104 5414 3947 5466
rect 3999 5414 4011 5466
rect 4063 5414 4075 5466
rect 4127 5414 4139 5466
rect 4191 5414 9878 5466
rect 9930 5414 9942 5466
rect 9994 5414 10006 5466
rect 10058 5414 10070 5466
rect 10122 5414 15808 5466
rect 15860 5414 15872 5466
rect 15924 5414 15936 5466
rect 15988 5414 16000 5466
rect 16052 5414 18860 5466
rect 1104 5392 18860 5414
rect 3510 5312 3516 5364
rect 3568 5352 3574 5364
rect 7282 5352 7288 5364
rect 3568 5324 7288 5352
rect 3568 5312 3574 5324
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 7558 5312 7564 5364
rect 7616 5352 7622 5364
rect 8665 5355 8723 5361
rect 8665 5352 8677 5355
rect 7616 5324 8677 5352
rect 7616 5312 7622 5324
rect 8665 5321 8677 5324
rect 8711 5321 8723 5355
rect 9674 5352 9680 5364
rect 9635 5324 9680 5352
rect 8665 5315 8723 5321
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 10594 5312 10600 5364
rect 10652 5352 10658 5364
rect 10689 5355 10747 5361
rect 10689 5352 10701 5355
rect 10652 5324 10701 5352
rect 10652 5312 10658 5324
rect 10689 5321 10701 5324
rect 10735 5321 10747 5355
rect 10689 5315 10747 5321
rect 13538 5312 13544 5364
rect 13596 5352 13602 5364
rect 15289 5355 15347 5361
rect 15289 5352 15301 5355
rect 13596 5324 15301 5352
rect 13596 5312 13602 5324
rect 15289 5321 15301 5324
rect 15335 5321 15347 5355
rect 15289 5315 15347 5321
rect 15378 5312 15384 5364
rect 15436 5352 15442 5364
rect 15565 5355 15623 5361
rect 15565 5352 15577 5355
rect 15436 5324 15577 5352
rect 15436 5312 15442 5324
rect 15565 5321 15577 5324
rect 15611 5321 15623 5355
rect 15565 5315 15623 5321
rect 3050 5244 3056 5296
rect 3108 5284 3114 5296
rect 5258 5284 5264 5296
rect 3108 5256 5264 5284
rect 3108 5244 3114 5256
rect 4246 5216 4252 5228
rect 4207 5188 4252 5216
rect 4246 5176 4252 5188
rect 4304 5176 4310 5228
rect 4356 5225 4384 5256
rect 5258 5244 5264 5256
rect 5316 5284 5322 5296
rect 9398 5284 9404 5296
rect 5316 5256 5396 5284
rect 5316 5244 5322 5256
rect 5368 5225 5396 5256
rect 7208 5256 9404 5284
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5185 4399 5219
rect 4341 5179 4399 5185
rect 5353 5219 5411 5225
rect 5353 5185 5365 5219
rect 5399 5185 5411 5219
rect 5353 5179 5411 5185
rect 6454 5176 6460 5228
rect 6512 5216 6518 5228
rect 7208 5225 7236 5256
rect 9398 5244 9404 5256
rect 9456 5244 9462 5296
rect 9858 5244 9864 5296
rect 9916 5284 9922 5296
rect 13814 5284 13820 5296
rect 9916 5256 13820 5284
rect 9916 5244 9922 5256
rect 13814 5244 13820 5256
rect 13872 5244 13878 5296
rect 7193 5219 7251 5225
rect 6512 5188 7144 5216
rect 6512 5176 6518 5188
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 1486 5148 1492 5160
rect 1443 5120 1492 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 1486 5108 1492 5120
rect 1544 5108 1550 5160
rect 3053 5151 3111 5157
rect 3053 5117 3065 5151
rect 3099 5148 3111 5151
rect 3099 5120 4108 5148
rect 3099 5117 3111 5120
rect 3053 5111 3111 5117
rect 1664 5083 1722 5089
rect 1664 5049 1676 5083
rect 1710 5080 1722 5083
rect 2958 5080 2964 5092
rect 1710 5052 2964 5080
rect 1710 5049 1722 5052
rect 1664 5043 1722 5049
rect 2958 5040 2964 5052
rect 3016 5040 3022 5092
rect 3329 5083 3387 5089
rect 3329 5049 3341 5083
rect 3375 5080 3387 5083
rect 3510 5080 3516 5092
rect 3375 5052 3516 5080
rect 3375 5049 3387 5052
rect 3329 5043 3387 5049
rect 3510 5040 3516 5052
rect 3568 5040 3574 5092
rect 4080 5080 4108 5120
rect 4154 5108 4160 5160
rect 4212 5148 4218 5160
rect 4212 5120 4257 5148
rect 4212 5108 4218 5120
rect 4706 5108 4712 5160
rect 4764 5148 4770 5160
rect 5813 5151 5871 5157
rect 4764 5120 5120 5148
rect 4764 5108 4770 5120
rect 4982 5080 4988 5092
rect 4080 5052 4988 5080
rect 4982 5040 4988 5052
rect 5040 5040 5046 5092
rect 5092 5080 5120 5120
rect 5813 5117 5825 5151
rect 5859 5148 5871 5151
rect 5994 5148 6000 5160
rect 5859 5120 6000 5148
rect 5859 5117 5871 5120
rect 5813 5111 5871 5117
rect 5994 5108 6000 5120
rect 6052 5108 6058 5160
rect 6914 5148 6920 5160
rect 6875 5120 6920 5148
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7116 5148 7144 5188
rect 7193 5185 7205 5219
rect 7239 5185 7251 5219
rect 7193 5179 7251 5185
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 7742 5216 7748 5228
rect 7607 5188 7748 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 7742 5176 7748 5188
rect 7800 5176 7806 5228
rect 8018 5176 8024 5228
rect 8076 5216 8082 5228
rect 8205 5219 8263 5225
rect 8205 5216 8217 5219
rect 8076 5188 8217 5216
rect 8076 5176 8082 5188
rect 8205 5185 8217 5188
rect 8251 5185 8263 5219
rect 9122 5216 9128 5228
rect 9083 5188 9128 5216
rect 8205 5179 8263 5185
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 9309 5219 9367 5225
rect 9309 5185 9321 5219
rect 9355 5216 9367 5219
rect 10229 5219 10287 5225
rect 10229 5216 10241 5219
rect 9355 5188 10241 5216
rect 9355 5185 9367 5188
rect 9309 5179 9367 5185
rect 10229 5185 10241 5188
rect 10275 5216 10287 5219
rect 11241 5219 11299 5225
rect 11241 5216 11253 5219
rect 10275 5188 11253 5216
rect 10275 5185 10287 5188
rect 10229 5179 10287 5185
rect 11241 5185 11253 5188
rect 11287 5185 11299 5219
rect 11241 5179 11299 5185
rect 8113 5151 8171 5157
rect 8113 5148 8125 5151
rect 7116 5120 8125 5148
rect 8113 5117 8125 5120
rect 8159 5148 8171 5151
rect 8159 5120 9168 5148
rect 8159 5117 8171 5120
rect 8113 5111 8171 5117
rect 5261 5083 5319 5089
rect 5261 5080 5273 5083
rect 5092 5052 5273 5080
rect 5261 5049 5273 5052
rect 5307 5049 5319 5083
rect 5261 5043 5319 5049
rect 6089 5083 6147 5089
rect 6089 5049 6101 5083
rect 6135 5080 6147 5083
rect 6454 5080 6460 5092
rect 6135 5052 6460 5080
rect 6135 5049 6147 5052
rect 6089 5043 6147 5049
rect 2774 4972 2780 5024
rect 2832 5012 2838 5024
rect 2832 4984 2877 5012
rect 2832 4972 2838 4984
rect 3418 4972 3424 5024
rect 3476 5012 3482 5024
rect 3789 5015 3847 5021
rect 3789 5012 3801 5015
rect 3476 4984 3801 5012
rect 3476 4972 3482 4984
rect 3789 4981 3801 4984
rect 3835 4981 3847 5015
rect 3789 4975 3847 4981
rect 4430 4972 4436 5024
rect 4488 5012 4494 5024
rect 4614 5012 4620 5024
rect 4488 4984 4620 5012
rect 4488 4972 4494 4984
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 4798 5012 4804 5024
rect 4759 4984 4804 5012
rect 4798 4972 4804 4984
rect 4856 4972 4862 5024
rect 5166 5012 5172 5024
rect 5127 4984 5172 5012
rect 5166 4972 5172 4984
rect 5224 4972 5230 5024
rect 5276 5012 5304 5043
rect 6454 5040 6460 5052
rect 6512 5040 6518 5092
rect 9033 5083 9091 5089
rect 9033 5080 9045 5083
rect 7668 5052 9045 5080
rect 7668 5021 7696 5052
rect 9033 5049 9045 5052
rect 9079 5049 9091 5083
rect 9140 5080 9168 5120
rect 9214 5108 9220 5160
rect 9272 5148 9278 5160
rect 9324 5148 9352 5179
rect 11330 5176 11336 5228
rect 11388 5216 11394 5228
rect 13170 5216 13176 5228
rect 11388 5188 13176 5216
rect 11388 5176 11394 5188
rect 13170 5176 13176 5188
rect 13228 5176 13234 5228
rect 13538 5216 13544 5228
rect 13499 5188 13544 5216
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 15102 5176 15108 5228
rect 15160 5216 15166 5228
rect 16117 5219 16175 5225
rect 16117 5216 16129 5219
rect 15160 5188 16129 5216
rect 15160 5176 15166 5188
rect 16117 5185 16129 5188
rect 16163 5185 16175 5219
rect 16117 5179 16175 5185
rect 9272 5120 9352 5148
rect 9272 5108 9278 5120
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 10686 5148 10692 5160
rect 10100 5120 10692 5148
rect 10100 5108 10106 5120
rect 10686 5108 10692 5120
rect 10744 5108 10750 5160
rect 11054 5148 11060 5160
rect 11015 5120 11060 5148
rect 11054 5108 11060 5120
rect 11112 5108 11118 5160
rect 11149 5151 11207 5157
rect 11149 5117 11161 5151
rect 11195 5148 11207 5151
rect 11422 5148 11428 5160
rect 11195 5120 11428 5148
rect 11195 5117 11207 5120
rect 11149 5111 11207 5117
rect 11422 5108 11428 5120
rect 11480 5108 11486 5160
rect 11701 5151 11759 5157
rect 11701 5117 11713 5151
rect 11747 5148 11759 5151
rect 12250 5148 12256 5160
rect 11747 5120 12256 5148
rect 11747 5117 11759 5120
rect 11701 5111 11759 5117
rect 12250 5108 12256 5120
rect 12308 5108 12314 5160
rect 13906 5148 13912 5160
rect 13867 5120 13912 5148
rect 13906 5108 13912 5120
rect 13964 5108 13970 5160
rect 14176 5151 14234 5157
rect 14176 5117 14188 5151
rect 14222 5148 14234 5151
rect 15120 5148 15148 5176
rect 16022 5148 16028 5160
rect 14222 5120 15148 5148
rect 15935 5120 16028 5148
rect 14222 5117 14234 5120
rect 14176 5111 14234 5117
rect 16022 5108 16028 5120
rect 16080 5148 16086 5160
rect 16574 5148 16580 5160
rect 16080 5120 16580 5148
rect 16080 5108 16086 5120
rect 16574 5108 16580 5120
rect 16632 5108 16638 5160
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5117 18107 5151
rect 18049 5111 18107 5117
rect 12526 5080 12532 5092
rect 9140 5052 12532 5080
rect 9033 5043 9091 5049
rect 12526 5040 12532 5052
rect 12584 5080 12590 5092
rect 13170 5080 13176 5092
rect 12584 5052 13176 5080
rect 12584 5040 12590 5052
rect 13170 5040 13176 5052
rect 13228 5040 13234 5092
rect 13265 5083 13323 5089
rect 13265 5049 13277 5083
rect 13311 5080 13323 5083
rect 13998 5080 14004 5092
rect 13311 5052 14004 5080
rect 13311 5049 13323 5052
rect 13265 5043 13323 5049
rect 13998 5040 14004 5052
rect 14056 5040 14062 5092
rect 18064 5080 18092 5111
rect 14108 5052 18092 5080
rect 7561 5015 7619 5021
rect 7561 5012 7573 5015
rect 5276 4984 7573 5012
rect 7561 4981 7573 4984
rect 7607 4981 7619 5015
rect 7561 4975 7619 4981
rect 7653 5015 7711 5021
rect 7653 4981 7665 5015
rect 7699 4981 7711 5015
rect 7653 4975 7711 4981
rect 7742 4972 7748 5024
rect 7800 5012 7806 5024
rect 8021 5015 8079 5021
rect 8021 5012 8033 5015
rect 7800 4984 8033 5012
rect 7800 4972 7806 4984
rect 8021 4981 8033 4984
rect 8067 5012 8079 5015
rect 9674 5012 9680 5024
rect 8067 4984 9680 5012
rect 8067 4981 8079 4984
rect 8021 4975 8079 4981
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 9766 4972 9772 5024
rect 9824 5012 9830 5024
rect 10045 5015 10103 5021
rect 10045 5012 10057 5015
rect 9824 4984 10057 5012
rect 9824 4972 9830 4984
rect 10045 4981 10057 4984
rect 10091 4981 10103 5015
rect 10045 4975 10103 4981
rect 10137 5015 10195 5021
rect 10137 4981 10149 5015
rect 10183 5012 10195 5015
rect 10778 5012 10784 5024
rect 10183 4984 10784 5012
rect 10183 4981 10195 4984
rect 10137 4975 10195 4981
rect 10778 4972 10784 4984
rect 10836 4972 10842 5024
rect 11422 4972 11428 5024
rect 11480 5012 11486 5024
rect 12897 5015 12955 5021
rect 12897 5012 12909 5015
rect 11480 4984 12909 5012
rect 11480 4972 11486 4984
rect 12897 4981 12909 4984
rect 12943 4981 12955 5015
rect 12897 4975 12955 4981
rect 13357 5015 13415 5021
rect 13357 4981 13369 5015
rect 13403 5012 13415 5015
rect 13630 5012 13636 5024
rect 13403 4984 13636 5012
rect 13403 4981 13415 4984
rect 13357 4975 13415 4981
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 13722 4972 13728 5024
rect 13780 5012 13786 5024
rect 14108 5012 14136 5052
rect 13780 4984 14136 5012
rect 13780 4972 13786 4984
rect 15010 4972 15016 5024
rect 15068 5012 15074 5024
rect 15286 5012 15292 5024
rect 15068 4984 15292 5012
rect 15068 4972 15074 4984
rect 15286 4972 15292 4984
rect 15344 4972 15350 5024
rect 15930 5012 15936 5024
rect 15891 4984 15936 5012
rect 15930 4972 15936 4984
rect 15988 4972 15994 5024
rect 18230 5012 18236 5024
rect 18191 4984 18236 5012
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 1104 4922 18860 4944
rect 1104 4870 6912 4922
rect 6964 4870 6976 4922
rect 7028 4870 7040 4922
rect 7092 4870 7104 4922
rect 7156 4870 12843 4922
rect 12895 4870 12907 4922
rect 12959 4870 12971 4922
rect 13023 4870 13035 4922
rect 13087 4870 18860 4922
rect 1104 4848 18860 4870
rect 2317 4811 2375 4817
rect 2317 4777 2329 4811
rect 2363 4808 2375 4811
rect 3142 4808 3148 4820
rect 2363 4780 3148 4808
rect 2363 4777 2375 4780
rect 2317 4771 2375 4777
rect 3142 4768 3148 4780
rect 3200 4768 3206 4820
rect 4706 4808 4712 4820
rect 3252 4780 4712 4808
rect 3252 4740 3280 4780
rect 4706 4768 4712 4780
rect 4764 4768 4770 4820
rect 5445 4811 5503 4817
rect 5445 4777 5457 4811
rect 5491 4808 5503 4811
rect 5534 4808 5540 4820
rect 5491 4780 5540 4808
rect 5491 4777 5503 4780
rect 5445 4771 5503 4777
rect 5534 4768 5540 4780
rect 5592 4768 5598 4820
rect 5902 4768 5908 4820
rect 5960 4808 5966 4820
rect 6733 4811 6791 4817
rect 6733 4808 6745 4811
rect 5960 4780 6745 4808
rect 5960 4768 5966 4780
rect 6733 4777 6745 4780
rect 6779 4777 6791 4811
rect 6733 4771 6791 4777
rect 7745 4811 7803 4817
rect 7745 4777 7757 4811
rect 7791 4808 7803 4811
rect 9122 4808 9128 4820
rect 7791 4780 9128 4808
rect 7791 4777 7803 4780
rect 7745 4771 7803 4777
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 9677 4811 9735 4817
rect 9677 4777 9689 4811
rect 9723 4808 9735 4811
rect 10226 4808 10232 4820
rect 9723 4780 10232 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 10226 4768 10232 4780
rect 10284 4768 10290 4820
rect 10502 4768 10508 4820
rect 10560 4808 10566 4820
rect 10689 4811 10747 4817
rect 10689 4808 10701 4811
rect 10560 4780 10701 4808
rect 10560 4768 10566 4780
rect 10689 4777 10701 4780
rect 10735 4777 10747 4811
rect 11422 4808 11428 4820
rect 11383 4780 11428 4808
rect 10689 4771 10747 4777
rect 11422 4768 11428 4780
rect 11480 4768 11486 4820
rect 13354 4808 13360 4820
rect 13315 4780 13360 4808
rect 13354 4768 13360 4780
rect 13412 4768 13418 4820
rect 13630 4808 13636 4820
rect 13591 4780 13636 4808
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 14645 4811 14703 4817
rect 14645 4777 14657 4811
rect 14691 4808 14703 4811
rect 15930 4808 15936 4820
rect 14691 4780 15936 4808
rect 14691 4777 14703 4780
rect 14645 4771 14703 4777
rect 15930 4768 15936 4780
rect 15988 4768 15994 4820
rect 1412 4712 3280 4740
rect 3329 4743 3387 4749
rect 1412 4681 1440 4712
rect 3329 4709 3341 4743
rect 3375 4740 3387 4743
rect 4798 4740 4804 4752
rect 3375 4712 4804 4740
rect 3375 4709 3387 4712
rect 3329 4703 3387 4709
rect 4798 4700 4804 4712
rect 4856 4700 4862 4752
rect 5258 4700 5264 4752
rect 5316 4740 5322 4752
rect 8110 4740 8116 4752
rect 5316 4712 6408 4740
rect 5316 4700 5322 4712
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4641 1455 4675
rect 1397 4635 1455 4641
rect 2409 4675 2467 4681
rect 2409 4641 2421 4675
rect 2455 4672 2467 4675
rect 3234 4672 3240 4684
rect 2455 4644 3240 4672
rect 2455 4641 2467 4644
rect 2409 4635 2467 4641
rect 3234 4632 3240 4644
rect 3292 4632 3298 4684
rect 3418 4632 3424 4684
rect 3476 4672 3482 4684
rect 4338 4681 4344 4684
rect 4332 4672 4344 4681
rect 3476 4644 3521 4672
rect 4299 4644 4344 4672
rect 3476 4632 3482 4644
rect 4332 4635 4344 4644
rect 4338 4632 4344 4635
rect 4396 4632 4402 4684
rect 4614 4632 4620 4684
rect 4672 4672 4678 4684
rect 4672 4644 5764 4672
rect 4672 4632 4678 4644
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4604 2651 4607
rect 2958 4604 2964 4616
rect 2639 4576 2964 4604
rect 2639 4573 2651 4576
rect 2593 4567 2651 4573
rect 2958 4564 2964 4576
rect 3016 4604 3022 4616
rect 3513 4607 3571 4613
rect 3513 4604 3525 4607
rect 3016 4576 3525 4604
rect 3016 4564 3022 4576
rect 3513 4573 3525 4576
rect 3559 4573 3571 4607
rect 3513 4567 3571 4573
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 1949 4539 2007 4545
rect 1949 4505 1961 4539
rect 1995 4536 2007 4539
rect 3050 4536 3056 4548
rect 1995 4508 3056 4536
rect 1995 4505 2007 4508
rect 1949 4499 2007 4505
rect 3050 4496 3056 4508
rect 3108 4496 3114 4548
rect 3418 4496 3424 4548
rect 3476 4536 3482 4548
rect 4080 4536 4108 4567
rect 3476 4508 4108 4536
rect 5736 4536 5764 4644
rect 5810 4632 5816 4684
rect 5868 4672 5874 4684
rect 6089 4675 6147 4681
rect 6089 4672 6101 4675
rect 5868 4644 6101 4672
rect 5868 4632 5874 4644
rect 6089 4641 6101 4644
rect 6135 4641 6147 4675
rect 6089 4635 6147 4641
rect 6178 4632 6184 4684
rect 6236 4672 6242 4684
rect 6236 4644 6281 4672
rect 6236 4632 6242 4644
rect 6380 4613 6408 4712
rect 7024 4712 8116 4740
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 7024 4536 7052 4712
rect 8110 4700 8116 4712
rect 8168 4700 8174 4752
rect 9214 4700 9220 4752
rect 9272 4740 9278 4752
rect 11330 4740 11336 4752
rect 9272 4712 10180 4740
rect 11291 4712 11336 4740
rect 9272 4700 9278 4712
rect 7101 4675 7159 4681
rect 7101 4641 7113 4675
rect 7147 4672 7159 4675
rect 7147 4644 7880 4672
rect 7147 4641 7159 4644
rect 7101 4635 7159 4641
rect 7190 4604 7196 4616
rect 7151 4576 7196 4604
rect 7190 4564 7196 4576
rect 7248 4564 7254 4616
rect 7282 4564 7288 4616
rect 7340 4604 7346 4616
rect 7340 4576 7385 4604
rect 7340 4564 7346 4576
rect 5736 4508 7052 4536
rect 7852 4536 7880 4644
rect 8018 4632 8024 4684
rect 8076 4672 8082 4684
rect 8757 4675 8815 4681
rect 8076 4644 8340 4672
rect 8076 4632 8082 4644
rect 7926 4564 7932 4616
rect 7984 4604 7990 4616
rect 8202 4604 8208 4616
rect 7984 4576 8208 4604
rect 7984 4564 7990 4576
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 8312 4613 8340 4644
rect 8757 4641 8769 4675
rect 8803 4672 8815 4675
rect 9858 4672 9864 4684
rect 8803 4644 9864 4672
rect 8803 4641 8815 4644
rect 8757 4635 8815 4641
rect 9858 4632 9864 4644
rect 9916 4632 9922 4684
rect 10042 4672 10048 4684
rect 10003 4644 10048 4672
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 10152 4672 10180 4712
rect 11330 4700 11336 4712
rect 11388 4700 11394 4752
rect 12222 4743 12280 4749
rect 12222 4740 12234 4743
rect 11624 4712 12234 4740
rect 10873 4675 10931 4681
rect 10152 4644 10272 4672
rect 8297 4607 8355 4613
rect 8297 4573 8309 4607
rect 8343 4573 8355 4607
rect 8297 4567 8355 4573
rect 8478 4564 8484 4616
rect 8536 4604 8542 4616
rect 8941 4607 8999 4613
rect 8941 4604 8953 4607
rect 8536 4576 8953 4604
rect 8536 4564 8542 4576
rect 8941 4573 8953 4576
rect 8987 4573 8999 4607
rect 8941 4567 8999 4573
rect 9122 4564 9128 4616
rect 9180 4604 9186 4616
rect 10244 4613 10272 4644
rect 10873 4641 10885 4675
rect 10919 4672 10931 4675
rect 11514 4672 11520 4684
rect 10919 4644 11520 4672
rect 10919 4641 10931 4644
rect 10873 4635 10931 4641
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 11624 4613 11652 4712
rect 12222 4709 12234 4712
rect 12268 4740 12280 4743
rect 12618 4740 12624 4752
rect 12268 4712 12624 4740
rect 12268 4709 12280 4712
rect 12222 4703 12280 4709
rect 12618 4700 12624 4712
rect 12676 4700 12682 4752
rect 15194 4740 15200 4752
rect 13832 4712 15200 4740
rect 13832 4672 13860 4712
rect 15194 4700 15200 4712
rect 15252 4700 15258 4752
rect 15562 4740 15568 4752
rect 15304 4712 15568 4740
rect 14001 4675 14059 4681
rect 14001 4672 14013 4675
rect 11716 4644 13860 4672
rect 13924 4644 14013 4672
rect 10137 4607 10195 4613
rect 10137 4604 10149 4607
rect 9180 4576 10149 4604
rect 9180 4564 9186 4576
rect 10137 4573 10149 4576
rect 10183 4573 10195 4607
rect 10137 4567 10195 4573
rect 10229 4607 10287 4613
rect 10229 4573 10241 4607
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 11609 4607 11667 4613
rect 11609 4573 11621 4607
rect 11655 4573 11667 4607
rect 11609 4567 11667 4573
rect 8386 4536 8392 4548
rect 7852 4508 8392 4536
rect 3476 4496 3482 4508
rect 8386 4496 8392 4508
rect 8444 4496 8450 4548
rect 8662 4496 8668 4548
rect 8720 4536 8726 4548
rect 11716 4536 11744 4644
rect 11974 4604 11980 4616
rect 11935 4576 11980 4604
rect 11974 4564 11980 4576
rect 12032 4564 12038 4616
rect 13170 4564 13176 4616
rect 13228 4604 13234 4616
rect 13924 4604 13952 4644
rect 14001 4641 14013 4644
rect 14047 4672 14059 4675
rect 15304 4672 15332 4712
rect 15562 4700 15568 4712
rect 15620 4700 15626 4752
rect 15746 4740 15752 4752
rect 15707 4712 15752 4740
rect 15746 4700 15752 4712
rect 15804 4700 15810 4752
rect 15654 4672 15660 4684
rect 14047 4644 15332 4672
rect 15615 4644 15660 4672
rect 14047 4641 14059 4644
rect 14001 4635 14059 4641
rect 15654 4632 15660 4644
rect 15712 4672 15718 4684
rect 17034 4672 17040 4684
rect 15712 4644 17040 4672
rect 15712 4632 15718 4644
rect 17034 4632 17040 4644
rect 17092 4632 17098 4684
rect 17218 4632 17224 4684
rect 17276 4672 17282 4684
rect 17313 4675 17371 4681
rect 17313 4672 17325 4675
rect 17276 4644 17325 4672
rect 17276 4632 17282 4644
rect 17313 4641 17325 4644
rect 17359 4641 17371 4675
rect 17862 4672 17868 4684
rect 17823 4644 17868 4672
rect 17313 4635 17371 4641
rect 17862 4632 17868 4644
rect 17920 4632 17926 4684
rect 14090 4604 14096 4616
rect 13228 4576 13952 4604
rect 14051 4576 14096 4604
rect 13228 4564 13234 4576
rect 14090 4564 14096 4576
rect 14148 4564 14154 4616
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4604 14335 4607
rect 15102 4604 15108 4616
rect 14323 4576 15108 4604
rect 14323 4573 14335 4576
rect 14277 4567 14335 4573
rect 15102 4564 15108 4576
rect 15160 4564 15166 4616
rect 15841 4607 15899 4613
rect 15841 4573 15853 4607
rect 15887 4573 15899 4607
rect 15841 4567 15899 4573
rect 8720 4508 11744 4536
rect 8720 4496 8726 4508
rect 13906 4496 13912 4548
rect 13964 4536 13970 4548
rect 15856 4536 15884 4567
rect 13964 4508 15884 4536
rect 13964 4496 13970 4508
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 2958 4468 2964 4480
rect 2919 4440 2964 4468
rect 2958 4428 2964 4440
rect 3016 4428 3022 4480
rect 3234 4428 3240 4480
rect 3292 4468 3298 4480
rect 5721 4471 5779 4477
rect 5721 4468 5733 4471
rect 3292 4440 5733 4468
rect 3292 4428 3298 4440
rect 5721 4437 5733 4440
rect 5767 4437 5779 4471
rect 5721 4431 5779 4437
rect 9674 4428 9680 4480
rect 9732 4468 9738 4480
rect 10870 4468 10876 4480
rect 9732 4440 10876 4468
rect 9732 4428 9738 4440
rect 10870 4428 10876 4440
rect 10928 4428 10934 4480
rect 10965 4471 11023 4477
rect 10965 4437 10977 4471
rect 11011 4468 11023 4471
rect 11422 4468 11428 4480
rect 11011 4440 11428 4468
rect 11011 4437 11023 4440
rect 10965 4431 11023 4437
rect 11422 4428 11428 4440
rect 11480 4428 11486 4480
rect 11974 4428 11980 4480
rect 12032 4468 12038 4480
rect 13354 4468 13360 4480
rect 12032 4440 13360 4468
rect 12032 4428 12038 4440
rect 13354 4428 13360 4440
rect 13412 4468 13418 4480
rect 13814 4468 13820 4480
rect 13412 4440 13820 4468
rect 13412 4428 13418 4440
rect 13814 4428 13820 4440
rect 13872 4428 13878 4480
rect 15286 4468 15292 4480
rect 15247 4440 15292 4468
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 17494 4468 17500 4480
rect 17455 4440 17500 4468
rect 17494 4428 17500 4440
rect 17552 4428 17558 4480
rect 17862 4428 17868 4480
rect 17920 4468 17926 4480
rect 18049 4471 18107 4477
rect 18049 4468 18061 4471
rect 17920 4440 18061 4468
rect 17920 4428 17926 4440
rect 18049 4437 18061 4440
rect 18095 4437 18107 4471
rect 18049 4431 18107 4437
rect 1104 4378 18860 4400
rect 1104 4326 3947 4378
rect 3999 4326 4011 4378
rect 4063 4326 4075 4378
rect 4127 4326 4139 4378
rect 4191 4326 9878 4378
rect 9930 4326 9942 4378
rect 9994 4326 10006 4378
rect 10058 4326 10070 4378
rect 10122 4326 15808 4378
rect 15860 4326 15872 4378
rect 15924 4326 15936 4378
rect 15988 4326 16000 4378
rect 16052 4326 18860 4378
rect 1104 4304 18860 4326
rect 4982 4224 4988 4276
rect 5040 4264 5046 4276
rect 5718 4264 5724 4276
rect 5040 4236 5724 4264
rect 5040 4224 5046 4236
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 5994 4224 6000 4276
rect 6052 4264 6058 4276
rect 9125 4267 9183 4273
rect 6052 4236 8708 4264
rect 6052 4224 6058 4236
rect 7282 4196 7288 4208
rect 5920 4168 7288 4196
rect 5920 4137 5948 4168
rect 7282 4156 7288 4168
rect 7340 4156 7346 4208
rect 8680 4196 8708 4236
rect 9125 4233 9137 4267
rect 9171 4264 9183 4267
rect 9214 4264 9220 4276
rect 9171 4236 9220 4264
rect 9171 4233 9183 4236
rect 9125 4227 9183 4233
rect 9214 4224 9220 4236
rect 9272 4224 9278 4276
rect 10318 4264 10324 4276
rect 9324 4236 10324 4264
rect 9324 4196 9352 4236
rect 10318 4224 10324 4236
rect 10376 4224 10382 4276
rect 10870 4224 10876 4276
rect 10928 4264 10934 4276
rect 10928 4236 12572 4264
rect 10928 4224 10934 4236
rect 12158 4196 12164 4208
rect 8680 4168 9352 4196
rect 11900 4168 12164 4196
rect 5169 4131 5227 4137
rect 5169 4097 5181 4131
rect 5215 4128 5227 4131
rect 5905 4131 5963 4137
rect 5905 4128 5917 4131
rect 5215 4100 5917 4128
rect 5215 4097 5227 4100
rect 5169 4091 5227 4097
rect 5905 4097 5917 4100
rect 5951 4097 5963 4131
rect 7374 4128 7380 4140
rect 5905 4091 5963 4097
rect 6012 4100 7380 4128
rect 1489 4063 1547 4069
rect 1489 4029 1501 4063
rect 1535 4060 1547 4063
rect 1670 4060 1676 4072
rect 1535 4032 1676 4060
rect 1535 4029 1547 4032
rect 1489 4023 1547 4029
rect 1670 4020 1676 4032
rect 1728 4060 1734 4072
rect 1946 4060 1952 4072
rect 1728 4032 1952 4060
rect 1728 4020 1734 4032
rect 1946 4020 1952 4032
rect 2004 4020 2010 4072
rect 2041 4063 2099 4069
rect 2041 4029 2053 4063
rect 2087 4060 2099 4063
rect 3418 4060 3424 4072
rect 2087 4032 3424 4060
rect 2087 4029 2099 4032
rect 2041 4023 2099 4029
rect 3418 4020 3424 4032
rect 3476 4060 3482 4072
rect 3694 4060 3700 4072
rect 3476 4032 3700 4060
rect 3476 4020 3482 4032
rect 3694 4020 3700 4032
rect 3752 4020 3758 4072
rect 6012 4060 6040 4100
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 7650 4088 7656 4140
rect 7708 4128 7714 4140
rect 7745 4131 7803 4137
rect 7745 4128 7757 4131
rect 7708 4100 7757 4128
rect 7708 4088 7714 4100
rect 7745 4097 7757 4100
rect 7791 4097 7803 4131
rect 7745 4091 7803 4097
rect 11054 4088 11060 4140
rect 11112 4128 11118 4140
rect 11606 4128 11612 4140
rect 11112 4100 11612 4128
rect 11112 4088 11118 4100
rect 11606 4088 11612 4100
rect 11664 4128 11670 4140
rect 11900 4137 11928 4168
rect 12158 4156 12164 4168
rect 12216 4156 12222 4208
rect 11793 4131 11851 4137
rect 11793 4128 11805 4131
rect 11664 4100 11805 4128
rect 11664 4088 11670 4100
rect 11793 4097 11805 4100
rect 11839 4097 11851 4131
rect 11793 4091 11851 4097
rect 11885 4131 11943 4137
rect 11885 4097 11897 4131
rect 11931 4097 11943 4131
rect 12544 4128 12572 4236
rect 13998 4224 14004 4276
rect 14056 4264 14062 4276
rect 15013 4267 15071 4273
rect 15013 4264 15025 4267
rect 14056 4236 15025 4264
rect 14056 4224 14062 4236
rect 15013 4233 15025 4236
rect 15059 4233 15071 4267
rect 15013 4227 15071 4233
rect 14737 4199 14795 4205
rect 14737 4165 14749 4199
rect 14783 4196 14795 4199
rect 15102 4196 15108 4208
rect 14783 4168 15108 4196
rect 14783 4165 14795 4168
rect 14737 4159 14795 4165
rect 15102 4156 15108 4168
rect 15160 4196 15166 4208
rect 15160 4168 15608 4196
rect 15160 4156 15166 4168
rect 12544 4100 13492 4128
rect 11885 4091 11943 4097
rect 4080 4032 6040 4060
rect 4080 4004 4108 4032
rect 6730 4020 6736 4072
rect 6788 4060 6794 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6788 4032 6837 4060
rect 6788 4020 6794 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 9677 4063 9735 4069
rect 9677 4029 9689 4063
rect 9723 4060 9735 4063
rect 10502 4060 10508 4072
rect 9723 4032 10508 4060
rect 9723 4029 9735 4032
rect 9677 4023 9735 4029
rect 10502 4020 10508 4032
rect 10560 4020 10566 4072
rect 12066 4020 12072 4072
rect 12124 4060 12130 4072
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 12124 4032 12449 4060
rect 12124 4020 12130 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 13354 4060 13360 4072
rect 13315 4032 13360 4060
rect 12437 4023 12495 4029
rect 13354 4020 13360 4032
rect 13412 4020 13418 4072
rect 13464 4060 13492 4100
rect 14458 4088 14464 4140
rect 14516 4128 14522 4140
rect 14918 4128 14924 4140
rect 14516 4100 14924 4128
rect 14516 4088 14522 4100
rect 14918 4088 14924 4100
rect 14976 4088 14982 4140
rect 15580 4137 15608 4168
rect 15565 4131 15623 4137
rect 15565 4097 15577 4131
rect 15611 4097 15623 4131
rect 15565 4091 15623 4097
rect 15473 4063 15531 4069
rect 15473 4060 15485 4063
rect 13464 4032 15485 4060
rect 15473 4029 15485 4032
rect 15519 4029 15531 4063
rect 15473 4023 15531 4029
rect 17405 4063 17463 4069
rect 17405 4029 17417 4063
rect 17451 4029 17463 4063
rect 17405 4023 17463 4029
rect 18049 4063 18107 4069
rect 18049 4029 18061 4063
rect 18095 4060 18107 4063
rect 18138 4060 18144 4072
rect 18095 4032 18144 4060
rect 18095 4029 18107 4032
rect 18049 4023 18107 4029
rect 2308 3995 2366 4001
rect 2308 3961 2320 3995
rect 2354 3992 2366 3995
rect 2774 3992 2780 4004
rect 2354 3964 2780 3992
rect 2354 3961 2366 3964
rect 2308 3955 2366 3961
rect 2774 3952 2780 3964
rect 2832 3952 2838 4004
rect 3942 3995 4000 4001
rect 3942 3992 3954 3995
rect 3436 3964 3954 3992
rect 3436 3936 3464 3964
rect 3942 3961 3954 3964
rect 3988 3961 4000 3995
rect 3942 3955 4000 3961
rect 4062 3952 4068 4004
rect 4120 3952 4126 4004
rect 4890 3952 4896 4004
rect 4948 3992 4954 4004
rect 8018 4001 8024 4004
rect 7101 3995 7159 4001
rect 7101 3992 7113 3995
rect 4948 3964 7113 3992
rect 4948 3952 4954 3964
rect 7101 3961 7113 3964
rect 7147 3961 7159 3995
rect 8012 3992 8024 4001
rect 7979 3964 8024 3992
rect 7101 3955 7159 3961
rect 8012 3955 8024 3964
rect 8018 3952 8024 3955
rect 8076 3952 8082 4004
rect 8110 3952 8116 4004
rect 8168 3992 8174 4004
rect 9944 3995 10002 4001
rect 8168 3964 9904 3992
rect 8168 3952 8174 3964
rect 1670 3924 1676 3936
rect 1631 3896 1676 3924
rect 1670 3884 1676 3896
rect 1728 3884 1734 3936
rect 3418 3924 3424 3936
rect 3379 3896 3424 3924
rect 3418 3884 3424 3896
rect 3476 3884 3482 3936
rect 4338 3884 4344 3936
rect 4396 3924 4402 3936
rect 5077 3927 5135 3933
rect 5077 3924 5089 3927
rect 4396 3896 5089 3924
rect 4396 3884 4402 3896
rect 5077 3893 5089 3896
rect 5123 3924 5135 3927
rect 5169 3927 5227 3933
rect 5169 3924 5181 3927
rect 5123 3896 5181 3924
rect 5123 3893 5135 3896
rect 5077 3887 5135 3893
rect 5169 3893 5181 3896
rect 5215 3893 5227 3927
rect 5350 3924 5356 3936
rect 5311 3896 5356 3924
rect 5169 3887 5227 3893
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 5626 3884 5632 3936
rect 5684 3924 5690 3936
rect 5721 3927 5779 3933
rect 5721 3924 5733 3927
rect 5684 3896 5733 3924
rect 5684 3884 5690 3896
rect 5721 3893 5733 3896
rect 5767 3893 5779 3927
rect 5721 3887 5779 3893
rect 5813 3927 5871 3933
rect 5813 3893 5825 3927
rect 5859 3924 5871 3927
rect 5994 3924 6000 3936
rect 5859 3896 6000 3924
rect 5859 3893 5871 3896
rect 5813 3887 5871 3893
rect 5994 3884 6000 3896
rect 6052 3884 6058 3936
rect 6086 3884 6092 3936
rect 6144 3924 6150 3936
rect 9674 3924 9680 3936
rect 6144 3896 9680 3924
rect 6144 3884 6150 3896
rect 9674 3884 9680 3896
rect 9732 3884 9738 3936
rect 9876 3924 9904 3964
rect 9944 3961 9956 3995
rect 9990 3992 10002 3995
rect 10042 3992 10048 4004
rect 9990 3964 10048 3992
rect 9990 3961 10002 3964
rect 9944 3955 10002 3961
rect 10042 3952 10048 3964
rect 10100 3952 10106 4004
rect 10143 3964 11744 3992
rect 10143 3924 10171 3964
rect 11054 3924 11060 3936
rect 9876 3896 10171 3924
rect 11015 3896 11060 3924
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 11330 3924 11336 3936
rect 11291 3896 11336 3924
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 11716 3933 11744 3964
rect 12158 3952 12164 4004
rect 12216 3992 12222 4004
rect 13630 4001 13636 4004
rect 12713 3995 12771 4001
rect 12713 3992 12725 3995
rect 12216 3964 12725 3992
rect 12216 3952 12222 3964
rect 12713 3961 12725 3964
rect 12759 3961 12771 3995
rect 13624 3992 13636 4001
rect 13591 3964 13636 3992
rect 12713 3955 12771 3961
rect 13624 3955 13636 3964
rect 13630 3952 13636 3955
rect 13688 3952 13694 4004
rect 14366 3952 14372 4004
rect 14424 3992 14430 4004
rect 14734 3992 14740 4004
rect 14424 3964 14740 3992
rect 14424 3952 14430 3964
rect 14734 3952 14740 3964
rect 14792 3952 14798 4004
rect 15378 3992 15384 4004
rect 15291 3964 15384 3992
rect 15378 3952 15384 3964
rect 15436 3992 15442 4004
rect 17420 3992 17448 4023
rect 18138 4020 18144 4032
rect 18196 4020 18202 4072
rect 15436 3964 17448 3992
rect 15436 3952 15442 3964
rect 11701 3927 11759 3933
rect 11701 3893 11713 3927
rect 11747 3924 11759 3927
rect 11882 3924 11888 3936
rect 11747 3896 11888 3924
rect 11747 3893 11759 3896
rect 11701 3887 11759 3893
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 12250 3884 12256 3936
rect 12308 3924 12314 3936
rect 13722 3924 13728 3936
rect 12308 3896 13728 3924
rect 12308 3884 12314 3896
rect 13722 3884 13728 3896
rect 13780 3884 13786 3936
rect 14274 3884 14280 3936
rect 14332 3924 14338 3936
rect 14826 3924 14832 3936
rect 14332 3896 14832 3924
rect 14332 3884 14338 3896
rect 14826 3884 14832 3896
rect 14884 3884 14890 3936
rect 17586 3924 17592 3936
rect 17547 3896 17592 3924
rect 17586 3884 17592 3896
rect 17644 3884 17650 3936
rect 17770 3884 17776 3936
rect 17828 3924 17834 3936
rect 18233 3927 18291 3933
rect 18233 3924 18245 3927
rect 17828 3896 18245 3924
rect 17828 3884 17834 3896
rect 18233 3893 18245 3896
rect 18279 3893 18291 3927
rect 18233 3887 18291 3893
rect 1104 3834 18860 3856
rect 1104 3782 6912 3834
rect 6964 3782 6976 3834
rect 7028 3782 7040 3834
rect 7092 3782 7104 3834
rect 7156 3782 12843 3834
rect 12895 3782 12907 3834
rect 12959 3782 12971 3834
rect 13023 3782 13035 3834
rect 13087 3782 18860 3834
rect 1104 3760 18860 3782
rect 2685 3723 2743 3729
rect 2685 3720 2697 3723
rect 1964 3692 2697 3720
rect 1964 3593 1992 3692
rect 2685 3689 2697 3692
rect 2731 3689 2743 3723
rect 2685 3683 2743 3689
rect 2774 3680 2780 3732
rect 2832 3720 2838 3732
rect 2832 3692 2912 3720
rect 2832 3680 2838 3692
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3553 1455 3587
rect 1397 3547 1455 3553
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3553 2007 3587
rect 2884 3584 2912 3692
rect 2958 3680 2964 3732
rect 3016 3720 3022 3732
rect 3145 3723 3203 3729
rect 3145 3720 3157 3723
rect 3016 3692 3157 3720
rect 3016 3680 3022 3692
rect 3145 3689 3157 3692
rect 3191 3689 3203 3723
rect 3145 3683 3203 3689
rect 3234 3680 3240 3732
rect 3292 3720 3298 3732
rect 4065 3723 4123 3729
rect 4065 3720 4077 3723
rect 3292 3692 4077 3720
rect 3292 3680 3298 3692
rect 4065 3689 4077 3692
rect 4111 3689 4123 3723
rect 4522 3720 4528 3732
rect 4483 3692 4528 3720
rect 4065 3683 4123 3689
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 5994 3680 6000 3732
rect 6052 3720 6058 3732
rect 6638 3720 6644 3732
rect 6052 3692 6644 3720
rect 6052 3680 6058 3692
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 6825 3723 6883 3729
rect 6825 3689 6837 3723
rect 6871 3689 6883 3723
rect 6825 3683 6883 3689
rect 3050 3652 3056 3664
rect 3011 3624 3056 3652
rect 3050 3612 3056 3624
rect 3108 3612 3114 3664
rect 3694 3612 3700 3664
rect 3752 3652 3758 3664
rect 5074 3652 5080 3664
rect 3752 3624 5080 3652
rect 3752 3612 3758 3624
rect 5074 3612 5080 3624
rect 5132 3652 5138 3664
rect 5132 3624 5488 3652
rect 5132 3612 5138 3624
rect 4430 3584 4436 3596
rect 2884 3556 3280 3584
rect 4391 3556 4436 3584
rect 1949 3547 2007 3553
rect 1412 3448 1440 3547
rect 2225 3519 2283 3525
rect 2225 3485 2237 3519
rect 2271 3516 2283 3519
rect 3050 3516 3056 3528
rect 2271 3488 3056 3516
rect 2271 3485 2283 3488
rect 2225 3479 2283 3485
rect 3050 3476 3056 3488
rect 3108 3476 3114 3528
rect 3252 3525 3280 3556
rect 4430 3544 4436 3556
rect 4488 3544 4494 3596
rect 5460 3593 5488 3624
rect 5534 3612 5540 3664
rect 5592 3652 5598 3664
rect 5690 3655 5748 3661
rect 5690 3652 5702 3655
rect 5592 3624 5702 3652
rect 5592 3612 5598 3624
rect 5690 3621 5702 3624
rect 5736 3621 5748 3655
rect 5690 3615 5748 3621
rect 5810 3612 5816 3664
rect 5868 3652 5874 3664
rect 6454 3652 6460 3664
rect 5868 3624 6460 3652
rect 5868 3612 5874 3624
rect 6454 3612 6460 3624
rect 6512 3612 6518 3664
rect 6840 3652 6868 3683
rect 8018 3680 8024 3732
rect 8076 3720 8082 3732
rect 8481 3723 8539 3729
rect 8481 3720 8493 3723
rect 8076 3692 8493 3720
rect 8076 3680 8082 3692
rect 8481 3689 8493 3692
rect 8527 3689 8539 3723
rect 8481 3683 8539 3689
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 11698 3720 11704 3732
rect 10100 3692 11704 3720
rect 10100 3680 10106 3692
rect 11698 3680 11704 3692
rect 11756 3680 11762 3732
rect 11793 3723 11851 3729
rect 11793 3689 11805 3723
rect 11839 3689 11851 3723
rect 11793 3683 11851 3689
rect 13725 3723 13783 3729
rect 13725 3689 13737 3723
rect 13771 3720 13783 3723
rect 14090 3720 14096 3732
rect 13771 3692 14096 3720
rect 13771 3689 13783 3692
rect 13725 3683 13783 3689
rect 7374 3661 7380 3664
rect 7346 3655 7380 3661
rect 7346 3652 7358 3655
rect 6840 3624 7358 3652
rect 7346 3621 7358 3624
rect 7432 3652 7438 3664
rect 7432 3624 7494 3652
rect 7346 3615 7380 3621
rect 7374 3612 7380 3615
rect 7432 3612 7438 3624
rect 7558 3612 7564 3664
rect 7616 3652 7622 3664
rect 9953 3655 10011 3661
rect 9953 3652 9965 3655
rect 7616 3624 9965 3652
rect 7616 3612 7622 3624
rect 9953 3621 9965 3624
rect 9999 3621 10011 3655
rect 11808 3652 11836 3683
rect 14090 3680 14096 3692
rect 14148 3680 14154 3732
rect 14182 3680 14188 3732
rect 14240 3720 14246 3732
rect 14240 3692 17724 3720
rect 14240 3680 14246 3692
rect 12314 3655 12372 3661
rect 12314 3652 12326 3655
rect 11808 3624 12326 3652
rect 9953 3615 10011 3621
rect 12314 3621 12326 3624
rect 12360 3652 12372 3655
rect 12360 3624 15884 3652
rect 12360 3621 12372 3624
rect 12314 3615 12372 3621
rect 5445 3587 5503 3593
rect 5445 3553 5457 3587
rect 5491 3553 5503 3587
rect 5445 3547 5503 3553
rect 7101 3587 7159 3593
rect 7101 3553 7113 3587
rect 7147 3584 7159 3587
rect 7650 3584 7656 3596
rect 7147 3556 7656 3584
rect 7147 3553 7159 3556
rect 7101 3547 7159 3553
rect 7650 3544 7656 3556
rect 7708 3544 7714 3596
rect 8294 3544 8300 3596
rect 8352 3584 8358 3596
rect 8757 3587 8815 3593
rect 8757 3584 8769 3587
rect 8352 3556 8769 3584
rect 8352 3544 8358 3556
rect 8757 3553 8769 3556
rect 8803 3553 8815 3587
rect 9674 3584 9680 3596
rect 9635 3556 9680 3584
rect 8757 3547 8815 3553
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 10413 3587 10471 3593
rect 10413 3553 10425 3587
rect 10459 3584 10471 3587
rect 10502 3584 10508 3596
rect 10459 3556 10508 3584
rect 10459 3553 10471 3556
rect 10413 3547 10471 3553
rect 10502 3544 10508 3556
rect 10560 3544 10566 3596
rect 10680 3587 10738 3593
rect 10680 3553 10692 3587
rect 10726 3584 10738 3587
rect 11054 3584 11060 3596
rect 10726 3556 11060 3584
rect 10726 3553 10738 3556
rect 10680 3547 10738 3553
rect 11054 3544 11060 3556
rect 11112 3584 11118 3596
rect 13998 3584 14004 3596
rect 11112 3556 14004 3584
rect 11112 3544 11118 3556
rect 13998 3544 14004 3556
rect 14056 3544 14062 3596
rect 14090 3544 14096 3596
rect 14148 3584 14154 3596
rect 14826 3584 14832 3596
rect 14148 3556 14832 3584
rect 14148 3544 14154 3556
rect 14826 3544 14832 3556
rect 14884 3544 14890 3596
rect 14918 3544 14924 3596
rect 14976 3584 14982 3596
rect 15657 3587 15715 3593
rect 15657 3584 15669 3587
rect 14976 3556 15669 3584
rect 14976 3544 14982 3556
rect 15657 3553 15669 3556
rect 15703 3553 15715 3587
rect 15657 3547 15715 3553
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3485 3295 3519
rect 3237 3479 3295 3485
rect 4709 3519 4767 3525
rect 4709 3485 4721 3519
rect 4755 3516 4767 3519
rect 5258 3516 5264 3528
rect 4755 3488 5264 3516
rect 4755 3485 4767 3488
rect 4709 3479 4767 3485
rect 5258 3476 5264 3488
rect 5316 3476 5322 3528
rect 8941 3519 8999 3525
rect 8941 3485 8953 3519
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 4246 3448 4252 3460
rect 1412 3420 4252 3448
rect 4246 3408 4252 3420
rect 4304 3408 4310 3460
rect 1581 3383 1639 3389
rect 1581 3349 1593 3383
rect 1627 3380 1639 3383
rect 2866 3380 2872 3392
rect 1627 3352 2872 3380
rect 1627 3349 1639 3352
rect 1581 3343 1639 3349
rect 2866 3340 2872 3352
rect 2924 3340 2930 3392
rect 3234 3340 3240 3392
rect 3292 3380 3298 3392
rect 3602 3380 3608 3392
rect 3292 3352 3608 3380
rect 3292 3340 3298 3352
rect 3602 3340 3608 3352
rect 3660 3340 3666 3392
rect 6730 3340 6736 3392
rect 6788 3380 6794 3392
rect 8956 3380 8984 3479
rect 11974 3476 11980 3528
rect 12032 3516 12038 3528
rect 12069 3519 12127 3525
rect 12069 3516 12081 3519
rect 12032 3488 12081 3516
rect 12032 3476 12038 3488
rect 12069 3485 12081 3488
rect 12115 3485 12127 3519
rect 12069 3479 12127 3485
rect 14369 3519 14427 3525
rect 14369 3485 14381 3519
rect 14415 3485 14427 3519
rect 14369 3479 14427 3485
rect 13449 3451 13507 3457
rect 13449 3417 13461 3451
rect 13495 3448 13507 3451
rect 13630 3448 13636 3460
rect 13495 3420 13636 3448
rect 13495 3417 13507 3420
rect 13449 3411 13507 3417
rect 13630 3408 13636 3420
rect 13688 3448 13694 3460
rect 14384 3448 14412 3479
rect 14458 3476 14464 3528
rect 14516 3516 14522 3528
rect 15856 3525 15884 3624
rect 16574 3544 16580 3596
rect 16632 3584 16638 3596
rect 17696 3593 17724 3692
rect 17129 3587 17187 3593
rect 17129 3584 17141 3587
rect 16632 3556 17141 3584
rect 16632 3544 16638 3556
rect 17129 3553 17141 3556
rect 17175 3553 17187 3587
rect 17129 3547 17187 3553
rect 17681 3587 17739 3593
rect 17681 3553 17693 3587
rect 17727 3553 17739 3587
rect 17681 3547 17739 3553
rect 15749 3519 15807 3525
rect 15749 3516 15761 3519
rect 14516 3488 15761 3516
rect 14516 3476 14522 3488
rect 15749 3485 15761 3488
rect 15795 3485 15807 3519
rect 15749 3479 15807 3485
rect 15841 3519 15899 3525
rect 15841 3485 15853 3519
rect 15887 3485 15899 3519
rect 15841 3479 15899 3485
rect 13688 3420 14412 3448
rect 13688 3408 13694 3420
rect 15194 3408 15200 3460
rect 15252 3448 15258 3460
rect 15289 3451 15347 3457
rect 15289 3448 15301 3451
rect 15252 3420 15301 3448
rect 15252 3408 15258 3420
rect 15289 3417 15301 3420
rect 15335 3417 15347 3451
rect 15289 3411 15347 3417
rect 16482 3408 16488 3460
rect 16540 3448 16546 3460
rect 17865 3451 17923 3457
rect 17865 3448 17877 3451
rect 16540 3420 17877 3448
rect 16540 3408 16546 3420
rect 17865 3417 17877 3420
rect 17911 3417 17923 3451
rect 17865 3411 17923 3417
rect 6788 3352 8984 3380
rect 6788 3340 6794 3352
rect 11606 3340 11612 3392
rect 11664 3380 11670 3392
rect 14182 3380 14188 3392
rect 11664 3352 14188 3380
rect 11664 3340 11670 3352
rect 14182 3340 14188 3352
rect 14240 3340 14246 3392
rect 17310 3380 17316 3392
rect 17271 3352 17316 3380
rect 17310 3340 17316 3352
rect 17368 3340 17374 3392
rect 1104 3290 18860 3312
rect 1104 3238 3947 3290
rect 3999 3238 4011 3290
rect 4063 3238 4075 3290
rect 4127 3238 4139 3290
rect 4191 3238 9878 3290
rect 9930 3238 9942 3290
rect 9994 3238 10006 3290
rect 10058 3238 10070 3290
rect 10122 3238 15808 3290
rect 15860 3238 15872 3290
rect 15924 3238 15936 3290
rect 15988 3238 16000 3290
rect 16052 3238 18860 3290
rect 1104 3216 18860 3238
rect 7837 3179 7895 3185
rect 7837 3145 7849 3179
rect 7883 3176 7895 3179
rect 9122 3176 9128 3188
rect 7883 3148 9128 3176
rect 7883 3145 7895 3148
rect 7837 3139 7895 3145
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 12253 3179 12311 3185
rect 10428 3148 11468 3176
rect 2133 3111 2191 3117
rect 2133 3077 2145 3111
rect 2179 3108 2191 3111
rect 3326 3108 3332 3120
rect 2179 3080 3332 3108
rect 2179 3077 2191 3080
rect 2133 3071 2191 3077
rect 3326 3068 3332 3080
rect 3384 3068 3390 3120
rect 4338 3068 4344 3120
rect 4396 3108 4402 3120
rect 6825 3111 6883 3117
rect 4396 3080 6040 3108
rect 4396 3068 4402 3080
rect 2685 3043 2743 3049
rect 2685 3009 2697 3043
rect 2731 3040 2743 3043
rect 3418 3040 3424 3052
rect 2731 3012 3424 3040
rect 2731 3009 2743 3012
rect 2685 3003 2743 3009
rect 3418 3000 3424 3012
rect 3476 3040 3482 3052
rect 6012 3049 6040 3080
rect 6825 3077 6837 3111
rect 6871 3108 6883 3111
rect 7282 3108 7288 3120
rect 6871 3080 7288 3108
rect 6871 3077 6883 3080
rect 6825 3071 6883 3077
rect 7282 3068 7288 3080
rect 7340 3068 7346 3120
rect 3789 3043 3847 3049
rect 3789 3040 3801 3043
rect 3476 3012 3801 3040
rect 3476 3000 3482 3012
rect 3789 3009 3801 3012
rect 3835 3040 3847 3043
rect 4985 3043 5043 3049
rect 4985 3040 4997 3043
rect 3835 3012 4997 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 4985 3009 4997 3012
rect 5031 3009 5043 3043
rect 4985 3003 5043 3009
rect 5997 3043 6055 3049
rect 5997 3009 6009 3043
rect 6043 3009 6055 3043
rect 7374 3040 7380 3052
rect 7335 3012 7380 3040
rect 5997 3003 6055 3009
rect 7374 3000 7380 3012
rect 7432 3000 7438 3052
rect 8018 3000 8024 3052
rect 8076 3040 8082 3052
rect 8389 3043 8447 3049
rect 8389 3040 8401 3043
rect 8076 3012 8401 3040
rect 8076 3000 8082 3012
rect 8389 3009 8401 3012
rect 8435 3009 8447 3043
rect 9306 3040 9312 3052
rect 9267 3012 9312 3040
rect 8389 3003 8447 3009
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 9490 3040 9496 3052
rect 9451 3012 9496 3040
rect 9490 3000 9496 3012
rect 9548 3040 9554 3052
rect 10428 3040 10456 3148
rect 10873 3111 10931 3117
rect 10873 3077 10885 3111
rect 10919 3108 10931 3111
rect 11330 3108 11336 3120
rect 10919 3080 11336 3108
rect 10919 3077 10931 3080
rect 10873 3071 10931 3077
rect 11330 3068 11336 3080
rect 11388 3068 11394 3120
rect 10597 3043 10655 3049
rect 10597 3040 10609 3043
rect 9548 3012 10609 3040
rect 9548 3000 9554 3012
rect 10597 3009 10609 3012
rect 10643 3009 10655 3043
rect 10597 3003 10655 3009
rect 11146 3000 11152 3052
rect 11204 3000 11210 3052
rect 11440 3040 11468 3148
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 14274 3176 14280 3188
rect 12299 3148 14280 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 14458 3176 14464 3188
rect 14419 3148 14464 3176
rect 14458 3136 14464 3148
rect 14516 3136 14522 3188
rect 14734 3136 14740 3188
rect 14792 3176 14798 3188
rect 14792 3148 18092 3176
rect 14792 3136 14798 3148
rect 12437 3111 12495 3117
rect 12437 3077 12449 3111
rect 12483 3108 12495 3111
rect 14918 3108 14924 3120
rect 12483 3080 14924 3108
rect 12483 3077 12495 3080
rect 12437 3071 12495 3077
rect 14918 3068 14924 3080
rect 14976 3068 14982 3120
rect 15562 3068 15568 3120
rect 15620 3108 15626 3120
rect 15620 3080 16988 3108
rect 15620 3068 15626 3080
rect 11609 3043 11667 3049
rect 11609 3040 11621 3043
rect 11440 3012 11621 3040
rect 11609 3009 11621 3012
rect 11655 3009 11667 3043
rect 11609 3003 11667 3009
rect 11698 3000 11704 3052
rect 11756 3040 11762 3052
rect 13081 3043 13139 3049
rect 13081 3040 13093 3043
rect 11756 3012 13093 3040
rect 11756 3000 11762 3012
rect 13081 3009 13093 3012
rect 13127 3040 13139 3043
rect 13446 3040 13452 3052
rect 13127 3012 13452 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 13446 3000 13452 3012
rect 13504 3040 13510 3052
rect 13906 3040 13912 3052
rect 13504 3012 13912 3040
rect 13504 3000 13510 3012
rect 13906 3000 13912 3012
rect 13964 3040 13970 3052
rect 14001 3043 14059 3049
rect 14001 3040 14013 3043
rect 13964 3012 14013 3040
rect 13964 3000 13970 3012
rect 14001 3009 14013 3012
rect 14047 3009 14059 3043
rect 14001 3003 14059 3009
rect 14090 3000 14096 3052
rect 14148 3040 14154 3052
rect 15013 3043 15071 3049
rect 15013 3040 15025 3043
rect 14148 3012 15025 3040
rect 14148 3000 14154 3012
rect 15013 3009 15025 3012
rect 15059 3009 15071 3043
rect 15657 3043 15715 3049
rect 15657 3040 15669 3043
rect 15013 3003 15071 3009
rect 15120 3012 15669 3040
rect 1394 2972 1400 2984
rect 1355 2944 1400 2972
rect 1394 2932 1400 2944
rect 1452 2932 1458 2984
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2972 1731 2975
rect 2130 2972 2136 2984
rect 1719 2944 2136 2972
rect 1719 2941 1731 2944
rect 1673 2935 1731 2941
rect 2130 2932 2136 2944
rect 2188 2932 2194 2984
rect 2406 2932 2412 2984
rect 2464 2972 2470 2984
rect 3605 2975 3663 2981
rect 3605 2972 3617 2975
rect 2464 2944 3617 2972
rect 2464 2932 2470 2944
rect 3605 2941 3617 2944
rect 3651 2941 3663 2975
rect 4798 2972 4804 2984
rect 4759 2944 4804 2972
rect 3605 2935 3663 2941
rect 4798 2932 4804 2944
rect 4856 2932 4862 2984
rect 4893 2975 4951 2981
rect 4893 2941 4905 2975
rect 4939 2972 4951 2975
rect 5442 2972 5448 2984
rect 4939 2944 5448 2972
rect 4939 2941 4951 2944
rect 4893 2935 4951 2941
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 5813 2975 5871 2981
rect 5813 2941 5825 2975
rect 5859 2972 5871 2975
rect 6270 2972 6276 2984
rect 5859 2944 6276 2972
rect 5859 2941 5871 2944
rect 5813 2935 5871 2941
rect 6270 2932 6276 2944
rect 6328 2932 6334 2984
rect 7193 2975 7251 2981
rect 7193 2941 7205 2975
rect 7239 2972 7251 2975
rect 7466 2972 7472 2984
rect 7239 2944 7472 2972
rect 7239 2941 7251 2944
rect 7193 2935 7251 2941
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 7834 2932 7840 2984
rect 7892 2972 7898 2984
rect 8110 2972 8116 2984
rect 7892 2944 8116 2972
rect 7892 2932 7898 2944
rect 8110 2932 8116 2944
rect 8168 2972 8174 2984
rect 8297 2975 8355 2981
rect 8297 2972 8309 2975
rect 8168 2944 8309 2972
rect 8168 2932 8174 2944
rect 8297 2941 8309 2944
rect 8343 2941 8355 2975
rect 8297 2935 8355 2941
rect 1946 2864 1952 2916
rect 2004 2904 2010 2916
rect 2501 2907 2559 2913
rect 2501 2904 2513 2907
rect 2004 2876 2513 2904
rect 2004 2864 2010 2876
rect 2501 2873 2513 2876
rect 2547 2873 2559 2907
rect 2501 2867 2559 2873
rect 2593 2907 2651 2913
rect 2593 2873 2605 2907
rect 2639 2904 2651 2907
rect 2682 2904 2688 2916
rect 2639 2876 2688 2904
rect 2639 2873 2651 2876
rect 2593 2867 2651 2873
rect 2682 2864 2688 2876
rect 2740 2864 2746 2916
rect 3513 2907 3571 2913
rect 3513 2873 3525 2907
rect 3559 2904 3571 2907
rect 3878 2904 3884 2916
rect 3559 2876 3884 2904
rect 3559 2873 3571 2876
rect 3513 2867 3571 2873
rect 3878 2864 3884 2876
rect 3936 2864 3942 2916
rect 5905 2907 5963 2913
rect 5905 2904 5917 2907
rect 4448 2876 5917 2904
rect 1394 2796 1400 2848
rect 1452 2836 1458 2848
rect 1762 2836 1768 2848
rect 1452 2808 1768 2836
rect 1452 2796 1458 2808
rect 1762 2796 1768 2808
rect 1820 2796 1826 2848
rect 3142 2836 3148 2848
rect 3103 2808 3148 2836
rect 3142 2796 3148 2808
rect 3200 2796 3206 2848
rect 4448 2845 4476 2876
rect 5905 2873 5917 2876
rect 5951 2873 5963 2907
rect 5905 2867 5963 2873
rect 5994 2864 6000 2916
rect 6052 2904 6058 2916
rect 7285 2907 7343 2913
rect 7285 2904 7297 2907
rect 6052 2876 7297 2904
rect 6052 2864 6058 2876
rect 7285 2873 7297 2876
rect 7331 2873 7343 2907
rect 7285 2867 7343 2873
rect 9306 2864 9312 2916
rect 9364 2904 9370 2916
rect 9508 2904 9536 3000
rect 10413 2975 10471 2981
rect 10413 2941 10425 2975
rect 10459 2972 10471 2975
rect 11164 2972 11192 3000
rect 10459 2944 11192 2972
rect 11425 2975 11483 2981
rect 10459 2941 10471 2944
rect 10413 2935 10471 2941
rect 11425 2941 11437 2975
rect 11471 2972 11483 2975
rect 11790 2972 11796 2984
rect 11471 2944 11796 2972
rect 11471 2941 11483 2944
rect 11425 2935 11483 2941
rect 11790 2932 11796 2944
rect 11848 2932 11854 2984
rect 13814 2932 13820 2984
rect 13872 2972 13878 2984
rect 13872 2944 14136 2972
rect 13872 2932 13878 2944
rect 9364 2876 9536 2904
rect 10505 2907 10563 2913
rect 9364 2864 9370 2876
rect 10505 2873 10517 2907
rect 10551 2904 10563 2907
rect 10873 2907 10931 2913
rect 10873 2904 10885 2907
rect 10551 2876 10885 2904
rect 10551 2873 10563 2876
rect 10505 2867 10563 2873
rect 10873 2873 10885 2876
rect 10919 2873 10931 2907
rect 10873 2867 10931 2873
rect 11146 2864 11152 2916
rect 11204 2904 11210 2916
rect 12897 2907 12955 2913
rect 12897 2904 12909 2907
rect 11204 2876 12909 2904
rect 11204 2864 11210 2876
rect 12897 2873 12909 2876
rect 12943 2873 12955 2907
rect 13998 2904 14004 2916
rect 12897 2867 12955 2873
rect 13464 2876 14004 2904
rect 4433 2839 4491 2845
rect 4433 2805 4445 2839
rect 4479 2805 4491 2839
rect 5442 2836 5448 2848
rect 5403 2808 5448 2836
rect 4433 2799 4491 2805
rect 5442 2796 5448 2808
rect 5500 2796 5506 2848
rect 6362 2796 6368 2848
rect 6420 2836 6426 2848
rect 8205 2839 8263 2845
rect 8205 2836 8217 2839
rect 6420 2808 8217 2836
rect 6420 2796 6426 2808
rect 8205 2805 8217 2808
rect 8251 2805 8263 2839
rect 8846 2836 8852 2848
rect 8807 2808 8852 2836
rect 8205 2799 8263 2805
rect 8846 2796 8852 2808
rect 8904 2796 8910 2848
rect 9217 2839 9275 2845
rect 9217 2805 9229 2839
rect 9263 2836 9275 2839
rect 9582 2836 9588 2848
rect 9263 2808 9588 2836
rect 9263 2805 9275 2808
rect 9217 2799 9275 2805
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 10042 2836 10048 2848
rect 10003 2808 10048 2836
rect 10042 2796 10048 2808
rect 10100 2796 10106 2848
rect 11054 2836 11060 2848
rect 11015 2808 11060 2836
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 11517 2839 11575 2845
rect 11517 2805 11529 2839
rect 11563 2836 11575 2839
rect 12253 2839 12311 2845
rect 12253 2836 12265 2839
rect 11563 2808 12265 2836
rect 11563 2805 11575 2808
rect 11517 2799 11575 2805
rect 12253 2805 12265 2808
rect 12299 2805 12311 2839
rect 12253 2799 12311 2805
rect 12805 2839 12863 2845
rect 12805 2805 12817 2839
rect 12851 2836 12863 2839
rect 13262 2836 13268 2848
rect 12851 2808 13268 2836
rect 12851 2805 12863 2808
rect 12805 2799 12863 2805
rect 13262 2796 13268 2808
rect 13320 2796 13326 2848
rect 13464 2845 13492 2876
rect 13998 2864 14004 2876
rect 14056 2864 14062 2916
rect 14108 2904 14136 2944
rect 14182 2932 14188 2984
rect 14240 2972 14246 2984
rect 14734 2972 14740 2984
rect 14240 2944 14740 2972
rect 14240 2932 14246 2944
rect 14734 2932 14740 2944
rect 14792 2932 14798 2984
rect 14826 2932 14832 2984
rect 14884 2972 14890 2984
rect 15120 2972 15148 3012
rect 15657 3009 15669 3012
rect 15703 3009 15715 3043
rect 15657 3003 15715 3009
rect 15470 2972 15476 2984
rect 14884 2944 15148 2972
rect 15431 2944 15476 2972
rect 14884 2932 14890 2944
rect 15470 2932 15476 2944
rect 15528 2932 15534 2984
rect 15562 2932 15568 2984
rect 15620 2972 15626 2984
rect 16960 2981 16988 3080
rect 18064 2981 18092 3148
rect 16393 2975 16451 2981
rect 16393 2972 16405 2975
rect 15620 2944 16405 2972
rect 15620 2932 15626 2944
rect 16393 2941 16405 2944
rect 16439 2941 16451 2975
rect 16393 2935 16451 2941
rect 16945 2975 17003 2981
rect 16945 2941 16957 2975
rect 16991 2941 17003 2975
rect 16945 2935 17003 2941
rect 18049 2975 18107 2981
rect 18049 2941 18061 2975
rect 18095 2941 18107 2975
rect 18049 2935 18107 2941
rect 14918 2904 14924 2916
rect 14108 2876 14780 2904
rect 14879 2876 14924 2904
rect 13449 2839 13507 2845
rect 13449 2805 13461 2839
rect 13495 2805 13507 2839
rect 13449 2799 13507 2805
rect 13722 2796 13728 2848
rect 13780 2836 13786 2848
rect 13817 2839 13875 2845
rect 13817 2836 13829 2839
rect 13780 2808 13829 2836
rect 13780 2796 13786 2808
rect 13817 2805 13829 2808
rect 13863 2805 13875 2839
rect 13817 2799 13875 2805
rect 13909 2839 13967 2845
rect 13909 2805 13921 2839
rect 13955 2836 13967 2839
rect 14642 2836 14648 2848
rect 13955 2808 14648 2836
rect 13955 2805 13967 2808
rect 13909 2799 13967 2805
rect 14642 2796 14648 2808
rect 14700 2796 14706 2848
rect 14752 2836 14780 2876
rect 14918 2864 14924 2876
rect 14976 2864 14982 2916
rect 16666 2904 16672 2916
rect 16408 2876 16672 2904
rect 16408 2848 16436 2876
rect 16666 2864 16672 2876
rect 16724 2864 16730 2916
rect 14829 2839 14887 2845
rect 14829 2836 14841 2839
rect 14752 2808 14841 2836
rect 14829 2805 14841 2808
rect 14875 2805 14887 2839
rect 14829 2799 14887 2805
rect 16390 2796 16396 2848
rect 16448 2796 16454 2848
rect 16574 2836 16580 2848
rect 16535 2808 16580 2836
rect 16574 2796 16580 2808
rect 16632 2796 16638 2848
rect 17129 2839 17187 2845
rect 17129 2805 17141 2839
rect 17175 2836 17187 2839
rect 17218 2836 17224 2848
rect 17175 2808 17224 2836
rect 17175 2805 17187 2808
rect 17129 2799 17187 2805
rect 17218 2796 17224 2808
rect 17276 2796 17282 2848
rect 18230 2836 18236 2848
rect 18191 2808 18236 2836
rect 18230 2796 18236 2808
rect 18288 2796 18294 2848
rect 1104 2746 18860 2768
rect 1104 2694 6912 2746
rect 6964 2694 6976 2746
rect 7028 2694 7040 2746
rect 7092 2694 7104 2746
rect 7156 2694 12843 2746
rect 12895 2694 12907 2746
rect 12959 2694 12971 2746
rect 13023 2694 13035 2746
rect 13087 2694 18860 2746
rect 1104 2672 18860 2694
rect 3326 2632 3332 2644
rect 3287 2604 3332 2632
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 4065 2635 4123 2641
rect 4065 2601 4077 2635
rect 4111 2632 4123 2635
rect 4430 2632 4436 2644
rect 4111 2604 4436 2632
rect 4111 2601 4123 2604
rect 4065 2595 4123 2601
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 4525 2635 4583 2641
rect 4525 2601 4537 2635
rect 4571 2601 4583 2635
rect 4525 2595 4583 2601
rect 4893 2635 4951 2641
rect 4893 2601 4905 2635
rect 4939 2632 4951 2635
rect 5442 2632 5448 2644
rect 4939 2604 5448 2632
rect 4939 2601 4951 2604
rect 4893 2595 4951 2601
rect 3142 2524 3148 2576
rect 3200 2564 3206 2576
rect 3421 2567 3479 2573
rect 3421 2564 3433 2567
rect 3200 2536 3433 2564
rect 3200 2524 3206 2536
rect 3421 2533 3433 2536
rect 3467 2533 3479 2567
rect 4540 2564 4568 2595
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 8665 2635 8723 2641
rect 8665 2632 8677 2635
rect 8067 2604 8677 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 8665 2601 8677 2604
rect 8711 2601 8723 2635
rect 9030 2632 9036 2644
rect 8991 2604 9036 2632
rect 8665 2595 8723 2601
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 10137 2635 10195 2641
rect 10137 2601 10149 2635
rect 10183 2632 10195 2635
rect 11054 2632 11060 2644
rect 10183 2604 11060 2632
rect 10183 2601 10195 2604
rect 10137 2595 10195 2601
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 11149 2635 11207 2641
rect 11149 2601 11161 2635
rect 11195 2632 11207 2635
rect 12342 2632 12348 2644
rect 11195 2604 12348 2632
rect 11195 2601 11207 2604
rect 11149 2595 11207 2601
rect 12342 2592 12348 2604
rect 12400 2592 12406 2644
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 12989 2635 13047 2641
rect 12989 2632 13001 2635
rect 12492 2604 13001 2632
rect 12492 2592 12498 2604
rect 12989 2601 13001 2604
rect 13035 2632 13047 2635
rect 13354 2632 13360 2644
rect 13035 2604 13360 2632
rect 13035 2601 13047 2604
rect 12989 2595 13047 2601
rect 13354 2592 13360 2604
rect 13412 2592 13418 2644
rect 13633 2635 13691 2641
rect 13633 2601 13645 2635
rect 13679 2601 13691 2635
rect 13998 2632 14004 2644
rect 13959 2604 14004 2632
rect 13633 2595 13691 2601
rect 5994 2564 6000 2576
rect 4540 2536 6000 2564
rect 3421 2527 3479 2533
rect 5994 2524 6000 2536
rect 6052 2524 6058 2576
rect 6365 2567 6423 2573
rect 6365 2533 6377 2567
rect 6411 2564 6423 2567
rect 6546 2564 6552 2576
rect 6411 2536 6552 2564
rect 6411 2533 6423 2536
rect 6365 2527 6423 2533
rect 6546 2524 6552 2536
rect 6604 2524 6610 2576
rect 8113 2567 8171 2573
rect 8113 2533 8125 2567
rect 8159 2564 8171 2567
rect 8846 2564 8852 2576
rect 8159 2536 8852 2564
rect 8159 2533 8171 2536
rect 8113 2527 8171 2533
rect 8846 2524 8852 2536
rect 8904 2524 8910 2576
rect 10042 2524 10048 2576
rect 10100 2564 10106 2576
rect 10229 2567 10287 2573
rect 10229 2564 10241 2567
rect 10100 2536 10241 2564
rect 10100 2524 10106 2536
rect 10229 2533 10241 2536
rect 10275 2533 10287 2567
rect 10229 2527 10287 2533
rect 10318 2524 10324 2576
rect 10376 2564 10382 2576
rect 12069 2567 12127 2573
rect 12069 2564 12081 2567
rect 10376 2536 12081 2564
rect 10376 2524 10382 2536
rect 12069 2533 12081 2536
rect 12115 2533 12127 2567
rect 13078 2564 13084 2576
rect 13039 2536 13084 2564
rect 12069 2527 12127 2533
rect 13078 2524 13084 2536
rect 13136 2524 13142 2576
rect 13538 2564 13544 2576
rect 13188 2536 13544 2564
rect 1394 2456 1400 2508
rect 1452 2496 1458 2508
rect 1581 2499 1639 2505
rect 1581 2496 1593 2499
rect 1452 2468 1593 2496
rect 1452 2456 1458 2468
rect 1581 2465 1593 2468
rect 1627 2465 1639 2499
rect 1581 2459 1639 2465
rect 2409 2499 2467 2505
rect 2409 2465 2421 2499
rect 2455 2496 2467 2499
rect 3878 2496 3884 2508
rect 2455 2468 3884 2496
rect 2455 2465 2467 2468
rect 2409 2459 2467 2465
rect 3878 2456 3884 2468
rect 3936 2456 3942 2508
rect 5718 2496 5724 2508
rect 5679 2468 5724 2496
rect 5718 2456 5724 2468
rect 5776 2456 5782 2508
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 7282 2496 7288 2508
rect 6963 2468 7288 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 7282 2456 7288 2468
rect 7340 2456 7346 2508
rect 8662 2456 8668 2508
rect 8720 2496 8726 2508
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 8720 2468 9137 2496
rect 8720 2456 8726 2468
rect 9125 2465 9137 2468
rect 9171 2465 9183 2499
rect 9125 2459 9183 2465
rect 10962 2456 10968 2508
rect 11020 2496 11026 2508
rect 11020 2468 11376 2496
rect 11020 2456 11026 2468
rect 1210 2388 1216 2440
rect 1268 2428 1274 2440
rect 1765 2431 1823 2437
rect 1765 2428 1777 2431
rect 1268 2400 1777 2428
rect 1268 2388 1274 2400
rect 1765 2397 1777 2400
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2428 3663 2431
rect 4338 2428 4344 2440
rect 3651 2400 4344 2428
rect 3651 2397 3663 2400
rect 3605 2391 3663 2397
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2397 5043 2431
rect 4985 2391 5043 2397
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2428 5227 2431
rect 5534 2428 5540 2440
rect 5215 2400 5540 2428
rect 5215 2397 5227 2400
rect 5169 2391 5227 2397
rect 2961 2363 3019 2369
rect 2961 2329 2973 2363
rect 3007 2360 3019 2363
rect 5000 2360 5028 2391
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 5626 2388 5632 2440
rect 5684 2428 5690 2440
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 5684 2400 7113 2428
rect 5684 2388 5690 2400
rect 7101 2397 7113 2400
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 8205 2431 8263 2437
rect 8205 2397 8217 2431
rect 8251 2397 8263 2431
rect 9306 2428 9312 2440
rect 9267 2400 9312 2428
rect 8205 2391 8263 2397
rect 3007 2332 5028 2360
rect 8220 2360 8248 2391
rect 9306 2388 9312 2400
rect 9364 2388 9370 2440
rect 11348 2437 11376 2468
rect 11422 2456 11428 2508
rect 11480 2496 11486 2508
rect 11793 2499 11851 2505
rect 11793 2496 11805 2499
rect 11480 2468 11805 2496
rect 11480 2456 11486 2468
rect 11793 2465 11805 2468
rect 11839 2465 11851 2499
rect 11793 2459 11851 2465
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 11241 2431 11299 2437
rect 11241 2397 11253 2431
rect 11287 2397 11299 2431
rect 11241 2391 11299 2397
rect 11333 2431 11391 2437
rect 11333 2397 11345 2431
rect 11379 2397 11391 2431
rect 13188 2428 13216 2536
rect 13538 2524 13544 2536
rect 13596 2524 13602 2576
rect 13648 2564 13676 2595
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 14093 2635 14151 2641
rect 14093 2601 14105 2635
rect 14139 2632 14151 2635
rect 15286 2632 15292 2644
rect 14139 2604 15292 2632
rect 14139 2601 14151 2604
rect 14093 2595 14151 2601
rect 15286 2592 15292 2604
rect 15344 2592 15350 2644
rect 14366 2564 14372 2576
rect 13648 2536 14372 2564
rect 14366 2524 14372 2536
rect 14424 2524 14430 2576
rect 16390 2564 16396 2576
rect 15488 2536 16396 2564
rect 13630 2456 13636 2508
rect 13688 2496 13694 2508
rect 13688 2468 14320 2496
rect 13688 2456 13694 2468
rect 11333 2391 11391 2397
rect 12544 2400 13216 2428
rect 13265 2431 13323 2437
rect 8754 2360 8760 2372
rect 8220 2332 8760 2360
rect 3007 2329 3019 2332
rect 2961 2323 3019 2329
rect 8754 2320 8760 2332
rect 8812 2360 8818 2372
rect 10336 2360 10364 2391
rect 8812 2332 10364 2360
rect 10781 2363 10839 2369
rect 8812 2320 8818 2332
rect 10781 2329 10793 2363
rect 10827 2360 10839 2363
rect 11146 2360 11152 2372
rect 10827 2332 11152 2360
rect 10827 2329 10839 2332
rect 10781 2323 10839 2329
rect 11146 2320 11152 2332
rect 11204 2320 11210 2372
rect 2593 2295 2651 2301
rect 2593 2261 2605 2295
rect 2639 2292 2651 2295
rect 2774 2292 2780 2304
rect 2639 2264 2780 2292
rect 2639 2261 2651 2264
rect 2593 2255 2651 2261
rect 2774 2252 2780 2264
rect 2832 2252 2838 2304
rect 7650 2292 7656 2304
rect 7611 2264 7656 2292
rect 7650 2252 7656 2264
rect 7708 2252 7714 2304
rect 9769 2295 9827 2301
rect 9769 2261 9781 2295
rect 9815 2292 9827 2295
rect 10410 2292 10416 2304
rect 9815 2264 10416 2292
rect 9815 2261 9827 2264
rect 9769 2255 9827 2261
rect 10410 2252 10416 2264
rect 10468 2252 10474 2304
rect 11256 2292 11284 2391
rect 12544 2292 12572 2400
rect 13265 2397 13277 2431
rect 13311 2428 13323 2431
rect 13446 2428 13452 2440
rect 13311 2400 13452 2428
rect 13311 2397 13323 2400
rect 13265 2391 13323 2397
rect 13446 2388 13452 2400
rect 13504 2388 13510 2440
rect 14182 2428 14188 2440
rect 14143 2400 14188 2428
rect 14182 2388 14188 2400
rect 14240 2388 14246 2440
rect 14292 2428 14320 2468
rect 14550 2456 14556 2508
rect 14608 2496 14614 2508
rect 15488 2505 15516 2536
rect 16390 2524 16396 2536
rect 16448 2524 16454 2576
rect 14645 2499 14703 2505
rect 14645 2496 14657 2499
rect 14608 2468 14657 2496
rect 14608 2456 14614 2468
rect 14645 2465 14657 2468
rect 14691 2465 14703 2499
rect 14645 2459 14703 2465
rect 15473 2499 15531 2505
rect 15473 2465 15485 2499
rect 15519 2465 15531 2499
rect 16206 2496 16212 2508
rect 16167 2468 16212 2496
rect 15473 2459 15531 2465
rect 16206 2456 16212 2468
rect 16264 2456 16270 2508
rect 16666 2456 16672 2508
rect 16724 2496 16730 2508
rect 16945 2499 17003 2505
rect 16945 2496 16957 2499
rect 16724 2468 16957 2496
rect 16724 2456 16730 2468
rect 16945 2465 16957 2468
rect 16991 2496 17003 2499
rect 17126 2496 17132 2508
rect 16991 2468 17132 2496
rect 16991 2465 17003 2468
rect 16945 2459 17003 2465
rect 17126 2456 17132 2468
rect 17184 2456 17190 2508
rect 17678 2496 17684 2508
rect 17639 2468 17684 2496
rect 17678 2456 17684 2468
rect 17736 2456 17742 2508
rect 14829 2431 14887 2437
rect 14829 2428 14841 2431
rect 14292 2400 14841 2428
rect 14829 2397 14841 2400
rect 14875 2397 14887 2431
rect 14829 2391 14887 2397
rect 15197 2431 15255 2437
rect 15197 2397 15209 2431
rect 15243 2428 15255 2431
rect 15657 2431 15715 2437
rect 15657 2428 15669 2431
rect 15243 2400 15669 2428
rect 15243 2397 15255 2400
rect 15197 2391 15255 2397
rect 15657 2397 15669 2400
rect 15703 2397 15715 2431
rect 15657 2391 15715 2397
rect 16393 2431 16451 2437
rect 16393 2397 16405 2431
rect 16439 2397 16451 2431
rect 16393 2391 16451 2397
rect 12621 2363 12679 2369
rect 12621 2329 12633 2363
rect 12667 2360 12679 2363
rect 13814 2360 13820 2372
rect 12667 2332 13820 2360
rect 12667 2329 12679 2332
rect 12621 2323 12679 2329
rect 13814 2320 13820 2332
rect 13872 2320 13878 2372
rect 13906 2320 13912 2372
rect 13964 2360 13970 2372
rect 16408 2360 16436 2391
rect 13964 2332 16436 2360
rect 13964 2320 13970 2332
rect 11256 2264 12572 2292
rect 13078 2252 13084 2304
rect 13136 2292 13142 2304
rect 15197 2295 15255 2301
rect 15197 2292 15209 2295
rect 13136 2264 15209 2292
rect 13136 2252 13142 2264
rect 15197 2261 15209 2264
rect 15243 2261 15255 2295
rect 17126 2292 17132 2304
rect 17087 2264 17132 2292
rect 15197 2255 15255 2261
rect 17126 2252 17132 2264
rect 17184 2252 17190 2304
rect 17862 2292 17868 2304
rect 17823 2264 17868 2292
rect 17862 2252 17868 2264
rect 17920 2252 17926 2304
rect 1104 2202 18860 2224
rect 1104 2150 3947 2202
rect 3999 2150 4011 2202
rect 4063 2150 4075 2202
rect 4127 2150 4139 2202
rect 4191 2150 9878 2202
rect 9930 2150 9942 2202
rect 9994 2150 10006 2202
rect 10058 2150 10070 2202
rect 10122 2150 15808 2202
rect 15860 2150 15872 2202
rect 15924 2150 15936 2202
rect 15988 2150 16000 2202
rect 16052 2150 18860 2202
rect 1104 2128 18860 2150
rect 382 2048 388 2100
rect 440 2088 446 2100
rect 17126 2088 17132 2100
rect 440 2060 17132 2088
rect 440 2048 446 2060
rect 17126 2048 17132 2060
rect 17184 2048 17190 2100
rect 7650 1912 7656 1964
rect 7708 1952 7714 1964
rect 7708 1924 12572 1952
rect 7708 1912 7714 1924
rect 12544 1816 12572 1924
rect 16298 1816 16304 1828
rect 12544 1788 16304 1816
rect 16298 1776 16304 1788
rect 16356 1776 16362 1828
rect 3970 1368 3976 1420
rect 4028 1408 4034 1420
rect 5626 1408 5632 1420
rect 4028 1380 5632 1408
rect 4028 1368 4034 1380
rect 5626 1368 5632 1380
rect 5684 1368 5690 1420
rect 11238 1368 11244 1420
rect 11296 1408 11302 1420
rect 13630 1408 13636 1420
rect 11296 1380 13636 1408
rect 11296 1368 11302 1380
rect 13630 1368 13636 1380
rect 13688 1368 13694 1420
<< via1 >>
rect 3976 15308 4028 15360
rect 6368 15308 6420 15360
rect 4068 15240 4120 15292
rect 8852 15240 8904 15292
rect 3516 14968 3568 15020
rect 6276 14968 6328 15020
rect 9036 14832 9088 14884
rect 18236 14832 18288 14884
rect 3700 14764 3752 14816
rect 11520 14764 11572 14816
rect 6912 14662 6964 14714
rect 6976 14662 7028 14714
rect 7040 14662 7092 14714
rect 7104 14662 7156 14714
rect 12843 14662 12895 14714
rect 12907 14662 12959 14714
rect 12971 14662 13023 14714
rect 13035 14662 13087 14714
rect 3792 14492 3844 14544
rect 8576 14492 8628 14544
rect 15476 14560 15528 14612
rect 11336 14492 11388 14544
rect 14372 14492 14424 14544
rect 8668 14424 8720 14476
rect 9588 14424 9640 14476
rect 11428 14424 11480 14476
rect 11980 14424 12032 14476
rect 12440 14424 12492 14476
rect 14740 14467 14792 14476
rect 14740 14433 14749 14467
rect 14749 14433 14783 14467
rect 14783 14433 14792 14467
rect 14740 14424 14792 14433
rect 8208 14399 8260 14408
rect 8208 14365 8217 14399
rect 8217 14365 8251 14399
rect 8251 14365 8260 14399
rect 8208 14356 8260 14365
rect 10600 14399 10652 14408
rect 10600 14365 10609 14399
rect 10609 14365 10643 14399
rect 10643 14365 10652 14399
rect 10600 14356 10652 14365
rect 10784 14399 10836 14408
rect 10784 14365 10793 14399
rect 10793 14365 10827 14399
rect 10827 14365 10836 14399
rect 10784 14356 10836 14365
rect 11060 14356 11112 14408
rect 12532 14356 12584 14408
rect 14924 14399 14976 14408
rect 13728 14288 13780 14340
rect 14924 14365 14933 14399
rect 14933 14365 14967 14399
rect 14967 14365 14976 14399
rect 14924 14356 14976 14365
rect 14188 14288 14240 14340
rect 15108 14424 15160 14476
rect 18788 14492 18840 14544
rect 15660 14356 15712 14408
rect 5724 14220 5776 14272
rect 9772 14220 9824 14272
rect 11152 14263 11204 14272
rect 11152 14229 11161 14263
rect 11161 14229 11195 14263
rect 11195 14229 11204 14263
rect 11152 14220 11204 14229
rect 13544 14220 13596 14272
rect 16212 14220 16264 14272
rect 3947 14118 3999 14170
rect 4011 14118 4063 14170
rect 4075 14118 4127 14170
rect 4139 14118 4191 14170
rect 9878 14118 9930 14170
rect 9942 14118 9994 14170
rect 10006 14118 10058 14170
rect 10070 14118 10122 14170
rect 15808 14118 15860 14170
rect 15872 14118 15924 14170
rect 15936 14118 15988 14170
rect 16000 14118 16052 14170
rect 3424 14016 3476 14068
rect 3332 13948 3384 14000
rect 8300 13948 8352 14000
rect 8668 14016 8720 14068
rect 9588 14059 9640 14068
rect 9588 14025 9597 14059
rect 9597 14025 9631 14059
rect 9631 14025 9640 14059
rect 9588 14016 9640 14025
rect 10600 14059 10652 14068
rect 10600 14025 10609 14059
rect 10609 14025 10643 14059
rect 10643 14025 10652 14059
rect 10600 14016 10652 14025
rect 12072 14016 12124 14068
rect 5448 13880 5500 13932
rect 8760 13880 8812 13932
rect 8944 13880 8996 13932
rect 9680 13880 9732 13932
rect 10784 13880 10836 13932
rect 10876 13880 10928 13932
rect 12164 13880 12216 13932
rect 14372 13880 14424 13932
rect 15936 13880 15988 13932
rect 16580 13880 16632 13932
rect 17132 13923 17184 13932
rect 17132 13889 17141 13923
rect 17141 13889 17175 13923
rect 17175 13889 17184 13923
rect 17132 13880 17184 13889
rect 8116 13812 8168 13864
rect 8668 13744 8720 13796
rect 9312 13812 9364 13864
rect 10508 13812 10560 13864
rect 11612 13855 11664 13864
rect 11612 13821 11621 13855
rect 11621 13821 11655 13855
rect 11655 13821 11664 13855
rect 11612 13812 11664 13821
rect 13176 13812 13228 13864
rect 13452 13855 13504 13864
rect 13452 13821 13461 13855
rect 13461 13821 13495 13855
rect 13495 13821 13504 13855
rect 13452 13812 13504 13821
rect 17408 13855 17460 13864
rect 10232 13744 10284 13796
rect 17408 13821 17417 13855
rect 17417 13821 17451 13855
rect 17451 13821 17460 13855
rect 17408 13812 17460 13821
rect 18512 13948 18564 14000
rect 15568 13744 15620 13796
rect 16212 13787 16264 13796
rect 16212 13753 16221 13787
rect 16221 13753 16255 13787
rect 16255 13753 16264 13787
rect 16212 13744 16264 13753
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 5632 13719 5684 13728
rect 5632 13685 5641 13719
rect 5641 13685 5675 13719
rect 5675 13685 5684 13719
rect 5632 13676 5684 13685
rect 6368 13676 6420 13728
rect 9496 13676 9548 13728
rect 9956 13719 10008 13728
rect 9956 13685 9965 13719
rect 9965 13685 9999 13719
rect 9999 13685 10008 13719
rect 9956 13676 10008 13685
rect 10324 13676 10376 13728
rect 10600 13676 10652 13728
rect 11244 13676 11296 13728
rect 11704 13676 11756 13728
rect 13912 13676 13964 13728
rect 15200 13676 15252 13728
rect 17592 13719 17644 13728
rect 17592 13685 17601 13719
rect 17601 13685 17635 13719
rect 17635 13685 17644 13719
rect 17592 13676 17644 13685
rect 6912 13574 6964 13626
rect 6976 13574 7028 13626
rect 7040 13574 7092 13626
rect 7104 13574 7156 13626
rect 12843 13574 12895 13626
rect 12907 13574 12959 13626
rect 12971 13574 13023 13626
rect 13035 13574 13087 13626
rect 5540 13472 5592 13524
rect 5080 13336 5132 13388
rect 6460 13336 6512 13388
rect 4068 13268 4120 13320
rect 5816 13268 5868 13320
rect 6184 13268 6236 13320
rect 8576 13515 8628 13524
rect 8576 13481 8585 13515
rect 8585 13481 8619 13515
rect 8619 13481 8628 13515
rect 8576 13472 8628 13481
rect 8944 13472 8996 13524
rect 9956 13472 10008 13524
rect 11244 13472 11296 13524
rect 12532 13472 12584 13524
rect 7840 13404 7892 13456
rect 11888 13404 11940 13456
rect 14648 13447 14700 13456
rect 7472 13336 7524 13388
rect 8852 13336 8904 13388
rect 9404 13336 9456 13388
rect 9496 13336 9548 13388
rect 14648 13413 14657 13447
rect 14657 13413 14691 13447
rect 14691 13413 14700 13447
rect 14648 13404 14700 13413
rect 14832 13404 14884 13456
rect 16304 13404 16356 13456
rect 18328 13404 18380 13456
rect 12440 13336 12492 13388
rect 13268 13336 13320 13388
rect 13912 13336 13964 13388
rect 16580 13336 16632 13388
rect 17868 13379 17920 13388
rect 7656 13268 7708 13320
rect 9680 13268 9732 13320
rect 10968 13311 11020 13320
rect 10968 13277 10977 13311
rect 10977 13277 11011 13311
rect 11011 13277 11020 13311
rect 10968 13268 11020 13277
rect 10692 13200 10744 13252
rect 10876 13200 10928 13252
rect 12900 13268 12952 13320
rect 13636 13311 13688 13320
rect 13636 13277 13645 13311
rect 13645 13277 13679 13311
rect 13679 13277 13688 13311
rect 13636 13268 13688 13277
rect 13820 13311 13872 13320
rect 13820 13277 13829 13311
rect 13829 13277 13863 13311
rect 13863 13277 13872 13311
rect 13820 13268 13872 13277
rect 14924 13268 14976 13320
rect 15936 13268 15988 13320
rect 17040 13311 17092 13320
rect 17040 13277 17049 13311
rect 17049 13277 17083 13311
rect 17083 13277 17092 13311
rect 17040 13268 17092 13277
rect 11888 13200 11940 13252
rect 14648 13200 14700 13252
rect 17868 13345 17877 13379
rect 17877 13345 17911 13379
rect 17911 13345 17920 13379
rect 17868 13336 17920 13345
rect 18328 13268 18380 13320
rect 6920 13132 6972 13184
rect 9128 13132 9180 13184
rect 10232 13132 10284 13184
rect 11796 13132 11848 13184
rect 14556 13132 14608 13184
rect 17224 13132 17276 13184
rect 3947 13030 3999 13082
rect 4011 13030 4063 13082
rect 4075 13030 4127 13082
rect 4139 13030 4191 13082
rect 9878 13030 9930 13082
rect 9942 13030 9994 13082
rect 10006 13030 10058 13082
rect 10070 13030 10122 13082
rect 15808 13030 15860 13082
rect 15872 13030 15924 13082
rect 15936 13030 15988 13082
rect 16000 13030 16052 13082
rect 3516 12928 3568 12980
rect 5632 12928 5684 12980
rect 6092 12860 6144 12912
rect 6736 12860 6788 12912
rect 5080 12835 5132 12844
rect 5080 12801 5089 12835
rect 5089 12801 5123 12835
rect 5123 12801 5132 12835
rect 5080 12792 5132 12801
rect 6000 12835 6052 12844
rect 6000 12801 6009 12835
rect 6009 12801 6043 12835
rect 6043 12801 6052 12835
rect 6000 12792 6052 12801
rect 6184 12835 6236 12844
rect 6184 12801 6193 12835
rect 6193 12801 6227 12835
rect 6227 12801 6236 12835
rect 6184 12792 6236 12801
rect 6644 12792 6696 12844
rect 3700 12724 3752 12776
rect 3976 12724 4028 12776
rect 8024 12928 8076 12980
rect 10324 12971 10376 12980
rect 10324 12937 10333 12971
rect 10333 12937 10367 12971
rect 10367 12937 10376 12971
rect 10324 12928 10376 12937
rect 12348 12928 12400 12980
rect 10692 12860 10744 12912
rect 13452 12928 13504 12980
rect 10416 12792 10468 12844
rect 10876 12835 10928 12844
rect 10876 12801 10885 12835
rect 10885 12801 10919 12835
rect 10919 12801 10928 12835
rect 10876 12792 10928 12801
rect 6920 12767 6972 12776
rect 6920 12733 6929 12767
rect 6929 12733 6963 12767
rect 6963 12733 6972 12767
rect 6920 12724 6972 12733
rect 7748 12724 7800 12776
rect 5448 12656 5500 12708
rect 6368 12656 6420 12708
rect 9680 12724 9732 12776
rect 10232 12724 10284 12776
rect 14556 12860 14608 12912
rect 11796 12835 11848 12844
rect 11796 12801 11805 12835
rect 11805 12801 11839 12835
rect 11839 12801 11848 12835
rect 11796 12792 11848 12801
rect 7932 12656 7984 12708
rect 16672 12792 16724 12844
rect 14924 12767 14976 12776
rect 2504 12631 2556 12640
rect 2504 12597 2513 12631
rect 2513 12597 2547 12631
rect 2547 12597 2556 12631
rect 2504 12588 2556 12597
rect 4160 12588 4212 12640
rect 7748 12588 7800 12640
rect 10876 12656 10928 12708
rect 11428 12656 11480 12708
rect 14924 12733 14933 12767
rect 14933 12733 14967 12767
rect 14967 12733 14976 12767
rect 14924 12724 14976 12733
rect 15016 12724 15068 12776
rect 16948 12724 17000 12776
rect 17224 12767 17276 12776
rect 17224 12733 17233 12767
rect 17233 12733 17267 12767
rect 17267 12733 17276 12767
rect 17224 12724 17276 12733
rect 8208 12588 8260 12640
rect 12532 12656 12584 12708
rect 12808 12656 12860 12708
rect 12900 12656 12952 12708
rect 16580 12656 16632 12708
rect 17592 12656 17644 12708
rect 13544 12588 13596 12640
rect 13636 12588 13688 12640
rect 16856 12631 16908 12640
rect 16856 12597 16865 12631
rect 16865 12597 16899 12631
rect 16899 12597 16908 12631
rect 16856 12588 16908 12597
rect 17316 12631 17368 12640
rect 17316 12597 17325 12631
rect 17325 12597 17359 12631
rect 17359 12597 17368 12631
rect 17316 12588 17368 12597
rect 6912 12486 6964 12538
rect 6976 12486 7028 12538
rect 7040 12486 7092 12538
rect 7104 12486 7156 12538
rect 12843 12486 12895 12538
rect 12907 12486 12959 12538
rect 12971 12486 13023 12538
rect 13035 12486 13087 12538
rect 3332 12427 3384 12436
rect 3332 12393 3341 12427
rect 3341 12393 3375 12427
rect 3375 12393 3384 12427
rect 3332 12384 3384 12393
rect 8116 12427 8168 12436
rect 8116 12393 8125 12427
rect 8125 12393 8159 12427
rect 8159 12393 8168 12427
rect 8116 12384 8168 12393
rect 9220 12384 9272 12436
rect 10324 12384 10376 12436
rect 10784 12384 10836 12436
rect 12164 12384 12216 12436
rect 13820 12384 13872 12436
rect 6184 12316 6236 12368
rect 7840 12316 7892 12368
rect 2228 12291 2280 12300
rect 2228 12257 2237 12291
rect 2237 12257 2271 12291
rect 2271 12257 2280 12291
rect 2228 12248 2280 12257
rect 2320 12223 2372 12232
rect 2320 12189 2329 12223
rect 2329 12189 2363 12223
rect 2363 12189 2372 12223
rect 2320 12180 2372 12189
rect 2596 12180 2648 12232
rect 4160 12248 4212 12300
rect 6828 12248 6880 12300
rect 6920 12248 6972 12300
rect 10232 12248 10284 12300
rect 10416 12316 10468 12368
rect 13360 12316 13412 12368
rect 13636 12316 13688 12368
rect 13728 12316 13780 12368
rect 14740 12384 14792 12436
rect 15568 12384 15620 12436
rect 18052 12384 18104 12436
rect 16948 12316 17000 12368
rect 11612 12248 11664 12300
rect 15568 12248 15620 12300
rect 16120 12291 16172 12300
rect 16120 12257 16129 12291
rect 16129 12257 16163 12291
rect 16163 12257 16172 12291
rect 16120 12248 16172 12257
rect 16764 12291 16816 12300
rect 16764 12257 16773 12291
rect 16773 12257 16807 12291
rect 16807 12257 16816 12291
rect 16764 12248 16816 12257
rect 17040 12291 17092 12300
rect 17040 12257 17074 12291
rect 17074 12257 17092 12291
rect 17040 12248 17092 12257
rect 2964 12155 3016 12164
rect 2964 12121 2973 12155
rect 2973 12121 3007 12155
rect 3007 12121 3016 12155
rect 2964 12112 3016 12121
rect 1860 12087 1912 12096
rect 1860 12053 1869 12087
rect 1869 12053 1903 12087
rect 1903 12053 1912 12087
rect 1860 12044 1912 12053
rect 3700 12180 3752 12232
rect 6552 12223 6604 12232
rect 6552 12189 6561 12223
rect 6561 12189 6595 12223
rect 6595 12189 6604 12223
rect 6552 12180 6604 12189
rect 7012 12180 7064 12232
rect 8576 12223 8628 12232
rect 8576 12189 8585 12223
rect 8585 12189 8619 12223
rect 8619 12189 8628 12223
rect 8576 12180 8628 12189
rect 8944 12180 8996 12232
rect 5448 12087 5500 12096
rect 5448 12053 5457 12087
rect 5457 12053 5491 12087
rect 5491 12053 5500 12087
rect 5448 12044 5500 12053
rect 6644 12112 6696 12164
rect 8484 12112 8536 12164
rect 8852 12112 8904 12164
rect 7196 12044 7248 12096
rect 9312 12044 9364 12096
rect 12808 12180 12860 12232
rect 13176 12180 13228 12232
rect 12532 12112 12584 12164
rect 14556 12180 14608 12232
rect 15016 12180 15068 12232
rect 14280 12112 14332 12164
rect 15108 12112 15160 12164
rect 10508 12044 10560 12096
rect 12072 12044 12124 12096
rect 12716 12044 12768 12096
rect 13636 12044 13688 12096
rect 14004 12044 14056 12096
rect 16212 12223 16264 12232
rect 16212 12189 16221 12223
rect 16221 12189 16255 12223
rect 16255 12189 16264 12223
rect 16212 12180 16264 12189
rect 16580 12180 16632 12232
rect 15660 12044 15712 12096
rect 3947 11942 3999 11994
rect 4011 11942 4063 11994
rect 4075 11942 4127 11994
rect 4139 11942 4191 11994
rect 9878 11942 9930 11994
rect 9942 11942 9994 11994
rect 10006 11942 10058 11994
rect 10070 11942 10122 11994
rect 15808 11942 15860 11994
rect 15872 11942 15924 11994
rect 15936 11942 15988 11994
rect 16000 11942 16052 11994
rect 2228 11883 2280 11892
rect 2228 11849 2237 11883
rect 2237 11849 2271 11883
rect 2271 11849 2280 11883
rect 2228 11840 2280 11849
rect 6828 11883 6880 11892
rect 6828 11849 6837 11883
rect 6837 11849 6871 11883
rect 6871 11849 6880 11883
rect 6828 11840 6880 11849
rect 6920 11772 6972 11824
rect 2412 11704 2464 11756
rect 6184 11704 6236 11756
rect 6644 11704 6696 11756
rect 9772 11772 9824 11824
rect 12256 11840 12308 11892
rect 13360 11840 13412 11892
rect 14740 11840 14792 11892
rect 15292 11840 15344 11892
rect 16120 11840 16172 11892
rect 11704 11772 11756 11824
rect 15568 11772 15620 11824
rect 18236 11772 18288 11824
rect 7472 11747 7524 11756
rect 1676 11679 1728 11688
rect 1676 11645 1685 11679
rect 1685 11645 1719 11679
rect 1719 11645 1728 11679
rect 1676 11636 1728 11645
rect 2504 11636 2556 11688
rect 2688 11611 2740 11620
rect 2688 11577 2697 11611
rect 2697 11577 2731 11611
rect 2731 11577 2740 11611
rect 2688 11568 2740 11577
rect 3700 11636 3752 11688
rect 3884 11636 3936 11688
rect 5080 11636 5132 11688
rect 1492 11500 1544 11552
rect 2964 11500 3016 11552
rect 4252 11568 4304 11620
rect 7104 11636 7156 11688
rect 7472 11713 7481 11747
rect 7481 11713 7515 11747
rect 7515 11713 7524 11747
rect 7472 11704 7524 11713
rect 8944 11704 8996 11756
rect 11888 11704 11940 11756
rect 12164 11704 12216 11756
rect 7656 11636 7708 11688
rect 8024 11636 8076 11688
rect 8208 11679 8260 11688
rect 8208 11645 8242 11679
rect 8242 11645 8260 11679
rect 8208 11636 8260 11645
rect 6828 11568 6880 11620
rect 12348 11636 12400 11688
rect 14096 11704 14148 11756
rect 15660 11747 15712 11756
rect 15660 11713 15669 11747
rect 15669 11713 15703 11747
rect 15703 11713 15712 11747
rect 15660 11704 15712 11713
rect 16120 11704 16172 11756
rect 16764 11747 16816 11756
rect 16764 11713 16773 11747
rect 16773 11713 16807 11747
rect 16807 11713 16816 11747
rect 16764 11704 16816 11713
rect 9496 11568 9548 11620
rect 11980 11568 12032 11620
rect 16304 11636 16356 11688
rect 17224 11636 17276 11688
rect 14464 11611 14516 11620
rect 5172 11543 5224 11552
rect 5172 11509 5181 11543
rect 5181 11509 5215 11543
rect 5215 11509 5224 11543
rect 5172 11500 5224 11509
rect 6000 11500 6052 11552
rect 6736 11500 6788 11552
rect 8668 11500 8720 11552
rect 9680 11500 9732 11552
rect 10600 11500 10652 11552
rect 14464 11577 14473 11611
rect 14473 11577 14507 11611
rect 14507 11577 14516 11611
rect 14464 11568 14516 11577
rect 16856 11568 16908 11620
rect 13176 11500 13228 11552
rect 13728 11500 13780 11552
rect 14372 11500 14424 11552
rect 15200 11543 15252 11552
rect 15200 11509 15209 11543
rect 15209 11509 15243 11543
rect 15243 11509 15252 11543
rect 15200 11500 15252 11509
rect 16948 11500 17000 11552
rect 6912 11398 6964 11450
rect 6976 11398 7028 11450
rect 7040 11398 7092 11450
rect 7104 11398 7156 11450
rect 12843 11398 12895 11450
rect 12907 11398 12959 11450
rect 12971 11398 13023 11450
rect 13035 11398 13087 11450
rect 2136 11296 2188 11348
rect 6368 11296 6420 11348
rect 6552 11339 6604 11348
rect 6552 11305 6561 11339
rect 6561 11305 6595 11339
rect 6595 11305 6604 11339
rect 6552 11296 6604 11305
rect 6736 11296 6788 11348
rect 8116 11296 8168 11348
rect 9496 11296 9548 11348
rect 9680 11339 9732 11348
rect 9680 11305 9689 11339
rect 9689 11305 9723 11339
rect 9723 11305 9732 11339
rect 9680 11296 9732 11305
rect 9864 11296 9916 11348
rect 13636 11296 13688 11348
rect 13912 11296 13964 11348
rect 14372 11296 14424 11348
rect 16212 11339 16264 11348
rect 16212 11305 16221 11339
rect 16221 11305 16255 11339
rect 16255 11305 16264 11339
rect 16212 11296 16264 11305
rect 17316 11296 17368 11348
rect 17500 11296 17552 11348
rect 18788 11296 18840 11348
rect 2688 11228 2740 11280
rect 2504 11203 2556 11212
rect 2504 11169 2538 11203
rect 2538 11169 2556 11203
rect 2504 11160 2556 11169
rect 5172 11160 5224 11212
rect 7840 11228 7892 11280
rect 10968 11228 11020 11280
rect 11888 11228 11940 11280
rect 6552 11160 6604 11212
rect 6920 11203 6972 11212
rect 6920 11169 6929 11203
rect 6929 11169 6963 11203
rect 6963 11169 6972 11203
rect 6920 11160 6972 11169
rect 7748 11160 7800 11212
rect 7932 11203 7984 11212
rect 7932 11169 7941 11203
rect 7941 11169 7975 11203
rect 7975 11169 7984 11203
rect 7932 11160 7984 11169
rect 8392 11160 8444 11212
rect 1308 11092 1360 11144
rect 3700 11092 3752 11144
rect 9220 11160 9272 11212
rect 9680 11160 9732 11212
rect 11704 11203 11756 11212
rect 1400 11024 1452 11076
rect 3240 11024 3292 11076
rect 5448 11067 5500 11076
rect 5448 11033 5457 11067
rect 5457 11033 5491 11067
rect 5491 11033 5500 11067
rect 5448 11024 5500 11033
rect 7472 11024 7524 11076
rect 3516 10956 3568 11008
rect 5264 10956 5316 11008
rect 5356 10956 5408 11008
rect 8852 11024 8904 11076
rect 9312 11092 9364 11144
rect 10324 11092 10376 11144
rect 10600 11092 10652 11144
rect 11704 11169 11713 11203
rect 11713 11169 11747 11203
rect 11747 11169 11756 11203
rect 11704 11160 11756 11169
rect 12348 11203 12400 11212
rect 12348 11169 12357 11203
rect 12357 11169 12391 11203
rect 12391 11169 12400 11203
rect 12348 11160 12400 11169
rect 12624 11203 12676 11212
rect 12624 11169 12658 11203
rect 12658 11169 12676 11203
rect 12624 11160 12676 11169
rect 14372 11203 14424 11212
rect 14372 11169 14381 11203
rect 14381 11169 14415 11203
rect 14415 11169 14424 11203
rect 14372 11160 14424 11169
rect 15660 11160 15712 11212
rect 17960 11228 18012 11280
rect 17592 11160 17644 11212
rect 11796 11135 11848 11144
rect 11428 11024 11480 11076
rect 11796 11101 11805 11135
rect 11805 11101 11839 11135
rect 11839 11101 11848 11135
rect 11796 11092 11848 11101
rect 11980 11135 12032 11144
rect 11980 11101 11989 11135
rect 11989 11101 12023 11135
rect 12023 11101 12032 11135
rect 11980 11092 12032 11101
rect 14004 11092 14056 11144
rect 14280 11092 14332 11144
rect 15292 11135 15344 11144
rect 8392 10956 8444 11008
rect 9588 10956 9640 11008
rect 10508 10956 10560 11008
rect 14096 11024 14148 11076
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 16672 11135 16724 11144
rect 16672 11101 16681 11135
rect 16681 11101 16715 11135
rect 16715 11101 16724 11135
rect 16672 11092 16724 11101
rect 16764 11092 16816 11144
rect 18328 11092 18380 11144
rect 13452 10956 13504 11008
rect 13544 10956 13596 11008
rect 17592 10956 17644 11008
rect 18052 10956 18104 11008
rect 3947 10854 3999 10906
rect 4011 10854 4063 10906
rect 4075 10854 4127 10906
rect 4139 10854 4191 10906
rect 9878 10854 9930 10906
rect 9942 10854 9994 10906
rect 10006 10854 10058 10906
rect 10070 10854 10122 10906
rect 15808 10854 15860 10906
rect 15872 10854 15924 10906
rect 15936 10854 15988 10906
rect 16000 10854 16052 10906
rect 2320 10752 2372 10804
rect 4804 10752 4856 10804
rect 6828 10752 6880 10804
rect 3332 10684 3384 10736
rect 2504 10616 2556 10668
rect 5172 10616 5224 10668
rect 5356 10616 5408 10668
rect 5448 10616 5500 10668
rect 8024 10752 8076 10804
rect 8760 10795 8812 10804
rect 8760 10761 8769 10795
rect 8769 10761 8803 10795
rect 8803 10761 8812 10795
rect 8760 10752 8812 10761
rect 10416 10795 10468 10804
rect 10416 10761 10425 10795
rect 10425 10761 10459 10795
rect 10459 10761 10468 10795
rect 10416 10752 10468 10761
rect 11704 10752 11756 10804
rect 14464 10752 14516 10804
rect 14556 10752 14608 10804
rect 12716 10684 12768 10736
rect 14280 10684 14332 10736
rect 5540 10548 5592 10600
rect 2780 10480 2832 10532
rect 4068 10480 4120 10532
rect 3424 10455 3476 10464
rect 3424 10421 3433 10455
rect 3433 10421 3467 10455
rect 3467 10421 3476 10455
rect 3424 10412 3476 10421
rect 3792 10455 3844 10464
rect 3792 10421 3801 10455
rect 3801 10421 3835 10455
rect 3835 10421 3844 10455
rect 3792 10412 3844 10421
rect 4344 10412 4396 10464
rect 6736 10480 6788 10532
rect 8944 10548 8996 10600
rect 12624 10616 12676 10668
rect 13176 10616 13228 10668
rect 8024 10480 8076 10532
rect 9588 10548 9640 10600
rect 12348 10548 12400 10600
rect 14096 10548 14148 10600
rect 14556 10616 14608 10668
rect 14924 10752 14976 10804
rect 14464 10548 14516 10600
rect 4804 10455 4856 10464
rect 4804 10421 4813 10455
rect 4813 10421 4847 10455
rect 4847 10421 4856 10455
rect 4804 10412 4856 10421
rect 5264 10412 5316 10464
rect 5448 10455 5500 10464
rect 5448 10421 5457 10455
rect 5457 10421 5491 10455
rect 5491 10421 5500 10455
rect 5448 10412 5500 10421
rect 5816 10455 5868 10464
rect 5816 10421 5825 10455
rect 5825 10421 5859 10455
rect 5859 10421 5868 10455
rect 5816 10412 5868 10421
rect 6184 10412 6236 10464
rect 7288 10412 7340 10464
rect 7932 10412 7984 10464
rect 13912 10480 13964 10532
rect 15292 10548 15344 10600
rect 16120 10752 16172 10804
rect 17040 10752 17092 10804
rect 15752 10548 15804 10600
rect 17500 10480 17552 10532
rect 9220 10412 9272 10464
rect 10968 10412 11020 10464
rect 11704 10455 11756 10464
rect 11704 10421 11713 10455
rect 11713 10421 11747 10455
rect 11747 10421 11756 10455
rect 11704 10412 11756 10421
rect 12716 10412 12768 10464
rect 13360 10412 13412 10464
rect 13820 10412 13872 10464
rect 14740 10412 14792 10464
rect 16580 10412 16632 10464
rect 6912 10310 6964 10362
rect 6976 10310 7028 10362
rect 7040 10310 7092 10362
rect 7104 10310 7156 10362
rect 12843 10310 12895 10362
rect 12907 10310 12959 10362
rect 12971 10310 13023 10362
rect 13035 10310 13087 10362
rect 1308 10208 1360 10260
rect 3700 10208 3752 10260
rect 3792 10208 3844 10260
rect 4988 10208 5040 10260
rect 5540 10251 5592 10260
rect 2596 10140 2648 10192
rect 3240 10140 3292 10192
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 6092 10208 6144 10260
rect 8576 10208 8628 10260
rect 11888 10208 11940 10260
rect 14464 10208 14516 10260
rect 17500 10251 17552 10260
rect 17500 10217 17509 10251
rect 17509 10217 17543 10251
rect 17543 10217 17552 10251
rect 17500 10208 17552 10217
rect 17868 10251 17920 10260
rect 17868 10217 17877 10251
rect 17877 10217 17911 10251
rect 17911 10217 17920 10251
rect 17868 10208 17920 10217
rect 1308 10004 1360 10056
rect 4896 10115 4948 10124
rect 4896 10081 4905 10115
rect 4905 10081 4939 10115
rect 4939 10081 4948 10115
rect 9772 10140 9824 10192
rect 12992 10140 13044 10192
rect 13176 10140 13228 10192
rect 5724 10115 5776 10124
rect 4896 10072 4948 10081
rect 5724 10081 5733 10115
rect 5733 10081 5767 10115
rect 5767 10081 5776 10115
rect 5724 10072 5776 10081
rect 8852 10072 8904 10124
rect 4620 10004 4672 10056
rect 5172 10004 5224 10056
rect 4804 9936 4856 9988
rect 5540 9936 5592 9988
rect 2780 9911 2832 9920
rect 2780 9877 2789 9911
rect 2789 9877 2823 9911
rect 2823 9877 2832 9911
rect 2780 9868 2832 9877
rect 3056 9868 3108 9920
rect 7196 10004 7248 10056
rect 7932 10047 7984 10056
rect 7932 10013 7941 10047
rect 7941 10013 7975 10047
rect 7975 10013 7984 10047
rect 7932 10004 7984 10013
rect 8024 10047 8076 10056
rect 8024 10013 8033 10047
rect 8033 10013 8067 10047
rect 8067 10013 8076 10047
rect 10416 10072 10468 10124
rect 10508 10072 10560 10124
rect 10876 10072 10928 10124
rect 12348 10072 12400 10124
rect 8024 10004 8076 10013
rect 10784 10004 10836 10056
rect 13820 10072 13872 10124
rect 11060 9979 11112 9988
rect 11060 9945 11069 9979
rect 11069 9945 11103 9979
rect 11103 9945 11112 9979
rect 11060 9936 11112 9945
rect 12256 9936 12308 9988
rect 6184 9868 6236 9920
rect 6736 9868 6788 9920
rect 7932 9868 7984 9920
rect 10876 9868 10928 9920
rect 12440 9868 12492 9920
rect 16212 10072 16264 10124
rect 16764 10140 16816 10192
rect 17776 10140 17828 10192
rect 17224 10072 17276 10124
rect 12716 9936 12768 9988
rect 15752 9936 15804 9988
rect 14372 9868 14424 9920
rect 17868 9868 17920 9920
rect 3947 9766 3999 9818
rect 4011 9766 4063 9818
rect 4075 9766 4127 9818
rect 4139 9766 4191 9818
rect 9878 9766 9930 9818
rect 9942 9766 9994 9818
rect 10006 9766 10058 9818
rect 10070 9766 10122 9818
rect 15808 9766 15860 9818
rect 15872 9766 15924 9818
rect 15936 9766 15988 9818
rect 16000 9766 16052 9818
rect 3608 9664 3660 9716
rect 5356 9664 5408 9716
rect 5816 9664 5868 9716
rect 9772 9664 9824 9716
rect 10784 9664 10836 9716
rect 10968 9664 11020 9716
rect 16488 9664 16540 9716
rect 4344 9596 4396 9648
rect 1308 9528 1360 9580
rect 4068 9528 4120 9580
rect 2780 9460 2832 9512
rect 4528 9460 4580 9512
rect 5172 9528 5224 9580
rect 6368 9571 6420 9580
rect 6368 9537 6377 9571
rect 6377 9537 6411 9571
rect 6411 9537 6420 9571
rect 6368 9528 6420 9537
rect 6736 9528 6788 9580
rect 7196 9460 7248 9512
rect 8576 9528 8628 9580
rect 12716 9596 12768 9648
rect 13452 9639 13504 9648
rect 9680 9528 9732 9580
rect 10876 9528 10928 9580
rect 8116 9460 8168 9512
rect 10416 9460 10468 9512
rect 5908 9392 5960 9444
rect 3148 9324 3200 9376
rect 3516 9367 3568 9376
rect 3516 9333 3525 9367
rect 3525 9333 3559 9367
rect 3559 9333 3568 9367
rect 3516 9324 3568 9333
rect 3608 9324 3660 9376
rect 4712 9324 4764 9376
rect 5816 9324 5868 9376
rect 6092 9367 6144 9376
rect 6092 9333 6101 9367
rect 6101 9333 6135 9367
rect 6135 9333 6144 9367
rect 6092 9324 6144 9333
rect 6184 9367 6236 9376
rect 6184 9333 6193 9367
rect 6193 9333 6227 9367
rect 6227 9333 6236 9367
rect 11060 9460 11112 9512
rect 13452 9605 13461 9639
rect 13461 9605 13495 9639
rect 13495 9605 13504 9639
rect 13452 9596 13504 9605
rect 13820 9596 13872 9648
rect 16672 9596 16724 9648
rect 13176 9528 13228 9580
rect 13912 9528 13964 9580
rect 14188 9571 14240 9580
rect 14188 9537 14197 9571
rect 14197 9537 14231 9571
rect 14231 9537 14240 9571
rect 14188 9528 14240 9537
rect 17408 9571 17460 9580
rect 17408 9537 17417 9571
rect 17417 9537 17451 9571
rect 17451 9537 17460 9571
rect 17408 9528 17460 9537
rect 14464 9435 14516 9444
rect 14464 9401 14498 9435
rect 14498 9401 14516 9435
rect 14464 9392 14516 9401
rect 6184 9324 6236 9333
rect 7656 9367 7708 9376
rect 7656 9333 7665 9367
rect 7665 9333 7699 9367
rect 7699 9333 7708 9367
rect 7656 9324 7708 9333
rect 8208 9367 8260 9376
rect 8208 9333 8217 9367
rect 8217 9333 8251 9367
rect 8251 9333 8260 9367
rect 8208 9324 8260 9333
rect 8392 9324 8444 9376
rect 9496 9324 9548 9376
rect 12532 9324 12584 9376
rect 15292 9392 15344 9444
rect 15384 9324 15436 9376
rect 17316 9324 17368 9376
rect 6912 9222 6964 9274
rect 6976 9222 7028 9274
rect 7040 9222 7092 9274
rect 7104 9222 7156 9274
rect 12843 9222 12895 9274
rect 12907 9222 12959 9274
rect 12971 9222 13023 9274
rect 13035 9222 13087 9274
rect 1860 9120 1912 9172
rect 3424 9163 3476 9172
rect 3424 9129 3433 9163
rect 3433 9129 3467 9163
rect 3467 9129 3476 9163
rect 3424 9120 3476 9129
rect 5908 9120 5960 9172
rect 6276 9120 6328 9172
rect 6460 9120 6512 9172
rect 3516 9052 3568 9104
rect 5816 9052 5868 9104
rect 5448 8984 5500 9036
rect 6276 8984 6328 9036
rect 6828 8984 6880 9036
rect 8024 9052 8076 9104
rect 8208 9120 8260 9172
rect 11520 9120 11572 9172
rect 11796 9120 11848 9172
rect 12532 9163 12584 9172
rect 12532 9129 12541 9163
rect 12541 9129 12575 9163
rect 12575 9129 12584 9163
rect 12532 9120 12584 9129
rect 14188 9120 14240 9172
rect 14556 9120 14608 9172
rect 12348 9052 12400 9104
rect 12440 9095 12492 9104
rect 12440 9061 12449 9095
rect 12449 9061 12483 9095
rect 12483 9061 12492 9095
rect 17776 9120 17828 9172
rect 12440 9052 12492 9061
rect 16212 9052 16264 9104
rect 13728 8984 13780 9036
rect 13820 8984 13872 9036
rect 16396 8984 16448 9036
rect 17408 8984 17460 9036
rect 2780 8916 2832 8968
rect 3240 8916 3292 8968
rect 3700 8916 3752 8968
rect 1768 8780 1820 8832
rect 4988 8780 5040 8832
rect 7288 8916 7340 8968
rect 9036 8959 9088 8968
rect 9036 8925 9045 8959
rect 9045 8925 9079 8959
rect 9079 8925 9088 8959
rect 9036 8916 9088 8925
rect 12624 8959 12676 8968
rect 12624 8925 12633 8959
rect 12633 8925 12667 8959
rect 12667 8925 12676 8959
rect 12624 8916 12676 8925
rect 14188 8916 14240 8968
rect 16212 8916 16264 8968
rect 6828 8780 6880 8832
rect 12808 8848 12860 8900
rect 8852 8780 8904 8832
rect 10324 8780 10376 8832
rect 16304 8848 16356 8900
rect 14464 8823 14516 8832
rect 14464 8789 14473 8823
rect 14473 8789 14507 8823
rect 14507 8789 14516 8823
rect 14464 8780 14516 8789
rect 3947 8678 3999 8730
rect 4011 8678 4063 8730
rect 4075 8678 4127 8730
rect 4139 8678 4191 8730
rect 9878 8678 9930 8730
rect 9942 8678 9994 8730
rect 10006 8678 10058 8730
rect 10070 8678 10122 8730
rect 15808 8678 15860 8730
rect 15872 8678 15924 8730
rect 15936 8678 15988 8730
rect 16000 8678 16052 8730
rect 5724 8576 5776 8628
rect 6184 8576 6236 8628
rect 3424 8508 3476 8560
rect 5356 8508 5408 8560
rect 1308 8440 1360 8492
rect 3516 8440 3568 8492
rect 4988 8483 5040 8492
rect 4988 8449 4997 8483
rect 4997 8449 5031 8483
rect 5031 8449 5040 8483
rect 4988 8440 5040 8449
rect 2504 8372 2556 8424
rect 2688 8304 2740 8356
rect 4252 8372 4304 8424
rect 4804 8415 4856 8424
rect 4804 8381 4813 8415
rect 4813 8381 4847 8415
rect 4847 8381 4856 8415
rect 4804 8372 4856 8381
rect 6460 8440 6512 8492
rect 6736 8440 6788 8492
rect 7196 8372 7248 8424
rect 4068 8304 4120 8356
rect 4436 8304 4488 8356
rect 5724 8304 5776 8356
rect 7288 8304 7340 8356
rect 2872 8236 2924 8288
rect 3332 8279 3384 8288
rect 3332 8245 3341 8279
rect 3341 8245 3375 8279
rect 3375 8245 3384 8279
rect 3332 8236 3384 8245
rect 3976 8236 4028 8288
rect 6460 8236 6512 8288
rect 6552 8236 6604 8288
rect 10968 8551 11020 8560
rect 10968 8517 10977 8551
rect 10977 8517 11011 8551
rect 11011 8517 11020 8551
rect 10968 8508 11020 8517
rect 12716 8576 12768 8628
rect 12808 8576 12860 8628
rect 12348 8508 12400 8560
rect 13912 8576 13964 8628
rect 11612 8483 11664 8492
rect 11612 8449 11621 8483
rect 11621 8449 11655 8483
rect 11655 8449 11664 8483
rect 11612 8440 11664 8449
rect 14464 8440 14516 8492
rect 13912 8372 13964 8424
rect 8392 8304 8444 8356
rect 12532 8304 12584 8356
rect 14740 8347 14792 8356
rect 14740 8313 14749 8347
rect 14749 8313 14783 8347
rect 14783 8313 14792 8347
rect 14740 8304 14792 8313
rect 14924 8304 14976 8356
rect 16396 8576 16448 8628
rect 17408 8619 17460 8628
rect 17408 8585 17417 8619
rect 17417 8585 17451 8619
rect 17451 8585 17460 8619
rect 17408 8576 17460 8585
rect 16028 8483 16080 8492
rect 16028 8449 16037 8483
rect 16037 8449 16071 8483
rect 16071 8449 16080 8483
rect 16028 8440 16080 8449
rect 15936 8372 15988 8424
rect 16304 8415 16356 8424
rect 16304 8381 16338 8415
rect 16338 8381 16356 8415
rect 16304 8372 16356 8381
rect 18052 8415 18104 8424
rect 18052 8381 18061 8415
rect 18061 8381 18095 8415
rect 18095 8381 18104 8415
rect 18052 8372 18104 8381
rect 16488 8304 16540 8356
rect 7656 8236 7708 8288
rect 8208 8236 8260 8288
rect 8760 8236 8812 8288
rect 8944 8236 8996 8288
rect 11060 8236 11112 8288
rect 11336 8279 11388 8288
rect 11336 8245 11345 8279
rect 11345 8245 11379 8279
rect 11379 8245 11388 8279
rect 11336 8236 11388 8245
rect 12440 8236 12492 8288
rect 13176 8236 13228 8288
rect 14372 8279 14424 8288
rect 14372 8245 14381 8279
rect 14381 8245 14415 8279
rect 14415 8245 14424 8279
rect 14372 8236 14424 8245
rect 15660 8236 15712 8288
rect 16580 8236 16632 8288
rect 18236 8279 18288 8288
rect 18236 8245 18245 8279
rect 18245 8245 18279 8279
rect 18279 8245 18288 8279
rect 18236 8236 18288 8245
rect 6912 8134 6964 8186
rect 6976 8134 7028 8186
rect 7040 8134 7092 8186
rect 7104 8134 7156 8186
rect 12843 8134 12895 8186
rect 12907 8134 12959 8186
rect 12971 8134 13023 8186
rect 13035 8134 13087 8186
rect 3332 8032 3384 8084
rect 6092 8032 6144 8084
rect 6460 8032 6512 8084
rect 4804 7964 4856 8016
rect 2320 7939 2372 7948
rect 2320 7905 2329 7939
rect 2329 7905 2363 7939
rect 2363 7905 2372 7939
rect 2320 7896 2372 7905
rect 2688 7896 2740 7948
rect 2872 7828 2924 7880
rect 3332 7939 3384 7948
rect 3332 7905 3341 7939
rect 3341 7905 3375 7939
rect 3375 7905 3384 7939
rect 3332 7896 3384 7905
rect 3976 7896 4028 7948
rect 4252 7828 4304 7880
rect 2780 7760 2832 7812
rect 1952 7735 2004 7744
rect 1952 7701 1961 7735
rect 1961 7701 1995 7735
rect 1995 7701 2004 7735
rect 1952 7692 2004 7701
rect 2688 7692 2740 7744
rect 3332 7692 3384 7744
rect 3700 7692 3752 7744
rect 4896 7896 4948 7948
rect 6368 7896 6420 7948
rect 6644 7896 6696 7948
rect 7288 8032 7340 8084
rect 7472 8075 7524 8084
rect 7472 8041 7481 8075
rect 7481 8041 7515 8075
rect 7515 8041 7524 8075
rect 7472 8032 7524 8041
rect 8116 8075 8168 8084
rect 8116 8041 8125 8075
rect 8125 8041 8159 8075
rect 8159 8041 8168 8075
rect 8116 8032 8168 8041
rect 8484 8075 8536 8084
rect 8484 8041 8493 8075
rect 8493 8041 8527 8075
rect 8527 8041 8536 8075
rect 8484 8032 8536 8041
rect 8576 8032 8628 8084
rect 10232 8032 10284 8084
rect 10876 8032 10928 8084
rect 11612 8032 11664 8084
rect 12532 8032 12584 8084
rect 13820 8032 13872 8084
rect 14188 8075 14240 8084
rect 14188 8041 14197 8075
rect 14197 8041 14231 8075
rect 14231 8041 14240 8075
rect 14188 8032 14240 8041
rect 14372 8032 14424 8084
rect 15936 8032 15988 8084
rect 7564 8007 7616 8016
rect 7564 7973 7573 8007
rect 7573 7973 7607 8007
rect 7607 7973 7616 8007
rect 7564 7964 7616 7973
rect 7748 7964 7800 8016
rect 7840 7964 7892 8016
rect 8024 7964 8076 8016
rect 8944 7964 8996 8016
rect 10508 7964 10560 8016
rect 10968 7964 11020 8016
rect 11060 7964 11112 8016
rect 13636 7964 13688 8016
rect 14556 8007 14608 8016
rect 14556 7973 14565 8007
rect 14565 7973 14599 8007
rect 14599 7973 14608 8007
rect 14556 7964 14608 7973
rect 14832 7964 14884 8016
rect 16212 7964 16264 8016
rect 8484 7896 8536 7948
rect 9864 7896 9916 7948
rect 6828 7828 6880 7880
rect 7656 7871 7708 7880
rect 6000 7760 6052 7812
rect 6276 7760 6328 7812
rect 7656 7837 7665 7871
rect 7665 7837 7699 7871
rect 7699 7837 7708 7871
rect 7656 7828 7708 7837
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8576 7828 8628 7837
rect 8668 7760 8720 7812
rect 8852 7828 8904 7880
rect 8944 7760 8996 7812
rect 11520 7896 11572 7948
rect 13268 7896 13320 7948
rect 16028 7939 16080 7948
rect 10508 7871 10560 7880
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10508 7828 10560 7837
rect 11612 7828 11664 7880
rect 12164 7735 12216 7744
rect 12164 7701 12173 7735
rect 12173 7701 12207 7735
rect 12207 7701 12216 7735
rect 12164 7692 12216 7701
rect 12348 7760 12400 7812
rect 13452 7828 13504 7880
rect 13728 7828 13780 7880
rect 15384 7828 15436 7880
rect 13912 7760 13964 7812
rect 15660 7692 15712 7744
rect 16028 7905 16037 7939
rect 16037 7905 16071 7939
rect 16071 7905 16080 7939
rect 16028 7896 16080 7905
rect 17868 7939 17920 7948
rect 17868 7905 17877 7939
rect 17877 7905 17911 7939
rect 17911 7905 17920 7939
rect 17868 7896 17920 7905
rect 17500 7692 17552 7744
rect 18052 7735 18104 7744
rect 18052 7701 18061 7735
rect 18061 7701 18095 7735
rect 18095 7701 18104 7735
rect 18052 7692 18104 7701
rect 3947 7590 3999 7642
rect 4011 7590 4063 7642
rect 4075 7590 4127 7642
rect 4139 7590 4191 7642
rect 9878 7590 9930 7642
rect 9942 7590 9994 7642
rect 10006 7590 10058 7642
rect 10070 7590 10122 7642
rect 15808 7590 15860 7642
rect 15872 7590 15924 7642
rect 15936 7590 15988 7642
rect 16000 7590 16052 7642
rect 2320 7488 2372 7540
rect 2596 7420 2648 7472
rect 4804 7488 4856 7540
rect 6368 7531 6420 7540
rect 4252 7420 4304 7472
rect 4988 7420 5040 7472
rect 6368 7497 6377 7531
rect 6377 7497 6411 7531
rect 6411 7497 6420 7531
rect 6368 7488 6420 7497
rect 6000 7352 6052 7404
rect 7564 7352 7616 7404
rect 8116 7395 8168 7404
rect 8116 7361 8125 7395
rect 8125 7361 8159 7395
rect 8159 7361 8168 7395
rect 8116 7352 8168 7361
rect 11336 7488 11388 7540
rect 11520 7488 11572 7540
rect 14280 7488 14332 7540
rect 14648 7488 14700 7540
rect 15016 7488 15068 7540
rect 10140 7352 10192 7404
rect 12164 7420 12216 7472
rect 10968 7395 11020 7404
rect 10968 7361 10977 7395
rect 10977 7361 11011 7395
rect 11011 7361 11020 7395
rect 10968 7352 11020 7361
rect 11244 7352 11296 7404
rect 12348 7420 12400 7472
rect 12532 7420 12584 7472
rect 14740 7420 14792 7472
rect 13084 7395 13136 7404
rect 13084 7361 13093 7395
rect 13093 7361 13127 7395
rect 13127 7361 13136 7395
rect 13084 7352 13136 7361
rect 1676 7284 1728 7336
rect 2872 7216 2924 7268
rect 3332 7216 3384 7268
rect 2320 7148 2372 7200
rect 2964 7191 3016 7200
rect 2964 7157 2973 7191
rect 2973 7157 3007 7191
rect 3007 7157 3016 7191
rect 2964 7148 3016 7157
rect 3792 7284 3844 7336
rect 4436 7284 4488 7336
rect 4896 7284 4948 7336
rect 5540 7284 5592 7336
rect 6368 7284 6420 7336
rect 8392 7284 8444 7336
rect 8576 7327 8628 7336
rect 8576 7293 8585 7327
rect 8585 7293 8619 7327
rect 8619 7293 8628 7327
rect 8576 7284 8628 7293
rect 6736 7216 6788 7268
rect 10600 7284 10652 7336
rect 13176 7284 13228 7336
rect 13912 7352 13964 7404
rect 14648 7352 14700 7404
rect 15660 7488 15712 7540
rect 16212 7488 16264 7540
rect 16856 7531 16908 7540
rect 16856 7497 16865 7531
rect 16865 7497 16899 7531
rect 16899 7497 16908 7531
rect 16856 7488 16908 7497
rect 17592 7531 17644 7540
rect 17592 7497 17601 7531
rect 17601 7497 17635 7531
rect 17635 7497 17644 7531
rect 17592 7488 17644 7497
rect 14096 7327 14148 7336
rect 14096 7293 14105 7327
rect 14105 7293 14139 7327
rect 14139 7293 14148 7327
rect 14096 7284 14148 7293
rect 14556 7284 14608 7336
rect 17500 7284 17552 7336
rect 8852 7259 8904 7268
rect 8852 7225 8886 7259
rect 8886 7225 8904 7259
rect 8852 7216 8904 7225
rect 8944 7216 8996 7268
rect 6644 7148 6696 7200
rect 7288 7148 7340 7200
rect 7472 7191 7524 7200
rect 7472 7157 7481 7191
rect 7481 7157 7515 7191
rect 7515 7157 7524 7191
rect 7472 7148 7524 7157
rect 9680 7148 9732 7200
rect 9772 7148 9824 7200
rect 10784 7148 10836 7200
rect 11336 7191 11388 7200
rect 11336 7157 11345 7191
rect 11345 7157 11379 7191
rect 11379 7157 11388 7191
rect 11336 7148 11388 7157
rect 11428 7148 11480 7200
rect 11796 7191 11848 7200
rect 11796 7157 11805 7191
rect 11805 7157 11839 7191
rect 11839 7157 11848 7191
rect 11796 7148 11848 7157
rect 11980 7148 12032 7200
rect 13268 7148 13320 7200
rect 13452 7148 13504 7200
rect 15384 7216 15436 7268
rect 13820 7148 13872 7200
rect 14740 7191 14792 7200
rect 14740 7157 14749 7191
rect 14749 7157 14783 7191
rect 14783 7157 14792 7191
rect 14740 7148 14792 7157
rect 15200 7148 15252 7200
rect 16212 7148 16264 7200
rect 18236 7191 18288 7200
rect 18236 7157 18245 7191
rect 18245 7157 18279 7191
rect 18279 7157 18288 7191
rect 18236 7148 18288 7157
rect 6912 7046 6964 7098
rect 6976 7046 7028 7098
rect 7040 7046 7092 7098
rect 7104 7046 7156 7098
rect 12843 7046 12895 7098
rect 12907 7046 12959 7098
rect 12971 7046 13023 7098
rect 13035 7046 13087 7098
rect 2872 6944 2924 6996
rect 10232 6944 10284 6996
rect 11796 6944 11848 6996
rect 7472 6876 7524 6928
rect 1860 6808 1912 6860
rect 2964 6808 3016 6860
rect 3792 6808 3844 6860
rect 4252 6808 4304 6860
rect 5632 6808 5684 6860
rect 7288 6808 7340 6860
rect 8576 6876 8628 6928
rect 8852 6876 8904 6928
rect 9312 6876 9364 6928
rect 2320 6783 2372 6792
rect 2320 6749 2329 6783
rect 2329 6749 2363 6783
rect 2363 6749 2372 6783
rect 2320 6740 2372 6749
rect 4620 6740 4672 6792
rect 4988 6740 5040 6792
rect 6644 6740 6696 6792
rect 3516 6604 3568 6656
rect 3700 6647 3752 6656
rect 3700 6613 3709 6647
rect 3709 6613 3743 6647
rect 3743 6613 3752 6647
rect 3700 6604 3752 6613
rect 5080 6647 5132 6656
rect 5080 6613 5089 6647
rect 5089 6613 5123 6647
rect 5123 6613 5132 6647
rect 5080 6604 5132 6613
rect 6736 6604 6788 6656
rect 6920 6604 6972 6656
rect 7196 6740 7248 6792
rect 8208 6808 8260 6860
rect 10508 6876 10560 6928
rect 11244 6876 11296 6928
rect 11336 6876 11388 6928
rect 12256 6876 12308 6928
rect 10968 6808 11020 6860
rect 8392 6740 8444 6792
rect 8668 6672 8720 6724
rect 11888 6740 11940 6792
rect 12348 6740 12400 6792
rect 13176 6783 13228 6792
rect 13176 6749 13185 6783
rect 13185 6749 13219 6783
rect 13219 6749 13228 6783
rect 13176 6740 13228 6749
rect 14096 6783 14148 6792
rect 14096 6749 14105 6783
rect 14105 6749 14139 6783
rect 14139 6749 14148 6783
rect 14096 6740 14148 6749
rect 14372 6808 14424 6860
rect 14832 6944 14884 6996
rect 15660 6987 15712 6996
rect 15660 6953 15669 6987
rect 15669 6953 15703 6987
rect 15703 6953 15712 6987
rect 15660 6944 15712 6953
rect 16304 6987 16356 6996
rect 16304 6953 16313 6987
rect 16313 6953 16347 6987
rect 16347 6953 16356 6987
rect 16304 6944 16356 6953
rect 14924 6876 14976 6928
rect 14832 6851 14884 6860
rect 14832 6817 14841 6851
rect 14841 6817 14875 6851
rect 14875 6817 14884 6851
rect 14832 6808 14884 6817
rect 15384 6808 15436 6860
rect 15016 6740 15068 6792
rect 16304 6808 16356 6860
rect 13452 6672 13504 6724
rect 16856 6783 16908 6792
rect 16856 6749 16865 6783
rect 16865 6749 16899 6783
rect 16899 6749 16908 6783
rect 16856 6740 16908 6749
rect 8116 6604 8168 6656
rect 8484 6604 8536 6656
rect 9312 6604 9364 6656
rect 12256 6604 12308 6656
rect 12716 6604 12768 6656
rect 13912 6604 13964 6656
rect 14556 6604 14608 6656
rect 18052 6647 18104 6656
rect 18052 6613 18061 6647
rect 18061 6613 18095 6647
rect 18095 6613 18104 6647
rect 18052 6604 18104 6613
rect 3947 6502 3999 6554
rect 4011 6502 4063 6554
rect 4075 6502 4127 6554
rect 4139 6502 4191 6554
rect 9878 6502 9930 6554
rect 9942 6502 9994 6554
rect 10006 6502 10058 6554
rect 10070 6502 10122 6554
rect 15808 6502 15860 6554
rect 15872 6502 15924 6554
rect 15936 6502 15988 6554
rect 16000 6502 16052 6554
rect 4252 6400 4304 6452
rect 7472 6400 7524 6452
rect 7564 6400 7616 6452
rect 8208 6443 8260 6452
rect 4896 6332 4948 6384
rect 6828 6332 6880 6384
rect 8208 6409 8217 6443
rect 8217 6409 8251 6443
rect 8251 6409 8260 6443
rect 8208 6400 8260 6409
rect 11888 6400 11940 6452
rect 12440 6400 12492 6452
rect 13452 6400 13504 6452
rect 14648 6443 14700 6452
rect 11520 6332 11572 6384
rect 12992 6375 13044 6384
rect 12992 6341 13001 6375
rect 13001 6341 13035 6375
rect 13035 6341 13044 6375
rect 12992 6332 13044 6341
rect 13176 6332 13228 6384
rect 14648 6409 14657 6443
rect 14657 6409 14691 6443
rect 14691 6409 14700 6443
rect 14648 6400 14700 6409
rect 14924 6443 14976 6452
rect 14924 6409 14933 6443
rect 14933 6409 14967 6443
rect 14967 6409 14976 6443
rect 14924 6400 14976 6409
rect 1952 6264 2004 6316
rect 2964 6264 3016 6316
rect 3332 6264 3384 6316
rect 3700 6264 3752 6316
rect 2872 6196 2924 6248
rect 5540 6264 5592 6316
rect 6644 6264 6696 6316
rect 4160 6239 4212 6248
rect 4160 6205 4183 6239
rect 4183 6205 4212 6239
rect 2320 6128 2372 6180
rect 1400 6060 1452 6112
rect 3424 6128 3476 6180
rect 4160 6196 4212 6205
rect 5356 6196 5408 6248
rect 3976 6128 4028 6180
rect 7656 6196 7708 6248
rect 8484 6239 8536 6248
rect 8484 6205 8493 6239
rect 8493 6205 8527 6239
rect 8527 6205 8536 6239
rect 8484 6196 8536 6205
rect 8668 6264 8720 6316
rect 11244 6264 11296 6316
rect 10416 6196 10468 6248
rect 12716 6264 12768 6316
rect 15384 6332 15436 6384
rect 17224 6332 17276 6384
rect 12624 6196 12676 6248
rect 4988 6060 5040 6112
rect 5264 6103 5316 6112
rect 5264 6069 5273 6103
rect 5273 6069 5307 6103
rect 5307 6069 5316 6103
rect 5264 6060 5316 6069
rect 5908 6103 5960 6112
rect 5908 6069 5917 6103
rect 5917 6069 5951 6103
rect 5951 6069 5960 6103
rect 5908 6060 5960 6069
rect 7196 6128 7248 6180
rect 9772 6128 9824 6180
rect 11612 6128 11664 6180
rect 11980 6128 12032 6180
rect 12900 6128 12952 6180
rect 13360 6196 13412 6248
rect 14740 6196 14792 6248
rect 15568 6196 15620 6248
rect 13912 6128 13964 6180
rect 17040 6196 17092 6248
rect 17960 6196 18012 6248
rect 10416 6103 10468 6112
rect 10416 6069 10425 6103
rect 10425 6069 10459 6103
rect 10459 6069 10468 6103
rect 10416 6060 10468 6069
rect 11060 6060 11112 6112
rect 11336 6103 11388 6112
rect 11336 6069 11345 6103
rect 11345 6069 11379 6103
rect 11379 6069 11388 6103
rect 11336 6060 11388 6069
rect 12164 6060 12216 6112
rect 14832 6060 14884 6112
rect 16396 6060 16448 6112
rect 17592 6103 17644 6112
rect 17592 6069 17601 6103
rect 17601 6069 17635 6103
rect 17635 6069 17644 6103
rect 17592 6060 17644 6069
rect 17868 6060 17920 6112
rect 6912 5958 6964 6010
rect 6976 5958 7028 6010
rect 7040 5958 7092 6010
rect 7104 5958 7156 6010
rect 12843 5958 12895 6010
rect 12907 5958 12959 6010
rect 12971 5958 13023 6010
rect 13035 5958 13087 6010
rect 4344 5856 4396 5908
rect 6644 5856 6696 5908
rect 8116 5856 8168 5908
rect 11612 5856 11664 5908
rect 16304 5856 16356 5908
rect 1492 5720 1544 5772
rect 2320 5788 2372 5840
rect 5080 5788 5132 5840
rect 3056 5720 3108 5772
rect 4436 5763 4488 5772
rect 4436 5729 4445 5763
rect 4445 5729 4479 5763
rect 4479 5729 4488 5763
rect 4436 5720 4488 5729
rect 4712 5720 4764 5772
rect 7656 5720 7708 5772
rect 8576 5788 8628 5840
rect 4160 5652 4212 5704
rect 4896 5584 4948 5636
rect 2964 5559 3016 5568
rect 2964 5525 2973 5559
rect 2973 5525 3007 5559
rect 3007 5525 3016 5559
rect 2964 5516 3016 5525
rect 3792 5516 3844 5568
rect 4252 5516 4304 5568
rect 5080 5559 5132 5568
rect 5080 5525 5089 5559
rect 5089 5525 5123 5559
rect 5123 5525 5132 5559
rect 5080 5516 5132 5525
rect 7656 5627 7708 5636
rect 7656 5593 7665 5627
rect 7665 5593 7699 5627
rect 7699 5593 7708 5627
rect 9220 5720 9272 5772
rect 10508 5788 10560 5840
rect 10416 5720 10468 5772
rect 10968 5720 11020 5772
rect 15384 5788 15436 5840
rect 16304 5720 16356 5772
rect 17316 5763 17368 5772
rect 17316 5729 17325 5763
rect 17325 5729 17359 5763
rect 17359 5729 17368 5763
rect 17316 5720 17368 5729
rect 17408 5720 17460 5772
rect 7656 5584 7708 5593
rect 6644 5516 6696 5568
rect 7380 5516 7432 5568
rect 7748 5516 7800 5568
rect 9772 5516 9824 5568
rect 13544 5652 13596 5704
rect 14280 5652 14332 5704
rect 15108 5652 15160 5704
rect 15752 5695 15804 5704
rect 15752 5661 15761 5695
rect 15761 5661 15795 5695
rect 15795 5661 15804 5695
rect 15752 5652 15804 5661
rect 17500 5627 17552 5636
rect 17500 5593 17509 5627
rect 17509 5593 17543 5627
rect 17543 5593 17552 5627
rect 17500 5584 17552 5593
rect 11704 5516 11756 5568
rect 12624 5516 12676 5568
rect 13176 5559 13228 5568
rect 13176 5525 13185 5559
rect 13185 5525 13219 5559
rect 13219 5525 13228 5559
rect 13176 5516 13228 5525
rect 13820 5516 13872 5568
rect 17776 5516 17828 5568
rect 3947 5414 3999 5466
rect 4011 5414 4063 5466
rect 4075 5414 4127 5466
rect 4139 5414 4191 5466
rect 9878 5414 9930 5466
rect 9942 5414 9994 5466
rect 10006 5414 10058 5466
rect 10070 5414 10122 5466
rect 15808 5414 15860 5466
rect 15872 5414 15924 5466
rect 15936 5414 15988 5466
rect 16000 5414 16052 5466
rect 3516 5312 3568 5364
rect 7288 5312 7340 5364
rect 7564 5312 7616 5364
rect 9680 5355 9732 5364
rect 9680 5321 9689 5355
rect 9689 5321 9723 5355
rect 9723 5321 9732 5355
rect 9680 5312 9732 5321
rect 10600 5312 10652 5364
rect 13544 5312 13596 5364
rect 15384 5312 15436 5364
rect 3056 5244 3108 5296
rect 4252 5219 4304 5228
rect 4252 5185 4261 5219
rect 4261 5185 4295 5219
rect 4295 5185 4304 5219
rect 4252 5176 4304 5185
rect 5264 5244 5316 5296
rect 6460 5176 6512 5228
rect 9404 5244 9456 5296
rect 9864 5244 9916 5296
rect 13820 5244 13872 5296
rect 1492 5108 1544 5160
rect 2964 5040 3016 5092
rect 3516 5040 3568 5092
rect 4160 5151 4212 5160
rect 4160 5117 4169 5151
rect 4169 5117 4203 5151
rect 4203 5117 4212 5151
rect 4160 5108 4212 5117
rect 4712 5108 4764 5160
rect 4988 5040 5040 5092
rect 6000 5108 6052 5160
rect 6920 5151 6972 5160
rect 6920 5117 6929 5151
rect 6929 5117 6963 5151
rect 6963 5117 6972 5151
rect 6920 5108 6972 5117
rect 7748 5176 7800 5228
rect 8024 5176 8076 5228
rect 9128 5219 9180 5228
rect 9128 5185 9137 5219
rect 9137 5185 9171 5219
rect 9171 5185 9180 5219
rect 9128 5176 9180 5185
rect 2780 5015 2832 5024
rect 2780 4981 2789 5015
rect 2789 4981 2823 5015
rect 2823 4981 2832 5015
rect 2780 4972 2832 4981
rect 3424 4972 3476 5024
rect 4436 4972 4488 5024
rect 4620 4972 4672 5024
rect 4804 5015 4856 5024
rect 4804 4981 4813 5015
rect 4813 4981 4847 5015
rect 4847 4981 4856 5015
rect 4804 4972 4856 4981
rect 5172 5015 5224 5024
rect 5172 4981 5181 5015
rect 5181 4981 5215 5015
rect 5215 4981 5224 5015
rect 5172 4972 5224 4981
rect 6460 5040 6512 5092
rect 9220 5108 9272 5160
rect 11336 5176 11388 5228
rect 13176 5176 13228 5228
rect 13544 5219 13596 5228
rect 13544 5185 13553 5219
rect 13553 5185 13587 5219
rect 13587 5185 13596 5219
rect 13544 5176 13596 5185
rect 15108 5176 15160 5228
rect 10048 5108 10100 5160
rect 10692 5108 10744 5160
rect 11060 5151 11112 5160
rect 11060 5117 11069 5151
rect 11069 5117 11103 5151
rect 11103 5117 11112 5151
rect 11060 5108 11112 5117
rect 11428 5108 11480 5160
rect 12256 5108 12308 5160
rect 13912 5151 13964 5160
rect 13912 5117 13921 5151
rect 13921 5117 13955 5151
rect 13955 5117 13964 5151
rect 13912 5108 13964 5117
rect 16028 5151 16080 5160
rect 16028 5117 16037 5151
rect 16037 5117 16071 5151
rect 16071 5117 16080 5151
rect 16028 5108 16080 5117
rect 16580 5108 16632 5160
rect 12532 5040 12584 5092
rect 13176 5040 13228 5092
rect 14004 5040 14056 5092
rect 7748 4972 7800 5024
rect 9680 4972 9732 5024
rect 9772 4972 9824 5024
rect 10784 4972 10836 5024
rect 11428 4972 11480 5024
rect 13636 4972 13688 5024
rect 13728 4972 13780 5024
rect 15016 4972 15068 5024
rect 15292 4972 15344 5024
rect 15936 5015 15988 5024
rect 15936 4981 15945 5015
rect 15945 4981 15979 5015
rect 15979 4981 15988 5015
rect 15936 4972 15988 4981
rect 18236 5015 18288 5024
rect 18236 4981 18245 5015
rect 18245 4981 18279 5015
rect 18279 4981 18288 5015
rect 18236 4972 18288 4981
rect 6912 4870 6964 4922
rect 6976 4870 7028 4922
rect 7040 4870 7092 4922
rect 7104 4870 7156 4922
rect 12843 4870 12895 4922
rect 12907 4870 12959 4922
rect 12971 4870 13023 4922
rect 13035 4870 13087 4922
rect 3148 4768 3200 4820
rect 4712 4768 4764 4820
rect 5540 4768 5592 4820
rect 5908 4768 5960 4820
rect 9128 4768 9180 4820
rect 10232 4768 10284 4820
rect 10508 4768 10560 4820
rect 11428 4811 11480 4820
rect 11428 4777 11437 4811
rect 11437 4777 11471 4811
rect 11471 4777 11480 4811
rect 11428 4768 11480 4777
rect 13360 4811 13412 4820
rect 13360 4777 13369 4811
rect 13369 4777 13403 4811
rect 13403 4777 13412 4811
rect 13360 4768 13412 4777
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 15936 4768 15988 4820
rect 4804 4700 4856 4752
rect 5264 4700 5316 4752
rect 8116 4743 8168 4752
rect 3240 4632 3292 4684
rect 3424 4675 3476 4684
rect 3424 4641 3433 4675
rect 3433 4641 3467 4675
rect 3467 4641 3476 4675
rect 4344 4675 4396 4684
rect 3424 4632 3476 4641
rect 4344 4641 4378 4675
rect 4378 4641 4396 4675
rect 4344 4632 4396 4641
rect 4620 4632 4672 4684
rect 2964 4564 3016 4616
rect 3056 4496 3108 4548
rect 3424 4496 3476 4548
rect 5816 4632 5868 4684
rect 6184 4675 6236 4684
rect 6184 4641 6193 4675
rect 6193 4641 6227 4675
rect 6227 4641 6236 4675
rect 6184 4632 6236 4641
rect 8116 4709 8125 4743
rect 8125 4709 8159 4743
rect 8159 4709 8168 4743
rect 8116 4700 8168 4709
rect 9220 4700 9272 4752
rect 11336 4743 11388 4752
rect 7196 4607 7248 4616
rect 7196 4573 7205 4607
rect 7205 4573 7239 4607
rect 7239 4573 7248 4607
rect 7196 4564 7248 4573
rect 7288 4607 7340 4616
rect 7288 4573 7297 4607
rect 7297 4573 7331 4607
rect 7331 4573 7340 4607
rect 7288 4564 7340 4573
rect 8024 4632 8076 4684
rect 7932 4564 7984 4616
rect 8208 4607 8260 4616
rect 8208 4573 8217 4607
rect 8217 4573 8251 4607
rect 8251 4573 8260 4607
rect 8208 4564 8260 4573
rect 9864 4632 9916 4684
rect 10048 4675 10100 4684
rect 10048 4641 10057 4675
rect 10057 4641 10091 4675
rect 10091 4641 10100 4675
rect 10048 4632 10100 4641
rect 11336 4709 11345 4743
rect 11345 4709 11379 4743
rect 11379 4709 11388 4743
rect 11336 4700 11388 4709
rect 8484 4564 8536 4616
rect 9128 4564 9180 4616
rect 11520 4632 11572 4684
rect 12624 4700 12676 4752
rect 15200 4700 15252 4752
rect 8392 4496 8444 4548
rect 8668 4496 8720 4548
rect 11980 4607 12032 4616
rect 11980 4573 11989 4607
rect 11989 4573 12023 4607
rect 12023 4573 12032 4607
rect 11980 4564 12032 4573
rect 13176 4564 13228 4616
rect 15568 4700 15620 4752
rect 15752 4743 15804 4752
rect 15752 4709 15761 4743
rect 15761 4709 15795 4743
rect 15795 4709 15804 4743
rect 15752 4700 15804 4709
rect 15660 4675 15712 4684
rect 15660 4641 15669 4675
rect 15669 4641 15703 4675
rect 15703 4641 15712 4675
rect 15660 4632 15712 4641
rect 17040 4632 17092 4684
rect 17224 4632 17276 4684
rect 17868 4675 17920 4684
rect 17868 4641 17877 4675
rect 17877 4641 17911 4675
rect 17911 4641 17920 4675
rect 17868 4632 17920 4641
rect 14096 4607 14148 4616
rect 14096 4573 14105 4607
rect 14105 4573 14139 4607
rect 14139 4573 14148 4607
rect 14096 4564 14148 4573
rect 15108 4564 15160 4616
rect 13912 4496 13964 4548
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 2964 4471 3016 4480
rect 2964 4437 2973 4471
rect 2973 4437 3007 4471
rect 3007 4437 3016 4471
rect 2964 4428 3016 4437
rect 3240 4428 3292 4480
rect 9680 4428 9732 4480
rect 10876 4428 10928 4480
rect 11428 4428 11480 4480
rect 11980 4428 12032 4480
rect 13360 4428 13412 4480
rect 13820 4428 13872 4480
rect 15292 4471 15344 4480
rect 15292 4437 15301 4471
rect 15301 4437 15335 4471
rect 15335 4437 15344 4471
rect 15292 4428 15344 4437
rect 17500 4471 17552 4480
rect 17500 4437 17509 4471
rect 17509 4437 17543 4471
rect 17543 4437 17552 4471
rect 17500 4428 17552 4437
rect 17868 4428 17920 4480
rect 3947 4326 3999 4378
rect 4011 4326 4063 4378
rect 4075 4326 4127 4378
rect 4139 4326 4191 4378
rect 9878 4326 9930 4378
rect 9942 4326 9994 4378
rect 10006 4326 10058 4378
rect 10070 4326 10122 4378
rect 15808 4326 15860 4378
rect 15872 4326 15924 4378
rect 15936 4326 15988 4378
rect 16000 4326 16052 4378
rect 4988 4224 5040 4276
rect 5724 4224 5776 4276
rect 6000 4224 6052 4276
rect 7288 4156 7340 4208
rect 9220 4224 9272 4276
rect 10324 4224 10376 4276
rect 10876 4224 10928 4276
rect 1676 4020 1728 4072
rect 1952 4020 2004 4072
rect 3424 4020 3476 4072
rect 3700 4063 3752 4072
rect 3700 4029 3709 4063
rect 3709 4029 3743 4063
rect 3743 4029 3752 4063
rect 3700 4020 3752 4029
rect 7380 4088 7432 4140
rect 7656 4088 7708 4140
rect 11060 4088 11112 4140
rect 11612 4088 11664 4140
rect 12164 4156 12216 4208
rect 14004 4224 14056 4276
rect 15108 4156 15160 4208
rect 6736 4020 6788 4072
rect 10508 4020 10560 4072
rect 12072 4020 12124 4072
rect 13360 4063 13412 4072
rect 13360 4029 13369 4063
rect 13369 4029 13403 4063
rect 13403 4029 13412 4063
rect 13360 4020 13412 4029
rect 14464 4088 14516 4140
rect 14924 4088 14976 4140
rect 2780 3952 2832 4004
rect 4068 3952 4120 4004
rect 4896 3952 4948 4004
rect 8024 3995 8076 4004
rect 8024 3961 8058 3995
rect 8058 3961 8076 3995
rect 8024 3952 8076 3961
rect 8116 3952 8168 4004
rect 1676 3927 1728 3936
rect 1676 3893 1685 3927
rect 1685 3893 1719 3927
rect 1719 3893 1728 3927
rect 1676 3884 1728 3893
rect 3424 3927 3476 3936
rect 3424 3893 3433 3927
rect 3433 3893 3467 3927
rect 3467 3893 3476 3927
rect 3424 3884 3476 3893
rect 4344 3884 4396 3936
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 5632 3884 5684 3936
rect 6000 3884 6052 3936
rect 6092 3884 6144 3936
rect 9680 3884 9732 3936
rect 10048 3952 10100 4004
rect 11060 3927 11112 3936
rect 11060 3893 11069 3927
rect 11069 3893 11103 3927
rect 11103 3893 11112 3927
rect 11060 3884 11112 3893
rect 11336 3927 11388 3936
rect 11336 3893 11345 3927
rect 11345 3893 11379 3927
rect 11379 3893 11388 3927
rect 11336 3884 11388 3893
rect 12164 3952 12216 4004
rect 13636 3995 13688 4004
rect 13636 3961 13670 3995
rect 13670 3961 13688 3995
rect 13636 3952 13688 3961
rect 14372 3952 14424 4004
rect 14740 3952 14792 4004
rect 15384 3995 15436 4004
rect 15384 3961 15393 3995
rect 15393 3961 15427 3995
rect 15427 3961 15436 3995
rect 18144 4020 18196 4072
rect 15384 3952 15436 3961
rect 11888 3884 11940 3936
rect 12256 3884 12308 3936
rect 13728 3884 13780 3936
rect 14280 3884 14332 3936
rect 14832 3884 14884 3936
rect 17592 3927 17644 3936
rect 17592 3893 17601 3927
rect 17601 3893 17635 3927
rect 17635 3893 17644 3927
rect 17592 3884 17644 3893
rect 17776 3884 17828 3936
rect 6912 3782 6964 3834
rect 6976 3782 7028 3834
rect 7040 3782 7092 3834
rect 7104 3782 7156 3834
rect 12843 3782 12895 3834
rect 12907 3782 12959 3834
rect 12971 3782 13023 3834
rect 13035 3782 13087 3834
rect 2780 3680 2832 3732
rect 2964 3680 3016 3732
rect 3240 3680 3292 3732
rect 4528 3723 4580 3732
rect 4528 3689 4537 3723
rect 4537 3689 4571 3723
rect 4571 3689 4580 3723
rect 4528 3680 4580 3689
rect 6000 3680 6052 3732
rect 6644 3680 6696 3732
rect 3056 3655 3108 3664
rect 3056 3621 3065 3655
rect 3065 3621 3099 3655
rect 3099 3621 3108 3655
rect 3056 3612 3108 3621
rect 3700 3612 3752 3664
rect 5080 3612 5132 3664
rect 4436 3587 4488 3596
rect 3056 3476 3108 3528
rect 4436 3553 4445 3587
rect 4445 3553 4479 3587
rect 4479 3553 4488 3587
rect 4436 3544 4488 3553
rect 5540 3612 5592 3664
rect 5816 3612 5868 3664
rect 6460 3612 6512 3664
rect 8024 3680 8076 3732
rect 10048 3680 10100 3732
rect 11704 3680 11756 3732
rect 7380 3655 7432 3664
rect 7380 3621 7392 3655
rect 7392 3621 7432 3655
rect 7380 3612 7432 3621
rect 7564 3612 7616 3664
rect 14096 3680 14148 3732
rect 14188 3723 14240 3732
rect 14188 3689 14197 3723
rect 14197 3689 14231 3723
rect 14231 3689 14240 3723
rect 14188 3680 14240 3689
rect 7656 3544 7708 3596
rect 8300 3544 8352 3596
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 10508 3544 10560 3596
rect 11060 3544 11112 3596
rect 14004 3544 14056 3596
rect 14096 3587 14148 3596
rect 14096 3553 14105 3587
rect 14105 3553 14139 3587
rect 14139 3553 14148 3587
rect 14096 3544 14148 3553
rect 14832 3544 14884 3596
rect 14924 3544 14976 3596
rect 5264 3476 5316 3528
rect 4252 3408 4304 3460
rect 2872 3340 2924 3392
rect 3240 3340 3292 3392
rect 3608 3340 3660 3392
rect 6736 3340 6788 3392
rect 11980 3476 12032 3528
rect 13636 3408 13688 3460
rect 14464 3476 14516 3528
rect 16580 3544 16632 3596
rect 15200 3408 15252 3460
rect 16488 3408 16540 3460
rect 11612 3340 11664 3392
rect 14188 3340 14240 3392
rect 17316 3383 17368 3392
rect 17316 3349 17325 3383
rect 17325 3349 17359 3383
rect 17359 3349 17368 3383
rect 17316 3340 17368 3349
rect 3947 3238 3999 3290
rect 4011 3238 4063 3290
rect 4075 3238 4127 3290
rect 4139 3238 4191 3290
rect 9878 3238 9930 3290
rect 9942 3238 9994 3290
rect 10006 3238 10058 3290
rect 10070 3238 10122 3290
rect 15808 3238 15860 3290
rect 15872 3238 15924 3290
rect 15936 3238 15988 3290
rect 16000 3238 16052 3290
rect 9128 3136 9180 3188
rect 3332 3068 3384 3120
rect 4344 3068 4396 3120
rect 3424 3000 3476 3052
rect 7288 3068 7340 3120
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 8024 3000 8076 3052
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 9496 3043 9548 3052
rect 9496 3009 9505 3043
rect 9505 3009 9539 3043
rect 9539 3009 9548 3043
rect 11336 3068 11388 3120
rect 9496 3000 9548 3009
rect 11152 3000 11204 3052
rect 14280 3136 14332 3188
rect 14464 3179 14516 3188
rect 14464 3145 14473 3179
rect 14473 3145 14507 3179
rect 14507 3145 14516 3179
rect 14464 3136 14516 3145
rect 14740 3136 14792 3188
rect 14924 3068 14976 3120
rect 15568 3068 15620 3120
rect 11704 3000 11756 3052
rect 13452 3000 13504 3052
rect 13912 3000 13964 3052
rect 14096 3000 14148 3052
rect 1400 2975 1452 2984
rect 1400 2941 1409 2975
rect 1409 2941 1443 2975
rect 1443 2941 1452 2975
rect 1400 2932 1452 2941
rect 2136 2932 2188 2984
rect 2412 2932 2464 2984
rect 4804 2975 4856 2984
rect 4804 2941 4813 2975
rect 4813 2941 4847 2975
rect 4847 2941 4856 2975
rect 4804 2932 4856 2941
rect 5448 2932 5500 2984
rect 6276 2932 6328 2984
rect 7472 2932 7524 2984
rect 7840 2932 7892 2984
rect 8116 2932 8168 2984
rect 1952 2864 2004 2916
rect 2688 2864 2740 2916
rect 3884 2864 3936 2916
rect 1400 2796 1452 2848
rect 1768 2796 1820 2848
rect 3148 2839 3200 2848
rect 3148 2805 3157 2839
rect 3157 2805 3191 2839
rect 3191 2805 3200 2839
rect 3148 2796 3200 2805
rect 6000 2864 6052 2916
rect 9312 2864 9364 2916
rect 11796 2932 11848 2984
rect 13820 2932 13872 2984
rect 11152 2864 11204 2916
rect 5448 2839 5500 2848
rect 5448 2805 5457 2839
rect 5457 2805 5491 2839
rect 5491 2805 5500 2839
rect 5448 2796 5500 2805
rect 6368 2796 6420 2848
rect 8852 2839 8904 2848
rect 8852 2805 8861 2839
rect 8861 2805 8895 2839
rect 8895 2805 8904 2839
rect 8852 2796 8904 2805
rect 9588 2796 9640 2848
rect 10048 2839 10100 2848
rect 10048 2805 10057 2839
rect 10057 2805 10091 2839
rect 10091 2805 10100 2839
rect 10048 2796 10100 2805
rect 11060 2839 11112 2848
rect 11060 2805 11069 2839
rect 11069 2805 11103 2839
rect 11103 2805 11112 2839
rect 11060 2796 11112 2805
rect 13268 2796 13320 2848
rect 14004 2864 14056 2916
rect 14188 2932 14240 2984
rect 14740 2932 14792 2984
rect 14832 2932 14884 2984
rect 15476 2975 15528 2984
rect 15476 2941 15485 2975
rect 15485 2941 15519 2975
rect 15519 2941 15528 2975
rect 15476 2932 15528 2941
rect 15568 2932 15620 2984
rect 14924 2907 14976 2916
rect 13728 2796 13780 2848
rect 14648 2796 14700 2848
rect 14924 2873 14933 2907
rect 14933 2873 14967 2907
rect 14967 2873 14976 2907
rect 14924 2864 14976 2873
rect 16672 2864 16724 2916
rect 16396 2796 16448 2848
rect 16580 2839 16632 2848
rect 16580 2805 16589 2839
rect 16589 2805 16623 2839
rect 16623 2805 16632 2839
rect 16580 2796 16632 2805
rect 17224 2796 17276 2848
rect 18236 2839 18288 2848
rect 18236 2805 18245 2839
rect 18245 2805 18279 2839
rect 18279 2805 18288 2839
rect 18236 2796 18288 2805
rect 6912 2694 6964 2746
rect 6976 2694 7028 2746
rect 7040 2694 7092 2746
rect 7104 2694 7156 2746
rect 12843 2694 12895 2746
rect 12907 2694 12959 2746
rect 12971 2694 13023 2746
rect 13035 2694 13087 2746
rect 3332 2635 3384 2644
rect 3332 2601 3341 2635
rect 3341 2601 3375 2635
rect 3375 2601 3384 2635
rect 3332 2592 3384 2601
rect 4436 2592 4488 2644
rect 3148 2524 3200 2576
rect 5448 2592 5500 2644
rect 9036 2635 9088 2644
rect 9036 2601 9045 2635
rect 9045 2601 9079 2635
rect 9079 2601 9088 2635
rect 9036 2592 9088 2601
rect 11060 2592 11112 2644
rect 12348 2592 12400 2644
rect 12440 2592 12492 2644
rect 13360 2592 13412 2644
rect 14004 2635 14056 2644
rect 6000 2524 6052 2576
rect 6552 2524 6604 2576
rect 8852 2524 8904 2576
rect 10048 2524 10100 2576
rect 10324 2524 10376 2576
rect 13084 2567 13136 2576
rect 13084 2533 13093 2567
rect 13093 2533 13127 2567
rect 13127 2533 13136 2567
rect 13084 2524 13136 2533
rect 1400 2456 1452 2508
rect 3884 2456 3936 2508
rect 5724 2499 5776 2508
rect 5724 2465 5733 2499
rect 5733 2465 5767 2499
rect 5767 2465 5776 2499
rect 5724 2456 5776 2465
rect 7288 2456 7340 2508
rect 8668 2456 8720 2508
rect 10968 2456 11020 2508
rect 1216 2388 1268 2440
rect 4344 2388 4396 2440
rect 5540 2388 5592 2440
rect 5632 2388 5684 2440
rect 9312 2431 9364 2440
rect 9312 2397 9321 2431
rect 9321 2397 9355 2431
rect 9355 2397 9364 2431
rect 9312 2388 9364 2397
rect 11428 2456 11480 2508
rect 13544 2524 13596 2576
rect 14004 2601 14013 2635
rect 14013 2601 14047 2635
rect 14047 2601 14056 2635
rect 14004 2592 14056 2601
rect 15292 2592 15344 2644
rect 14372 2524 14424 2576
rect 13636 2456 13688 2508
rect 8760 2320 8812 2372
rect 11152 2320 11204 2372
rect 2780 2252 2832 2304
rect 7656 2295 7708 2304
rect 7656 2261 7665 2295
rect 7665 2261 7699 2295
rect 7699 2261 7708 2295
rect 7656 2252 7708 2261
rect 10416 2252 10468 2304
rect 13452 2388 13504 2440
rect 14188 2431 14240 2440
rect 14188 2397 14197 2431
rect 14197 2397 14231 2431
rect 14231 2397 14240 2431
rect 14188 2388 14240 2397
rect 14556 2456 14608 2508
rect 16396 2524 16448 2576
rect 16212 2499 16264 2508
rect 16212 2465 16221 2499
rect 16221 2465 16255 2499
rect 16255 2465 16264 2499
rect 16212 2456 16264 2465
rect 16672 2456 16724 2508
rect 17132 2456 17184 2508
rect 17684 2499 17736 2508
rect 17684 2465 17693 2499
rect 17693 2465 17727 2499
rect 17727 2465 17736 2499
rect 17684 2456 17736 2465
rect 13820 2320 13872 2372
rect 13912 2320 13964 2372
rect 13084 2252 13136 2304
rect 17132 2295 17184 2304
rect 17132 2261 17141 2295
rect 17141 2261 17175 2295
rect 17175 2261 17184 2295
rect 17132 2252 17184 2261
rect 17868 2295 17920 2304
rect 17868 2261 17877 2295
rect 17877 2261 17911 2295
rect 17911 2261 17920 2295
rect 17868 2252 17920 2261
rect 3947 2150 3999 2202
rect 4011 2150 4063 2202
rect 4075 2150 4127 2202
rect 4139 2150 4191 2202
rect 9878 2150 9930 2202
rect 9942 2150 9994 2202
rect 10006 2150 10058 2202
rect 10070 2150 10122 2202
rect 15808 2150 15860 2202
rect 15872 2150 15924 2202
rect 15936 2150 15988 2202
rect 16000 2150 16052 2202
rect 388 2048 440 2100
rect 17132 2048 17184 2100
rect 7656 1912 7708 1964
rect 16304 1776 16356 1828
rect 3976 1368 4028 1420
rect 5632 1368 5684 1420
rect 11244 1368 11296 1420
rect 13636 1368 13688 1420
<< metal2 >>
rect 1122 16200 1178 17000
rect 3330 16200 3386 17000
rect 4066 16280 4122 16289
rect 4066 16215 4122 16224
rect 1136 12753 1164 16200
rect 2778 15872 2834 15881
rect 2778 15807 2834 15816
rect 1122 12744 1178 12753
rect 1122 12679 1178 12688
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 2134 12200 2190 12209
rect 2134 12135 2190 12144
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 1492 11552 1544 11558
rect 1492 11494 1544 11500
rect 1308 11144 1360 11150
rect 1308 11086 1360 11092
rect 1320 10266 1348 11086
rect 1400 11076 1452 11082
rect 1400 11018 1452 11024
rect 1308 10260 1360 10266
rect 1308 10202 1360 10208
rect 1320 10062 1348 10202
rect 1308 10056 1360 10062
rect 1308 9998 1360 10004
rect 1320 9586 1348 9998
rect 1308 9580 1360 9586
rect 1308 9522 1360 9528
rect 1320 8498 1348 9522
rect 1308 8492 1360 8498
rect 1308 8434 1360 8440
rect 1412 7585 1440 11018
rect 1504 7993 1532 11494
rect 1688 11257 1716 11630
rect 1674 11248 1730 11257
rect 1674 11183 1730 11192
rect 1872 9178 1900 12038
rect 2148 11354 2176 12135
rect 2240 11898 2268 12242
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2332 10810 2360 12174
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2424 11370 2452 11698
rect 2516 11694 2544 12582
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2424 11342 2544 11370
rect 2516 11218 2544 11342
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2516 10674 2544 11154
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2608 10198 2636 12174
rect 2686 11656 2742 11665
rect 2686 11591 2688 11600
rect 2740 11591 2742 11600
rect 2688 11562 2740 11568
rect 2700 11286 2728 11562
rect 2688 11280 2740 11286
rect 2688 11222 2740 11228
rect 2792 10538 2820 15807
rect 3344 14090 3372 16200
rect 3974 15464 4030 15473
rect 3974 15399 4030 15408
rect 3988 15366 4016 15399
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 4080 15298 4108 16215
rect 5538 16200 5594 17000
rect 7746 16200 7802 17000
rect 8390 16688 8446 16697
rect 8390 16623 8446 16632
rect 4068 15292 4120 15298
rect 4068 15234 4120 15240
rect 3514 15056 3570 15065
rect 3514 14991 3516 15000
rect 3568 14991 3570 15000
rect 3516 14962 3568 14968
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3712 14249 3740 14758
rect 4434 14648 4490 14657
rect 4434 14583 4490 14592
rect 3792 14544 3844 14550
rect 3792 14486 3844 14492
rect 3698 14240 3754 14249
rect 3698 14175 3754 14184
rect 3344 14074 3464 14090
rect 3344 14068 3476 14074
rect 3344 14062 3424 14068
rect 3424 14010 3476 14016
rect 3332 14000 3384 14006
rect 3332 13942 3384 13948
rect 3344 12442 3372 13942
rect 3804 13841 3832 14486
rect 3921 14172 4217 14192
rect 3977 14170 4001 14172
rect 4057 14170 4081 14172
rect 4137 14170 4161 14172
rect 3999 14118 4001 14170
rect 4063 14118 4075 14170
rect 4137 14118 4139 14170
rect 3977 14116 4001 14118
rect 4057 14116 4081 14118
rect 4137 14116 4161 14118
rect 3921 14096 4217 14116
rect 3790 13832 3846 13841
rect 3790 13767 3846 13776
rect 4066 13424 4122 13433
rect 4066 13359 4122 13368
rect 4080 13326 4108 13359
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 3921 13084 4217 13104
rect 3977 13082 4001 13084
rect 4057 13082 4081 13084
rect 4137 13082 4161 13084
rect 3999 13030 4001 13082
rect 4063 13030 4075 13082
rect 4137 13030 4139 13082
rect 3977 13028 4001 13030
rect 4057 13028 4081 13030
rect 4137 13028 4161 13030
rect 3514 13016 3570 13025
rect 3921 13008 4217 13028
rect 3514 12951 3516 12960
rect 3568 12951 3570 12960
rect 3516 12922 3568 12928
rect 3700 12776 3752 12782
rect 3700 12718 3752 12724
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 3712 12238 3740 12718
rect 3988 12617 4016 12718
rect 4160 12640 4212 12646
rect 3974 12608 4030 12617
rect 4160 12582 4212 12588
rect 3974 12543 4030 12552
rect 4172 12306 4200 12582
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 3700 12232 3752 12238
rect 2962 12200 3018 12209
rect 3700 12174 3752 12180
rect 2962 12135 2964 12144
rect 3016 12135 3018 12144
rect 2964 12106 3016 12112
rect 3712 11694 3740 12174
rect 4172 12084 4200 12242
rect 4172 12056 4292 12084
rect 3921 11996 4217 12016
rect 3977 11994 4001 11996
rect 4057 11994 4081 11996
rect 4137 11994 4161 11996
rect 3999 11942 4001 11994
rect 4063 11942 4075 11994
rect 4137 11942 4139 11994
rect 3977 11940 4001 11942
rect 4057 11940 4081 11942
rect 4137 11940 4161 11942
rect 3921 11920 4217 11940
rect 3882 11792 3938 11801
rect 3882 11727 3938 11736
rect 3896 11694 3924 11727
rect 3700 11688 3752 11694
rect 3700 11630 3752 11636
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2780 10532 2832 10538
rect 2780 10474 2832 10480
rect 2596 10192 2648 10198
rect 2596 10134 2648 10140
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2792 9518 2820 9862
rect 2870 9752 2926 9761
rect 2870 9687 2926 9696
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 2792 8974 2820 9454
rect 2780 8968 2832 8974
rect 2502 8936 2558 8945
rect 2780 8910 2832 8916
rect 2502 8871 2558 8880
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1490 7984 1546 7993
rect 1490 7919 1546 7928
rect 1398 7576 1454 7585
rect 1398 7511 1454 7520
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1412 2990 1440 6054
rect 1492 5772 1544 5778
rect 1492 5714 1544 5720
rect 1504 5166 1532 5714
rect 1492 5160 1544 5166
rect 1492 5102 1544 5108
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1400 2984 1452 2990
rect 1400 2926 1452 2932
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1412 2514 1440 2790
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1216 2440 1268 2446
rect 1216 2382 1268 2388
rect 388 2100 440 2106
rect 388 2042 440 2048
rect 400 800 428 2042
rect 1228 800 1256 2382
rect 1596 1873 1624 4422
rect 1688 4078 1716 7278
rect 1676 4072 1728 4078
rect 1676 4014 1728 4020
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1582 1864 1638 1873
rect 1582 1799 1638 1808
rect 1688 1465 1716 3878
rect 1780 2854 1808 8774
rect 2516 8430 2544 8871
rect 2884 8480 2912 9687
rect 2608 8452 2912 8480
rect 2504 8424 2556 8430
rect 2424 8384 2504 8412
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1858 7032 1914 7041
rect 1858 6967 1914 6976
rect 1872 6866 1900 6967
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 1964 6322 1992 7686
rect 2332 7546 2360 7890
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 2332 6798 2360 7142
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 2332 6186 2360 6734
rect 2320 6180 2372 6186
rect 2320 6122 2372 6128
rect 2332 5846 2360 6122
rect 2320 5840 2372 5846
rect 2320 5782 2372 5788
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 1964 2922 1992 4014
rect 2424 2990 2452 8384
rect 2504 8366 2556 8372
rect 2608 7732 2636 8452
rect 2976 8401 3004 11494
rect 3712 11150 3740 11630
rect 4264 11626 4292 12056
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 3790 11384 3846 11393
rect 3790 11319 3846 11328
rect 3700 11144 3752 11150
rect 3700 11086 3752 11092
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3252 10198 3280 11018
rect 3516 11008 3568 11014
rect 3514 10976 3516 10985
rect 3568 10976 3570 10985
rect 3514 10911 3570 10920
rect 3332 10736 3384 10742
rect 3332 10678 3384 10684
rect 3240 10192 3292 10198
rect 3240 10134 3292 10140
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 2962 8392 3018 8401
rect 2688 8356 2740 8362
rect 2962 8327 3018 8336
rect 2688 8298 2740 8304
rect 2700 7954 2728 8298
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2884 7886 2912 8230
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2780 7812 2832 7818
rect 2780 7754 2832 7760
rect 2688 7744 2740 7750
rect 2608 7704 2688 7732
rect 2688 7686 2740 7692
rect 2596 7472 2648 7478
rect 2516 7432 2596 7460
rect 2516 3505 2544 7432
rect 2596 7414 2648 7420
rect 2594 6896 2650 6905
rect 2594 6831 2650 6840
rect 2502 3496 2558 3505
rect 2502 3431 2558 3440
rect 2608 3097 2636 6831
rect 2594 3088 2650 3097
rect 2594 3023 2650 3032
rect 2136 2984 2188 2990
rect 2136 2926 2188 2932
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 1952 2916 2004 2922
rect 1952 2858 2004 2864
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 1674 1456 1730 1465
rect 1674 1391 1730 1400
rect 2148 800 2176 2926
rect 2700 2922 2728 7686
rect 2792 6905 2820 7754
rect 2884 7274 2912 7822
rect 2872 7268 2924 7274
rect 2872 7210 2924 7216
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 2778 6896 2834 6905
rect 2778 6831 2834 6840
rect 2884 6254 2912 6938
rect 2976 6866 3004 7142
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2976 6322 3004 6802
rect 3068 6361 3096 9862
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3054 6352 3110 6361
rect 2964 6316 3016 6322
rect 3054 6287 3110 6296
rect 2964 6258 3016 6264
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 3160 5794 3188 9318
rect 3252 8974 3280 10134
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3344 8378 3372 10678
rect 3606 10568 3662 10577
rect 3606 10503 3662 10512
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3436 9178 3464 10406
rect 3620 9722 3648 10503
rect 3712 10266 3740 11086
rect 3804 10554 3832 11319
rect 3921 10908 4217 10928
rect 3977 10906 4001 10908
rect 4057 10906 4081 10908
rect 4137 10906 4161 10908
rect 3999 10854 4001 10906
rect 4063 10854 4075 10906
rect 4137 10854 4139 10906
rect 3977 10852 4001 10854
rect 4057 10852 4081 10854
rect 4137 10852 4161 10854
rect 3921 10832 4217 10852
rect 4066 10704 4122 10713
rect 4066 10639 4122 10648
rect 3804 10526 3924 10554
rect 4080 10538 4108 10639
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3804 10266 3832 10406
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 3608 9716 3660 9722
rect 3608 9658 3660 9664
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3528 9110 3556 9318
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3424 8560 3476 8566
rect 3424 8502 3476 8508
rect 3252 8350 3372 8378
rect 3252 5930 3280 8350
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3344 8090 3372 8230
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3344 7750 3372 7890
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3332 7268 3384 7274
rect 3332 7210 3384 7216
rect 3344 6322 3372 7210
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3436 6186 3464 8502
rect 3528 8498 3556 9046
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3620 6769 3648 9318
rect 3712 8974 3740 10202
rect 3896 9908 3924 10526
rect 4068 10532 4120 10538
rect 4068 10474 4120 10480
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 3804 9880 3924 9908
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3606 6760 3662 6769
rect 3712 6746 3740 7686
rect 3804 7342 3832 9880
rect 3921 9820 4217 9840
rect 3977 9818 4001 9820
rect 4057 9818 4081 9820
rect 4137 9818 4161 9820
rect 3999 9766 4001 9818
rect 4063 9766 4075 9818
rect 4137 9766 4139 9818
rect 3977 9764 4001 9766
rect 4057 9764 4081 9766
rect 4137 9764 4161 9766
rect 3921 9744 4217 9764
rect 4356 9654 4384 10406
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 4080 9353 4108 9522
rect 4066 9344 4122 9353
rect 4066 9279 4122 9288
rect 4080 8922 4108 9279
rect 4080 8894 4384 8922
rect 3921 8732 4217 8752
rect 3977 8730 4001 8732
rect 4057 8730 4081 8732
rect 4137 8730 4161 8732
rect 3999 8678 4001 8730
rect 4063 8678 4075 8730
rect 4137 8678 4139 8730
rect 3977 8676 4001 8678
rect 4057 8676 4081 8678
rect 4137 8676 4161 8678
rect 3921 8656 4217 8676
rect 4250 8528 4306 8537
rect 4250 8463 4306 8472
rect 4264 8430 4292 8463
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3988 7954 4016 8230
rect 4080 7993 4108 8298
rect 4066 7984 4122 7993
rect 3976 7948 4028 7954
rect 4066 7919 4122 7928
rect 3976 7890 4028 7896
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 3921 7644 4217 7664
rect 3977 7642 4001 7644
rect 4057 7642 4081 7644
rect 4137 7642 4161 7644
rect 3999 7590 4001 7642
rect 4063 7590 4075 7642
rect 4137 7590 4139 7642
rect 3977 7588 4001 7590
rect 4057 7588 4081 7590
rect 4137 7588 4161 7590
rect 3921 7568 4217 7588
rect 4264 7478 4292 7822
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3804 6866 3832 7278
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 3712 6718 3832 6746
rect 3606 6695 3662 6704
rect 3516 6656 3568 6662
rect 3700 6656 3752 6662
rect 3568 6616 3648 6644
rect 3516 6598 3568 6604
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3252 5902 3464 5930
rect 3056 5772 3108 5778
rect 3160 5766 3372 5794
rect 3056 5714 3108 5720
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2976 5098 3004 5510
rect 3068 5302 3096 5714
rect 3056 5296 3108 5302
rect 3056 5238 3108 5244
rect 2964 5092 3016 5098
rect 2964 5034 3016 5040
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2792 4010 2820 4966
rect 2976 4622 3004 5034
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2780 4004 2832 4010
rect 2780 3946 2832 3952
rect 2792 3738 2820 3946
rect 2976 3738 3004 4422
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 3068 3670 3096 4490
rect 3160 3720 3188 4762
rect 3344 4729 3372 5766
rect 3436 5137 3464 5902
rect 3514 5536 3570 5545
rect 3514 5471 3570 5480
rect 3528 5370 3556 5471
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3422 5128 3478 5137
rect 3422 5063 3478 5072
rect 3516 5092 3568 5098
rect 3516 5034 3568 5040
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3330 4720 3386 4729
rect 3240 4684 3292 4690
rect 3436 4690 3464 4966
rect 3330 4655 3386 4664
rect 3424 4684 3476 4690
rect 3240 4626 3292 4632
rect 3424 4626 3476 4632
rect 3252 4486 3280 4626
rect 3424 4548 3476 4554
rect 3424 4490 3476 4496
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3436 4078 3464 4490
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 3240 3732 3292 3738
rect 3160 3692 3240 3720
rect 3240 3674 3292 3680
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 2688 2916 2740 2922
rect 2688 2858 2740 2864
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 386 0 442 800
rect 1214 0 1270 800
rect 2134 0 2190 800
rect 2792 649 2820 2246
rect 2884 1057 2912 3334
rect 2870 1048 2926 1057
rect 2870 983 2926 992
rect 3068 800 3096 3470
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 3160 2582 3188 2790
rect 3252 2689 3280 3334
rect 3332 3120 3384 3126
rect 3332 3062 3384 3068
rect 3238 2680 3294 2689
rect 3344 2650 3372 3062
rect 3436 3058 3464 3878
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 3238 2615 3294 2624
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3148 2576 3200 2582
rect 3148 2518 3200 2524
rect 2778 640 2834 649
rect 2778 575 2834 584
rect 3054 0 3110 800
rect 3528 241 3556 5034
rect 3620 3398 3648 6616
rect 3700 6598 3752 6604
rect 3712 6322 3740 6598
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3804 5658 3832 6718
rect 3921 6556 4217 6576
rect 3977 6554 4001 6556
rect 4057 6554 4081 6556
rect 4137 6554 4161 6556
rect 3999 6502 4001 6554
rect 4063 6502 4075 6554
rect 4137 6502 4139 6554
rect 3977 6500 4001 6502
rect 4057 6500 4081 6502
rect 4137 6500 4161 6502
rect 3921 6480 4217 6500
rect 4264 6458 4292 6802
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 3988 5953 4016 6122
rect 3974 5944 4030 5953
rect 3974 5879 4030 5888
rect 4172 5710 4200 6190
rect 4356 5914 4384 8894
rect 4448 8362 4476 14583
rect 5552 14498 5580 16200
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6276 15020 6328 15026
rect 6276 14962 6328 14968
rect 5552 14470 5948 14498
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5080 13388 5132 13394
rect 5080 13330 5132 13336
rect 5092 12850 5120 13330
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 5460 12714 5488 13874
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5552 13530 5580 13670
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5644 12986 5672 13670
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5460 12102 5488 12650
rect 5448 12096 5500 12102
rect 5446 12064 5448 12073
rect 5500 12064 5502 12073
rect 5446 11999 5502 12008
rect 5736 11914 5764 14214
rect 5816 13320 5868 13326
rect 5920 13297 5948 14470
rect 6184 13320 6236 13326
rect 5816 13262 5868 13268
rect 5906 13288 5962 13297
rect 5644 11886 5764 11914
rect 5080 11688 5132 11694
rect 5080 11630 5132 11636
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4816 10470 4844 10746
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4434 7440 4490 7449
rect 4434 7375 4490 7384
rect 4448 7342 4476 7375
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 3712 5630 3832 5658
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 3712 4321 3740 5630
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 3698 4312 3754 4321
rect 3698 4247 3754 4256
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3712 3670 3740 4014
rect 3700 3664 3752 3670
rect 3700 3606 3752 3612
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3698 2272 3754 2281
rect 3804 2258 3832 5510
rect 3921 5468 4217 5488
rect 3977 5466 4001 5468
rect 4057 5466 4081 5468
rect 4137 5466 4161 5468
rect 3999 5414 4001 5466
rect 4063 5414 4075 5466
rect 4137 5414 4139 5466
rect 3977 5412 4001 5414
rect 4057 5412 4081 5414
rect 4137 5412 4161 5414
rect 3921 5392 4217 5412
rect 4158 5264 4214 5273
rect 4264 5234 4292 5510
rect 4158 5199 4214 5208
rect 4252 5228 4304 5234
rect 4172 5166 4200 5199
rect 4252 5170 4304 5176
rect 4160 5160 4212 5166
rect 4448 5114 4476 5714
rect 4160 5102 4212 5108
rect 4264 5086 4476 5114
rect 3921 4380 4217 4400
rect 3977 4378 4001 4380
rect 4057 4378 4081 4380
rect 4137 4378 4161 4380
rect 3999 4326 4001 4378
rect 4063 4326 4075 4378
rect 4137 4326 4139 4378
rect 3977 4324 4001 4326
rect 4057 4324 4081 4326
rect 4137 4324 4161 4326
rect 3921 4304 4217 4324
rect 4068 4004 4120 4010
rect 4068 3946 4120 3952
rect 4080 3913 4108 3946
rect 4066 3904 4122 3913
rect 4066 3839 4122 3848
rect 4264 3466 4292 5086
rect 4448 5030 4476 5086
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4540 4729 4568 9454
rect 4632 6798 4660 9998
rect 4816 9994 4844 10406
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 4894 10160 4950 10169
rect 4894 10095 4896 10104
rect 4948 10095 4950 10104
rect 4896 10066 4948 10072
rect 5000 10033 5028 10202
rect 4986 10024 5042 10033
rect 4804 9988 4856 9994
rect 4986 9959 5042 9968
rect 4804 9930 4856 9936
rect 4710 9888 4766 9897
rect 4710 9823 4766 9832
rect 4724 9382 4752 9823
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4632 5681 4660 6734
rect 4724 5778 4752 9318
rect 5092 9081 5120 11630
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 5184 11218 5212 11494
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5184 10674 5212 11154
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5184 10062 5212 10610
rect 5276 10470 5304 10950
rect 5368 10674 5396 10950
rect 5460 10674 5488 11018
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5184 9586 5212 9998
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5078 9072 5134 9081
rect 5078 9007 5134 9016
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 5000 8498 5028 8774
rect 5092 8616 5120 9007
rect 5092 8588 5212 8616
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 4816 8022 4844 8366
rect 4804 8016 4856 8022
rect 4804 7958 4856 7964
rect 4816 7546 4844 7958
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 4908 7342 4936 7890
rect 5000 7478 5028 8434
rect 4988 7472 5040 7478
rect 4988 7414 5040 7420
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4908 6644 4936 7278
rect 5000 6798 5028 7414
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 5080 6656 5132 6662
rect 4908 6616 5028 6644
rect 4896 6384 4948 6390
rect 4896 6326 4948 6332
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4618 5672 4674 5681
rect 4908 5642 4936 6326
rect 5000 6118 5028 6616
rect 5080 6598 5132 6604
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4618 5607 4674 5616
rect 4896 5636 4948 5642
rect 4896 5578 4948 5584
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4526 4720 4582 4729
rect 4344 4684 4396 4690
rect 4632 4690 4660 4966
rect 4724 4826 4752 5102
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4816 4758 4844 4966
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4526 4655 4582 4664
rect 4620 4684 4672 4690
rect 4344 4626 4396 4632
rect 4356 3942 4384 4626
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4252 3460 4304 3466
rect 4252 3402 4304 3408
rect 3921 3292 4217 3312
rect 3977 3290 4001 3292
rect 4057 3290 4081 3292
rect 4137 3290 4161 3292
rect 3999 3238 4001 3290
rect 4063 3238 4075 3290
rect 4137 3238 4139 3290
rect 3977 3236 4001 3238
rect 4057 3236 4081 3238
rect 4137 3236 4161 3238
rect 3921 3216 4217 3236
rect 4356 3126 4384 3878
rect 4540 3738 4568 4655
rect 4620 4626 4672 4632
rect 4908 4570 4936 5578
rect 5000 5556 5028 6054
rect 5092 5846 5120 6598
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 5080 5568 5132 5574
rect 5000 5528 5080 5556
rect 5080 5510 5132 5516
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 4816 4542 4936 4570
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 3882 2952 3938 2961
rect 3882 2887 3884 2896
rect 3936 2887 3938 2896
rect 3884 2858 3936 2864
rect 3896 2514 3924 2858
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 4356 2446 4384 3062
rect 4448 2650 4476 3538
rect 4816 2990 4844 4542
rect 5000 4282 5028 5034
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 3754 2230 3832 2258
rect 3698 2207 3754 2216
rect 3921 2204 4217 2224
rect 3977 2202 4001 2204
rect 4057 2202 4081 2204
rect 4137 2202 4161 2204
rect 3999 2150 4001 2202
rect 4063 2150 4075 2202
rect 4137 2150 4139 2202
rect 3977 2148 4001 2150
rect 4057 2148 4081 2150
rect 4137 2148 4161 2150
rect 3921 2128 4217 2148
rect 3976 1420 4028 1426
rect 3976 1362 4028 1368
rect 3988 800 4016 1362
rect 4908 800 4936 3946
rect 5092 3670 5120 5510
rect 5184 5030 5212 8588
rect 5276 7721 5304 10406
rect 5354 10160 5410 10169
rect 5354 10095 5410 10104
rect 5368 9722 5396 10095
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5368 8922 5396 9658
rect 5460 9042 5488 10406
rect 5552 10266 5580 10542
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5368 8894 5488 8922
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 5262 7712 5318 7721
rect 5262 7647 5318 7656
rect 5368 7177 5396 8502
rect 5354 7168 5410 7177
rect 5354 7103 5410 7112
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5276 5302 5304 6054
rect 5264 5296 5316 5302
rect 5264 5238 5316 5244
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5276 4758 5304 5238
rect 5264 4752 5316 4758
rect 5264 4694 5316 4700
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 5276 3534 5304 4694
rect 5368 3942 5396 6190
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5460 2990 5488 8894
rect 5552 7342 5580 9930
rect 5644 8809 5672 11886
rect 5828 10470 5856 13262
rect 6184 13262 6236 13268
rect 5906 13223 5962 13232
rect 6092 12912 6144 12918
rect 5998 12880 6054 12889
rect 6092 12854 6144 12860
rect 5920 12824 5998 12832
rect 5920 12804 6000 12824
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5724 10124 5776 10130
rect 5724 10066 5776 10072
rect 5630 8800 5686 8809
rect 5630 8735 5686 8744
rect 5736 8634 5764 10066
rect 5828 9722 5856 10406
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5920 9489 5948 12804
rect 6052 12815 6054 12824
rect 6000 12786 6052 12792
rect 6000 11552 6052 11558
rect 6104 11540 6132 12854
rect 6196 12850 6224 13262
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 6196 12374 6224 12786
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 6196 11762 6224 12310
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6052 11512 6132 11540
rect 6000 11494 6052 11500
rect 5906 9480 5962 9489
rect 5906 9415 5908 9424
rect 5960 9415 5962 9424
rect 5908 9386 5960 9392
rect 5816 9376 5868 9382
rect 5920 9355 5948 9386
rect 5816 9318 5868 9324
rect 5828 9110 5856 9318
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5920 8922 5948 9114
rect 5828 8894 5948 8922
rect 5724 8628 5776 8634
rect 5644 8588 5724 8616
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5552 7041 5580 7278
rect 5538 7032 5594 7041
rect 5538 6967 5594 6976
rect 5644 6866 5672 8588
rect 5724 8570 5776 8576
rect 5724 8356 5776 8362
rect 5724 8298 5776 8304
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5552 4826 5580 6258
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5552 3670 5580 4762
rect 5630 4584 5686 4593
rect 5736 4570 5764 8298
rect 5828 5545 5856 8894
rect 5906 8800 5962 8809
rect 5906 8735 5962 8744
rect 5920 7936 5948 8735
rect 6012 8129 6040 11494
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6104 9897 6132 10202
rect 6196 9926 6224 10406
rect 6184 9920 6236 9926
rect 6090 9888 6146 9897
rect 6184 9862 6236 9868
rect 6090 9823 6146 9832
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 5998 8120 6054 8129
rect 6104 8090 6132 9318
rect 6196 8634 6224 9318
rect 6288 9178 6316 14962
rect 6380 13734 6408 15302
rect 6886 14716 7182 14736
rect 6942 14714 6966 14716
rect 7022 14714 7046 14716
rect 7102 14714 7126 14716
rect 6964 14662 6966 14714
rect 7028 14662 7040 14714
rect 7102 14662 7104 14714
rect 6942 14660 6966 14662
rect 7022 14660 7046 14662
rect 7102 14660 7126 14662
rect 6886 14640 7182 14660
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6380 12714 6408 13670
rect 6886 13628 7182 13648
rect 6942 13626 6966 13628
rect 7022 13626 7046 13628
rect 7102 13626 7126 13628
rect 6964 13574 6966 13626
rect 7028 13574 7040 13626
rect 7102 13574 7104 13626
rect 6942 13572 6966 13574
rect 7022 13572 7046 13574
rect 7102 13572 7126 13574
rect 6886 13552 7182 13572
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 6368 12708 6420 12714
rect 6368 12650 6420 12656
rect 6366 12336 6422 12345
rect 6366 12271 6422 12280
rect 6380 11354 6408 12271
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6182 8528 6238 8537
rect 6182 8463 6238 8472
rect 5998 8055 6054 8064
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 5920 7908 6132 7936
rect 6000 7812 6052 7818
rect 6000 7754 6052 7760
rect 6012 7410 6040 7754
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5814 5536 5870 5545
rect 5814 5471 5870 5480
rect 5828 4690 5856 5471
rect 5920 4826 5948 6054
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5686 4542 5764 4570
rect 5630 4519 5686 4528
rect 5644 3942 5672 4519
rect 6012 4282 6040 5102
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5460 2650 5488 2790
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5552 2446 5580 3606
rect 5736 3505 5764 4218
rect 6104 3942 6132 7908
rect 6196 7426 6224 8463
rect 6288 7818 6316 8978
rect 6380 7954 6408 9522
rect 6472 9178 6500 13330
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6564 11354 6592 12174
rect 6656 12170 6684 12786
rect 6644 12164 6696 12170
rect 6644 12106 6696 12112
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6472 8498 6500 9114
rect 6564 8537 6592 11154
rect 6550 8528 6606 8537
rect 6460 8492 6512 8498
rect 6550 8463 6606 8472
rect 6460 8434 6512 8440
rect 6458 8392 6514 8401
rect 6458 8327 6514 8336
rect 6472 8294 6500 8327
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6458 8120 6514 8129
rect 6458 8055 6460 8064
rect 6512 8055 6514 8064
rect 6460 8026 6512 8032
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6276 7812 6328 7818
rect 6276 7754 6328 7760
rect 6380 7546 6408 7890
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 6196 7398 6316 7426
rect 6182 7304 6238 7313
rect 6182 7239 6238 7248
rect 6196 4690 6224 7239
rect 6288 5137 6316 7398
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6274 5128 6330 5137
rect 6274 5063 6330 5072
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6012 3738 6040 3878
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5816 3664 5868 3670
rect 5816 3606 5868 3612
rect 5722 3496 5778 3505
rect 5722 3431 5778 3440
rect 5736 2514 5764 3431
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 5644 1426 5672 2382
rect 5632 1420 5684 1426
rect 5632 1362 5684 1368
rect 5828 800 5856 3606
rect 6288 2990 6316 5063
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 6000 2916 6052 2922
rect 6000 2858 6052 2864
rect 6012 2582 6040 2858
rect 6380 2854 6408 7278
rect 6458 5264 6514 5273
rect 6458 5199 6460 5208
rect 6512 5199 6514 5208
rect 6460 5170 6512 5176
rect 6460 5092 6512 5098
rect 6460 5034 6512 5040
rect 6472 3670 6500 5034
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 6564 2582 6592 8230
rect 6656 7954 6684 11698
rect 6748 11642 6776 12854
rect 6932 12782 6960 13126
rect 7484 13025 7512 13330
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7470 13016 7526 13025
rect 7470 12951 7526 12960
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 6886 12540 7182 12560
rect 6942 12538 6966 12540
rect 7022 12538 7046 12540
rect 7102 12538 7126 12540
rect 6964 12486 6966 12538
rect 7028 12486 7040 12538
rect 7102 12486 7104 12538
rect 6942 12484 6966 12486
rect 7022 12484 7046 12486
rect 7102 12484 7126 12486
rect 6886 12464 7182 12484
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6840 11898 6868 12242
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 6932 11830 6960 12242
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 7024 12073 7052 12174
rect 7196 12096 7248 12102
rect 7010 12064 7066 12073
rect 7010 11999 7066 12008
rect 7116 12056 7196 12084
rect 6920 11824 6972 11830
rect 6920 11766 6972 11772
rect 7116 11694 7144 12056
rect 7196 12038 7248 12044
rect 7484 11762 7512 12951
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7104 11688 7156 11694
rect 6748 11626 6868 11642
rect 7104 11630 7156 11636
rect 6748 11620 6880 11626
rect 6748 11614 6828 11620
rect 6828 11562 6880 11568
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6748 11354 6776 11494
rect 6886 11452 7182 11472
rect 6942 11450 6966 11452
rect 7022 11450 7046 11452
rect 7102 11450 7126 11452
rect 6964 11398 6966 11450
rect 7028 11398 7040 11450
rect 7102 11398 7104 11450
rect 6942 11396 6966 11398
rect 7022 11396 7046 11398
rect 7102 11396 7126 11398
rect 6886 11376 7182 11396
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6932 11121 6960 11154
rect 6918 11112 6974 11121
rect 7484 11082 7512 11698
rect 7668 11694 7696 13262
rect 7760 12782 7788 16200
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 7840 13456 7892 13462
rect 7840 13398 7892 13404
rect 7852 12889 7880 13398
rect 8022 13016 8078 13025
rect 8022 12951 8024 12960
rect 8076 12951 8078 12960
rect 8024 12922 8076 12928
rect 7838 12880 7894 12889
rect 7838 12815 7894 12824
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7932 12708 7984 12714
rect 7932 12650 7984 12656
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7656 11688 7708 11694
rect 7576 11648 7656 11676
rect 6918 11047 6974 11056
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7470 10976 7526 10985
rect 7470 10911 7526 10920
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6840 10577 6868 10746
rect 6826 10568 6882 10577
rect 6736 10532 6788 10538
rect 6826 10503 6882 10512
rect 6736 10474 6788 10480
rect 6748 9926 6776 10474
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 6886 10364 7182 10384
rect 6942 10362 6966 10364
rect 7022 10362 7046 10364
rect 7102 10362 7126 10364
rect 6964 10310 6966 10362
rect 7028 10310 7040 10362
rect 7102 10310 7104 10362
rect 6942 10308 6966 10310
rect 7022 10308 7046 10310
rect 7102 10308 7126 10310
rect 6886 10288 7182 10308
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6748 8498 6776 9522
rect 7208 9518 7236 9998
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 6886 9276 7182 9296
rect 6942 9274 6966 9276
rect 7022 9274 7046 9276
rect 7102 9274 7126 9276
rect 6964 9222 6966 9274
rect 7028 9222 7040 9274
rect 7102 9222 7104 9274
rect 6942 9220 6966 9222
rect 7022 9220 7046 9222
rect 7102 9220 7126 9222
rect 6886 9200 7182 9220
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6840 8838 6868 8978
rect 7300 8974 7328 10406
rect 7288 8968 7340 8974
rect 7208 8928 7288 8956
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6656 7206 6684 7890
rect 6748 7868 6776 8434
rect 7208 8430 7236 8928
rect 7288 8910 7340 8916
rect 7484 8673 7512 10911
rect 7470 8664 7526 8673
rect 7470 8599 7526 8608
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 6886 8188 7182 8208
rect 6942 8186 6966 8188
rect 7022 8186 7046 8188
rect 7102 8186 7126 8188
rect 6964 8134 6966 8186
rect 7028 8134 7040 8186
rect 7102 8134 7104 8186
rect 6942 8132 6966 8134
rect 7022 8132 7046 8134
rect 7102 8132 7126 8134
rect 6886 8112 7182 8132
rect 7300 8090 7328 8298
rect 7484 8090 7512 8599
rect 7576 8401 7604 11648
rect 7656 11630 7708 11636
rect 7654 11248 7710 11257
rect 7760 11218 7788 12582
rect 7840 12368 7892 12374
rect 7840 12310 7892 12316
rect 7852 12209 7880 12310
rect 7838 12200 7894 12209
rect 7838 12135 7894 12144
rect 7944 11676 7972 12650
rect 8128 12442 8156 13806
rect 8220 12646 8248 14350
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 8116 12436 8168 12442
rect 8116 12378 8168 12384
rect 8220 11694 8248 12582
rect 8024 11688 8076 11694
rect 7838 11656 7894 11665
rect 7944 11648 8024 11676
rect 8024 11630 8076 11636
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 7838 11591 7894 11600
rect 7852 11286 7880 11591
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 7654 11183 7710 11192
rect 7748 11212 7800 11218
rect 7668 9382 7696 11183
rect 7748 11154 7800 11160
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7562 8392 7618 8401
rect 7562 8327 7618 8336
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7564 8016 7616 8022
rect 7562 7984 7564 7993
rect 7616 7984 7618 7993
rect 7562 7919 7618 7928
rect 7668 7886 7696 8230
rect 7760 8022 7788 11154
rect 7944 10470 7972 11154
rect 8036 10810 8064 11630
rect 8114 11384 8170 11393
rect 8114 11319 8116 11328
rect 8168 11319 8170 11328
rect 8116 11290 8168 11296
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 8036 10538 8064 10746
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 7932 10464 7984 10470
rect 7852 10424 7932 10452
rect 7852 8022 7880 10424
rect 7932 10406 7984 10412
rect 8128 10169 8156 11290
rect 8114 10160 8170 10169
rect 8114 10095 8170 10104
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 7944 9926 7972 9998
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7840 8016 7892 8022
rect 7840 7958 7892 7964
rect 6828 7880 6880 7886
rect 6748 7840 6828 7868
rect 6748 7274 6776 7840
rect 6828 7822 6880 7828
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7746 7712 7802 7721
rect 7746 7647 7802 7656
rect 7760 7426 7788 7647
rect 7564 7404 7616 7410
rect 7760 7398 7880 7426
rect 7564 7346 7616 7352
rect 7576 7313 7604 7346
rect 7562 7304 7618 7313
rect 6736 7268 6788 7274
rect 7562 7239 7618 7248
rect 6736 7210 6788 7216
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 6886 7100 7182 7120
rect 6942 7098 6966 7100
rect 7022 7098 7046 7100
rect 7102 7098 7126 7100
rect 6964 7046 6966 7098
rect 7028 7046 7040 7098
rect 7102 7046 7104 7098
rect 6942 7044 6966 7046
rect 7022 7044 7046 7046
rect 7102 7044 7126 7046
rect 6886 7024 7182 7044
rect 7300 7018 7328 7142
rect 7300 6990 7420 7018
rect 7288 6860 7340 6866
rect 7288 6802 7340 6808
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 6656 6322 6684 6734
rect 6736 6656 6788 6662
rect 6920 6656 6972 6662
rect 6736 6598 6788 6604
rect 6918 6624 6920 6633
rect 6972 6624 6974 6633
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6656 5914 6684 6258
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6656 3738 6684 5510
rect 6748 4078 6776 6598
rect 6918 6559 6974 6568
rect 6918 6488 6974 6497
rect 6840 6446 6918 6474
rect 6840 6390 6868 6446
rect 6918 6423 6974 6432
rect 6828 6384 6880 6390
rect 6828 6326 6880 6332
rect 7208 6186 7236 6734
rect 7196 6180 7248 6186
rect 7196 6122 7248 6128
rect 6886 6012 7182 6032
rect 6942 6010 6966 6012
rect 7022 6010 7046 6012
rect 7102 6010 7126 6012
rect 6964 5958 6966 6010
rect 7028 5958 7040 6010
rect 7102 5958 7104 6010
rect 6942 5956 6966 5958
rect 7022 5956 7046 5958
rect 7102 5956 7126 5958
rect 6886 5936 7182 5956
rect 7300 5817 7328 6802
rect 7286 5808 7342 5817
rect 7286 5743 7342 5752
rect 7194 5672 7250 5681
rect 7392 5658 7420 6990
rect 7484 6934 7512 7142
rect 7472 6928 7524 6934
rect 7472 6870 7524 6876
rect 7562 6624 7618 6633
rect 7562 6559 7618 6568
rect 7576 6458 7604 6559
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7194 5607 7250 5616
rect 7300 5630 7420 5658
rect 6918 5264 6974 5273
rect 7208 5250 7236 5607
rect 7300 5370 7328 5630
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7208 5222 7328 5250
rect 6918 5199 6974 5208
rect 6932 5166 6960 5199
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6886 4924 7182 4944
rect 6942 4922 6966 4924
rect 7022 4922 7046 4924
rect 7102 4922 7126 4924
rect 6964 4870 6966 4922
rect 7028 4870 7040 4922
rect 7102 4870 7104 4922
rect 6942 4868 6966 4870
rect 7022 4868 7046 4870
rect 7102 4868 7126 4870
rect 6886 4848 7182 4868
rect 7300 4808 7328 5222
rect 7208 4780 7328 4808
rect 7208 4622 7236 4780
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7208 4185 7236 4558
rect 7300 4214 7328 4558
rect 7288 4208 7340 4214
rect 7194 4176 7250 4185
rect 7288 4150 7340 4156
rect 7392 4146 7420 5510
rect 7194 4111 7250 4120
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6886 3836 7182 3856
rect 6942 3834 6966 3836
rect 7022 3834 7046 3836
rect 7102 3834 7126 3836
rect 6964 3782 6966 3834
rect 7028 3782 7040 3834
rect 7102 3782 7104 3834
rect 6942 3780 6966 3782
rect 7022 3780 7046 3782
rect 7102 3780 7126 3782
rect 6886 3760 7182 3780
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 7380 3664 7432 3670
rect 7380 3606 7432 3612
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6000 2576 6052 2582
rect 6000 2518 6052 2524
rect 6552 2576 6604 2582
rect 6552 2518 6604 2524
rect 6748 800 6776 3334
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 6886 2748 7182 2768
rect 6942 2746 6966 2748
rect 7022 2746 7046 2748
rect 7102 2746 7126 2748
rect 6964 2694 6966 2746
rect 7028 2694 7040 2746
rect 7102 2694 7104 2746
rect 6942 2692 6966 2694
rect 7022 2692 7046 2694
rect 7102 2692 7126 2694
rect 6886 2672 7182 2692
rect 7300 2514 7328 3062
rect 7392 3058 7420 3606
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7484 2990 7512 6394
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7562 5808 7618 5817
rect 7668 5778 7696 6190
rect 7562 5743 7618 5752
rect 7656 5772 7708 5778
rect 7576 5370 7604 5743
rect 7656 5714 7708 5720
rect 7656 5636 7708 5642
rect 7656 5578 7708 5584
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7668 4146 7696 5578
rect 7748 5568 7800 5574
rect 7746 5536 7748 5545
rect 7800 5536 7802 5545
rect 7746 5471 7802 5480
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 7760 5030 7788 5170
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7576 800 7604 3606
rect 7668 3602 7696 4082
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7852 2990 7880 7398
rect 7944 4622 7972 9862
rect 8036 9110 8064 9998
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 8128 8090 8156 9454
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8220 9178 8248 9318
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8116 8084 8168 8090
rect 8116 8026 8168 8032
rect 8024 8016 8076 8022
rect 8024 7958 8076 7964
rect 8036 6497 8064 7958
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8128 6662 8156 7346
rect 8220 6866 8248 8230
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8022 6488 8078 6497
rect 8022 6423 8078 6432
rect 8128 5914 8156 6598
rect 8220 6458 8248 6802
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 8036 4690 8064 5170
rect 8116 4752 8168 4758
rect 8116 4694 8168 4700
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 8036 4010 8064 4626
rect 8128 4010 8156 4694
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8220 4049 8248 4558
rect 8206 4040 8262 4049
rect 8024 4004 8076 4010
rect 8024 3946 8076 3952
rect 8116 4004 8168 4010
rect 8206 3975 8262 3984
rect 8116 3946 8168 3952
rect 8036 3738 8064 3946
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 8036 3058 8064 3674
rect 8312 3602 8340 13942
rect 8404 11218 8432 16623
rect 9954 16200 10010 17000
rect 12162 16200 12218 17000
rect 14370 16200 14426 17000
rect 16578 16200 16634 17000
rect 18326 16688 18382 16697
rect 18326 16623 18382 16632
rect 18234 16280 18290 16289
rect 18234 16215 18290 16224
rect 8852 15292 8904 15298
rect 8852 15234 8904 15240
rect 8576 14544 8628 14550
rect 8576 14486 8628 14492
rect 8588 13530 8616 14486
rect 8668 14476 8720 14482
rect 8668 14418 8720 14424
rect 8680 14074 8708 14418
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8668 13796 8720 13802
rect 8668 13738 8720 13744
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8392 11212 8444 11218
rect 8392 11154 8444 11160
rect 8404 11014 8432 11154
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8404 8362 8432 9318
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8496 8090 8524 12106
rect 8588 10266 8616 12174
rect 8680 11558 8708 13738
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8772 10810 8800 13874
rect 8864 13394 8892 15234
rect 9036 14884 9088 14890
rect 9036 14826 9088 14832
rect 9048 14056 9076 14826
rect 9968 14498 9996 16200
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11336 14544 11388 14550
rect 9588 14476 9640 14482
rect 9968 14470 10272 14498
rect 11336 14486 11388 14492
rect 9588 14418 9640 14424
rect 9600 14074 9628 14418
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9588 14068 9640 14074
rect 9048 14028 9352 14056
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 8956 13530 8984 13874
rect 8944 13524 8996 13530
rect 8944 13466 8996 13472
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 8864 12170 8892 13330
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8852 12164 8904 12170
rect 8852 12106 8904 12112
rect 8956 11762 8984 12174
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 8852 11076 8904 11082
rect 8852 11018 8904 11024
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8864 10130 8892 11018
rect 8956 10606 8984 11698
rect 9048 11257 9076 14028
rect 9324 13870 9352 14028
rect 9588 14010 9640 14016
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9402 13424 9458 13433
rect 9508 13394 9536 13670
rect 9402 13359 9404 13368
rect 9456 13359 9458 13368
rect 9496 13388 9548 13394
rect 9404 13330 9456 13336
rect 9496 13330 9548 13336
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 9034 11248 9090 11257
rect 9034 11183 9090 11192
rect 9140 11121 9168 13126
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9232 11218 9260 12378
rect 9310 12200 9366 12209
rect 9310 12135 9366 12144
rect 9324 12102 9352 12135
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9324 11150 9352 12038
rect 9312 11144 9364 11150
rect 9126 11112 9182 11121
rect 9312 11086 9364 11092
rect 9126 11047 9182 11056
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 9218 10568 9274 10577
rect 9218 10503 9274 10512
rect 9232 10470 9260 10503
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8588 8090 8616 9522
rect 8666 9480 8722 9489
rect 8666 9415 8722 9424
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8496 7954 8524 8026
rect 8680 7970 8708 9415
rect 8864 8838 8892 10066
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 8588 7942 8708 7970
rect 8588 7886 8616 7942
rect 8576 7880 8628 7886
rect 8390 7848 8446 7857
rect 8576 7822 8628 7828
rect 8390 7783 8446 7792
rect 8668 7812 8720 7818
rect 8404 7342 8432 7783
rect 8668 7754 8720 7760
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8588 6934 8616 7278
rect 8576 6928 8628 6934
rect 8576 6870 8628 6876
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8404 4554 8432 6734
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8496 6254 8524 6598
rect 8588 6304 8616 6870
rect 8680 6730 8708 7754
rect 8772 7732 8800 8230
rect 8864 7886 8892 8774
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 8956 8022 8984 8230
rect 8944 8016 8996 8022
rect 8944 7958 8996 7964
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8944 7812 8996 7818
rect 8944 7754 8996 7760
rect 8772 7704 8892 7732
rect 8864 7274 8892 7704
rect 8956 7449 8984 7754
rect 8942 7440 8998 7449
rect 8942 7375 8998 7384
rect 8942 7304 8998 7313
rect 8852 7268 8904 7274
rect 8942 7239 8944 7248
rect 8852 7210 8904 7216
rect 8996 7239 8998 7248
rect 8944 7210 8996 7216
rect 8864 7154 8892 7210
rect 8864 7126 8984 7154
rect 8852 6928 8904 6934
rect 8852 6870 8904 6876
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8668 6316 8720 6322
rect 8588 6276 8668 6304
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8588 5846 8616 6276
rect 8668 6258 8720 6264
rect 8576 5840 8628 5846
rect 8576 5782 8628 5788
rect 8666 5264 8722 5273
rect 8666 5199 8722 5208
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7840 2984 7892 2990
rect 8116 2984 8168 2990
rect 7840 2926 7892 2932
rect 8114 2952 8116 2961
rect 8168 2952 8170 2961
rect 8114 2887 8170 2896
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 7668 1970 7696 2246
rect 7656 1964 7708 1970
rect 7656 1906 7708 1912
rect 8496 800 8524 4558
rect 8680 4554 8708 5199
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8864 3618 8892 6870
rect 8680 3590 8892 3618
rect 8680 2514 8708 3590
rect 8956 3482 8984 7126
rect 8772 3454 8984 3482
rect 8668 2508 8720 2514
rect 8668 2450 8720 2456
rect 8772 2378 8800 3454
rect 8852 2848 8904 2854
rect 8852 2790 8904 2796
rect 8864 2582 8892 2790
rect 9048 2650 9076 8910
rect 9324 6934 9352 11086
rect 9416 7857 9444 13330
rect 9692 13326 9720 13874
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9692 12782 9720 13262
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9784 11830 9812 14214
rect 9852 14172 10148 14192
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 9930 14118 9932 14170
rect 9994 14118 10006 14170
rect 10068 14118 10070 14170
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 9852 14096 10148 14116
rect 10244 13802 10272 14470
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 10612 14074 10640 14350
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10796 13938 10824 14350
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10508 13864 10560 13870
rect 10508 13806 10560 13812
rect 10232 13796 10284 13802
rect 10232 13738 10284 13744
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 9968 13530 9996 13670
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 9852 13084 10148 13104
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 9930 13030 9932 13082
rect 9994 13030 10006 13082
rect 10068 13030 10070 13082
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 9852 13008 10148 13028
rect 10244 12889 10272 13126
rect 10336 12986 10364 13670
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10230 12880 10286 12889
rect 10230 12815 10286 12824
rect 10416 12844 10468 12850
rect 10244 12782 10272 12815
rect 10416 12786 10468 12792
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 9852 11996 10148 12016
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 9930 11942 9932 11994
rect 9994 11942 10006 11994
rect 10068 11942 10070 11994
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 9852 11920 10148 11940
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 9496 11620 9548 11626
rect 9496 11562 9548 11568
rect 9508 11354 9536 11562
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9692 11354 9720 11494
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9600 10606 9628 10950
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9402 7848 9458 7857
rect 9402 7783 9458 7792
rect 9312 6928 9364 6934
rect 9312 6870 9364 6876
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9220 5772 9272 5778
rect 9220 5714 9272 5720
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9140 4826 9168 5170
rect 9232 5166 9260 5714
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9232 4758 9260 5102
rect 9220 4752 9272 4758
rect 9220 4694 9272 4700
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9140 3194 9168 4558
rect 9232 4282 9260 4694
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9324 3058 9352 6598
rect 9404 5296 9456 5302
rect 9404 5238 9456 5244
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9312 2916 9364 2922
rect 9312 2858 9364 2864
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 8852 2576 8904 2582
rect 8852 2518 8904 2524
rect 9324 2446 9352 2858
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 8760 2372 8812 2378
rect 8760 2314 8812 2320
rect 9416 800 9444 5238
rect 9508 3058 9536 9318
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 9600 2854 9628 10542
rect 9692 9586 9720 11154
rect 9784 10198 9812 11766
rect 9862 11384 9918 11393
rect 9862 11319 9864 11328
rect 9916 11319 9918 11328
rect 9864 11290 9916 11296
rect 9852 10908 10148 10928
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 9930 10854 9932 10906
rect 9994 10854 10006 10906
rect 10068 10854 10070 10906
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 9852 10832 10148 10852
rect 9772 10192 9824 10198
rect 9772 10134 9824 10140
rect 9852 9820 10148 9840
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 9930 9766 9932 9818
rect 9994 9766 10006 9818
rect 10068 9766 10070 9818
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 9852 9744 10148 9764
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9784 7970 9812 9658
rect 9852 8732 10148 8752
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 9930 8678 9932 8730
rect 9994 8678 10006 8730
rect 10068 8678 10070 8730
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 9852 8656 10148 8676
rect 10244 8090 10272 12242
rect 10336 11801 10364 12378
rect 10428 12374 10456 12786
rect 10416 12368 10468 12374
rect 10520 12345 10548 13806
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10416 12310 10468 12316
rect 10506 12336 10562 12345
rect 10322 11792 10378 11801
rect 10322 11727 10378 11736
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10336 9364 10364 11086
rect 10428 10810 10456 12310
rect 10506 12271 10562 12280
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10520 11014 10548 12038
rect 10612 11558 10640 13670
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10704 13161 10732 13194
rect 10690 13152 10746 13161
rect 10690 13087 10746 13096
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10612 11150 10640 11494
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10520 10690 10548 10950
rect 10428 10662 10548 10690
rect 10428 10130 10456 10662
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10428 9518 10456 10066
rect 10520 10033 10548 10066
rect 10506 10024 10562 10033
rect 10506 9959 10562 9968
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10336 9336 10456 9364
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 9784 7954 9904 7970
rect 9784 7948 9916 7954
rect 9784 7942 9864 7948
rect 9864 7890 9916 7896
rect 9852 7644 10148 7664
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 9930 7590 9932 7642
rect 9994 7590 10006 7642
rect 10068 7590 10070 7642
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 9852 7568 10148 7588
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9692 5370 9720 7142
rect 9784 6186 9812 7142
rect 10152 7041 10180 7346
rect 10138 7032 10194 7041
rect 10138 6967 10194 6976
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 9852 6556 10148 6576
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 9930 6502 9932 6554
rect 9994 6502 10006 6554
rect 10068 6502 10070 6554
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 9852 6480 10148 6500
rect 9772 6180 9824 6186
rect 9772 6122 9824 6128
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9784 5030 9812 5510
rect 9852 5468 10148 5488
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 9930 5414 9932 5466
rect 9994 5414 10006 5466
rect 10068 5414 10070 5466
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 9852 5392 10148 5412
rect 9864 5296 9916 5302
rect 9864 5238 9916 5244
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9692 4486 9720 4966
rect 9876 4690 9904 5238
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 10060 4690 10088 5102
rect 10244 4826 10272 6938
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9852 4380 10148 4400
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 9930 4326 9932 4378
rect 9994 4326 10006 4378
rect 10068 4326 10070 4378
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 9852 4304 10148 4324
rect 10336 4282 10364 8774
rect 10428 6254 10456 9336
rect 10520 8022 10548 9959
rect 10508 8016 10560 8022
rect 10508 7958 10560 7964
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10520 6934 10548 7822
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10508 6928 10560 6934
rect 10508 6870 10560 6876
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10428 5778 10456 6054
rect 10520 5846 10548 6870
rect 10508 5840 10560 5846
rect 10508 5782 10560 5788
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10414 5672 10470 5681
rect 10414 5607 10470 5616
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9692 3602 9720 3878
rect 10060 3738 10088 3946
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9852 3292 10148 3312
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 9930 3238 9932 3290
rect 9994 3238 10006 3290
rect 10068 3238 10070 3290
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 9852 3216 10148 3236
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10060 2582 10088 2790
rect 10048 2576 10100 2582
rect 10048 2518 10100 2524
rect 10324 2576 10376 2582
rect 10324 2518 10376 2524
rect 9852 2204 10148 2224
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 9930 2150 9932 2202
rect 9994 2150 10006 2202
rect 10068 2150 10070 2202
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 9852 2128 10148 2148
rect 10336 800 10364 2518
rect 10428 2310 10456 5607
rect 10520 4826 10548 5782
rect 10612 5370 10640 7278
rect 10704 6225 10732 12854
rect 10796 12442 10824 13874
rect 10888 13258 10916 13874
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10888 12850 10916 13194
rect 10980 13161 11008 13262
rect 10966 13152 11022 13161
rect 10966 13087 11022 13096
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 10888 10130 10916 12650
rect 10968 11280 11020 11286
rect 10966 11248 10968 11257
rect 11020 11248 11022 11257
rect 10966 11183 11022 11192
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10796 9722 10824 9998
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10888 9586 10916 9862
rect 10980 9722 11008 10406
rect 11072 9994 11100 14350
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 11072 9518 11100 9930
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 10980 8401 11008 8502
rect 10966 8392 11022 8401
rect 10966 8327 11022 8336
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10782 7304 10838 7313
rect 10782 7239 10838 7248
rect 10796 7206 10824 7239
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10690 6216 10746 6225
rect 10690 6151 10746 6160
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10704 5166 10732 6151
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10796 5030 10824 7142
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10520 4078 10548 4762
rect 10888 4486 10916 8026
rect 11072 8022 11100 8230
rect 10968 8016 11020 8022
rect 10968 7958 11020 7964
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 10980 7410 11008 7958
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10980 6866 11008 7346
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 10888 4282 10916 4422
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10520 3602 10548 4014
rect 10508 3596 10560 3602
rect 10508 3538 10560 3544
rect 10980 2514 11008 5714
rect 11072 5166 11100 6054
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 11072 4049 11100 4082
rect 11058 4040 11114 4049
rect 11058 3975 11114 3984
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11072 3602 11100 3878
rect 11060 3596 11112 3602
rect 11060 3538 11112 3544
rect 11164 3058 11192 14214
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 11256 13530 11284 13670
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 11348 13410 11376 14486
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 11256 13382 11376 13410
rect 11256 8378 11284 13382
rect 11440 12714 11468 14418
rect 11428 12708 11480 12714
rect 11428 12650 11480 12656
rect 11426 11656 11482 11665
rect 11426 11591 11482 11600
rect 11440 11082 11468 11591
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 11532 10452 11560 14758
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 11624 12306 11652 13806
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11716 11830 11744 13670
rect 11888 13456 11940 13462
rect 11888 13398 11940 13404
rect 11900 13258 11928 13398
rect 11888 13252 11940 13258
rect 11888 13194 11940 13200
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11808 12850 11836 13126
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11992 12288 12020 14418
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 11808 12260 12020 12288
rect 11704 11824 11756 11830
rect 11704 11766 11756 11772
rect 11808 11234 11836 12260
rect 12084 12186 12112 14010
rect 12176 13938 12204 16200
rect 12817 14716 13113 14736
rect 12873 14714 12897 14716
rect 12953 14714 12977 14716
rect 13033 14714 13057 14716
rect 12895 14662 12897 14714
rect 12959 14662 12971 14714
rect 13033 14662 13035 14714
rect 12873 14660 12897 14662
rect 12953 14660 12977 14662
rect 13033 14660 13057 14662
rect 12817 14640 13113 14660
rect 14384 14550 14412 16200
rect 15290 15872 15346 15881
rect 15290 15807 15346 15816
rect 15106 15464 15162 15473
rect 15106 15399 15162 15408
rect 14372 14544 14424 14550
rect 14372 14486 14424 14492
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12452 13546 12480 14418
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12360 13518 12480 13546
rect 12544 13530 12572 14350
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 14188 14340 14240 14346
rect 14188 14282 14240 14288
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 12817 13628 13113 13648
rect 12873 13626 12897 13628
rect 12953 13626 12977 13628
rect 13033 13626 13057 13628
rect 12895 13574 12897 13626
rect 12959 13574 12971 13626
rect 13033 13574 13035 13626
rect 12873 13572 12897 13574
rect 12953 13572 12977 13574
rect 13033 13572 13057 13574
rect 12817 13552 13113 13572
rect 12532 13524 12584 13530
rect 12360 12986 12388 13518
rect 12532 13466 12584 13472
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12348 12980 12400 12986
rect 12348 12922 12400 12928
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 11900 12158 12112 12186
rect 11900 11762 11928 12158
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11980 11620 12032 11626
rect 11980 11562 12032 11568
rect 11900 11286 11928 11317
rect 11888 11280 11940 11286
rect 11808 11228 11888 11234
rect 11808 11222 11940 11228
rect 11704 11212 11756 11218
rect 11808 11206 11928 11222
rect 11704 11154 11756 11160
rect 11716 10810 11744 11154
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11704 10464 11756 10470
rect 11532 10424 11704 10452
rect 11704 10406 11756 10412
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11256 8350 11468 8378
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11348 7546 11376 8230
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 11440 7449 11468 8350
rect 11532 8129 11560 9114
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11518 8120 11574 8129
rect 11624 8090 11652 8434
rect 11518 8055 11574 8064
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11532 7546 11560 7890
rect 11612 7880 11664 7886
rect 11610 7848 11612 7857
rect 11664 7848 11666 7857
rect 11610 7783 11666 7792
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11426 7440 11482 7449
rect 11244 7404 11296 7410
rect 11426 7375 11482 7384
rect 11244 7346 11296 7352
rect 11256 6934 11284 7346
rect 11440 7206 11468 7375
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11348 6934 11376 7142
rect 11244 6928 11296 6934
rect 11244 6870 11296 6876
rect 11336 6928 11388 6934
rect 11336 6870 11388 6876
rect 11256 6322 11284 6870
rect 11334 6488 11390 6497
rect 11334 6423 11390 6432
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11348 6118 11376 6423
rect 11520 6384 11572 6390
rect 11520 6326 11572 6332
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11242 5128 11298 5137
rect 11242 5063 11298 5072
rect 11256 4729 11284 5063
rect 11348 4758 11376 5170
rect 11428 5160 11480 5166
rect 11426 5128 11428 5137
rect 11480 5128 11482 5137
rect 11426 5063 11482 5072
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 11440 4826 11468 4966
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11336 4752 11388 4758
rect 11242 4720 11298 4729
rect 11336 4694 11388 4700
rect 11532 4690 11560 6326
rect 11612 6180 11664 6186
rect 11612 6122 11664 6128
rect 11624 5914 11652 6122
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11716 5794 11744 10406
rect 11808 9178 11836 11086
rect 11900 10266 11928 11206
rect 11992 11150 12020 11562
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11808 7002 11836 7142
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 11900 6458 11928 6734
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11992 6186 12020 7142
rect 11980 6180 12032 6186
rect 11980 6122 12032 6128
rect 11794 5808 11850 5817
rect 11716 5766 11794 5794
rect 11794 5743 11850 5752
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11242 4655 11298 4664
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11428 4480 11480 4486
rect 11428 4422 11480 4428
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11348 3126 11376 3878
rect 11336 3120 11388 3126
rect 11336 3062 11388 3068
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 11072 2650 11100 2790
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 11164 2378 11192 2858
rect 11440 2514 11468 4422
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 11624 3398 11652 4082
rect 11716 3738 11744 5510
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11716 3058 11744 3674
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11808 2990 11836 5743
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11992 4486 12020 4558
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11900 3641 11928 3878
rect 11886 3632 11942 3641
rect 11886 3567 11942 3576
rect 11992 3534 12020 4422
rect 12084 4078 12112 12038
rect 12176 11762 12204 12378
rect 12452 11914 12480 13330
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12728 12714 12848 12730
rect 12912 12714 12940 13262
rect 13188 12753 13216 13806
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13174 12744 13230 12753
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12728 12708 12860 12714
rect 12728 12702 12808 12708
rect 12544 12170 12572 12650
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12268 11898 12480 11914
rect 12256 11892 12480 11898
rect 12308 11886 12480 11892
rect 12256 11834 12308 11840
rect 12544 11812 12572 12106
rect 12728 12102 12756 12702
rect 12808 12650 12860 12656
rect 12900 12708 12952 12714
rect 13174 12679 13230 12688
rect 12900 12650 12952 12656
rect 12817 12540 13113 12560
rect 12873 12538 12897 12540
rect 12953 12538 12977 12540
rect 13033 12538 13057 12540
rect 12895 12486 12897 12538
rect 12959 12486 12971 12538
rect 13033 12486 13035 12538
rect 12873 12484 12897 12486
rect 12953 12484 12977 12486
rect 13033 12484 13057 12486
rect 12817 12464 13113 12484
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12360 11784 12572 11812
rect 12164 11756 12216 11762
rect 12164 11698 12216 11704
rect 12360 11694 12388 11784
rect 12348 11688 12400 11694
rect 12820 11665 12848 12174
rect 12348 11630 12400 11636
rect 12806 11656 12862 11665
rect 12360 11218 12388 11630
rect 12806 11591 12862 11600
rect 13188 11558 13216 12174
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 12817 11452 13113 11472
rect 12873 11450 12897 11452
rect 12953 11450 12977 11452
rect 13033 11450 13057 11452
rect 12895 11398 12897 11450
rect 12959 11398 12971 11450
rect 13033 11398 13035 11450
rect 12873 11396 12897 11398
rect 12953 11396 12977 11398
rect 13033 11396 13057 11398
rect 12817 11376 13113 11396
rect 12348 11212 12400 11218
rect 12624 11212 12676 11218
rect 12400 11172 12480 11200
rect 12348 11154 12400 11160
rect 12346 11112 12402 11121
rect 12346 11047 12402 11056
rect 12360 10606 12388 11047
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12360 10033 12388 10066
rect 12346 10024 12402 10033
rect 12256 9988 12308 9994
rect 12452 10010 12480 11172
rect 12624 11154 12676 11160
rect 12636 10674 12664 11154
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12636 10248 12664 10610
rect 12728 10470 12756 10678
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12817 10364 13113 10384
rect 12873 10362 12897 10364
rect 12953 10362 12977 10364
rect 13033 10362 13057 10364
rect 12895 10310 12897 10362
rect 12959 10310 12971 10362
rect 13033 10310 13035 10362
rect 12873 10308 12897 10310
rect 12953 10308 12977 10310
rect 13033 10308 13057 10310
rect 12817 10288 13113 10308
rect 12636 10220 12848 10248
rect 12452 9994 12756 10010
rect 12452 9988 12768 9994
rect 12452 9982 12716 9988
rect 12346 9959 12402 9968
rect 12256 9930 12308 9936
rect 12716 9930 12768 9936
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 12176 7478 12204 7686
rect 12164 7472 12216 7478
rect 12164 7414 12216 7420
rect 12268 7290 12296 9930
rect 12440 9920 12492 9926
rect 12820 9874 12848 10220
rect 13188 10198 13216 10610
rect 12992 10192 13044 10198
rect 12992 10134 13044 10140
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 12440 9862 12492 9868
rect 12452 9110 12480 9862
rect 12636 9846 12848 9874
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12544 9178 12572 9318
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12348 9104 12400 9110
rect 12348 9046 12400 9052
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 12360 8945 12388 9046
rect 12636 8974 12664 9846
rect 12716 9648 12768 9654
rect 12716 9590 12768 9596
rect 12624 8968 12676 8974
rect 12346 8936 12402 8945
rect 12624 8910 12676 8916
rect 12346 8871 12402 8880
rect 12728 8786 12756 9590
rect 13004 9364 13032 10134
rect 13188 9586 13216 10134
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13004 9336 13216 9364
rect 12817 9276 13113 9296
rect 12873 9274 12897 9276
rect 12953 9274 12977 9276
rect 13033 9274 13057 9276
rect 12895 9222 12897 9274
rect 12959 9222 12971 9274
rect 13033 9222 13035 9274
rect 12873 9220 12897 9222
rect 12953 9220 12977 9222
rect 13033 9220 13057 9222
rect 12817 9200 13113 9220
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12452 8758 12756 8786
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 12360 8378 12388 8502
rect 12452 8378 12480 8758
rect 12360 8350 12480 8378
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12348 7812 12400 7818
rect 12348 7754 12400 7760
rect 12360 7478 12388 7754
rect 12348 7472 12400 7478
rect 12348 7414 12400 7420
rect 12176 7262 12296 7290
rect 12176 6118 12204 7262
rect 12254 7032 12310 7041
rect 12254 6967 12310 6976
rect 12268 6934 12296 6967
rect 12256 6928 12308 6934
rect 12256 6870 12308 6876
rect 12346 6896 12402 6905
rect 12346 6831 12402 6840
rect 12360 6798 12388 6831
rect 12348 6792 12400 6798
rect 12254 6760 12310 6769
rect 12452 6780 12480 8230
rect 12544 8090 12572 8298
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12544 6905 12572 7414
rect 12530 6896 12586 6905
rect 12530 6831 12586 6840
rect 12452 6752 12572 6780
rect 12348 6734 12400 6740
rect 12254 6695 12310 6704
rect 12268 6662 12296 6695
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12176 4214 12204 6054
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 12164 4208 12216 4214
rect 12164 4150 12216 4156
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 12164 4004 12216 4010
rect 12164 3946 12216 3952
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 11152 2372 11204 2378
rect 11152 2314 11204 2320
rect 10416 2304 10468 2310
rect 10416 2246 10468 2252
rect 11244 1420 11296 1426
rect 11244 1362 11296 1368
rect 11256 800 11284 1362
rect 12176 800 12204 3946
rect 12268 3942 12296 5102
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12360 2650 12388 6734
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12452 2650 12480 6394
rect 12544 5098 12572 6752
rect 12636 6254 12664 8758
rect 12820 8634 12848 8842
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12728 6905 12756 8570
rect 13188 8294 13216 9336
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 12817 8188 13113 8208
rect 12873 8186 12897 8188
rect 12953 8186 12977 8188
rect 13033 8186 13057 8188
rect 12895 8134 12897 8186
rect 12959 8134 12971 8186
rect 13033 8134 13035 8186
rect 12873 8132 12897 8134
rect 12953 8132 12977 8134
rect 13033 8132 13057 8134
rect 12817 8112 13113 8132
rect 13280 7954 13308 13330
rect 13464 12986 13492 13806
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13556 12646 13584 14214
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13648 12753 13676 13262
rect 13634 12744 13690 12753
rect 13634 12679 13690 12688
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13648 12374 13676 12582
rect 13740 12374 13768 14282
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 13924 13394 13952 13670
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13832 12442 13860 13262
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13360 12368 13412 12374
rect 13360 12310 13412 12316
rect 13636 12368 13688 12374
rect 13636 12310 13688 12316
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13372 11898 13400 12310
rect 13636 12096 13688 12102
rect 13740 12084 13768 12310
rect 13688 12056 13768 12084
rect 13636 12038 13688 12044
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13924 11744 13952 13330
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 13556 11716 13952 11744
rect 13556 11234 13584 11716
rect 14016 11642 14044 12038
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 13648 11614 14044 11642
rect 13648 11354 13676 11614
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13556 11206 13676 11234
rect 13542 11112 13598 11121
rect 13542 11047 13598 11056
rect 13556 11014 13584 11047
rect 13452 11008 13504 11014
rect 13452 10950 13504 10956
rect 13544 11008 13596 11014
rect 13544 10950 13596 10956
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 13372 9466 13400 10406
rect 13464 9654 13492 10950
rect 13452 9648 13504 9654
rect 13452 9590 13504 9596
rect 13648 9489 13676 11206
rect 13634 9480 13690 9489
rect 13372 9438 13584 9466
rect 13556 9081 13584 9438
rect 13634 9415 13690 9424
rect 13542 9072 13598 9081
rect 13542 9007 13598 9016
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13082 7576 13138 7585
rect 13082 7511 13138 7520
rect 13096 7410 13124 7511
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 12817 7100 13113 7120
rect 12873 7098 12897 7100
rect 12953 7098 12977 7100
rect 13033 7098 13057 7100
rect 12895 7046 12897 7098
rect 12959 7046 12971 7098
rect 13033 7046 13035 7098
rect 12873 7044 12897 7046
rect 12953 7044 12977 7046
rect 13033 7044 13057 7046
rect 12817 7024 13113 7044
rect 12714 6896 12770 6905
rect 12714 6831 12770 6840
rect 13188 6798 13216 7278
rect 13464 7206 13492 7822
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12990 6624 13046 6633
rect 12728 6322 12756 6598
rect 12990 6559 13046 6568
rect 13004 6390 13032 6559
rect 13188 6390 13216 6734
rect 12992 6384 13044 6390
rect 12898 6352 12954 6361
rect 12716 6316 12768 6322
rect 12992 6326 13044 6332
rect 13176 6384 13228 6390
rect 13176 6326 13228 6332
rect 12898 6287 12954 6296
rect 12716 6258 12768 6264
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12912 6186 12940 6287
rect 12900 6180 12952 6186
rect 12900 6122 12952 6128
rect 12817 6012 13113 6032
rect 12873 6010 12897 6012
rect 12953 6010 12977 6012
rect 13033 6010 13057 6012
rect 12895 5958 12897 6010
rect 12959 5958 12971 6010
rect 13033 5958 13035 6010
rect 12873 5956 12897 5958
rect 12953 5956 12977 5958
rect 13033 5956 13057 5958
rect 12817 5936 13113 5956
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 12636 4758 12664 5510
rect 13188 5234 13216 5510
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 13176 5092 13228 5098
rect 13176 5034 13228 5040
rect 12817 4924 13113 4944
rect 12873 4922 12897 4924
rect 12953 4922 12977 4924
rect 13033 4922 13057 4924
rect 12895 4870 12897 4922
rect 12959 4870 12971 4922
rect 13033 4870 13035 4922
rect 12873 4868 12897 4870
rect 12953 4868 12977 4870
rect 13033 4868 13057 4870
rect 12817 4848 13113 4868
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 13188 4622 13216 5034
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 13280 4060 13308 7142
rect 13450 6896 13506 6905
rect 13450 6831 13506 6840
rect 13464 6730 13492 6831
rect 13452 6724 13504 6730
rect 13452 6666 13504 6672
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13360 6248 13412 6254
rect 13464 6225 13492 6394
rect 13360 6190 13412 6196
rect 13450 6216 13506 6225
rect 13372 4826 13400 6190
rect 13450 6151 13506 6160
rect 13556 6100 13584 9007
rect 13648 8106 13676 9415
rect 13740 9042 13768 11494
rect 14108 11370 14136 11698
rect 13924 11354 14136 11370
rect 13912 11348 14136 11354
rect 13964 11342 14136 11348
rect 13912 11290 13964 11296
rect 13818 11248 13874 11257
rect 13818 11183 13874 11192
rect 13832 10470 13860 11183
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 13820 10464 13872 10470
rect 13924 10441 13952 10474
rect 13820 10406 13872 10412
rect 13910 10432 13966 10441
rect 13910 10367 13966 10376
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13832 9654 13860 10066
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13648 8078 13768 8106
rect 13832 8090 13860 8978
rect 13924 8634 13952 9522
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 13464 6072 13584 6100
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 13372 4078 13400 4422
rect 13188 4032 13308 4060
rect 13360 4072 13412 4078
rect 12817 3836 13113 3856
rect 12873 3834 12897 3836
rect 12953 3834 12977 3836
rect 13033 3834 13057 3836
rect 12895 3782 12897 3834
rect 12959 3782 12971 3834
rect 13033 3782 13035 3834
rect 12873 3780 12897 3782
rect 12953 3780 12977 3782
rect 13033 3780 13057 3782
rect 12817 3760 13113 3780
rect 12817 2748 13113 2768
rect 12873 2746 12897 2748
rect 12953 2746 12977 2748
rect 13033 2746 13057 2748
rect 12895 2694 12897 2746
rect 12959 2694 12971 2746
rect 13033 2694 13035 2746
rect 12873 2692 12897 2694
rect 12953 2692 12977 2694
rect 13033 2692 13057 2694
rect 12817 2672 13113 2692
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 13084 2576 13136 2582
rect 13188 2564 13216 4032
rect 13464 4049 13492 6072
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13556 5370 13584 5646
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 13556 5234 13584 5306
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13648 5114 13676 7958
rect 13740 7886 13768 8078
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13924 7936 13952 8366
rect 13832 7908 13952 7936
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13832 7290 13860 7908
rect 13912 7812 13964 7818
rect 13912 7754 13964 7760
rect 13924 7410 13952 7754
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13832 7262 13952 7290
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13832 6361 13860 7142
rect 13924 6662 13952 7262
rect 14016 6769 14044 11086
rect 14096 11076 14148 11082
rect 14096 11018 14148 11024
rect 14108 10606 14136 11018
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14200 10146 14228 14282
rect 14384 13938 14412 14486
rect 15120 14482 15148 15399
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 15108 14476 15160 14482
rect 15108 14418 15160 14424
rect 14372 13932 14424 13938
rect 14372 13874 14424 13880
rect 14648 13456 14700 13462
rect 14648 13398 14700 13404
rect 14660 13258 14688 13398
rect 14648 13252 14700 13258
rect 14648 13194 14700 13200
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14568 12918 14596 13126
rect 14556 12912 14608 12918
rect 14556 12854 14608 12860
rect 14568 12238 14596 12854
rect 14646 12744 14702 12753
rect 14646 12679 14702 12688
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 14292 11150 14320 12106
rect 14554 11656 14610 11665
rect 14464 11620 14516 11626
rect 14554 11591 14610 11600
rect 14464 11562 14516 11568
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14384 11354 14412 11494
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14280 10736 14332 10742
rect 14384 10713 14412 11154
rect 14476 10810 14504 11562
rect 14568 10810 14596 11591
rect 14464 10804 14516 10810
rect 14464 10746 14516 10752
rect 14556 10804 14608 10810
rect 14556 10746 14608 10752
rect 14280 10678 14332 10684
rect 14370 10704 14426 10713
rect 14108 10118 14228 10146
rect 14108 8945 14136 10118
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14200 9178 14228 9522
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14188 8968 14240 8974
rect 14094 8936 14150 8945
rect 14188 8910 14240 8916
rect 14094 8871 14150 8880
rect 14108 7342 14136 8871
rect 14200 8090 14228 8910
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14292 7546 14320 10678
rect 14370 10639 14426 10648
rect 14556 10668 14608 10674
rect 14384 9926 14412 10639
rect 14556 10610 14608 10616
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14476 10266 14504 10542
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 14464 9444 14516 9450
rect 14464 9386 14516 9392
rect 14476 8838 14504 9386
rect 14568 9178 14596 10610
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14476 8498 14504 8774
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14462 8392 14518 8401
rect 14462 8327 14518 8336
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 14384 8090 14412 8230
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 14096 6792 14148 6798
rect 14002 6760 14058 6769
rect 14096 6734 14148 6740
rect 14002 6695 14058 6704
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13818 6352 13874 6361
rect 13818 6287 13874 6296
rect 13924 6186 13952 6598
rect 14108 6497 14136 6734
rect 14094 6488 14150 6497
rect 14094 6423 14150 6432
rect 13912 6180 13964 6186
rect 13912 6122 13964 6128
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13832 5302 13860 5510
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 13924 5166 13952 6122
rect 14292 5710 14320 7482
rect 14372 6860 14424 6866
rect 14372 6802 14424 6808
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 13912 5160 13964 5166
rect 13648 5086 13768 5114
rect 13912 5102 13964 5108
rect 13740 5030 13768 5086
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13728 5024 13780 5030
rect 13728 4966 13780 4972
rect 13648 4826 13676 4966
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13924 4706 13952 5102
rect 14004 5092 14056 5098
rect 14004 5034 14056 5040
rect 13832 4678 13952 4706
rect 13832 4486 13860 4678
rect 13912 4548 13964 4554
rect 13912 4490 13964 4496
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13360 4014 13412 4020
rect 13450 4040 13506 4049
rect 13450 3975 13506 3984
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 13648 3466 13676 3946
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13358 2816 13414 2825
rect 13136 2536 13216 2564
rect 13280 2553 13308 2790
rect 13358 2751 13414 2760
rect 13372 2650 13400 2751
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13266 2544 13322 2553
rect 13084 2518 13136 2524
rect 13266 2479 13322 2488
rect 13464 2446 13492 2994
rect 13740 2854 13768 3878
rect 13924 3058 13952 4490
rect 14016 4282 14044 5034
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 14108 3738 14136 4558
rect 14384 4010 14412 6802
rect 14476 4264 14504 8327
rect 14556 8016 14608 8022
rect 14556 7958 14608 7964
rect 14568 7585 14596 7958
rect 14554 7576 14610 7585
rect 14660 7546 14688 12679
rect 14752 12442 14780 14418
rect 14924 14408 14976 14414
rect 14924 14350 14976 14356
rect 15106 14376 15162 14385
rect 14832 13456 14884 13462
rect 14832 13398 14884 13404
rect 14844 13161 14872 13398
rect 14936 13326 14964 14350
rect 15106 14311 15162 14320
rect 14924 13320 14976 13326
rect 14924 13262 14976 13268
rect 14830 13152 14886 13161
rect 14936 13138 14964 13262
rect 14936 13110 15056 13138
rect 14830 13087 14886 13096
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14752 10470 14780 11834
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14738 8528 14794 8537
rect 14738 8463 14794 8472
rect 14752 8362 14780 8463
rect 14740 8356 14792 8362
rect 14740 8298 14792 8304
rect 14554 7511 14610 7520
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 14752 7478 14780 8298
rect 14844 8022 14872 13087
rect 15028 12782 15056 13110
rect 14924 12776 14976 12782
rect 14924 12718 14976 12724
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 14936 12617 14964 12718
rect 14922 12608 14978 12617
rect 14922 12543 14978 12552
rect 14936 10810 14964 12543
rect 15016 12232 15068 12238
rect 15016 12174 15068 12180
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 14924 8356 14976 8362
rect 15028 8344 15056 12174
rect 15120 12170 15148 14311
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 15108 12164 15160 12170
rect 15108 12106 15160 12112
rect 15212 11642 15240 13670
rect 15304 11898 15332 15807
rect 15382 14648 15438 14657
rect 15382 14583 15438 14592
rect 15476 14612 15528 14618
rect 15396 11937 15424 14583
rect 15476 14554 15528 14560
rect 15382 11928 15438 11937
rect 15292 11892 15344 11898
rect 15382 11863 15438 11872
rect 15292 11834 15344 11840
rect 15212 11614 15424 11642
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15106 11248 15162 11257
rect 15106 11183 15162 11192
rect 14976 8316 15056 8344
rect 14924 8298 14976 8304
rect 14832 8016 14884 8022
rect 14832 7958 14884 7964
rect 14936 7834 14964 8298
rect 14844 7806 14964 7834
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 14568 6662 14596 7278
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14660 6458 14688 7346
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14752 6254 14780 7142
rect 14844 7002 14872 7806
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 14832 6996 14884 7002
rect 14832 6938 14884 6944
rect 14924 6928 14976 6934
rect 14924 6870 14976 6876
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14844 6633 14872 6802
rect 14830 6624 14886 6633
rect 14830 6559 14886 6568
rect 14936 6458 14964 6870
rect 15028 6798 15056 7482
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 15120 6644 15148 11183
rect 15212 7206 15240 11494
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15304 10606 15332 11086
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15396 10441 15424 11614
rect 15382 10432 15438 10441
rect 15382 10367 15438 10376
rect 15292 9444 15344 9450
rect 15292 9386 15344 9392
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15028 6616 15148 6644
rect 14924 6452 14976 6458
rect 14924 6394 14976 6400
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 14646 5536 14702 5545
rect 14646 5471 14702 5480
rect 14476 4236 14596 4264
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14372 4004 14424 4010
rect 14372 3946 14424 3952
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14094 3632 14150 3641
rect 14004 3596 14056 3602
rect 14094 3567 14096 3576
rect 14004 3538 14056 3544
rect 14148 3567 14150 3576
rect 14096 3538 14148 3544
rect 14016 3074 14044 3538
rect 14200 3398 14228 3674
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 14292 3194 14320 3878
rect 14476 3618 14504 4082
rect 14384 3590 14504 3618
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14016 3058 14136 3074
rect 13912 3052 13964 3058
rect 14016 3052 14148 3058
rect 14016 3046 14096 3052
rect 13912 2994 13964 3000
rect 14096 2994 14148 3000
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 13542 2680 13598 2689
rect 13542 2615 13598 2624
rect 13556 2582 13584 2615
rect 13544 2576 13596 2582
rect 13544 2518 13596 2524
rect 13636 2508 13688 2514
rect 13636 2450 13688 2456
rect 13452 2440 13504 2446
rect 13452 2382 13504 2388
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 13096 800 13124 2246
rect 13648 1426 13676 2450
rect 13832 2378 13860 2926
rect 14004 2916 14056 2922
rect 14004 2858 14056 2864
rect 14016 2650 14044 2858
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14108 2564 14136 2994
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14200 2689 14228 2926
rect 14186 2680 14242 2689
rect 14186 2615 14242 2624
rect 14384 2582 14412 3590
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14476 3194 14504 3470
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 14372 2576 14424 2582
rect 14108 2536 14228 2564
rect 14200 2446 14228 2536
rect 14372 2518 14424 2524
rect 14568 2514 14596 4236
rect 14660 4185 14688 5471
rect 14646 4176 14702 4185
rect 14646 4111 14702 4120
rect 14660 2854 14688 4111
rect 14740 4004 14792 4010
rect 14740 3946 14792 3952
rect 14752 3194 14780 3946
rect 14844 3942 14872 6054
rect 15028 5273 15056 6616
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15014 5264 15070 5273
rect 15120 5234 15148 5646
rect 15014 5199 15070 5208
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14936 3602 14964 4082
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 14924 3596 14976 3602
rect 14924 3538 14976 3544
rect 14844 3482 14872 3538
rect 15028 3482 15056 4966
rect 15120 4622 15148 5170
rect 15304 5030 15332 9386
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15396 7886 15424 9318
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15396 7274 15424 7822
rect 15384 7268 15436 7274
rect 15384 7210 15436 7216
rect 15396 6866 15424 7210
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15396 6390 15424 6802
rect 15384 6384 15436 6390
rect 15384 6326 15436 6332
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 15396 5370 15424 5782
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 15200 4752 15252 4758
rect 15200 4694 15252 4700
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 15120 4214 15148 4558
rect 15108 4208 15160 4214
rect 15108 4150 15160 4156
rect 14844 3454 15056 3482
rect 15212 3466 15240 4694
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 15200 3460 15252 3466
rect 15200 3402 15252 3408
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 14752 2990 14780 3130
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14832 2984 14884 2990
rect 14832 2926 14884 2932
rect 14648 2848 14700 2854
rect 14648 2790 14700 2796
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 13912 2372 13964 2378
rect 13912 2314 13964 2320
rect 13636 1420 13688 1426
rect 13636 1362 13688 1368
rect 13924 800 13952 2314
rect 14844 800 14872 2926
rect 14936 2922 14964 3062
rect 14924 2916 14976 2922
rect 14924 2858 14976 2864
rect 15304 2650 15332 4422
rect 15382 4040 15438 4049
rect 15382 3975 15384 3984
rect 15436 3975 15438 3984
rect 15384 3946 15436 3952
rect 15488 2990 15516 14554
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15580 12442 15608 13738
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15580 12306 15608 12378
rect 15672 12345 15700 14350
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 15782 14172 16078 14192
rect 15838 14170 15862 14172
rect 15918 14170 15942 14172
rect 15998 14170 16022 14172
rect 15860 14118 15862 14170
rect 15924 14118 15936 14170
rect 15998 14118 16000 14170
rect 15838 14116 15862 14118
rect 15918 14116 15942 14118
rect 15998 14116 16022 14118
rect 15782 14096 16078 14116
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 15948 13326 15976 13874
rect 16224 13802 16252 14214
rect 16592 13938 16620 16200
rect 17958 15056 18014 15065
rect 17958 14991 18014 15000
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16304 13456 16356 13462
rect 16304 13398 16356 13404
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15782 13084 16078 13104
rect 15838 13082 15862 13084
rect 15918 13082 15942 13084
rect 15998 13082 16022 13084
rect 15860 13030 15862 13082
rect 15924 13030 15936 13082
rect 15998 13030 16000 13082
rect 15838 13028 15862 13030
rect 15918 13028 15942 13030
rect 15998 13028 16022 13030
rect 15782 13008 16078 13028
rect 15658 12336 15714 12345
rect 15568 12300 15620 12306
rect 15658 12271 15714 12280
rect 16120 12300 16172 12306
rect 15568 12242 15620 12248
rect 16120 12242 16172 12248
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15568 11824 15620 11830
rect 15568 11766 15620 11772
rect 15580 6254 15608 11766
rect 15672 11762 15700 12038
rect 15782 11996 16078 12016
rect 15838 11994 15862 11996
rect 15918 11994 15942 11996
rect 15998 11994 16022 11996
rect 15860 11942 15862 11994
rect 15924 11942 15936 11994
rect 15998 11942 16000 11994
rect 15838 11940 15862 11942
rect 15918 11940 15942 11942
rect 15998 11940 16022 11942
rect 15782 11920 16078 11940
rect 16132 11898 16160 12242
rect 16212 12232 16264 12238
rect 16316 12209 16344 13398
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 16592 12889 16620 13330
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 16578 12880 16634 12889
rect 16578 12815 16634 12824
rect 16672 12844 16724 12850
rect 16592 12714 16620 12815
rect 16672 12786 16724 12792
rect 16580 12708 16632 12714
rect 16580 12650 16632 12656
rect 16394 12336 16450 12345
rect 16684 12322 16712 12786
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16856 12640 16908 12646
rect 16762 12608 16818 12617
rect 16856 12582 16908 12588
rect 16762 12543 16818 12552
rect 16394 12271 16450 12280
rect 16592 12294 16712 12322
rect 16776 12306 16804 12543
rect 16764 12300 16816 12306
rect 16212 12174 16264 12180
rect 16302 12200 16358 12209
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15672 8294 15700 11154
rect 15782 10908 16078 10928
rect 15838 10906 15862 10908
rect 15918 10906 15942 10908
rect 15998 10906 16022 10908
rect 15860 10854 15862 10906
rect 15924 10854 15936 10906
rect 15998 10854 16000 10906
rect 15838 10852 15862 10854
rect 15918 10852 15942 10854
rect 15998 10852 16022 10854
rect 15782 10832 16078 10852
rect 16132 10810 16160 11698
rect 16224 11354 16252 12174
rect 16302 12135 16358 12144
rect 16302 12064 16358 12073
rect 16302 11999 16358 12008
rect 16316 11694 16344 11999
rect 16304 11688 16356 11694
rect 16304 11630 16356 11636
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16408 10690 16436 12271
rect 16592 12238 16620 12294
rect 16764 12242 16816 12248
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16486 10840 16542 10849
rect 16486 10775 16542 10784
rect 16132 10662 16436 10690
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 15764 9994 15792 10542
rect 15752 9988 15804 9994
rect 15752 9930 15804 9936
rect 15782 9820 16078 9840
rect 15838 9818 15862 9820
rect 15918 9818 15942 9820
rect 15998 9818 16022 9820
rect 15860 9766 15862 9818
rect 15924 9766 15936 9818
rect 15998 9766 16000 9818
rect 15838 9764 15862 9766
rect 15918 9764 15942 9766
rect 15998 9764 16022 9766
rect 15782 9744 16078 9764
rect 15782 8732 16078 8752
rect 15838 8730 15862 8732
rect 15918 8730 15942 8732
rect 15998 8730 16022 8732
rect 15860 8678 15862 8730
rect 15924 8678 15936 8730
rect 15998 8678 16000 8730
rect 15838 8676 15862 8678
rect 15918 8676 15942 8678
rect 15998 8676 16022 8678
rect 15782 8656 16078 8676
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 15936 8424 15988 8430
rect 15936 8366 15988 8372
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15948 8090 15976 8366
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 16040 7954 16068 8434
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15672 7546 15700 7686
rect 15782 7644 16078 7664
rect 15838 7642 15862 7644
rect 15918 7642 15942 7644
rect 15998 7642 16022 7644
rect 15860 7590 15862 7642
rect 15924 7590 15936 7642
rect 15998 7590 16000 7642
rect 15838 7588 15862 7590
rect 15918 7588 15942 7590
rect 15998 7588 16022 7590
rect 15782 7568 16078 7588
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15672 7002 15700 7482
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15782 6556 16078 6576
rect 15838 6554 15862 6556
rect 15918 6554 15942 6556
rect 15998 6554 16022 6556
rect 15860 6502 15862 6554
rect 15924 6502 15936 6554
rect 15998 6502 16000 6554
rect 15838 6500 15862 6502
rect 15918 6500 15942 6502
rect 15998 6500 16022 6502
rect 15782 6480 16078 6500
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15752 5704 15804 5710
rect 15750 5672 15752 5681
rect 15804 5672 15806 5681
rect 15750 5607 15806 5616
rect 15782 5468 16078 5488
rect 15838 5466 15862 5468
rect 15918 5466 15942 5468
rect 15998 5466 16022 5468
rect 15860 5414 15862 5466
rect 15924 5414 15936 5466
rect 15998 5414 16000 5466
rect 15838 5412 15862 5414
rect 15918 5412 15942 5414
rect 15998 5412 16022 5414
rect 15782 5392 16078 5412
rect 15750 5264 15806 5273
rect 15750 5199 15806 5208
rect 15764 4758 15792 5199
rect 16028 5160 16080 5166
rect 16026 5128 16028 5137
rect 16080 5128 16082 5137
rect 16026 5063 16082 5072
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 15948 4826 15976 4966
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 15568 4752 15620 4758
rect 15568 4694 15620 4700
rect 15752 4752 15804 4758
rect 15752 4694 15804 4700
rect 15580 3126 15608 4694
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15672 4593 15700 4626
rect 15658 4584 15714 4593
rect 15658 4519 15714 4528
rect 15782 4380 16078 4400
rect 15838 4378 15862 4380
rect 15918 4378 15942 4380
rect 15998 4378 16022 4380
rect 15860 4326 15862 4378
rect 15924 4326 15936 4378
rect 15998 4326 16000 4378
rect 15838 4324 15862 4326
rect 15918 4324 15942 4326
rect 15998 4324 16022 4326
rect 15782 4304 16078 4324
rect 15782 3292 16078 3312
rect 15838 3290 15862 3292
rect 15918 3290 15942 3292
rect 15998 3290 16022 3292
rect 15860 3238 15862 3290
rect 15924 3238 15936 3290
rect 15998 3238 16000 3290
rect 15838 3236 15862 3238
rect 15918 3236 15942 3238
rect 15998 3236 16022 3238
rect 15782 3216 16078 3236
rect 15568 3120 15620 3126
rect 15568 3062 15620 3068
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15580 2825 15608 2926
rect 15566 2816 15622 2825
rect 15566 2751 15622 2760
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 15782 2204 16078 2224
rect 15838 2202 15862 2204
rect 15918 2202 15942 2204
rect 15998 2202 16022 2204
rect 15860 2150 15862 2202
rect 15924 2150 15936 2202
rect 15998 2150 16000 2202
rect 15838 2148 15862 2150
rect 15918 2148 15942 2150
rect 15998 2148 16022 2150
rect 15782 2128 16078 2148
rect 16132 1442 16160 10662
rect 16394 10568 16450 10577
rect 16394 10503 16450 10512
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16224 9110 16252 10066
rect 16408 9194 16436 10503
rect 16500 9722 16528 10775
rect 16592 10470 16620 12174
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16776 11150 16804 11698
rect 16868 11626 16896 12582
rect 16960 12374 16988 12718
rect 16948 12368 17000 12374
rect 16948 12310 17000 12316
rect 17052 12306 17080 13262
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16488 9716 16540 9722
rect 16488 9658 16540 9664
rect 16684 9654 16712 11086
rect 16776 10198 16804 11086
rect 16764 10192 16816 10198
rect 16764 10134 16816 10140
rect 16960 9897 16988 11494
rect 17052 10810 17080 12242
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 16946 9888 17002 9897
rect 16946 9823 17002 9832
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16408 9166 16528 9194
rect 16212 9104 16264 9110
rect 16212 9046 16264 9052
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 16224 8022 16252 8910
rect 16304 8900 16356 8906
rect 16304 8842 16356 8848
rect 16316 8430 16344 8842
rect 16408 8634 16436 8978
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16500 8514 16528 9166
rect 16408 8486 16528 8514
rect 16304 8424 16356 8430
rect 16304 8366 16356 8372
rect 16212 8016 16264 8022
rect 16212 7958 16264 7964
rect 16302 7984 16358 7993
rect 16224 7546 16252 7958
rect 16302 7919 16358 7928
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16224 2514 16252 7142
rect 16316 7002 16344 7919
rect 16408 7313 16436 8486
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16394 7304 16450 7313
rect 16394 7239 16450 7248
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16316 5914 16344 6802
rect 16408 6118 16436 7239
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 16304 5772 16356 5778
rect 16304 5714 16356 5720
rect 16212 2508 16264 2514
rect 16212 2450 16264 2456
rect 16316 1834 16344 5714
rect 16500 3754 16528 8298
rect 16580 8288 16632 8294
rect 16580 8230 16632 8236
rect 16592 5166 16620 8230
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16868 6798 16896 7482
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 16580 5160 16632 5166
rect 16580 5102 16632 5108
rect 17052 4690 17080 6190
rect 17040 4684 17092 4690
rect 17040 4626 17092 4632
rect 16500 3726 16712 3754
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16488 3460 16540 3466
rect 16488 3402 16540 3408
rect 16396 2848 16448 2854
rect 16396 2790 16448 2796
rect 16408 2582 16436 2790
rect 16396 2576 16448 2582
rect 16396 2518 16448 2524
rect 16304 1828 16356 1834
rect 16304 1770 16356 1776
rect 15764 1414 16160 1442
rect 15764 800 15792 1414
rect 3514 232 3570 241
rect 3514 167 3570 176
rect 3974 0 4030 800
rect 4894 0 4950 800
rect 5814 0 5870 800
rect 6734 0 6790 800
rect 7562 0 7618 800
rect 8482 0 8538 800
rect 9402 0 9458 800
rect 10322 0 10378 800
rect 11242 0 11298 800
rect 12162 0 12218 800
rect 13082 0 13138 800
rect 13910 0 13966 800
rect 14830 0 14886 800
rect 15750 0 15806 800
rect 16500 649 16528 3402
rect 16592 2961 16620 3538
rect 16578 2952 16634 2961
rect 16684 2922 16712 3726
rect 16578 2887 16634 2896
rect 16672 2916 16724 2922
rect 16672 2858 16724 2864
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 16592 2689 16620 2790
rect 16578 2680 16634 2689
rect 16578 2615 16634 2624
rect 17144 2514 17172 13874
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 17236 12782 17264 13126
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 17236 10130 17264 11630
rect 17328 11354 17356 12582
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17420 10146 17448 13806
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17604 13433 17632 13670
rect 17590 13424 17646 13433
rect 17590 13359 17646 13368
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17592 12708 17644 12714
rect 17592 12650 17644 12656
rect 17498 11792 17554 11801
rect 17498 11727 17554 11736
rect 17512 11354 17540 11727
rect 17604 11370 17632 12650
rect 17500 11348 17552 11354
rect 17604 11342 17724 11370
rect 17500 11290 17552 11296
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17604 11014 17632 11154
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17696 10826 17724 11342
rect 17604 10798 17724 10826
rect 17500 10532 17552 10538
rect 17500 10474 17552 10480
rect 17512 10266 17540 10474
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17224 10124 17276 10130
rect 17420 10118 17540 10146
rect 17224 10066 17276 10072
rect 17236 8514 17264 10066
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17328 9081 17356 9318
rect 17314 9072 17370 9081
rect 17420 9042 17448 9522
rect 17314 9007 17370 9016
rect 17408 9036 17460 9042
rect 17408 8978 17460 8984
rect 17420 8634 17448 8978
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17236 8486 17448 8514
rect 17224 6384 17276 6390
rect 17224 6326 17276 6332
rect 17236 4690 17264 6326
rect 17314 5808 17370 5817
rect 17420 5778 17448 8486
rect 17512 7936 17540 10118
rect 17604 8673 17632 10798
rect 17880 10266 17908 13330
rect 17972 11286 18000 14991
rect 18248 14890 18276 16215
rect 18236 14884 18288 14890
rect 18236 14826 18288 14832
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 18064 12322 18092 12378
rect 18064 12294 18184 12322
rect 17960 11280 18012 11286
rect 17960 11222 18012 11228
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17776 10192 17828 10198
rect 17776 10134 17828 10140
rect 17788 9178 17816 10134
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17590 8664 17646 8673
rect 17590 8599 17646 8608
rect 17880 7954 17908 9862
rect 18064 8430 18092 10950
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 17868 7948 17920 7954
rect 17512 7908 17724 7936
rect 17590 7848 17646 7857
rect 17590 7783 17646 7792
rect 17500 7744 17552 7750
rect 17500 7686 17552 7692
rect 17512 7342 17540 7686
rect 17604 7546 17632 7783
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 17500 7336 17552 7342
rect 17500 7278 17552 7284
rect 17592 6112 17644 6118
rect 17590 6080 17592 6089
rect 17644 6080 17646 6089
rect 17590 6015 17646 6024
rect 17314 5743 17316 5752
rect 17368 5743 17370 5752
rect 17408 5772 17460 5778
rect 17316 5714 17368 5720
rect 17408 5714 17460 5720
rect 17498 5672 17554 5681
rect 17498 5607 17500 5616
rect 17552 5607 17554 5616
rect 17500 5578 17552 5584
rect 17224 4684 17276 4690
rect 17224 4626 17276 4632
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 17512 4049 17540 4422
rect 17498 4040 17554 4049
rect 17498 3975 17554 3984
rect 17592 3936 17644 3942
rect 17592 3878 17644 3884
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 17224 2848 17276 2854
rect 17224 2790 17276 2796
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 16684 800 16712 2450
rect 17132 2304 17184 2310
rect 17132 2246 17184 2252
rect 17144 2106 17172 2246
rect 17132 2100 17184 2106
rect 17132 2042 17184 2048
rect 17236 1465 17264 2790
rect 17328 2281 17356 3334
rect 17604 3097 17632 3878
rect 17590 3088 17646 3097
rect 17590 3023 17646 3032
rect 17696 2972 17724 7908
rect 17868 7890 17920 7896
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 18064 7449 18092 7686
rect 17866 7440 17922 7449
rect 18050 7440 18106 7449
rect 17922 7398 18000 7426
rect 17866 7375 17922 7384
rect 17972 6254 18000 7398
rect 18050 7375 18106 7384
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 18064 6497 18092 6598
rect 18050 6488 18106 6497
rect 18050 6423 18106 6432
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17788 4865 17816 5510
rect 17880 5273 17908 6054
rect 17866 5264 17922 5273
rect 17866 5199 17922 5208
rect 17774 4856 17830 4865
rect 17774 4791 17830 4800
rect 17866 4720 17922 4729
rect 17866 4655 17868 4664
rect 17920 4655 17922 4664
rect 17868 4626 17920 4632
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17604 2944 17724 2972
rect 17314 2272 17370 2281
rect 17314 2207 17370 2216
rect 17222 1456 17278 1465
rect 17222 1391 17278 1400
rect 17604 800 17632 2944
rect 17682 2544 17738 2553
rect 17682 2479 17684 2488
rect 17736 2479 17738 2488
rect 17684 2450 17736 2456
rect 17788 1873 17816 3878
rect 17880 3641 17908 4422
rect 18156 4078 18184 12294
rect 18248 11830 18276 14826
rect 18340 13462 18368 16623
rect 18786 16200 18842 17000
rect 18800 14550 18828 16200
rect 18788 14544 18840 14550
rect 18788 14486 18840 14492
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 18328 13456 18380 13462
rect 18328 13398 18380 13404
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18340 11150 18368 13262
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18236 8288 18288 8294
rect 18234 8256 18236 8265
rect 18288 8256 18290 8265
rect 18234 8191 18290 8200
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 18248 7041 18276 7142
rect 18234 7032 18290 7041
rect 18234 6967 18290 6976
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18248 4457 18276 4966
rect 18234 4448 18290 4457
rect 18234 4383 18290 4392
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 17866 3632 17922 3641
rect 17866 3567 17922 3576
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 17868 2304 17920 2310
rect 17868 2246 17920 2252
rect 17774 1864 17830 1873
rect 17774 1799 17830 1808
rect 17880 1057 17908 2246
rect 17866 1048 17922 1057
rect 17866 983 17922 992
rect 16486 640 16542 649
rect 16486 575 16542 584
rect 16670 0 16726 800
rect 17590 0 17646 800
rect 18248 241 18276 2790
rect 18524 800 18552 13942
rect 18786 13288 18842 13297
rect 18786 13223 18842 13232
rect 18800 11354 18828 13223
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 19430 3360 19486 3369
rect 19430 3295 19486 3304
rect 19444 800 19472 3295
rect 18234 232 18290 241
rect 18234 167 18290 176
rect 18510 0 18566 800
rect 19430 0 19486 800
<< via2 >>
rect 4066 16224 4122 16280
rect 2778 15816 2834 15872
rect 1122 12688 1178 12744
rect 2134 12144 2190 12200
rect 1674 11192 1730 11248
rect 2686 11620 2742 11656
rect 2686 11600 2688 11620
rect 2688 11600 2740 11620
rect 2740 11600 2742 11620
rect 3974 15408 4030 15464
rect 8390 16632 8446 16688
rect 3514 15020 3570 15056
rect 3514 15000 3516 15020
rect 3516 15000 3568 15020
rect 3568 15000 3570 15020
rect 4434 14592 4490 14648
rect 3698 14184 3754 14240
rect 3921 14170 3977 14172
rect 4001 14170 4057 14172
rect 4081 14170 4137 14172
rect 4161 14170 4217 14172
rect 3921 14118 3947 14170
rect 3947 14118 3977 14170
rect 4001 14118 4011 14170
rect 4011 14118 4057 14170
rect 4081 14118 4127 14170
rect 4127 14118 4137 14170
rect 4161 14118 4191 14170
rect 4191 14118 4217 14170
rect 3921 14116 3977 14118
rect 4001 14116 4057 14118
rect 4081 14116 4137 14118
rect 4161 14116 4217 14118
rect 3790 13776 3846 13832
rect 4066 13368 4122 13424
rect 3921 13082 3977 13084
rect 4001 13082 4057 13084
rect 4081 13082 4137 13084
rect 4161 13082 4217 13084
rect 3921 13030 3947 13082
rect 3947 13030 3977 13082
rect 4001 13030 4011 13082
rect 4011 13030 4057 13082
rect 4081 13030 4127 13082
rect 4127 13030 4137 13082
rect 4161 13030 4191 13082
rect 4191 13030 4217 13082
rect 3921 13028 3977 13030
rect 4001 13028 4057 13030
rect 4081 13028 4137 13030
rect 4161 13028 4217 13030
rect 3514 12980 3570 13016
rect 3514 12960 3516 12980
rect 3516 12960 3568 12980
rect 3568 12960 3570 12980
rect 3974 12552 4030 12608
rect 2962 12164 3018 12200
rect 2962 12144 2964 12164
rect 2964 12144 3016 12164
rect 3016 12144 3018 12164
rect 3921 11994 3977 11996
rect 4001 11994 4057 11996
rect 4081 11994 4137 11996
rect 4161 11994 4217 11996
rect 3921 11942 3947 11994
rect 3947 11942 3977 11994
rect 4001 11942 4011 11994
rect 4011 11942 4057 11994
rect 4081 11942 4127 11994
rect 4127 11942 4137 11994
rect 4161 11942 4191 11994
rect 4191 11942 4217 11994
rect 3921 11940 3977 11942
rect 4001 11940 4057 11942
rect 4081 11940 4137 11942
rect 4161 11940 4217 11942
rect 3882 11736 3938 11792
rect 2870 9696 2926 9752
rect 2502 8880 2558 8936
rect 1490 7928 1546 7984
rect 1398 7520 1454 7576
rect 1582 1808 1638 1864
rect 1858 6976 1914 7032
rect 3790 11328 3846 11384
rect 3514 10956 3516 10976
rect 3516 10956 3568 10976
rect 3568 10956 3570 10976
rect 3514 10920 3570 10956
rect 2962 8336 3018 8392
rect 2594 6840 2650 6896
rect 2502 3440 2558 3496
rect 2594 3032 2650 3088
rect 1674 1400 1730 1456
rect 2778 6840 2834 6896
rect 3054 6296 3110 6352
rect 3606 10512 3662 10568
rect 3921 10906 3977 10908
rect 4001 10906 4057 10908
rect 4081 10906 4137 10908
rect 4161 10906 4217 10908
rect 3921 10854 3947 10906
rect 3947 10854 3977 10906
rect 4001 10854 4011 10906
rect 4011 10854 4057 10906
rect 4081 10854 4127 10906
rect 4127 10854 4137 10906
rect 4161 10854 4191 10906
rect 4191 10854 4217 10906
rect 3921 10852 3977 10854
rect 4001 10852 4057 10854
rect 4081 10852 4137 10854
rect 4161 10852 4217 10854
rect 4066 10648 4122 10704
rect 3606 6704 3662 6760
rect 3921 9818 3977 9820
rect 4001 9818 4057 9820
rect 4081 9818 4137 9820
rect 4161 9818 4217 9820
rect 3921 9766 3947 9818
rect 3947 9766 3977 9818
rect 4001 9766 4011 9818
rect 4011 9766 4057 9818
rect 4081 9766 4127 9818
rect 4127 9766 4137 9818
rect 4161 9766 4191 9818
rect 4191 9766 4217 9818
rect 3921 9764 3977 9766
rect 4001 9764 4057 9766
rect 4081 9764 4137 9766
rect 4161 9764 4217 9766
rect 4066 9288 4122 9344
rect 3921 8730 3977 8732
rect 4001 8730 4057 8732
rect 4081 8730 4137 8732
rect 4161 8730 4217 8732
rect 3921 8678 3947 8730
rect 3947 8678 3977 8730
rect 4001 8678 4011 8730
rect 4011 8678 4057 8730
rect 4081 8678 4127 8730
rect 4127 8678 4137 8730
rect 4161 8678 4191 8730
rect 4191 8678 4217 8730
rect 3921 8676 3977 8678
rect 4001 8676 4057 8678
rect 4081 8676 4137 8678
rect 4161 8676 4217 8678
rect 4250 8472 4306 8528
rect 4066 7928 4122 7984
rect 3921 7642 3977 7644
rect 4001 7642 4057 7644
rect 4081 7642 4137 7644
rect 4161 7642 4217 7644
rect 3921 7590 3947 7642
rect 3947 7590 3977 7642
rect 4001 7590 4011 7642
rect 4011 7590 4057 7642
rect 4081 7590 4127 7642
rect 4127 7590 4137 7642
rect 4161 7590 4191 7642
rect 4191 7590 4217 7642
rect 3921 7588 3977 7590
rect 4001 7588 4057 7590
rect 4081 7588 4137 7590
rect 4161 7588 4217 7590
rect 3514 5480 3570 5536
rect 3422 5072 3478 5128
rect 3330 4664 3386 4720
rect 2870 992 2926 1048
rect 3238 2624 3294 2680
rect 2778 584 2834 640
rect 3921 6554 3977 6556
rect 4001 6554 4057 6556
rect 4081 6554 4137 6556
rect 4161 6554 4217 6556
rect 3921 6502 3947 6554
rect 3947 6502 3977 6554
rect 4001 6502 4011 6554
rect 4011 6502 4057 6554
rect 4081 6502 4127 6554
rect 4127 6502 4137 6554
rect 4161 6502 4191 6554
rect 4191 6502 4217 6554
rect 3921 6500 3977 6502
rect 4001 6500 4057 6502
rect 4081 6500 4137 6502
rect 4161 6500 4217 6502
rect 3974 5888 4030 5944
rect 5446 12044 5448 12064
rect 5448 12044 5500 12064
rect 5500 12044 5502 12064
rect 5446 12008 5502 12044
rect 4434 7384 4490 7440
rect 3698 4256 3754 4312
rect 3698 2216 3754 2272
rect 3921 5466 3977 5468
rect 4001 5466 4057 5468
rect 4081 5466 4137 5468
rect 4161 5466 4217 5468
rect 3921 5414 3947 5466
rect 3947 5414 3977 5466
rect 4001 5414 4011 5466
rect 4011 5414 4057 5466
rect 4081 5414 4127 5466
rect 4127 5414 4137 5466
rect 4161 5414 4191 5466
rect 4191 5414 4217 5466
rect 3921 5412 3977 5414
rect 4001 5412 4057 5414
rect 4081 5412 4137 5414
rect 4161 5412 4217 5414
rect 4158 5208 4214 5264
rect 3921 4378 3977 4380
rect 4001 4378 4057 4380
rect 4081 4378 4137 4380
rect 4161 4378 4217 4380
rect 3921 4326 3947 4378
rect 3947 4326 3977 4378
rect 4001 4326 4011 4378
rect 4011 4326 4057 4378
rect 4081 4326 4127 4378
rect 4127 4326 4137 4378
rect 4161 4326 4191 4378
rect 4191 4326 4217 4378
rect 3921 4324 3977 4326
rect 4001 4324 4057 4326
rect 4081 4324 4137 4326
rect 4161 4324 4217 4326
rect 4066 3848 4122 3904
rect 4894 10124 4950 10160
rect 4894 10104 4896 10124
rect 4896 10104 4948 10124
rect 4948 10104 4950 10124
rect 4986 9968 5042 10024
rect 4710 9832 4766 9888
rect 5078 9016 5134 9072
rect 4618 5616 4674 5672
rect 4526 4664 4582 4720
rect 3921 3290 3977 3292
rect 4001 3290 4057 3292
rect 4081 3290 4137 3292
rect 4161 3290 4217 3292
rect 3921 3238 3947 3290
rect 3947 3238 3977 3290
rect 4001 3238 4011 3290
rect 4011 3238 4057 3290
rect 4081 3238 4127 3290
rect 4127 3238 4137 3290
rect 4161 3238 4191 3290
rect 4191 3238 4217 3290
rect 3921 3236 3977 3238
rect 4001 3236 4057 3238
rect 4081 3236 4137 3238
rect 4161 3236 4217 3238
rect 3882 2916 3938 2952
rect 3882 2896 3884 2916
rect 3884 2896 3936 2916
rect 3936 2896 3938 2916
rect 3921 2202 3977 2204
rect 4001 2202 4057 2204
rect 4081 2202 4137 2204
rect 4161 2202 4217 2204
rect 3921 2150 3947 2202
rect 3947 2150 3977 2202
rect 4001 2150 4011 2202
rect 4011 2150 4057 2202
rect 4081 2150 4127 2202
rect 4127 2150 4137 2202
rect 4161 2150 4191 2202
rect 4191 2150 4217 2202
rect 3921 2148 3977 2150
rect 4001 2148 4057 2150
rect 4081 2148 4137 2150
rect 4161 2148 4217 2150
rect 5354 10104 5410 10160
rect 5262 7656 5318 7712
rect 5354 7112 5410 7168
rect 5906 13232 5962 13288
rect 5998 12844 6054 12880
rect 5998 12824 6000 12844
rect 6000 12824 6052 12844
rect 6052 12824 6054 12844
rect 5630 8744 5686 8800
rect 5906 9444 5962 9480
rect 5906 9424 5908 9444
rect 5908 9424 5960 9444
rect 5960 9424 5962 9444
rect 5538 6976 5594 7032
rect 5630 4528 5686 4584
rect 5906 8744 5962 8800
rect 6090 9832 6146 9888
rect 5998 8064 6054 8120
rect 6886 14714 6942 14716
rect 6966 14714 7022 14716
rect 7046 14714 7102 14716
rect 7126 14714 7182 14716
rect 6886 14662 6912 14714
rect 6912 14662 6942 14714
rect 6966 14662 6976 14714
rect 6976 14662 7022 14714
rect 7046 14662 7092 14714
rect 7092 14662 7102 14714
rect 7126 14662 7156 14714
rect 7156 14662 7182 14714
rect 6886 14660 6942 14662
rect 6966 14660 7022 14662
rect 7046 14660 7102 14662
rect 7126 14660 7182 14662
rect 6886 13626 6942 13628
rect 6966 13626 7022 13628
rect 7046 13626 7102 13628
rect 7126 13626 7182 13628
rect 6886 13574 6912 13626
rect 6912 13574 6942 13626
rect 6966 13574 6976 13626
rect 6976 13574 7022 13626
rect 7046 13574 7092 13626
rect 7092 13574 7102 13626
rect 7126 13574 7156 13626
rect 7156 13574 7182 13626
rect 6886 13572 6942 13574
rect 6966 13572 7022 13574
rect 7046 13572 7102 13574
rect 7126 13572 7182 13574
rect 6366 12280 6422 12336
rect 6182 8472 6238 8528
rect 5814 5480 5870 5536
rect 6550 8472 6606 8528
rect 6458 8336 6514 8392
rect 6458 8084 6514 8120
rect 6458 8064 6460 8084
rect 6460 8064 6512 8084
rect 6512 8064 6514 8084
rect 6182 7248 6238 7304
rect 6274 5072 6330 5128
rect 5722 3440 5778 3496
rect 6458 5228 6514 5264
rect 6458 5208 6460 5228
rect 6460 5208 6512 5228
rect 6512 5208 6514 5228
rect 7470 12960 7526 13016
rect 6886 12538 6942 12540
rect 6966 12538 7022 12540
rect 7046 12538 7102 12540
rect 7126 12538 7182 12540
rect 6886 12486 6912 12538
rect 6912 12486 6942 12538
rect 6966 12486 6976 12538
rect 6976 12486 7022 12538
rect 7046 12486 7092 12538
rect 7092 12486 7102 12538
rect 7126 12486 7156 12538
rect 7156 12486 7182 12538
rect 6886 12484 6942 12486
rect 6966 12484 7022 12486
rect 7046 12484 7102 12486
rect 7126 12484 7182 12486
rect 7010 12008 7066 12064
rect 6886 11450 6942 11452
rect 6966 11450 7022 11452
rect 7046 11450 7102 11452
rect 7126 11450 7182 11452
rect 6886 11398 6912 11450
rect 6912 11398 6942 11450
rect 6966 11398 6976 11450
rect 6976 11398 7022 11450
rect 7046 11398 7092 11450
rect 7092 11398 7102 11450
rect 7126 11398 7156 11450
rect 7156 11398 7182 11450
rect 6886 11396 6942 11398
rect 6966 11396 7022 11398
rect 7046 11396 7102 11398
rect 7126 11396 7182 11398
rect 6918 11056 6974 11112
rect 8022 12980 8078 13016
rect 8022 12960 8024 12980
rect 8024 12960 8076 12980
rect 8076 12960 8078 12980
rect 7838 12824 7894 12880
rect 7470 10920 7526 10976
rect 6826 10512 6882 10568
rect 6886 10362 6942 10364
rect 6966 10362 7022 10364
rect 7046 10362 7102 10364
rect 7126 10362 7182 10364
rect 6886 10310 6912 10362
rect 6912 10310 6942 10362
rect 6966 10310 6976 10362
rect 6976 10310 7022 10362
rect 7046 10310 7092 10362
rect 7092 10310 7102 10362
rect 7126 10310 7156 10362
rect 7156 10310 7182 10362
rect 6886 10308 6942 10310
rect 6966 10308 7022 10310
rect 7046 10308 7102 10310
rect 7126 10308 7182 10310
rect 6886 9274 6942 9276
rect 6966 9274 7022 9276
rect 7046 9274 7102 9276
rect 7126 9274 7182 9276
rect 6886 9222 6912 9274
rect 6912 9222 6942 9274
rect 6966 9222 6976 9274
rect 6976 9222 7022 9274
rect 7046 9222 7092 9274
rect 7092 9222 7102 9274
rect 7126 9222 7156 9274
rect 7156 9222 7182 9274
rect 6886 9220 6942 9222
rect 6966 9220 7022 9222
rect 7046 9220 7102 9222
rect 7126 9220 7182 9222
rect 7470 8608 7526 8664
rect 6886 8186 6942 8188
rect 6966 8186 7022 8188
rect 7046 8186 7102 8188
rect 7126 8186 7182 8188
rect 6886 8134 6912 8186
rect 6912 8134 6942 8186
rect 6966 8134 6976 8186
rect 6976 8134 7022 8186
rect 7046 8134 7092 8186
rect 7092 8134 7102 8186
rect 7126 8134 7156 8186
rect 7156 8134 7182 8186
rect 6886 8132 6942 8134
rect 6966 8132 7022 8134
rect 7046 8132 7102 8134
rect 7126 8132 7182 8134
rect 7654 11192 7710 11248
rect 7838 12144 7894 12200
rect 7838 11600 7894 11656
rect 7562 8336 7618 8392
rect 7562 7964 7564 7984
rect 7564 7964 7616 7984
rect 7616 7964 7618 7984
rect 7562 7928 7618 7964
rect 8114 11348 8170 11384
rect 8114 11328 8116 11348
rect 8116 11328 8168 11348
rect 8168 11328 8170 11348
rect 8114 10104 8170 10160
rect 7746 7656 7802 7712
rect 7562 7248 7618 7304
rect 6886 7098 6942 7100
rect 6966 7098 7022 7100
rect 7046 7098 7102 7100
rect 7126 7098 7182 7100
rect 6886 7046 6912 7098
rect 6912 7046 6942 7098
rect 6966 7046 6976 7098
rect 6976 7046 7022 7098
rect 7046 7046 7092 7098
rect 7092 7046 7102 7098
rect 7126 7046 7156 7098
rect 7156 7046 7182 7098
rect 6886 7044 6942 7046
rect 6966 7044 7022 7046
rect 7046 7044 7102 7046
rect 7126 7044 7182 7046
rect 6918 6604 6920 6624
rect 6920 6604 6972 6624
rect 6972 6604 6974 6624
rect 6918 6568 6974 6604
rect 6918 6432 6974 6488
rect 6886 6010 6942 6012
rect 6966 6010 7022 6012
rect 7046 6010 7102 6012
rect 7126 6010 7182 6012
rect 6886 5958 6912 6010
rect 6912 5958 6942 6010
rect 6966 5958 6976 6010
rect 6976 5958 7022 6010
rect 7046 5958 7092 6010
rect 7092 5958 7102 6010
rect 7126 5958 7156 6010
rect 7156 5958 7182 6010
rect 6886 5956 6942 5958
rect 6966 5956 7022 5958
rect 7046 5956 7102 5958
rect 7126 5956 7182 5958
rect 7286 5752 7342 5808
rect 7194 5616 7250 5672
rect 7562 6568 7618 6624
rect 6918 5208 6974 5264
rect 6886 4922 6942 4924
rect 6966 4922 7022 4924
rect 7046 4922 7102 4924
rect 7126 4922 7182 4924
rect 6886 4870 6912 4922
rect 6912 4870 6942 4922
rect 6966 4870 6976 4922
rect 6976 4870 7022 4922
rect 7046 4870 7092 4922
rect 7092 4870 7102 4922
rect 7126 4870 7156 4922
rect 7156 4870 7182 4922
rect 6886 4868 6942 4870
rect 6966 4868 7022 4870
rect 7046 4868 7102 4870
rect 7126 4868 7182 4870
rect 7194 4120 7250 4176
rect 6886 3834 6942 3836
rect 6966 3834 7022 3836
rect 7046 3834 7102 3836
rect 7126 3834 7182 3836
rect 6886 3782 6912 3834
rect 6912 3782 6942 3834
rect 6966 3782 6976 3834
rect 6976 3782 7022 3834
rect 7046 3782 7092 3834
rect 7092 3782 7102 3834
rect 7126 3782 7156 3834
rect 7156 3782 7182 3834
rect 6886 3780 6942 3782
rect 6966 3780 7022 3782
rect 7046 3780 7102 3782
rect 7126 3780 7182 3782
rect 6886 2746 6942 2748
rect 6966 2746 7022 2748
rect 7046 2746 7102 2748
rect 7126 2746 7182 2748
rect 6886 2694 6912 2746
rect 6912 2694 6942 2746
rect 6966 2694 6976 2746
rect 6976 2694 7022 2746
rect 7046 2694 7092 2746
rect 7092 2694 7102 2746
rect 7126 2694 7156 2746
rect 7156 2694 7182 2746
rect 6886 2692 6942 2694
rect 6966 2692 7022 2694
rect 7046 2692 7102 2694
rect 7126 2692 7182 2694
rect 7562 5752 7618 5808
rect 7746 5516 7748 5536
rect 7748 5516 7800 5536
rect 7800 5516 7802 5536
rect 7746 5480 7802 5516
rect 8022 6432 8078 6488
rect 8206 3984 8262 4040
rect 18326 16632 18382 16688
rect 18234 16224 18290 16280
rect 9402 13388 9458 13424
rect 9402 13368 9404 13388
rect 9404 13368 9456 13388
rect 9456 13368 9458 13388
rect 9034 11192 9090 11248
rect 9310 12144 9366 12200
rect 9126 11056 9182 11112
rect 9218 10512 9274 10568
rect 8666 9424 8722 9480
rect 8390 7792 8446 7848
rect 8942 7384 8998 7440
rect 8942 7268 8998 7304
rect 8942 7248 8944 7268
rect 8944 7248 8996 7268
rect 8996 7248 8998 7268
rect 8666 5208 8722 5264
rect 8114 2932 8116 2952
rect 8116 2932 8168 2952
rect 8168 2932 8170 2952
rect 8114 2896 8170 2932
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9878 14170
rect 9878 14118 9908 14170
rect 9932 14118 9942 14170
rect 9942 14118 9988 14170
rect 10012 14118 10058 14170
rect 10058 14118 10068 14170
rect 10092 14118 10122 14170
rect 10122 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9878 13082
rect 9878 13030 9908 13082
rect 9932 13030 9942 13082
rect 9942 13030 9988 13082
rect 10012 13030 10058 13082
rect 10058 13030 10068 13082
rect 10092 13030 10122 13082
rect 10122 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 10230 12824 10286 12880
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9878 11994
rect 9878 11942 9908 11994
rect 9932 11942 9942 11994
rect 9942 11942 9988 11994
rect 10012 11942 10058 11994
rect 10058 11942 10068 11994
rect 10092 11942 10122 11994
rect 10122 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 9402 7792 9458 7848
rect 9862 11348 9918 11384
rect 9862 11328 9864 11348
rect 9864 11328 9916 11348
rect 9916 11328 9918 11348
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9878 10906
rect 9878 10854 9908 10906
rect 9932 10854 9942 10906
rect 9942 10854 9988 10906
rect 10012 10854 10058 10906
rect 10058 10854 10068 10906
rect 10092 10854 10122 10906
rect 10122 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9878 9818
rect 9878 9766 9908 9818
rect 9932 9766 9942 9818
rect 9942 9766 9988 9818
rect 10012 9766 10058 9818
rect 10058 9766 10068 9818
rect 10092 9766 10122 9818
rect 10122 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9878 8730
rect 9878 8678 9908 8730
rect 9932 8678 9942 8730
rect 9942 8678 9988 8730
rect 10012 8678 10058 8730
rect 10058 8678 10068 8730
rect 10092 8678 10122 8730
rect 10122 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 10322 11736 10378 11792
rect 10506 12280 10562 12336
rect 10690 13096 10746 13152
rect 10506 9968 10562 10024
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9878 7642
rect 9878 7590 9908 7642
rect 9932 7590 9942 7642
rect 9942 7590 9988 7642
rect 10012 7590 10058 7642
rect 10058 7590 10068 7642
rect 10092 7590 10122 7642
rect 10122 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 10138 6976 10194 7032
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9878 6554
rect 9878 6502 9908 6554
rect 9932 6502 9942 6554
rect 9942 6502 9988 6554
rect 10012 6502 10058 6554
rect 10058 6502 10068 6554
rect 10092 6502 10122 6554
rect 10122 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9878 5466
rect 9878 5414 9908 5466
rect 9932 5414 9942 5466
rect 9942 5414 9988 5466
rect 10012 5414 10058 5466
rect 10058 5414 10068 5466
rect 10092 5414 10122 5466
rect 10122 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9878 4378
rect 9878 4326 9908 4378
rect 9932 4326 9942 4378
rect 9942 4326 9988 4378
rect 10012 4326 10058 4378
rect 10058 4326 10068 4378
rect 10092 4326 10122 4378
rect 10122 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 10414 5616 10470 5672
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9878 3290
rect 9878 3238 9908 3290
rect 9932 3238 9942 3290
rect 9942 3238 9988 3290
rect 10012 3238 10058 3290
rect 10058 3238 10068 3290
rect 10092 3238 10122 3290
rect 10122 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9878 2202
rect 9878 2150 9908 2202
rect 9932 2150 9942 2202
rect 9942 2150 9988 2202
rect 10012 2150 10058 2202
rect 10058 2150 10068 2202
rect 10092 2150 10122 2202
rect 10122 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 10966 13096 11022 13152
rect 10966 11228 10968 11248
rect 10968 11228 11020 11248
rect 11020 11228 11022 11248
rect 10966 11192 11022 11228
rect 10966 8336 11022 8392
rect 10782 7248 10838 7304
rect 10690 6160 10746 6216
rect 11058 3984 11114 4040
rect 11426 11600 11482 11656
rect 12817 14714 12873 14716
rect 12897 14714 12953 14716
rect 12977 14714 13033 14716
rect 13057 14714 13113 14716
rect 12817 14662 12843 14714
rect 12843 14662 12873 14714
rect 12897 14662 12907 14714
rect 12907 14662 12953 14714
rect 12977 14662 13023 14714
rect 13023 14662 13033 14714
rect 13057 14662 13087 14714
rect 13087 14662 13113 14714
rect 12817 14660 12873 14662
rect 12897 14660 12953 14662
rect 12977 14660 13033 14662
rect 13057 14660 13113 14662
rect 15290 15816 15346 15872
rect 15106 15408 15162 15464
rect 12817 13626 12873 13628
rect 12897 13626 12953 13628
rect 12977 13626 13033 13628
rect 13057 13626 13113 13628
rect 12817 13574 12843 13626
rect 12843 13574 12873 13626
rect 12897 13574 12907 13626
rect 12907 13574 12953 13626
rect 12977 13574 13023 13626
rect 13023 13574 13033 13626
rect 13057 13574 13087 13626
rect 13087 13574 13113 13626
rect 12817 13572 12873 13574
rect 12897 13572 12953 13574
rect 12977 13572 13033 13574
rect 13057 13572 13113 13574
rect 11518 8064 11574 8120
rect 11610 7828 11612 7848
rect 11612 7828 11664 7848
rect 11664 7828 11666 7848
rect 11610 7792 11666 7828
rect 11426 7384 11482 7440
rect 11334 6432 11390 6488
rect 11242 5072 11298 5128
rect 11426 5108 11428 5128
rect 11428 5108 11480 5128
rect 11480 5108 11482 5128
rect 11426 5072 11482 5108
rect 11242 4664 11298 4720
rect 11794 5752 11850 5808
rect 11886 3576 11942 3632
rect 13174 12688 13230 12744
rect 12817 12538 12873 12540
rect 12897 12538 12953 12540
rect 12977 12538 13033 12540
rect 13057 12538 13113 12540
rect 12817 12486 12843 12538
rect 12843 12486 12873 12538
rect 12897 12486 12907 12538
rect 12907 12486 12953 12538
rect 12977 12486 13023 12538
rect 13023 12486 13033 12538
rect 13057 12486 13087 12538
rect 13087 12486 13113 12538
rect 12817 12484 12873 12486
rect 12897 12484 12953 12486
rect 12977 12484 13033 12486
rect 13057 12484 13113 12486
rect 12806 11600 12862 11656
rect 12817 11450 12873 11452
rect 12897 11450 12953 11452
rect 12977 11450 13033 11452
rect 13057 11450 13113 11452
rect 12817 11398 12843 11450
rect 12843 11398 12873 11450
rect 12897 11398 12907 11450
rect 12907 11398 12953 11450
rect 12977 11398 13023 11450
rect 13023 11398 13033 11450
rect 13057 11398 13087 11450
rect 13087 11398 13113 11450
rect 12817 11396 12873 11398
rect 12897 11396 12953 11398
rect 12977 11396 13033 11398
rect 13057 11396 13113 11398
rect 12346 11056 12402 11112
rect 12346 9968 12402 10024
rect 12817 10362 12873 10364
rect 12897 10362 12953 10364
rect 12977 10362 13033 10364
rect 13057 10362 13113 10364
rect 12817 10310 12843 10362
rect 12843 10310 12873 10362
rect 12897 10310 12907 10362
rect 12907 10310 12953 10362
rect 12977 10310 13023 10362
rect 13023 10310 13033 10362
rect 13057 10310 13087 10362
rect 13087 10310 13113 10362
rect 12817 10308 12873 10310
rect 12897 10308 12953 10310
rect 12977 10308 13033 10310
rect 13057 10308 13113 10310
rect 12346 8880 12402 8936
rect 12817 9274 12873 9276
rect 12897 9274 12953 9276
rect 12977 9274 13033 9276
rect 13057 9274 13113 9276
rect 12817 9222 12843 9274
rect 12843 9222 12873 9274
rect 12897 9222 12907 9274
rect 12907 9222 12953 9274
rect 12977 9222 13023 9274
rect 13023 9222 13033 9274
rect 13057 9222 13087 9274
rect 13087 9222 13113 9274
rect 12817 9220 12873 9222
rect 12897 9220 12953 9222
rect 12977 9220 13033 9222
rect 13057 9220 13113 9222
rect 12254 6976 12310 7032
rect 12346 6840 12402 6896
rect 12254 6704 12310 6760
rect 12530 6840 12586 6896
rect 12817 8186 12873 8188
rect 12897 8186 12953 8188
rect 12977 8186 13033 8188
rect 13057 8186 13113 8188
rect 12817 8134 12843 8186
rect 12843 8134 12873 8186
rect 12897 8134 12907 8186
rect 12907 8134 12953 8186
rect 12977 8134 13023 8186
rect 13023 8134 13033 8186
rect 13057 8134 13087 8186
rect 13087 8134 13113 8186
rect 12817 8132 12873 8134
rect 12897 8132 12953 8134
rect 12977 8132 13033 8134
rect 13057 8132 13113 8134
rect 13634 12688 13690 12744
rect 13542 11056 13598 11112
rect 13634 9424 13690 9480
rect 13542 9016 13598 9072
rect 13082 7520 13138 7576
rect 12817 7098 12873 7100
rect 12897 7098 12953 7100
rect 12977 7098 13033 7100
rect 13057 7098 13113 7100
rect 12817 7046 12843 7098
rect 12843 7046 12873 7098
rect 12897 7046 12907 7098
rect 12907 7046 12953 7098
rect 12977 7046 13023 7098
rect 13023 7046 13033 7098
rect 13057 7046 13087 7098
rect 13087 7046 13113 7098
rect 12817 7044 12873 7046
rect 12897 7044 12953 7046
rect 12977 7044 13033 7046
rect 13057 7044 13113 7046
rect 12714 6840 12770 6896
rect 12990 6568 13046 6624
rect 12898 6296 12954 6352
rect 12817 6010 12873 6012
rect 12897 6010 12953 6012
rect 12977 6010 13033 6012
rect 13057 6010 13113 6012
rect 12817 5958 12843 6010
rect 12843 5958 12873 6010
rect 12897 5958 12907 6010
rect 12907 5958 12953 6010
rect 12977 5958 13023 6010
rect 13023 5958 13033 6010
rect 13057 5958 13087 6010
rect 13087 5958 13113 6010
rect 12817 5956 12873 5958
rect 12897 5956 12953 5958
rect 12977 5956 13033 5958
rect 13057 5956 13113 5958
rect 12817 4922 12873 4924
rect 12897 4922 12953 4924
rect 12977 4922 13033 4924
rect 13057 4922 13113 4924
rect 12817 4870 12843 4922
rect 12843 4870 12873 4922
rect 12897 4870 12907 4922
rect 12907 4870 12953 4922
rect 12977 4870 13023 4922
rect 13023 4870 13033 4922
rect 13057 4870 13087 4922
rect 13087 4870 13113 4922
rect 12817 4868 12873 4870
rect 12897 4868 12953 4870
rect 12977 4868 13033 4870
rect 13057 4868 13113 4870
rect 13450 6840 13506 6896
rect 13450 6160 13506 6216
rect 13818 11192 13874 11248
rect 13910 10376 13966 10432
rect 12817 3834 12873 3836
rect 12897 3834 12953 3836
rect 12977 3834 13033 3836
rect 13057 3834 13113 3836
rect 12817 3782 12843 3834
rect 12843 3782 12873 3834
rect 12897 3782 12907 3834
rect 12907 3782 12953 3834
rect 12977 3782 13023 3834
rect 13023 3782 13033 3834
rect 13057 3782 13087 3834
rect 13087 3782 13113 3834
rect 12817 3780 12873 3782
rect 12897 3780 12953 3782
rect 12977 3780 13033 3782
rect 13057 3780 13113 3782
rect 12817 2746 12873 2748
rect 12897 2746 12953 2748
rect 12977 2746 13033 2748
rect 13057 2746 13113 2748
rect 12817 2694 12843 2746
rect 12843 2694 12873 2746
rect 12897 2694 12907 2746
rect 12907 2694 12953 2746
rect 12977 2694 13023 2746
rect 13023 2694 13033 2746
rect 13057 2694 13087 2746
rect 13087 2694 13113 2746
rect 12817 2692 12873 2694
rect 12897 2692 12953 2694
rect 12977 2692 13033 2694
rect 13057 2692 13113 2694
rect 14646 12688 14702 12744
rect 14554 11600 14610 11656
rect 14094 8880 14150 8936
rect 14370 10648 14426 10704
rect 14462 8336 14518 8392
rect 14002 6704 14058 6760
rect 13818 6296 13874 6352
rect 14094 6432 14150 6488
rect 13450 3984 13506 4040
rect 13358 2760 13414 2816
rect 13266 2488 13322 2544
rect 14554 7520 14610 7576
rect 15106 14320 15162 14376
rect 14830 13096 14886 13152
rect 14738 8472 14794 8528
rect 14922 12552 14978 12608
rect 15382 14592 15438 14648
rect 15382 11872 15438 11928
rect 15106 11192 15162 11248
rect 14830 6568 14886 6624
rect 15382 10376 15438 10432
rect 14646 5480 14702 5536
rect 14094 3596 14150 3632
rect 14094 3576 14096 3596
rect 14096 3576 14148 3596
rect 14148 3576 14150 3596
rect 13542 2624 13598 2680
rect 14186 2624 14242 2680
rect 14646 4120 14702 4176
rect 15014 5208 15070 5264
rect 15382 4004 15438 4040
rect 15382 3984 15384 4004
rect 15384 3984 15436 4004
rect 15436 3984 15438 4004
rect 15782 14170 15838 14172
rect 15862 14170 15918 14172
rect 15942 14170 15998 14172
rect 16022 14170 16078 14172
rect 15782 14118 15808 14170
rect 15808 14118 15838 14170
rect 15862 14118 15872 14170
rect 15872 14118 15918 14170
rect 15942 14118 15988 14170
rect 15988 14118 15998 14170
rect 16022 14118 16052 14170
rect 16052 14118 16078 14170
rect 15782 14116 15838 14118
rect 15862 14116 15918 14118
rect 15942 14116 15998 14118
rect 16022 14116 16078 14118
rect 17958 15000 18014 15056
rect 15782 13082 15838 13084
rect 15862 13082 15918 13084
rect 15942 13082 15998 13084
rect 16022 13082 16078 13084
rect 15782 13030 15808 13082
rect 15808 13030 15838 13082
rect 15862 13030 15872 13082
rect 15872 13030 15918 13082
rect 15942 13030 15988 13082
rect 15988 13030 15998 13082
rect 16022 13030 16052 13082
rect 16052 13030 16078 13082
rect 15782 13028 15838 13030
rect 15862 13028 15918 13030
rect 15942 13028 15998 13030
rect 16022 13028 16078 13030
rect 15658 12280 15714 12336
rect 15782 11994 15838 11996
rect 15862 11994 15918 11996
rect 15942 11994 15998 11996
rect 16022 11994 16078 11996
rect 15782 11942 15808 11994
rect 15808 11942 15838 11994
rect 15862 11942 15872 11994
rect 15872 11942 15918 11994
rect 15942 11942 15988 11994
rect 15988 11942 15998 11994
rect 16022 11942 16052 11994
rect 16052 11942 16078 11994
rect 15782 11940 15838 11942
rect 15862 11940 15918 11942
rect 15942 11940 15998 11942
rect 16022 11940 16078 11942
rect 16578 12824 16634 12880
rect 16394 12280 16450 12336
rect 16762 12552 16818 12608
rect 15782 10906 15838 10908
rect 15862 10906 15918 10908
rect 15942 10906 15998 10908
rect 16022 10906 16078 10908
rect 15782 10854 15808 10906
rect 15808 10854 15838 10906
rect 15862 10854 15872 10906
rect 15872 10854 15918 10906
rect 15942 10854 15988 10906
rect 15988 10854 15998 10906
rect 16022 10854 16052 10906
rect 16052 10854 16078 10906
rect 15782 10852 15838 10854
rect 15862 10852 15918 10854
rect 15942 10852 15998 10854
rect 16022 10852 16078 10854
rect 16302 12144 16358 12200
rect 16302 12008 16358 12064
rect 16486 10784 16542 10840
rect 15782 9818 15838 9820
rect 15862 9818 15918 9820
rect 15942 9818 15998 9820
rect 16022 9818 16078 9820
rect 15782 9766 15808 9818
rect 15808 9766 15838 9818
rect 15862 9766 15872 9818
rect 15872 9766 15918 9818
rect 15942 9766 15988 9818
rect 15988 9766 15998 9818
rect 16022 9766 16052 9818
rect 16052 9766 16078 9818
rect 15782 9764 15838 9766
rect 15862 9764 15918 9766
rect 15942 9764 15998 9766
rect 16022 9764 16078 9766
rect 15782 8730 15838 8732
rect 15862 8730 15918 8732
rect 15942 8730 15998 8732
rect 16022 8730 16078 8732
rect 15782 8678 15808 8730
rect 15808 8678 15838 8730
rect 15862 8678 15872 8730
rect 15872 8678 15918 8730
rect 15942 8678 15988 8730
rect 15988 8678 15998 8730
rect 16022 8678 16052 8730
rect 16052 8678 16078 8730
rect 15782 8676 15838 8678
rect 15862 8676 15918 8678
rect 15942 8676 15998 8678
rect 16022 8676 16078 8678
rect 15782 7642 15838 7644
rect 15862 7642 15918 7644
rect 15942 7642 15998 7644
rect 16022 7642 16078 7644
rect 15782 7590 15808 7642
rect 15808 7590 15838 7642
rect 15862 7590 15872 7642
rect 15872 7590 15918 7642
rect 15942 7590 15988 7642
rect 15988 7590 15998 7642
rect 16022 7590 16052 7642
rect 16052 7590 16078 7642
rect 15782 7588 15838 7590
rect 15862 7588 15918 7590
rect 15942 7588 15998 7590
rect 16022 7588 16078 7590
rect 15782 6554 15838 6556
rect 15862 6554 15918 6556
rect 15942 6554 15998 6556
rect 16022 6554 16078 6556
rect 15782 6502 15808 6554
rect 15808 6502 15838 6554
rect 15862 6502 15872 6554
rect 15872 6502 15918 6554
rect 15942 6502 15988 6554
rect 15988 6502 15998 6554
rect 16022 6502 16052 6554
rect 16052 6502 16078 6554
rect 15782 6500 15838 6502
rect 15862 6500 15918 6502
rect 15942 6500 15998 6502
rect 16022 6500 16078 6502
rect 15750 5652 15752 5672
rect 15752 5652 15804 5672
rect 15804 5652 15806 5672
rect 15750 5616 15806 5652
rect 15782 5466 15838 5468
rect 15862 5466 15918 5468
rect 15942 5466 15998 5468
rect 16022 5466 16078 5468
rect 15782 5414 15808 5466
rect 15808 5414 15838 5466
rect 15862 5414 15872 5466
rect 15872 5414 15918 5466
rect 15942 5414 15988 5466
rect 15988 5414 15998 5466
rect 16022 5414 16052 5466
rect 16052 5414 16078 5466
rect 15782 5412 15838 5414
rect 15862 5412 15918 5414
rect 15942 5412 15998 5414
rect 16022 5412 16078 5414
rect 15750 5208 15806 5264
rect 16026 5108 16028 5128
rect 16028 5108 16080 5128
rect 16080 5108 16082 5128
rect 16026 5072 16082 5108
rect 15658 4528 15714 4584
rect 15782 4378 15838 4380
rect 15862 4378 15918 4380
rect 15942 4378 15998 4380
rect 16022 4378 16078 4380
rect 15782 4326 15808 4378
rect 15808 4326 15838 4378
rect 15862 4326 15872 4378
rect 15872 4326 15918 4378
rect 15942 4326 15988 4378
rect 15988 4326 15998 4378
rect 16022 4326 16052 4378
rect 16052 4326 16078 4378
rect 15782 4324 15838 4326
rect 15862 4324 15918 4326
rect 15942 4324 15998 4326
rect 16022 4324 16078 4326
rect 15782 3290 15838 3292
rect 15862 3290 15918 3292
rect 15942 3290 15998 3292
rect 16022 3290 16078 3292
rect 15782 3238 15808 3290
rect 15808 3238 15838 3290
rect 15862 3238 15872 3290
rect 15872 3238 15918 3290
rect 15942 3238 15988 3290
rect 15988 3238 15998 3290
rect 16022 3238 16052 3290
rect 16052 3238 16078 3290
rect 15782 3236 15838 3238
rect 15862 3236 15918 3238
rect 15942 3236 15998 3238
rect 16022 3236 16078 3238
rect 15566 2760 15622 2816
rect 15782 2202 15838 2204
rect 15862 2202 15918 2204
rect 15942 2202 15998 2204
rect 16022 2202 16078 2204
rect 15782 2150 15808 2202
rect 15808 2150 15838 2202
rect 15862 2150 15872 2202
rect 15872 2150 15918 2202
rect 15942 2150 15988 2202
rect 15988 2150 15998 2202
rect 16022 2150 16052 2202
rect 16052 2150 16078 2202
rect 15782 2148 15838 2150
rect 15862 2148 15918 2150
rect 15942 2148 15998 2150
rect 16022 2148 16078 2150
rect 16394 10512 16450 10568
rect 16946 9832 17002 9888
rect 16302 7928 16358 7984
rect 16394 7248 16450 7304
rect 3514 176 3570 232
rect 16578 2896 16634 2952
rect 16578 2624 16634 2680
rect 17590 13368 17646 13424
rect 17498 11736 17554 11792
rect 17314 9016 17370 9072
rect 17314 5772 17370 5808
rect 17590 8608 17646 8664
rect 17590 7792 17646 7848
rect 17590 6060 17592 6080
rect 17592 6060 17644 6080
rect 17644 6060 17646 6080
rect 17590 6024 17646 6060
rect 17314 5752 17316 5772
rect 17316 5752 17368 5772
rect 17368 5752 17370 5772
rect 17498 5636 17554 5672
rect 17498 5616 17500 5636
rect 17500 5616 17552 5636
rect 17552 5616 17554 5636
rect 17498 3984 17554 4040
rect 17590 3032 17646 3088
rect 17866 7384 17922 7440
rect 18050 7384 18106 7440
rect 18050 6432 18106 6488
rect 17866 5208 17922 5264
rect 17774 4800 17830 4856
rect 17866 4684 17922 4720
rect 17866 4664 17868 4684
rect 17868 4664 17920 4684
rect 17920 4664 17922 4684
rect 17314 2216 17370 2272
rect 17222 1400 17278 1456
rect 17682 2508 17738 2544
rect 17682 2488 17684 2508
rect 17684 2488 17736 2508
rect 17736 2488 17738 2508
rect 18234 8236 18236 8256
rect 18236 8236 18288 8256
rect 18288 8236 18290 8256
rect 18234 8200 18290 8236
rect 18234 6976 18290 7032
rect 18234 4392 18290 4448
rect 17866 3576 17922 3632
rect 17774 1808 17830 1864
rect 17866 992 17922 1048
rect 16486 584 16542 640
rect 18786 13232 18842 13288
rect 19430 3304 19486 3360
rect 18234 176 18290 232
<< metal3 >>
rect 0 16690 800 16720
rect 8385 16690 8451 16693
rect 0 16688 8451 16690
rect 0 16632 8390 16688
rect 8446 16632 8451 16688
rect 0 16630 8451 16632
rect 0 16600 800 16630
rect 8385 16627 8451 16630
rect 18321 16690 18387 16693
rect 19200 16690 20000 16720
rect 18321 16688 20000 16690
rect 18321 16632 18326 16688
rect 18382 16632 20000 16688
rect 18321 16630 20000 16632
rect 18321 16627 18387 16630
rect 19200 16600 20000 16630
rect 0 16282 800 16312
rect 4061 16282 4127 16285
rect 0 16280 4127 16282
rect 0 16224 4066 16280
rect 4122 16224 4127 16280
rect 0 16222 4127 16224
rect 0 16192 800 16222
rect 4061 16219 4127 16222
rect 18229 16282 18295 16285
rect 19200 16282 20000 16312
rect 18229 16280 20000 16282
rect 18229 16224 18234 16280
rect 18290 16224 20000 16280
rect 18229 16222 20000 16224
rect 18229 16219 18295 16222
rect 19200 16192 20000 16222
rect 0 15874 800 15904
rect 2773 15874 2839 15877
rect 0 15872 2839 15874
rect 0 15816 2778 15872
rect 2834 15816 2839 15872
rect 0 15814 2839 15816
rect 0 15784 800 15814
rect 2773 15811 2839 15814
rect 15285 15874 15351 15877
rect 19200 15874 20000 15904
rect 15285 15872 20000 15874
rect 15285 15816 15290 15872
rect 15346 15816 20000 15872
rect 15285 15814 20000 15816
rect 15285 15811 15351 15814
rect 19200 15784 20000 15814
rect 0 15466 800 15496
rect 3969 15466 4035 15469
rect 0 15464 4035 15466
rect 0 15408 3974 15464
rect 4030 15408 4035 15464
rect 0 15406 4035 15408
rect 0 15376 800 15406
rect 3969 15403 4035 15406
rect 15101 15466 15167 15469
rect 19200 15466 20000 15496
rect 15101 15464 20000 15466
rect 15101 15408 15106 15464
rect 15162 15408 20000 15464
rect 15101 15406 20000 15408
rect 15101 15403 15167 15406
rect 19200 15376 20000 15406
rect 0 15058 800 15088
rect 3509 15058 3575 15061
rect 0 15056 3575 15058
rect 0 15000 3514 15056
rect 3570 15000 3575 15056
rect 0 14998 3575 15000
rect 0 14968 800 14998
rect 3509 14995 3575 14998
rect 17953 15058 18019 15061
rect 19200 15058 20000 15088
rect 17953 15056 20000 15058
rect 17953 15000 17958 15056
rect 18014 15000 20000 15056
rect 17953 14998 20000 15000
rect 17953 14995 18019 14998
rect 19200 14968 20000 14998
rect 6874 14720 7194 14721
rect 0 14650 800 14680
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7194 14720
rect 6874 14655 7194 14656
rect 12805 14720 13125 14721
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 14655 13125 14656
rect 4429 14650 4495 14653
rect 0 14648 4495 14650
rect 0 14592 4434 14648
rect 4490 14592 4495 14648
rect 0 14590 4495 14592
rect 0 14560 800 14590
rect 4429 14587 4495 14590
rect 15377 14650 15443 14653
rect 19200 14650 20000 14680
rect 15377 14648 20000 14650
rect 15377 14592 15382 14648
rect 15438 14592 20000 14648
rect 15377 14590 20000 14592
rect 15377 14587 15443 14590
rect 19200 14560 20000 14590
rect 15101 14378 15167 14381
rect 15101 14376 16866 14378
rect 15101 14320 15106 14376
rect 15162 14320 16866 14376
rect 15101 14318 16866 14320
rect 15101 14315 15167 14318
rect 0 14242 800 14272
rect 3693 14242 3759 14245
rect 0 14240 3759 14242
rect 0 14184 3698 14240
rect 3754 14184 3759 14240
rect 0 14182 3759 14184
rect 16806 14242 16866 14318
rect 19200 14242 20000 14272
rect 16806 14182 20000 14242
rect 0 14152 800 14182
rect 3693 14179 3759 14182
rect 3909 14176 4229 14177
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 14111 4229 14112
rect 9840 14176 10160 14177
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14111 10160 14112
rect 15770 14176 16090 14177
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 19200 14152 20000 14182
rect 15770 14111 16090 14112
rect 0 13834 800 13864
rect 3785 13834 3851 13837
rect 19200 13834 20000 13864
rect 0 13832 3851 13834
rect 0 13776 3790 13832
rect 3846 13776 3851 13832
rect 0 13774 3851 13776
rect 0 13744 800 13774
rect 3785 13771 3851 13774
rect 15702 13774 20000 13834
rect 6874 13632 7194 13633
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7194 13632
rect 6874 13567 7194 13568
rect 12805 13632 13125 13633
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 13567 13125 13568
rect 0 13426 800 13456
rect 4061 13426 4127 13429
rect 0 13424 4127 13426
rect 0 13368 4066 13424
rect 4122 13368 4127 13424
rect 0 13366 4127 13368
rect 0 13336 800 13366
rect 4061 13363 4127 13366
rect 9397 13426 9463 13429
rect 15702 13426 15762 13774
rect 19200 13744 20000 13774
rect 17585 13426 17651 13429
rect 9397 13424 15762 13426
rect 9397 13368 9402 13424
rect 9458 13368 15762 13424
rect 9397 13366 15762 13368
rect 15886 13424 17651 13426
rect 15886 13368 17590 13424
rect 17646 13368 17651 13424
rect 15886 13366 17651 13368
rect 9397 13363 9463 13366
rect 5901 13290 5967 13293
rect 15886 13290 15946 13366
rect 17585 13363 17651 13366
rect 5901 13288 15946 13290
rect 5901 13232 5906 13288
rect 5962 13232 15946 13288
rect 5901 13230 15946 13232
rect 18781 13290 18847 13293
rect 19200 13290 20000 13320
rect 18781 13288 20000 13290
rect 18781 13232 18786 13288
rect 18842 13232 20000 13288
rect 18781 13230 20000 13232
rect 5901 13227 5967 13230
rect 18781 13227 18847 13230
rect 19200 13200 20000 13230
rect 10685 13154 10751 13157
rect 10961 13154 11027 13157
rect 14825 13154 14891 13157
rect 10685 13152 14891 13154
rect 10685 13096 10690 13152
rect 10746 13096 10966 13152
rect 11022 13096 14830 13152
rect 14886 13096 14891 13152
rect 10685 13094 14891 13096
rect 10685 13091 10751 13094
rect 10961 13091 11027 13094
rect 14825 13091 14891 13094
rect 3909 13088 4229 13089
rect 0 13018 800 13048
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 13023 4229 13024
rect 9840 13088 10160 13089
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 13023 10160 13024
rect 15770 13088 16090 13089
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15770 13023 16090 13024
rect 3509 13018 3575 13021
rect 0 13016 3575 13018
rect 0 12960 3514 13016
rect 3570 12960 3575 13016
rect 0 12958 3575 12960
rect 0 12928 800 12958
rect 3509 12955 3575 12958
rect 7465 13018 7531 13021
rect 8017 13018 8083 13021
rect 7465 13016 8083 13018
rect 7465 12960 7470 13016
rect 7526 12960 8022 13016
rect 8078 12960 8083 13016
rect 7465 12958 8083 12960
rect 7465 12955 7531 12958
rect 8017 12955 8083 12958
rect 5993 12882 6059 12885
rect 7833 12882 7899 12885
rect 5993 12880 7899 12882
rect 5993 12824 5998 12880
rect 6054 12824 7838 12880
rect 7894 12824 7899 12880
rect 5993 12822 7899 12824
rect 5993 12819 6059 12822
rect 7833 12819 7899 12822
rect 10225 12882 10291 12885
rect 16573 12882 16639 12885
rect 19200 12882 20000 12912
rect 10225 12880 16639 12882
rect 10225 12824 10230 12880
rect 10286 12824 16578 12880
rect 16634 12824 16639 12880
rect 10225 12822 16639 12824
rect 10225 12819 10291 12822
rect 16573 12819 16639 12822
rect 16806 12822 20000 12882
rect 1117 12746 1183 12749
rect 13169 12746 13235 12749
rect 1117 12744 13235 12746
rect 1117 12688 1122 12744
rect 1178 12688 13174 12744
rect 13230 12688 13235 12744
rect 1117 12686 13235 12688
rect 1117 12683 1183 12686
rect 13169 12683 13235 12686
rect 13629 12746 13695 12749
rect 14641 12746 14707 12749
rect 16806 12746 16866 12822
rect 19200 12792 20000 12822
rect 13629 12744 16866 12746
rect 13629 12688 13634 12744
rect 13690 12688 14646 12744
rect 14702 12688 16866 12744
rect 13629 12686 16866 12688
rect 13629 12683 13695 12686
rect 14641 12683 14707 12686
rect 0 12610 800 12640
rect 3969 12610 4035 12613
rect 0 12608 4035 12610
rect 0 12552 3974 12608
rect 4030 12552 4035 12608
rect 0 12550 4035 12552
rect 0 12520 800 12550
rect 3969 12547 4035 12550
rect 14917 12610 14983 12613
rect 16757 12610 16823 12613
rect 14917 12608 16823 12610
rect 14917 12552 14922 12608
rect 14978 12552 16762 12608
rect 16818 12552 16823 12608
rect 14917 12550 16823 12552
rect 14917 12547 14983 12550
rect 16757 12547 16823 12550
rect 6874 12544 7194 12545
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7194 12544
rect 6874 12479 7194 12480
rect 12805 12544 13125 12545
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 12479 13125 12480
rect 16246 12412 16252 12476
rect 16316 12474 16322 12476
rect 19200 12474 20000 12504
rect 16316 12414 20000 12474
rect 16316 12412 16322 12414
rect 19200 12384 20000 12414
rect 6361 12338 6427 12341
rect 10501 12338 10567 12341
rect 6361 12336 10567 12338
rect 6361 12280 6366 12336
rect 6422 12280 10506 12336
rect 10562 12280 10567 12336
rect 6361 12278 10567 12280
rect 6361 12275 6427 12278
rect 10501 12275 10567 12278
rect 15653 12338 15719 12341
rect 16389 12338 16455 12341
rect 15653 12336 16455 12338
rect 15653 12280 15658 12336
rect 15714 12280 16394 12336
rect 16450 12280 16455 12336
rect 15653 12278 16455 12280
rect 15653 12275 15719 12278
rect 16389 12275 16455 12278
rect 0 12202 800 12232
rect 2129 12202 2195 12205
rect 0 12200 2195 12202
rect 0 12144 2134 12200
rect 2190 12144 2195 12200
rect 0 12142 2195 12144
rect 0 12112 800 12142
rect 2129 12139 2195 12142
rect 2957 12202 3023 12205
rect 7833 12202 7899 12205
rect 2957 12200 7899 12202
rect 2957 12144 2962 12200
rect 3018 12144 7838 12200
rect 7894 12144 7899 12200
rect 2957 12142 7899 12144
rect 2957 12139 3023 12142
rect 7833 12139 7899 12142
rect 9305 12202 9371 12205
rect 16297 12202 16363 12205
rect 9305 12200 16363 12202
rect 9305 12144 9310 12200
rect 9366 12144 16302 12200
rect 16358 12144 16363 12200
rect 9305 12142 16363 12144
rect 9305 12139 9371 12142
rect 16297 12139 16363 12142
rect 5441 12066 5507 12069
rect 7005 12066 7071 12069
rect 5441 12064 7071 12066
rect 5441 12008 5446 12064
rect 5502 12008 7010 12064
rect 7066 12008 7071 12064
rect 5441 12006 7071 12008
rect 5441 12003 5507 12006
rect 7005 12003 7071 12006
rect 16297 12066 16363 12069
rect 19200 12066 20000 12096
rect 16297 12064 20000 12066
rect 16297 12008 16302 12064
rect 16358 12008 20000 12064
rect 16297 12006 20000 12008
rect 16297 12003 16363 12006
rect 3909 12000 4229 12001
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 11935 4229 11936
rect 9840 12000 10160 12001
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 11935 10160 11936
rect 15770 12000 16090 12001
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 19200 11976 20000 12006
rect 15770 11935 16090 11936
rect 15377 11932 15443 11933
rect 15326 11930 15332 11932
rect 15286 11870 15332 11930
rect 15396 11928 15443 11932
rect 15438 11872 15443 11928
rect 15326 11868 15332 11870
rect 15396 11868 15443 11872
rect 15377 11867 15443 11868
rect 0 11794 800 11824
rect 3877 11794 3943 11797
rect 0 11792 3943 11794
rect 0 11736 3882 11792
rect 3938 11736 3943 11792
rect 0 11734 3943 11736
rect 0 11704 800 11734
rect 3877 11731 3943 11734
rect 10317 11794 10383 11797
rect 17493 11794 17559 11797
rect 10317 11792 17559 11794
rect 10317 11736 10322 11792
rect 10378 11736 17498 11792
rect 17554 11736 17559 11792
rect 10317 11734 17559 11736
rect 10317 11731 10383 11734
rect 17493 11731 17559 11734
rect 2681 11658 2747 11661
rect 7833 11658 7899 11661
rect 2681 11656 7899 11658
rect 2681 11600 2686 11656
rect 2742 11600 7838 11656
rect 7894 11600 7899 11656
rect 2681 11598 7899 11600
rect 2681 11595 2747 11598
rect 7833 11595 7899 11598
rect 11421 11658 11487 11661
rect 12801 11658 12867 11661
rect 11421 11656 12867 11658
rect 11421 11600 11426 11656
rect 11482 11600 12806 11656
rect 12862 11600 12867 11656
rect 11421 11598 12867 11600
rect 11421 11595 11487 11598
rect 12801 11595 12867 11598
rect 14549 11658 14615 11661
rect 19200 11658 20000 11688
rect 14549 11656 20000 11658
rect 14549 11600 14554 11656
rect 14610 11600 20000 11656
rect 14549 11598 20000 11600
rect 14549 11595 14615 11598
rect 19200 11568 20000 11598
rect 6874 11456 7194 11457
rect 0 11386 800 11416
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7194 11456
rect 6874 11391 7194 11392
rect 12805 11456 13125 11457
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 11391 13125 11392
rect 3785 11386 3851 11389
rect 0 11384 3851 11386
rect 0 11328 3790 11384
rect 3846 11328 3851 11384
rect 0 11326 3851 11328
rect 0 11296 800 11326
rect 3785 11323 3851 11326
rect 8109 11386 8175 11389
rect 9857 11386 9923 11389
rect 8109 11384 9923 11386
rect 8109 11328 8114 11384
rect 8170 11328 9862 11384
rect 9918 11328 9923 11384
rect 8109 11326 9923 11328
rect 8109 11323 8175 11326
rect 9857 11323 9923 11326
rect 1669 11250 1735 11253
rect 7649 11250 7715 11253
rect 9029 11250 9095 11253
rect 1669 11248 9095 11250
rect 1669 11192 1674 11248
rect 1730 11192 7654 11248
rect 7710 11192 9034 11248
rect 9090 11192 9095 11248
rect 1669 11190 9095 11192
rect 1669 11187 1735 11190
rect 7649 11187 7715 11190
rect 9029 11187 9095 11190
rect 10961 11250 11027 11253
rect 13813 11250 13879 11253
rect 10961 11248 13879 11250
rect 10961 11192 10966 11248
rect 11022 11192 13818 11248
rect 13874 11192 13879 11248
rect 10961 11190 13879 11192
rect 10961 11187 11027 11190
rect 13813 11187 13879 11190
rect 15101 11250 15167 11253
rect 19200 11250 20000 11280
rect 15101 11248 20000 11250
rect 15101 11192 15106 11248
rect 15162 11192 20000 11248
rect 15101 11190 20000 11192
rect 15101 11187 15167 11190
rect 19200 11160 20000 11190
rect 6913 11114 6979 11117
rect 9121 11114 9187 11117
rect 6913 11112 9187 11114
rect 6913 11056 6918 11112
rect 6974 11056 9126 11112
rect 9182 11056 9187 11112
rect 6913 11054 9187 11056
rect 6913 11051 6979 11054
rect 0 10978 800 11008
rect 7468 10981 7528 11054
rect 9121 11051 9187 11054
rect 12341 11114 12407 11117
rect 13537 11114 13603 11117
rect 12341 11112 13603 11114
rect 12341 11056 12346 11112
rect 12402 11056 13542 11112
rect 13598 11056 13603 11112
rect 12341 11054 13603 11056
rect 12341 11051 12407 11054
rect 13537 11051 13603 11054
rect 3509 10978 3575 10981
rect 0 10976 3575 10978
rect 0 10920 3514 10976
rect 3570 10920 3575 10976
rect 0 10918 3575 10920
rect 0 10888 800 10918
rect 3509 10915 3575 10918
rect 7465 10976 7531 10981
rect 7465 10920 7470 10976
rect 7526 10920 7531 10976
rect 7465 10915 7531 10920
rect 3909 10912 4229 10913
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 10847 4229 10848
rect 9840 10912 10160 10913
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10847 10160 10848
rect 15770 10912 16090 10913
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 10847 16090 10848
rect 16481 10842 16547 10845
rect 19200 10842 20000 10872
rect 16481 10840 20000 10842
rect 16481 10784 16486 10840
rect 16542 10784 20000 10840
rect 16481 10782 20000 10784
rect 16481 10779 16547 10782
rect 19200 10752 20000 10782
rect 4061 10706 4127 10709
rect 14365 10706 14431 10709
rect 4061 10704 14431 10706
rect 4061 10648 4066 10704
rect 4122 10648 14370 10704
rect 14426 10648 14431 10704
rect 4061 10646 14431 10648
rect 4061 10643 4127 10646
rect 14365 10643 14431 10646
rect 0 10570 800 10600
rect 3601 10570 3667 10573
rect 0 10568 3667 10570
rect 0 10512 3606 10568
rect 3662 10512 3667 10568
rect 0 10510 3667 10512
rect 0 10480 800 10510
rect 3601 10507 3667 10510
rect 6821 10570 6887 10573
rect 9213 10570 9279 10573
rect 6821 10568 9279 10570
rect 6821 10512 6826 10568
rect 6882 10512 9218 10568
rect 9274 10512 9279 10568
rect 6821 10510 9279 10512
rect 6821 10507 6887 10510
rect 9213 10507 9279 10510
rect 16246 10508 16252 10572
rect 16316 10570 16322 10572
rect 16389 10570 16455 10573
rect 16316 10568 16455 10570
rect 16316 10512 16394 10568
rect 16450 10512 16455 10568
rect 16316 10510 16455 10512
rect 16316 10508 16322 10510
rect 16389 10507 16455 10510
rect 13905 10434 13971 10437
rect 15377 10434 15443 10437
rect 19200 10434 20000 10464
rect 13905 10432 20000 10434
rect 13905 10376 13910 10432
rect 13966 10376 15382 10432
rect 15438 10376 20000 10432
rect 13905 10374 20000 10376
rect 13905 10371 13971 10374
rect 15377 10371 15443 10374
rect 6874 10368 7194 10369
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7194 10368
rect 6874 10303 7194 10304
rect 12805 10368 13125 10369
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 19200 10344 20000 10374
rect 12805 10303 13125 10304
rect 0 10162 800 10192
rect 4889 10162 4955 10165
rect 0 10160 4955 10162
rect 0 10104 4894 10160
rect 4950 10104 4955 10160
rect 0 10102 4955 10104
rect 0 10072 800 10102
rect 4889 10099 4955 10102
rect 5349 10162 5415 10165
rect 8109 10162 8175 10165
rect 5349 10160 8175 10162
rect 5349 10104 5354 10160
rect 5410 10104 8114 10160
rect 8170 10104 8175 10160
rect 5349 10102 8175 10104
rect 5349 10099 5415 10102
rect 8109 10099 8175 10102
rect 4981 10026 5047 10029
rect 10501 10026 10567 10029
rect 4981 10024 10567 10026
rect 4981 9968 4986 10024
rect 5042 9968 10506 10024
rect 10562 9968 10567 10024
rect 4981 9966 10567 9968
rect 4981 9963 5047 9966
rect 10501 9963 10567 9966
rect 12341 10026 12407 10029
rect 12341 10024 17004 10026
rect 12341 9968 12346 10024
rect 12402 9968 17004 10024
rect 12341 9966 17004 9968
rect 12341 9963 12407 9966
rect 16944 9893 17004 9966
rect 4705 9890 4771 9893
rect 6085 9890 6151 9893
rect 4705 9888 6151 9890
rect 4705 9832 4710 9888
rect 4766 9832 6090 9888
rect 6146 9832 6151 9888
rect 4705 9830 6151 9832
rect 4705 9827 4771 9830
rect 6085 9827 6151 9830
rect 16941 9890 17007 9893
rect 19200 9890 20000 9920
rect 16941 9888 20000 9890
rect 16941 9832 16946 9888
rect 17002 9832 20000 9888
rect 16941 9830 20000 9832
rect 16941 9827 17007 9830
rect 3909 9824 4229 9825
rect 0 9754 800 9784
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 9759 4229 9760
rect 9840 9824 10160 9825
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 9759 10160 9760
rect 15770 9824 16090 9825
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 19200 9800 20000 9830
rect 15770 9759 16090 9760
rect 2865 9754 2931 9757
rect 0 9752 2931 9754
rect 0 9696 2870 9752
rect 2926 9696 2931 9752
rect 0 9694 2931 9696
rect 0 9664 800 9694
rect 2865 9691 2931 9694
rect 5901 9482 5967 9485
rect 8661 9482 8727 9485
rect 5901 9480 8727 9482
rect 5901 9424 5906 9480
rect 5962 9424 8666 9480
rect 8722 9424 8727 9480
rect 5901 9422 8727 9424
rect 5901 9419 5967 9422
rect 8661 9419 8727 9422
rect 13629 9482 13695 9485
rect 19200 9482 20000 9512
rect 13629 9480 20000 9482
rect 13629 9424 13634 9480
rect 13690 9424 20000 9480
rect 13629 9422 20000 9424
rect 13629 9419 13695 9422
rect 19200 9392 20000 9422
rect 0 9346 800 9376
rect 4061 9346 4127 9349
rect 0 9344 4127 9346
rect 0 9288 4066 9344
rect 4122 9288 4127 9344
rect 0 9286 4127 9288
rect 0 9256 800 9286
rect 4061 9283 4127 9286
rect 6874 9280 7194 9281
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7194 9280
rect 6874 9215 7194 9216
rect 12805 9280 13125 9281
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 9215 13125 9216
rect 5073 9074 5139 9077
rect 13537 9074 13603 9077
rect 5073 9072 13603 9074
rect 5073 9016 5078 9072
rect 5134 9016 13542 9072
rect 13598 9016 13603 9072
rect 5073 9014 13603 9016
rect 5073 9011 5139 9014
rect 13537 9011 13603 9014
rect 17309 9074 17375 9077
rect 19200 9074 20000 9104
rect 17309 9072 20000 9074
rect 17309 9016 17314 9072
rect 17370 9016 20000 9072
rect 17309 9014 20000 9016
rect 17309 9011 17375 9014
rect 19200 8984 20000 9014
rect 0 8938 800 8968
rect 2497 8938 2563 8941
rect 0 8936 2563 8938
rect 0 8880 2502 8936
rect 2558 8880 2563 8936
rect 0 8878 2563 8880
rect 0 8848 800 8878
rect 2497 8875 2563 8878
rect 12341 8938 12407 8941
rect 14089 8938 14155 8941
rect 12341 8936 14155 8938
rect 12341 8880 12346 8936
rect 12402 8880 14094 8936
rect 14150 8880 14155 8936
rect 12341 8878 14155 8880
rect 12341 8875 12407 8878
rect 14089 8875 14155 8878
rect 5625 8802 5691 8805
rect 5901 8802 5967 8805
rect 5625 8800 5967 8802
rect 5625 8744 5630 8800
rect 5686 8744 5906 8800
rect 5962 8744 5967 8800
rect 5625 8742 5967 8744
rect 5625 8739 5691 8742
rect 5901 8739 5967 8742
rect 3909 8736 4229 8737
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 8671 4229 8672
rect 9840 8736 10160 8737
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 8671 10160 8672
rect 15770 8736 16090 8737
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 15770 8671 16090 8672
rect 7465 8666 7531 8669
rect 17585 8666 17651 8669
rect 19200 8666 20000 8696
rect 4524 8664 7531 8666
rect 4524 8608 7470 8664
rect 7526 8608 7531 8664
rect 4524 8606 7531 8608
rect 4245 8532 4311 8533
rect 4245 8528 4292 8532
rect 4356 8530 4362 8532
rect 4524 8530 4584 8606
rect 7465 8603 7531 8606
rect 16254 8664 20000 8666
rect 16254 8608 17590 8664
rect 17646 8608 20000 8664
rect 16254 8606 20000 8608
rect 4245 8472 4250 8528
rect 4245 8468 4292 8472
rect 4356 8470 4584 8530
rect 6177 8530 6243 8533
rect 6545 8530 6611 8533
rect 6177 8528 6611 8530
rect 6177 8472 6182 8528
rect 6238 8472 6550 8528
rect 6606 8472 6611 8528
rect 6177 8470 6611 8472
rect 4356 8468 4362 8470
rect 4245 8467 4311 8468
rect 6177 8467 6243 8470
rect 6545 8467 6611 8470
rect 14733 8530 14799 8533
rect 16254 8530 16314 8606
rect 17585 8603 17651 8606
rect 19200 8576 20000 8606
rect 14733 8528 16314 8530
rect 14733 8472 14738 8528
rect 14794 8472 16314 8528
rect 14733 8470 16314 8472
rect 14733 8467 14799 8470
rect 0 8394 800 8424
rect 2957 8394 3023 8397
rect 0 8392 3023 8394
rect 0 8336 2962 8392
rect 3018 8336 3023 8392
rect 0 8334 3023 8336
rect 0 8304 800 8334
rect 2957 8331 3023 8334
rect 6453 8394 6519 8397
rect 7557 8394 7623 8397
rect 6453 8392 7623 8394
rect 6453 8336 6458 8392
rect 6514 8336 7562 8392
rect 7618 8336 7623 8392
rect 6453 8334 7623 8336
rect 6453 8331 6519 8334
rect 7557 8331 7623 8334
rect 10961 8394 11027 8397
rect 14457 8394 14523 8397
rect 10961 8392 14523 8394
rect 10961 8336 10966 8392
rect 11022 8336 14462 8392
rect 14518 8336 14523 8392
rect 10961 8334 14523 8336
rect 10961 8331 11027 8334
rect 14457 8331 14523 8334
rect 18229 8258 18295 8261
rect 19200 8258 20000 8288
rect 18229 8256 20000 8258
rect 18229 8200 18234 8256
rect 18290 8200 20000 8256
rect 18229 8198 20000 8200
rect 18229 8195 18295 8198
rect 6874 8192 7194 8193
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7194 8192
rect 6874 8127 7194 8128
rect 12805 8192 13125 8193
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 19200 8168 20000 8198
rect 12805 8127 13125 8128
rect 5993 8122 6059 8125
rect 6453 8122 6519 8125
rect 5993 8120 6519 8122
rect 5993 8064 5998 8120
rect 6054 8064 6458 8120
rect 6514 8064 6519 8120
rect 5993 8062 6519 8064
rect 5993 8059 6059 8062
rect 6453 8059 6519 8062
rect 11513 8122 11579 8125
rect 11513 8120 12634 8122
rect 11513 8064 11518 8120
rect 11574 8064 12634 8120
rect 11513 8062 12634 8064
rect 11513 8059 11579 8062
rect 0 7986 800 8016
rect 1485 7986 1551 7989
rect 0 7984 1551 7986
rect 0 7928 1490 7984
rect 1546 7928 1551 7984
rect 0 7926 1551 7928
rect 0 7896 800 7926
rect 1485 7923 1551 7926
rect 4061 7986 4127 7989
rect 7557 7986 7623 7989
rect 4061 7984 7623 7986
rect 4061 7928 4066 7984
rect 4122 7928 7562 7984
rect 7618 7928 7623 7984
rect 4061 7926 7623 7928
rect 12574 7986 12634 8062
rect 16297 7986 16363 7989
rect 12574 7984 16363 7986
rect 12574 7928 16302 7984
rect 16358 7928 16363 7984
rect 12574 7926 16363 7928
rect 4061 7923 4127 7926
rect 7557 7923 7623 7926
rect 16297 7923 16363 7926
rect 8385 7850 8451 7853
rect 9397 7850 9463 7853
rect 11605 7850 11671 7853
rect 8385 7848 11671 7850
rect 8385 7792 8390 7848
rect 8446 7792 9402 7848
rect 9458 7792 11610 7848
rect 11666 7792 11671 7848
rect 8385 7790 11671 7792
rect 8385 7787 8451 7790
rect 9397 7787 9463 7790
rect 11605 7787 11671 7790
rect 17585 7850 17651 7853
rect 19200 7850 20000 7880
rect 17585 7848 20000 7850
rect 17585 7792 17590 7848
rect 17646 7792 20000 7848
rect 17585 7790 20000 7792
rect 17585 7787 17651 7790
rect 19200 7760 20000 7790
rect 5257 7714 5323 7717
rect 7741 7714 7807 7717
rect 5257 7712 7807 7714
rect 5257 7656 5262 7712
rect 5318 7656 7746 7712
rect 7802 7656 7807 7712
rect 5257 7654 7807 7656
rect 5257 7651 5323 7654
rect 7741 7651 7807 7654
rect 3909 7648 4229 7649
rect 0 7578 800 7608
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 7583 4229 7584
rect 9840 7648 10160 7649
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 7583 10160 7584
rect 15770 7648 16090 7649
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 7583 16090 7584
rect 1393 7578 1459 7581
rect 0 7576 1459 7578
rect 0 7520 1398 7576
rect 1454 7520 1459 7576
rect 0 7518 1459 7520
rect 0 7488 800 7518
rect 1393 7515 1459 7518
rect 13077 7578 13143 7581
rect 13302 7578 13308 7580
rect 13077 7576 13308 7578
rect 13077 7520 13082 7576
rect 13138 7520 13308 7576
rect 13077 7518 13308 7520
rect 13077 7515 13143 7518
rect 13302 7516 13308 7518
rect 13372 7578 13378 7580
rect 14549 7578 14615 7581
rect 13372 7576 14615 7578
rect 13372 7520 14554 7576
rect 14610 7520 14615 7576
rect 13372 7518 14615 7520
rect 13372 7516 13378 7518
rect 14549 7515 14615 7518
rect 4429 7442 4495 7445
rect 8937 7442 9003 7445
rect 4429 7440 9003 7442
rect 4429 7384 4434 7440
rect 4490 7384 8942 7440
rect 8998 7384 9003 7440
rect 4429 7382 9003 7384
rect 4429 7379 4495 7382
rect 6180 7309 6240 7382
rect 8937 7379 9003 7382
rect 11421 7442 11487 7445
rect 17861 7442 17927 7445
rect 11421 7440 17927 7442
rect 11421 7384 11426 7440
rect 11482 7384 17866 7440
rect 17922 7384 17927 7440
rect 11421 7382 17927 7384
rect 11421 7379 11487 7382
rect 17861 7379 17927 7382
rect 18045 7442 18111 7445
rect 19200 7442 20000 7472
rect 18045 7440 20000 7442
rect 18045 7384 18050 7440
rect 18106 7384 20000 7440
rect 18045 7382 20000 7384
rect 18045 7379 18111 7382
rect 19200 7352 20000 7382
rect 6177 7304 6243 7309
rect 6177 7248 6182 7304
rect 6238 7248 6243 7304
rect 6177 7243 6243 7248
rect 7557 7306 7623 7309
rect 8937 7306 9003 7309
rect 7557 7304 9003 7306
rect 7557 7248 7562 7304
rect 7618 7248 8942 7304
rect 8998 7248 9003 7304
rect 7557 7246 9003 7248
rect 7557 7243 7623 7246
rect 8937 7243 9003 7246
rect 10777 7306 10843 7309
rect 16389 7306 16455 7309
rect 10777 7304 16455 7306
rect 10777 7248 10782 7304
rect 10838 7248 16394 7304
rect 16450 7248 16455 7304
rect 10777 7246 16455 7248
rect 10777 7243 10843 7246
rect 16389 7243 16455 7246
rect 0 7170 800 7200
rect 5349 7170 5415 7173
rect 0 7168 5415 7170
rect 0 7112 5354 7168
rect 5410 7112 5415 7168
rect 0 7110 5415 7112
rect 0 7080 800 7110
rect 5349 7107 5415 7110
rect 6874 7104 7194 7105
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7194 7104
rect 6874 7039 7194 7040
rect 12805 7104 13125 7105
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 7039 13125 7040
rect 1853 7034 1919 7037
rect 5533 7034 5599 7037
rect 1853 7032 5599 7034
rect 1853 6976 1858 7032
rect 1914 6976 5538 7032
rect 5594 6976 5599 7032
rect 1853 6974 5599 6976
rect 1853 6971 1919 6974
rect 5533 6971 5599 6974
rect 10133 7034 10199 7037
rect 12249 7034 12315 7037
rect 12382 7034 12388 7036
rect 10133 7032 12388 7034
rect 10133 6976 10138 7032
rect 10194 6976 12254 7032
rect 12310 6976 12388 7032
rect 10133 6974 12388 6976
rect 10133 6971 10199 6974
rect 12249 6971 12315 6974
rect 12382 6972 12388 6974
rect 12452 6972 12458 7036
rect 18229 7034 18295 7037
rect 19200 7034 20000 7064
rect 18229 7032 20000 7034
rect 18229 6976 18234 7032
rect 18290 6976 20000 7032
rect 18229 6974 20000 6976
rect 18229 6971 18295 6974
rect 19200 6944 20000 6974
rect 2589 6898 2655 6901
rect 2773 6898 2839 6901
rect 2589 6896 2839 6898
rect 2589 6840 2594 6896
rect 2650 6840 2778 6896
rect 2834 6840 2839 6896
rect 2589 6838 2839 6840
rect 2589 6835 2655 6838
rect 2773 6835 2839 6838
rect 12341 6898 12407 6901
rect 12525 6898 12591 6901
rect 12341 6896 12591 6898
rect 12341 6840 12346 6896
rect 12402 6840 12530 6896
rect 12586 6840 12591 6896
rect 12341 6838 12591 6840
rect 12341 6835 12407 6838
rect 12525 6835 12591 6838
rect 12709 6898 12775 6901
rect 13445 6898 13511 6901
rect 12709 6896 13511 6898
rect 12709 6840 12714 6896
rect 12770 6840 13450 6896
rect 13506 6840 13511 6896
rect 12709 6838 13511 6840
rect 12709 6835 12775 6838
rect 13445 6835 13511 6838
rect 0 6762 800 6792
rect 3601 6762 3667 6765
rect 0 6760 3667 6762
rect 0 6704 3606 6760
rect 3662 6704 3667 6760
rect 0 6702 3667 6704
rect 0 6672 800 6702
rect 3601 6699 3667 6702
rect 12249 6762 12315 6765
rect 13997 6762 14063 6765
rect 12249 6760 14063 6762
rect 12249 6704 12254 6760
rect 12310 6704 14002 6760
rect 14058 6704 14063 6760
rect 12249 6702 14063 6704
rect 12249 6699 12315 6702
rect 13997 6699 14063 6702
rect 6913 6626 6979 6629
rect 7557 6626 7623 6629
rect 6913 6624 7623 6626
rect 6913 6568 6918 6624
rect 6974 6568 7562 6624
rect 7618 6568 7623 6624
rect 6913 6566 7623 6568
rect 6913 6563 6979 6566
rect 7557 6563 7623 6566
rect 12985 6626 13051 6629
rect 14825 6626 14891 6629
rect 12985 6624 14891 6626
rect 12985 6568 12990 6624
rect 13046 6568 14830 6624
rect 14886 6568 14891 6624
rect 12985 6566 14891 6568
rect 12985 6563 13051 6566
rect 14825 6563 14891 6566
rect 3909 6560 4229 6561
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 6495 4229 6496
rect 9840 6560 10160 6561
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6495 10160 6496
rect 15770 6560 16090 6561
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 15770 6495 16090 6496
rect 6913 6490 6979 6493
rect 8017 6490 8083 6493
rect 6913 6488 8083 6490
rect 6913 6432 6918 6488
rect 6974 6432 8022 6488
rect 8078 6432 8083 6488
rect 6913 6430 8083 6432
rect 6913 6427 6979 6430
rect 8017 6427 8083 6430
rect 11329 6490 11395 6493
rect 14089 6490 14155 6493
rect 11329 6488 14155 6490
rect 11329 6432 11334 6488
rect 11390 6432 14094 6488
rect 14150 6432 14155 6488
rect 11329 6430 14155 6432
rect 11329 6427 11395 6430
rect 14089 6427 14155 6430
rect 18045 6490 18111 6493
rect 19200 6490 20000 6520
rect 18045 6488 20000 6490
rect 18045 6432 18050 6488
rect 18106 6432 20000 6488
rect 18045 6430 20000 6432
rect 18045 6427 18111 6430
rect 19200 6400 20000 6430
rect 0 6354 800 6384
rect 3049 6354 3115 6357
rect 0 6352 3115 6354
rect 0 6296 3054 6352
rect 3110 6296 3115 6352
rect 0 6294 3115 6296
rect 0 6264 800 6294
rect 3049 6291 3115 6294
rect 12893 6354 12959 6357
rect 13813 6354 13879 6357
rect 12893 6352 13879 6354
rect 12893 6296 12898 6352
rect 12954 6296 13818 6352
rect 13874 6296 13879 6352
rect 12893 6294 13879 6296
rect 12893 6291 12959 6294
rect 13813 6291 13879 6294
rect 10685 6218 10751 6221
rect 13445 6218 13511 6221
rect 10685 6216 13511 6218
rect 10685 6160 10690 6216
rect 10746 6160 13450 6216
rect 13506 6160 13511 6216
rect 10685 6158 13511 6160
rect 10685 6155 10751 6158
rect 13445 6155 13511 6158
rect 17585 6082 17651 6085
rect 19200 6082 20000 6112
rect 17585 6080 20000 6082
rect 17585 6024 17590 6080
rect 17646 6024 20000 6080
rect 17585 6022 20000 6024
rect 17585 6019 17651 6022
rect 6874 6016 7194 6017
rect 0 5946 800 5976
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7194 6016
rect 6874 5951 7194 5952
rect 12805 6016 13125 6017
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 19200 5992 20000 6022
rect 12805 5951 13125 5952
rect 3969 5946 4035 5949
rect 0 5944 4035 5946
rect 0 5888 3974 5944
rect 4030 5888 4035 5944
rect 0 5886 4035 5888
rect 0 5856 800 5886
rect 3969 5883 4035 5886
rect 7281 5810 7347 5813
rect 7557 5810 7623 5813
rect 7281 5808 7623 5810
rect 7281 5752 7286 5808
rect 7342 5752 7562 5808
rect 7618 5752 7623 5808
rect 7281 5750 7623 5752
rect 7281 5747 7347 5750
rect 7557 5747 7623 5750
rect 11789 5810 11855 5813
rect 17309 5810 17375 5813
rect 11789 5808 17375 5810
rect 11789 5752 11794 5808
rect 11850 5752 17314 5808
rect 17370 5752 17375 5808
rect 11789 5750 17375 5752
rect 11789 5747 11855 5750
rect 17309 5747 17375 5750
rect 4613 5674 4679 5677
rect 7189 5674 7255 5677
rect 4613 5672 7255 5674
rect 4613 5616 4618 5672
rect 4674 5616 7194 5672
rect 7250 5616 7255 5672
rect 4613 5614 7255 5616
rect 4613 5611 4679 5614
rect 7189 5611 7255 5614
rect 10409 5674 10475 5677
rect 15745 5674 15811 5677
rect 10409 5672 15811 5674
rect 10409 5616 10414 5672
rect 10470 5616 15750 5672
rect 15806 5616 15811 5672
rect 10409 5614 15811 5616
rect 10409 5611 10475 5614
rect 15745 5611 15811 5614
rect 17493 5674 17559 5677
rect 19200 5674 20000 5704
rect 17493 5672 20000 5674
rect 17493 5616 17498 5672
rect 17554 5616 20000 5672
rect 17493 5614 20000 5616
rect 17493 5611 17559 5614
rect 19200 5584 20000 5614
rect 0 5538 800 5568
rect 3509 5538 3575 5541
rect 0 5536 3575 5538
rect 0 5480 3514 5536
rect 3570 5480 3575 5536
rect 0 5478 3575 5480
rect 0 5448 800 5478
rect 3509 5475 3575 5478
rect 5809 5538 5875 5541
rect 7741 5538 7807 5541
rect 5809 5536 7807 5538
rect 5809 5480 5814 5536
rect 5870 5480 7746 5536
rect 7802 5480 7807 5536
rect 5809 5478 7807 5480
rect 5809 5475 5875 5478
rect 7741 5475 7807 5478
rect 14641 5538 14707 5541
rect 15326 5538 15332 5540
rect 14641 5536 15332 5538
rect 14641 5480 14646 5536
rect 14702 5480 15332 5536
rect 14641 5478 15332 5480
rect 14641 5475 14707 5478
rect 15326 5476 15332 5478
rect 15396 5476 15402 5540
rect 3909 5472 4229 5473
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 5407 4229 5408
rect 9840 5472 10160 5473
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 5407 10160 5408
rect 15770 5472 16090 5473
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15770 5407 16090 5408
rect 4153 5266 4219 5269
rect 6453 5266 6519 5269
rect 4153 5264 6519 5266
rect 4153 5208 4158 5264
rect 4214 5208 6458 5264
rect 6514 5208 6519 5264
rect 4153 5206 6519 5208
rect 4153 5203 4219 5206
rect 6453 5203 6519 5206
rect 6913 5266 6979 5269
rect 8661 5266 8727 5269
rect 6913 5264 8727 5266
rect 6913 5208 6918 5264
rect 6974 5208 8666 5264
rect 8722 5208 8727 5264
rect 6913 5206 8727 5208
rect 6913 5203 6979 5206
rect 8661 5203 8727 5206
rect 12382 5204 12388 5268
rect 12452 5266 12458 5268
rect 15009 5266 15075 5269
rect 15745 5266 15811 5269
rect 12452 5264 15811 5266
rect 12452 5208 15014 5264
rect 15070 5208 15750 5264
rect 15806 5208 15811 5264
rect 12452 5206 15811 5208
rect 12452 5204 12458 5206
rect 15009 5203 15075 5206
rect 15745 5203 15811 5206
rect 17861 5266 17927 5269
rect 19200 5266 20000 5296
rect 17861 5264 20000 5266
rect 17861 5208 17866 5264
rect 17922 5208 20000 5264
rect 17861 5206 20000 5208
rect 17861 5203 17927 5206
rect 19200 5176 20000 5206
rect 0 5130 800 5160
rect 3417 5130 3483 5133
rect 0 5128 3483 5130
rect 0 5072 3422 5128
rect 3478 5072 3483 5128
rect 0 5070 3483 5072
rect 0 5040 800 5070
rect 3417 5067 3483 5070
rect 6269 5130 6335 5133
rect 11237 5130 11303 5133
rect 11421 5130 11487 5133
rect 16021 5130 16087 5133
rect 6269 5128 11162 5130
rect 6269 5072 6274 5128
rect 6330 5072 11162 5128
rect 6269 5070 11162 5072
rect 6269 5067 6335 5070
rect 11102 4994 11162 5070
rect 11237 5128 16087 5130
rect 11237 5072 11242 5128
rect 11298 5072 11426 5128
rect 11482 5072 16026 5128
rect 16082 5072 16087 5128
rect 11237 5070 16087 5072
rect 11237 5067 11303 5070
rect 11421 5067 11487 5070
rect 16021 5067 16087 5070
rect 11102 4934 11530 4994
rect 6874 4928 7194 4929
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7194 4928
rect 6874 4863 7194 4864
rect 0 4722 800 4752
rect 3325 4722 3391 4725
rect 0 4720 3391 4722
rect 0 4664 3330 4720
rect 3386 4664 3391 4720
rect 0 4662 3391 4664
rect 0 4632 800 4662
rect 3325 4659 3391 4662
rect 4521 4722 4587 4725
rect 11237 4722 11303 4725
rect 4521 4720 11303 4722
rect 4521 4664 4526 4720
rect 4582 4664 11242 4720
rect 11298 4664 11303 4720
rect 4521 4662 11303 4664
rect 11470 4722 11530 4934
rect 12805 4928 13125 4929
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 4863 13125 4864
rect 17769 4858 17835 4861
rect 19200 4858 20000 4888
rect 17769 4856 20000 4858
rect 17769 4800 17774 4856
rect 17830 4800 20000 4856
rect 17769 4798 20000 4800
rect 17769 4795 17835 4798
rect 19200 4768 20000 4798
rect 17861 4722 17927 4725
rect 11470 4720 17927 4722
rect 11470 4664 17866 4720
rect 17922 4664 17927 4720
rect 11470 4662 17927 4664
rect 4521 4659 4587 4662
rect 11237 4659 11303 4662
rect 17861 4659 17927 4662
rect 5625 4586 5691 4589
rect 15653 4586 15719 4589
rect 5625 4584 15719 4586
rect 5625 4528 5630 4584
rect 5686 4528 15658 4584
rect 15714 4528 15719 4584
rect 5625 4526 15719 4528
rect 5625 4523 5691 4526
rect 15653 4523 15719 4526
rect 18229 4450 18295 4453
rect 19200 4450 20000 4480
rect 18229 4448 20000 4450
rect 18229 4392 18234 4448
rect 18290 4392 20000 4448
rect 18229 4390 20000 4392
rect 18229 4387 18295 4390
rect 3909 4384 4229 4385
rect 0 4314 800 4344
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 4319 4229 4320
rect 9840 4384 10160 4385
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 4319 10160 4320
rect 15770 4384 16090 4385
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 19200 4360 20000 4390
rect 15770 4319 16090 4320
rect 3693 4314 3759 4317
rect 0 4312 3759 4314
rect 0 4256 3698 4312
rect 3754 4256 3759 4312
rect 0 4254 3759 4256
rect 0 4224 800 4254
rect 3693 4251 3759 4254
rect 7189 4178 7255 4181
rect 14641 4178 14707 4181
rect 7189 4176 14707 4178
rect 7189 4120 7194 4176
rect 7250 4120 14646 4176
rect 14702 4120 14707 4176
rect 7189 4118 14707 4120
rect 7189 4115 7255 4118
rect 14641 4115 14707 4118
rect 8201 4042 8267 4045
rect 11053 4042 11119 4045
rect 8201 4040 11119 4042
rect 8201 3984 8206 4040
rect 8262 3984 11058 4040
rect 11114 3984 11119 4040
rect 8201 3982 11119 3984
rect 8201 3979 8267 3982
rect 11053 3979 11119 3982
rect 13445 4042 13511 4045
rect 15377 4042 15443 4045
rect 13445 4040 15443 4042
rect 13445 3984 13450 4040
rect 13506 3984 15382 4040
rect 15438 3984 15443 4040
rect 13445 3982 15443 3984
rect 13445 3979 13511 3982
rect 15377 3979 15443 3982
rect 17493 4042 17559 4045
rect 19200 4042 20000 4072
rect 17493 4040 20000 4042
rect 17493 3984 17498 4040
rect 17554 3984 20000 4040
rect 17493 3982 20000 3984
rect 17493 3979 17559 3982
rect 19200 3952 20000 3982
rect 0 3906 800 3936
rect 4061 3906 4127 3909
rect 0 3904 4127 3906
rect 0 3848 4066 3904
rect 4122 3848 4127 3904
rect 0 3846 4127 3848
rect 0 3816 800 3846
rect 4061 3843 4127 3846
rect 6874 3840 7194 3841
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7194 3840
rect 6874 3775 7194 3776
rect 12805 3840 13125 3841
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 3775 13125 3776
rect 11881 3634 11947 3637
rect 14089 3634 14155 3637
rect 11881 3632 14155 3634
rect 11881 3576 11886 3632
rect 11942 3576 14094 3632
rect 14150 3576 14155 3632
rect 11881 3574 14155 3576
rect 11881 3571 11947 3574
rect 14089 3571 14155 3574
rect 17861 3634 17927 3637
rect 19200 3634 20000 3664
rect 17861 3632 20000 3634
rect 17861 3576 17866 3632
rect 17922 3576 20000 3632
rect 17861 3574 20000 3576
rect 17861 3571 17927 3574
rect 19200 3544 20000 3574
rect 0 3498 800 3528
rect 2497 3498 2563 3501
rect 0 3496 2563 3498
rect 0 3440 2502 3496
rect 2558 3440 2563 3496
rect 0 3438 2563 3440
rect 0 3408 800 3438
rect 2497 3435 2563 3438
rect 5717 3498 5783 3501
rect 5717 3496 16314 3498
rect 5717 3440 5722 3496
rect 5778 3440 16314 3496
rect 5717 3438 16314 3440
rect 5717 3435 5783 3438
rect 16254 3362 16314 3438
rect 19425 3362 19491 3365
rect 16254 3360 19491 3362
rect 16254 3304 19430 3360
rect 19486 3304 19491 3360
rect 16254 3302 19491 3304
rect 19425 3299 19491 3302
rect 3909 3296 4229 3297
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 3231 4229 3232
rect 9840 3296 10160 3297
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 3231 10160 3232
rect 15770 3296 16090 3297
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 3231 16090 3232
rect 0 3090 800 3120
rect 2589 3090 2655 3093
rect 0 3088 2655 3090
rect 0 3032 2594 3088
rect 2650 3032 2655 3088
rect 0 3030 2655 3032
rect 0 3000 800 3030
rect 2589 3027 2655 3030
rect 17585 3090 17651 3093
rect 19200 3090 20000 3120
rect 17585 3088 20000 3090
rect 17585 3032 17590 3088
rect 17646 3032 20000 3088
rect 17585 3030 20000 3032
rect 17585 3027 17651 3030
rect 19200 3000 20000 3030
rect 3877 2954 3943 2957
rect 4286 2954 4292 2956
rect 3877 2952 4292 2954
rect 3877 2896 3882 2952
rect 3938 2896 4292 2952
rect 3877 2894 4292 2896
rect 3877 2891 3943 2894
rect 4286 2892 4292 2894
rect 4356 2892 4362 2956
rect 8109 2954 8175 2957
rect 16573 2954 16639 2957
rect 8109 2952 16639 2954
rect 8109 2896 8114 2952
rect 8170 2896 16578 2952
rect 16634 2896 16639 2952
rect 8109 2894 16639 2896
rect 8109 2891 8175 2894
rect 16573 2891 16639 2894
rect 13353 2818 13419 2821
rect 15561 2818 15627 2821
rect 13353 2816 15627 2818
rect 13353 2760 13358 2816
rect 13414 2760 15566 2816
rect 15622 2760 15627 2816
rect 13353 2758 15627 2760
rect 13353 2755 13419 2758
rect 15561 2755 15627 2758
rect 6874 2752 7194 2753
rect 0 2682 800 2712
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7194 2752
rect 6874 2687 7194 2688
rect 12805 2752 13125 2753
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2687 13125 2688
rect 3233 2682 3299 2685
rect 0 2680 3299 2682
rect 0 2624 3238 2680
rect 3294 2624 3299 2680
rect 0 2622 3299 2624
rect 0 2592 800 2622
rect 3233 2619 3299 2622
rect 13537 2682 13603 2685
rect 14181 2682 14247 2685
rect 13537 2680 14247 2682
rect 13537 2624 13542 2680
rect 13598 2624 14186 2680
rect 14242 2624 14247 2680
rect 13537 2622 14247 2624
rect 13537 2619 13603 2622
rect 14181 2619 14247 2622
rect 16573 2682 16639 2685
rect 19200 2682 20000 2712
rect 16573 2680 20000 2682
rect 16573 2624 16578 2680
rect 16634 2624 20000 2680
rect 16573 2622 20000 2624
rect 16573 2619 16639 2622
rect 19200 2592 20000 2622
rect 13261 2548 13327 2549
rect 13261 2546 13308 2548
rect 13180 2544 13308 2546
rect 13372 2546 13378 2548
rect 17677 2546 17743 2549
rect 13372 2544 17743 2546
rect 13180 2488 13266 2544
rect 13372 2488 17682 2544
rect 17738 2488 17743 2544
rect 13180 2486 13308 2488
rect 13261 2484 13308 2486
rect 13372 2486 17743 2488
rect 13372 2484 13378 2486
rect 13261 2483 13327 2484
rect 17677 2483 17743 2486
rect 0 2274 800 2304
rect 3693 2274 3759 2277
rect 0 2272 3759 2274
rect 0 2216 3698 2272
rect 3754 2216 3759 2272
rect 0 2214 3759 2216
rect 0 2184 800 2214
rect 3693 2211 3759 2214
rect 17309 2274 17375 2277
rect 19200 2274 20000 2304
rect 17309 2272 20000 2274
rect 17309 2216 17314 2272
rect 17370 2216 20000 2272
rect 17309 2214 20000 2216
rect 17309 2211 17375 2214
rect 3909 2208 4229 2209
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2143 4229 2144
rect 9840 2208 10160 2209
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2143 10160 2144
rect 15770 2208 16090 2209
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 19200 2184 20000 2214
rect 15770 2143 16090 2144
rect 0 1866 800 1896
rect 1577 1866 1643 1869
rect 0 1864 1643 1866
rect 0 1808 1582 1864
rect 1638 1808 1643 1864
rect 0 1806 1643 1808
rect 0 1776 800 1806
rect 1577 1803 1643 1806
rect 17769 1866 17835 1869
rect 19200 1866 20000 1896
rect 17769 1864 20000 1866
rect 17769 1808 17774 1864
rect 17830 1808 20000 1864
rect 17769 1806 20000 1808
rect 17769 1803 17835 1806
rect 19200 1776 20000 1806
rect 0 1458 800 1488
rect 1669 1458 1735 1461
rect 0 1456 1735 1458
rect 0 1400 1674 1456
rect 1730 1400 1735 1456
rect 0 1398 1735 1400
rect 0 1368 800 1398
rect 1669 1395 1735 1398
rect 17217 1458 17283 1461
rect 19200 1458 20000 1488
rect 17217 1456 20000 1458
rect 17217 1400 17222 1456
rect 17278 1400 20000 1456
rect 17217 1398 20000 1400
rect 17217 1395 17283 1398
rect 19200 1368 20000 1398
rect 0 1050 800 1080
rect 2865 1050 2931 1053
rect 0 1048 2931 1050
rect 0 992 2870 1048
rect 2926 992 2931 1048
rect 0 990 2931 992
rect 0 960 800 990
rect 2865 987 2931 990
rect 17861 1050 17927 1053
rect 19200 1050 20000 1080
rect 17861 1048 20000 1050
rect 17861 992 17866 1048
rect 17922 992 20000 1048
rect 17861 990 20000 992
rect 17861 987 17927 990
rect 19200 960 20000 990
rect 0 642 800 672
rect 2773 642 2839 645
rect 0 640 2839 642
rect 0 584 2778 640
rect 2834 584 2839 640
rect 0 582 2839 584
rect 0 552 800 582
rect 2773 579 2839 582
rect 16481 642 16547 645
rect 19200 642 20000 672
rect 16481 640 20000 642
rect 16481 584 16486 640
rect 16542 584 20000 640
rect 16481 582 20000 584
rect 16481 579 16547 582
rect 19200 552 20000 582
rect 0 234 800 264
rect 3509 234 3575 237
rect 0 232 3575 234
rect 0 176 3514 232
rect 3570 176 3575 232
rect 0 174 3575 176
rect 0 144 800 174
rect 3509 171 3575 174
rect 18229 234 18295 237
rect 19200 234 20000 264
rect 18229 232 20000 234
rect 18229 176 18234 232
rect 18290 176 20000 232
rect 18229 174 20000 176
rect 18229 171 18295 174
rect 19200 144 20000 174
<< via3 >>
rect 6882 14716 6946 14720
rect 6882 14660 6886 14716
rect 6886 14660 6942 14716
rect 6942 14660 6946 14716
rect 6882 14656 6946 14660
rect 6962 14716 7026 14720
rect 6962 14660 6966 14716
rect 6966 14660 7022 14716
rect 7022 14660 7026 14716
rect 6962 14656 7026 14660
rect 7042 14716 7106 14720
rect 7042 14660 7046 14716
rect 7046 14660 7102 14716
rect 7102 14660 7106 14716
rect 7042 14656 7106 14660
rect 7122 14716 7186 14720
rect 7122 14660 7126 14716
rect 7126 14660 7182 14716
rect 7182 14660 7186 14716
rect 7122 14656 7186 14660
rect 12813 14716 12877 14720
rect 12813 14660 12817 14716
rect 12817 14660 12873 14716
rect 12873 14660 12877 14716
rect 12813 14656 12877 14660
rect 12893 14716 12957 14720
rect 12893 14660 12897 14716
rect 12897 14660 12953 14716
rect 12953 14660 12957 14716
rect 12893 14656 12957 14660
rect 12973 14716 13037 14720
rect 12973 14660 12977 14716
rect 12977 14660 13033 14716
rect 13033 14660 13037 14716
rect 12973 14656 13037 14660
rect 13053 14716 13117 14720
rect 13053 14660 13057 14716
rect 13057 14660 13113 14716
rect 13113 14660 13117 14716
rect 13053 14656 13117 14660
rect 3917 14172 3981 14176
rect 3917 14116 3921 14172
rect 3921 14116 3977 14172
rect 3977 14116 3981 14172
rect 3917 14112 3981 14116
rect 3997 14172 4061 14176
rect 3997 14116 4001 14172
rect 4001 14116 4057 14172
rect 4057 14116 4061 14172
rect 3997 14112 4061 14116
rect 4077 14172 4141 14176
rect 4077 14116 4081 14172
rect 4081 14116 4137 14172
rect 4137 14116 4141 14172
rect 4077 14112 4141 14116
rect 4157 14172 4221 14176
rect 4157 14116 4161 14172
rect 4161 14116 4217 14172
rect 4217 14116 4221 14172
rect 4157 14112 4221 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 15778 14172 15842 14176
rect 15778 14116 15782 14172
rect 15782 14116 15838 14172
rect 15838 14116 15842 14172
rect 15778 14112 15842 14116
rect 15858 14172 15922 14176
rect 15858 14116 15862 14172
rect 15862 14116 15918 14172
rect 15918 14116 15922 14172
rect 15858 14112 15922 14116
rect 15938 14172 16002 14176
rect 15938 14116 15942 14172
rect 15942 14116 15998 14172
rect 15998 14116 16002 14172
rect 15938 14112 16002 14116
rect 16018 14172 16082 14176
rect 16018 14116 16022 14172
rect 16022 14116 16078 14172
rect 16078 14116 16082 14172
rect 16018 14112 16082 14116
rect 6882 13628 6946 13632
rect 6882 13572 6886 13628
rect 6886 13572 6942 13628
rect 6942 13572 6946 13628
rect 6882 13568 6946 13572
rect 6962 13628 7026 13632
rect 6962 13572 6966 13628
rect 6966 13572 7022 13628
rect 7022 13572 7026 13628
rect 6962 13568 7026 13572
rect 7042 13628 7106 13632
rect 7042 13572 7046 13628
rect 7046 13572 7102 13628
rect 7102 13572 7106 13628
rect 7042 13568 7106 13572
rect 7122 13628 7186 13632
rect 7122 13572 7126 13628
rect 7126 13572 7182 13628
rect 7182 13572 7186 13628
rect 7122 13568 7186 13572
rect 12813 13628 12877 13632
rect 12813 13572 12817 13628
rect 12817 13572 12873 13628
rect 12873 13572 12877 13628
rect 12813 13568 12877 13572
rect 12893 13628 12957 13632
rect 12893 13572 12897 13628
rect 12897 13572 12953 13628
rect 12953 13572 12957 13628
rect 12893 13568 12957 13572
rect 12973 13628 13037 13632
rect 12973 13572 12977 13628
rect 12977 13572 13033 13628
rect 13033 13572 13037 13628
rect 12973 13568 13037 13572
rect 13053 13628 13117 13632
rect 13053 13572 13057 13628
rect 13057 13572 13113 13628
rect 13113 13572 13117 13628
rect 13053 13568 13117 13572
rect 3917 13084 3981 13088
rect 3917 13028 3921 13084
rect 3921 13028 3977 13084
rect 3977 13028 3981 13084
rect 3917 13024 3981 13028
rect 3997 13084 4061 13088
rect 3997 13028 4001 13084
rect 4001 13028 4057 13084
rect 4057 13028 4061 13084
rect 3997 13024 4061 13028
rect 4077 13084 4141 13088
rect 4077 13028 4081 13084
rect 4081 13028 4137 13084
rect 4137 13028 4141 13084
rect 4077 13024 4141 13028
rect 4157 13084 4221 13088
rect 4157 13028 4161 13084
rect 4161 13028 4217 13084
rect 4217 13028 4221 13084
rect 4157 13024 4221 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 15778 13084 15842 13088
rect 15778 13028 15782 13084
rect 15782 13028 15838 13084
rect 15838 13028 15842 13084
rect 15778 13024 15842 13028
rect 15858 13084 15922 13088
rect 15858 13028 15862 13084
rect 15862 13028 15918 13084
rect 15918 13028 15922 13084
rect 15858 13024 15922 13028
rect 15938 13084 16002 13088
rect 15938 13028 15942 13084
rect 15942 13028 15998 13084
rect 15998 13028 16002 13084
rect 15938 13024 16002 13028
rect 16018 13084 16082 13088
rect 16018 13028 16022 13084
rect 16022 13028 16078 13084
rect 16078 13028 16082 13084
rect 16018 13024 16082 13028
rect 6882 12540 6946 12544
rect 6882 12484 6886 12540
rect 6886 12484 6942 12540
rect 6942 12484 6946 12540
rect 6882 12480 6946 12484
rect 6962 12540 7026 12544
rect 6962 12484 6966 12540
rect 6966 12484 7022 12540
rect 7022 12484 7026 12540
rect 6962 12480 7026 12484
rect 7042 12540 7106 12544
rect 7042 12484 7046 12540
rect 7046 12484 7102 12540
rect 7102 12484 7106 12540
rect 7042 12480 7106 12484
rect 7122 12540 7186 12544
rect 7122 12484 7126 12540
rect 7126 12484 7182 12540
rect 7182 12484 7186 12540
rect 7122 12480 7186 12484
rect 12813 12540 12877 12544
rect 12813 12484 12817 12540
rect 12817 12484 12873 12540
rect 12873 12484 12877 12540
rect 12813 12480 12877 12484
rect 12893 12540 12957 12544
rect 12893 12484 12897 12540
rect 12897 12484 12953 12540
rect 12953 12484 12957 12540
rect 12893 12480 12957 12484
rect 12973 12540 13037 12544
rect 12973 12484 12977 12540
rect 12977 12484 13033 12540
rect 13033 12484 13037 12540
rect 12973 12480 13037 12484
rect 13053 12540 13117 12544
rect 13053 12484 13057 12540
rect 13057 12484 13113 12540
rect 13113 12484 13117 12540
rect 13053 12480 13117 12484
rect 16252 12412 16316 12476
rect 3917 11996 3981 12000
rect 3917 11940 3921 11996
rect 3921 11940 3977 11996
rect 3977 11940 3981 11996
rect 3917 11936 3981 11940
rect 3997 11996 4061 12000
rect 3997 11940 4001 11996
rect 4001 11940 4057 11996
rect 4057 11940 4061 11996
rect 3997 11936 4061 11940
rect 4077 11996 4141 12000
rect 4077 11940 4081 11996
rect 4081 11940 4137 11996
rect 4137 11940 4141 11996
rect 4077 11936 4141 11940
rect 4157 11996 4221 12000
rect 4157 11940 4161 11996
rect 4161 11940 4217 11996
rect 4217 11940 4221 11996
rect 4157 11936 4221 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 15778 11996 15842 12000
rect 15778 11940 15782 11996
rect 15782 11940 15838 11996
rect 15838 11940 15842 11996
rect 15778 11936 15842 11940
rect 15858 11996 15922 12000
rect 15858 11940 15862 11996
rect 15862 11940 15918 11996
rect 15918 11940 15922 11996
rect 15858 11936 15922 11940
rect 15938 11996 16002 12000
rect 15938 11940 15942 11996
rect 15942 11940 15998 11996
rect 15998 11940 16002 11996
rect 15938 11936 16002 11940
rect 16018 11996 16082 12000
rect 16018 11940 16022 11996
rect 16022 11940 16078 11996
rect 16078 11940 16082 11996
rect 16018 11936 16082 11940
rect 15332 11928 15396 11932
rect 15332 11872 15382 11928
rect 15382 11872 15396 11928
rect 15332 11868 15396 11872
rect 6882 11452 6946 11456
rect 6882 11396 6886 11452
rect 6886 11396 6942 11452
rect 6942 11396 6946 11452
rect 6882 11392 6946 11396
rect 6962 11452 7026 11456
rect 6962 11396 6966 11452
rect 6966 11396 7022 11452
rect 7022 11396 7026 11452
rect 6962 11392 7026 11396
rect 7042 11452 7106 11456
rect 7042 11396 7046 11452
rect 7046 11396 7102 11452
rect 7102 11396 7106 11452
rect 7042 11392 7106 11396
rect 7122 11452 7186 11456
rect 7122 11396 7126 11452
rect 7126 11396 7182 11452
rect 7182 11396 7186 11452
rect 7122 11392 7186 11396
rect 12813 11452 12877 11456
rect 12813 11396 12817 11452
rect 12817 11396 12873 11452
rect 12873 11396 12877 11452
rect 12813 11392 12877 11396
rect 12893 11452 12957 11456
rect 12893 11396 12897 11452
rect 12897 11396 12953 11452
rect 12953 11396 12957 11452
rect 12893 11392 12957 11396
rect 12973 11452 13037 11456
rect 12973 11396 12977 11452
rect 12977 11396 13033 11452
rect 13033 11396 13037 11452
rect 12973 11392 13037 11396
rect 13053 11452 13117 11456
rect 13053 11396 13057 11452
rect 13057 11396 13113 11452
rect 13113 11396 13117 11452
rect 13053 11392 13117 11396
rect 3917 10908 3981 10912
rect 3917 10852 3921 10908
rect 3921 10852 3977 10908
rect 3977 10852 3981 10908
rect 3917 10848 3981 10852
rect 3997 10908 4061 10912
rect 3997 10852 4001 10908
rect 4001 10852 4057 10908
rect 4057 10852 4061 10908
rect 3997 10848 4061 10852
rect 4077 10908 4141 10912
rect 4077 10852 4081 10908
rect 4081 10852 4137 10908
rect 4137 10852 4141 10908
rect 4077 10848 4141 10852
rect 4157 10908 4221 10912
rect 4157 10852 4161 10908
rect 4161 10852 4217 10908
rect 4217 10852 4221 10908
rect 4157 10848 4221 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 15778 10908 15842 10912
rect 15778 10852 15782 10908
rect 15782 10852 15838 10908
rect 15838 10852 15842 10908
rect 15778 10848 15842 10852
rect 15858 10908 15922 10912
rect 15858 10852 15862 10908
rect 15862 10852 15918 10908
rect 15918 10852 15922 10908
rect 15858 10848 15922 10852
rect 15938 10908 16002 10912
rect 15938 10852 15942 10908
rect 15942 10852 15998 10908
rect 15998 10852 16002 10908
rect 15938 10848 16002 10852
rect 16018 10908 16082 10912
rect 16018 10852 16022 10908
rect 16022 10852 16078 10908
rect 16078 10852 16082 10908
rect 16018 10848 16082 10852
rect 16252 10508 16316 10572
rect 6882 10364 6946 10368
rect 6882 10308 6886 10364
rect 6886 10308 6942 10364
rect 6942 10308 6946 10364
rect 6882 10304 6946 10308
rect 6962 10364 7026 10368
rect 6962 10308 6966 10364
rect 6966 10308 7022 10364
rect 7022 10308 7026 10364
rect 6962 10304 7026 10308
rect 7042 10364 7106 10368
rect 7042 10308 7046 10364
rect 7046 10308 7102 10364
rect 7102 10308 7106 10364
rect 7042 10304 7106 10308
rect 7122 10364 7186 10368
rect 7122 10308 7126 10364
rect 7126 10308 7182 10364
rect 7182 10308 7186 10364
rect 7122 10304 7186 10308
rect 12813 10364 12877 10368
rect 12813 10308 12817 10364
rect 12817 10308 12873 10364
rect 12873 10308 12877 10364
rect 12813 10304 12877 10308
rect 12893 10364 12957 10368
rect 12893 10308 12897 10364
rect 12897 10308 12953 10364
rect 12953 10308 12957 10364
rect 12893 10304 12957 10308
rect 12973 10364 13037 10368
rect 12973 10308 12977 10364
rect 12977 10308 13033 10364
rect 13033 10308 13037 10364
rect 12973 10304 13037 10308
rect 13053 10364 13117 10368
rect 13053 10308 13057 10364
rect 13057 10308 13113 10364
rect 13113 10308 13117 10364
rect 13053 10304 13117 10308
rect 3917 9820 3981 9824
rect 3917 9764 3921 9820
rect 3921 9764 3977 9820
rect 3977 9764 3981 9820
rect 3917 9760 3981 9764
rect 3997 9820 4061 9824
rect 3997 9764 4001 9820
rect 4001 9764 4057 9820
rect 4057 9764 4061 9820
rect 3997 9760 4061 9764
rect 4077 9820 4141 9824
rect 4077 9764 4081 9820
rect 4081 9764 4137 9820
rect 4137 9764 4141 9820
rect 4077 9760 4141 9764
rect 4157 9820 4221 9824
rect 4157 9764 4161 9820
rect 4161 9764 4217 9820
rect 4217 9764 4221 9820
rect 4157 9760 4221 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 15778 9820 15842 9824
rect 15778 9764 15782 9820
rect 15782 9764 15838 9820
rect 15838 9764 15842 9820
rect 15778 9760 15842 9764
rect 15858 9820 15922 9824
rect 15858 9764 15862 9820
rect 15862 9764 15918 9820
rect 15918 9764 15922 9820
rect 15858 9760 15922 9764
rect 15938 9820 16002 9824
rect 15938 9764 15942 9820
rect 15942 9764 15998 9820
rect 15998 9764 16002 9820
rect 15938 9760 16002 9764
rect 16018 9820 16082 9824
rect 16018 9764 16022 9820
rect 16022 9764 16078 9820
rect 16078 9764 16082 9820
rect 16018 9760 16082 9764
rect 6882 9276 6946 9280
rect 6882 9220 6886 9276
rect 6886 9220 6942 9276
rect 6942 9220 6946 9276
rect 6882 9216 6946 9220
rect 6962 9276 7026 9280
rect 6962 9220 6966 9276
rect 6966 9220 7022 9276
rect 7022 9220 7026 9276
rect 6962 9216 7026 9220
rect 7042 9276 7106 9280
rect 7042 9220 7046 9276
rect 7046 9220 7102 9276
rect 7102 9220 7106 9276
rect 7042 9216 7106 9220
rect 7122 9276 7186 9280
rect 7122 9220 7126 9276
rect 7126 9220 7182 9276
rect 7182 9220 7186 9276
rect 7122 9216 7186 9220
rect 12813 9276 12877 9280
rect 12813 9220 12817 9276
rect 12817 9220 12873 9276
rect 12873 9220 12877 9276
rect 12813 9216 12877 9220
rect 12893 9276 12957 9280
rect 12893 9220 12897 9276
rect 12897 9220 12953 9276
rect 12953 9220 12957 9276
rect 12893 9216 12957 9220
rect 12973 9276 13037 9280
rect 12973 9220 12977 9276
rect 12977 9220 13033 9276
rect 13033 9220 13037 9276
rect 12973 9216 13037 9220
rect 13053 9276 13117 9280
rect 13053 9220 13057 9276
rect 13057 9220 13113 9276
rect 13113 9220 13117 9276
rect 13053 9216 13117 9220
rect 3917 8732 3981 8736
rect 3917 8676 3921 8732
rect 3921 8676 3977 8732
rect 3977 8676 3981 8732
rect 3917 8672 3981 8676
rect 3997 8732 4061 8736
rect 3997 8676 4001 8732
rect 4001 8676 4057 8732
rect 4057 8676 4061 8732
rect 3997 8672 4061 8676
rect 4077 8732 4141 8736
rect 4077 8676 4081 8732
rect 4081 8676 4137 8732
rect 4137 8676 4141 8732
rect 4077 8672 4141 8676
rect 4157 8732 4221 8736
rect 4157 8676 4161 8732
rect 4161 8676 4217 8732
rect 4217 8676 4221 8732
rect 4157 8672 4221 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 15778 8732 15842 8736
rect 15778 8676 15782 8732
rect 15782 8676 15838 8732
rect 15838 8676 15842 8732
rect 15778 8672 15842 8676
rect 15858 8732 15922 8736
rect 15858 8676 15862 8732
rect 15862 8676 15918 8732
rect 15918 8676 15922 8732
rect 15858 8672 15922 8676
rect 15938 8732 16002 8736
rect 15938 8676 15942 8732
rect 15942 8676 15998 8732
rect 15998 8676 16002 8732
rect 15938 8672 16002 8676
rect 16018 8732 16082 8736
rect 16018 8676 16022 8732
rect 16022 8676 16078 8732
rect 16078 8676 16082 8732
rect 16018 8672 16082 8676
rect 4292 8528 4356 8532
rect 4292 8472 4306 8528
rect 4306 8472 4356 8528
rect 4292 8468 4356 8472
rect 6882 8188 6946 8192
rect 6882 8132 6886 8188
rect 6886 8132 6942 8188
rect 6942 8132 6946 8188
rect 6882 8128 6946 8132
rect 6962 8188 7026 8192
rect 6962 8132 6966 8188
rect 6966 8132 7022 8188
rect 7022 8132 7026 8188
rect 6962 8128 7026 8132
rect 7042 8188 7106 8192
rect 7042 8132 7046 8188
rect 7046 8132 7102 8188
rect 7102 8132 7106 8188
rect 7042 8128 7106 8132
rect 7122 8188 7186 8192
rect 7122 8132 7126 8188
rect 7126 8132 7182 8188
rect 7182 8132 7186 8188
rect 7122 8128 7186 8132
rect 12813 8188 12877 8192
rect 12813 8132 12817 8188
rect 12817 8132 12873 8188
rect 12873 8132 12877 8188
rect 12813 8128 12877 8132
rect 12893 8188 12957 8192
rect 12893 8132 12897 8188
rect 12897 8132 12953 8188
rect 12953 8132 12957 8188
rect 12893 8128 12957 8132
rect 12973 8188 13037 8192
rect 12973 8132 12977 8188
rect 12977 8132 13033 8188
rect 13033 8132 13037 8188
rect 12973 8128 13037 8132
rect 13053 8188 13117 8192
rect 13053 8132 13057 8188
rect 13057 8132 13113 8188
rect 13113 8132 13117 8188
rect 13053 8128 13117 8132
rect 3917 7644 3981 7648
rect 3917 7588 3921 7644
rect 3921 7588 3977 7644
rect 3977 7588 3981 7644
rect 3917 7584 3981 7588
rect 3997 7644 4061 7648
rect 3997 7588 4001 7644
rect 4001 7588 4057 7644
rect 4057 7588 4061 7644
rect 3997 7584 4061 7588
rect 4077 7644 4141 7648
rect 4077 7588 4081 7644
rect 4081 7588 4137 7644
rect 4137 7588 4141 7644
rect 4077 7584 4141 7588
rect 4157 7644 4221 7648
rect 4157 7588 4161 7644
rect 4161 7588 4217 7644
rect 4217 7588 4221 7644
rect 4157 7584 4221 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 15778 7644 15842 7648
rect 15778 7588 15782 7644
rect 15782 7588 15838 7644
rect 15838 7588 15842 7644
rect 15778 7584 15842 7588
rect 15858 7644 15922 7648
rect 15858 7588 15862 7644
rect 15862 7588 15918 7644
rect 15918 7588 15922 7644
rect 15858 7584 15922 7588
rect 15938 7644 16002 7648
rect 15938 7588 15942 7644
rect 15942 7588 15998 7644
rect 15998 7588 16002 7644
rect 15938 7584 16002 7588
rect 16018 7644 16082 7648
rect 16018 7588 16022 7644
rect 16022 7588 16078 7644
rect 16078 7588 16082 7644
rect 16018 7584 16082 7588
rect 13308 7516 13372 7580
rect 6882 7100 6946 7104
rect 6882 7044 6886 7100
rect 6886 7044 6942 7100
rect 6942 7044 6946 7100
rect 6882 7040 6946 7044
rect 6962 7100 7026 7104
rect 6962 7044 6966 7100
rect 6966 7044 7022 7100
rect 7022 7044 7026 7100
rect 6962 7040 7026 7044
rect 7042 7100 7106 7104
rect 7042 7044 7046 7100
rect 7046 7044 7102 7100
rect 7102 7044 7106 7100
rect 7042 7040 7106 7044
rect 7122 7100 7186 7104
rect 7122 7044 7126 7100
rect 7126 7044 7182 7100
rect 7182 7044 7186 7100
rect 7122 7040 7186 7044
rect 12813 7100 12877 7104
rect 12813 7044 12817 7100
rect 12817 7044 12873 7100
rect 12873 7044 12877 7100
rect 12813 7040 12877 7044
rect 12893 7100 12957 7104
rect 12893 7044 12897 7100
rect 12897 7044 12953 7100
rect 12953 7044 12957 7100
rect 12893 7040 12957 7044
rect 12973 7100 13037 7104
rect 12973 7044 12977 7100
rect 12977 7044 13033 7100
rect 13033 7044 13037 7100
rect 12973 7040 13037 7044
rect 13053 7100 13117 7104
rect 13053 7044 13057 7100
rect 13057 7044 13113 7100
rect 13113 7044 13117 7100
rect 13053 7040 13117 7044
rect 12388 6972 12452 7036
rect 3917 6556 3981 6560
rect 3917 6500 3921 6556
rect 3921 6500 3977 6556
rect 3977 6500 3981 6556
rect 3917 6496 3981 6500
rect 3997 6556 4061 6560
rect 3997 6500 4001 6556
rect 4001 6500 4057 6556
rect 4057 6500 4061 6556
rect 3997 6496 4061 6500
rect 4077 6556 4141 6560
rect 4077 6500 4081 6556
rect 4081 6500 4137 6556
rect 4137 6500 4141 6556
rect 4077 6496 4141 6500
rect 4157 6556 4221 6560
rect 4157 6500 4161 6556
rect 4161 6500 4217 6556
rect 4217 6500 4221 6556
rect 4157 6496 4221 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 15778 6556 15842 6560
rect 15778 6500 15782 6556
rect 15782 6500 15838 6556
rect 15838 6500 15842 6556
rect 15778 6496 15842 6500
rect 15858 6556 15922 6560
rect 15858 6500 15862 6556
rect 15862 6500 15918 6556
rect 15918 6500 15922 6556
rect 15858 6496 15922 6500
rect 15938 6556 16002 6560
rect 15938 6500 15942 6556
rect 15942 6500 15998 6556
rect 15998 6500 16002 6556
rect 15938 6496 16002 6500
rect 16018 6556 16082 6560
rect 16018 6500 16022 6556
rect 16022 6500 16078 6556
rect 16078 6500 16082 6556
rect 16018 6496 16082 6500
rect 6882 6012 6946 6016
rect 6882 5956 6886 6012
rect 6886 5956 6942 6012
rect 6942 5956 6946 6012
rect 6882 5952 6946 5956
rect 6962 6012 7026 6016
rect 6962 5956 6966 6012
rect 6966 5956 7022 6012
rect 7022 5956 7026 6012
rect 6962 5952 7026 5956
rect 7042 6012 7106 6016
rect 7042 5956 7046 6012
rect 7046 5956 7102 6012
rect 7102 5956 7106 6012
rect 7042 5952 7106 5956
rect 7122 6012 7186 6016
rect 7122 5956 7126 6012
rect 7126 5956 7182 6012
rect 7182 5956 7186 6012
rect 7122 5952 7186 5956
rect 12813 6012 12877 6016
rect 12813 5956 12817 6012
rect 12817 5956 12873 6012
rect 12873 5956 12877 6012
rect 12813 5952 12877 5956
rect 12893 6012 12957 6016
rect 12893 5956 12897 6012
rect 12897 5956 12953 6012
rect 12953 5956 12957 6012
rect 12893 5952 12957 5956
rect 12973 6012 13037 6016
rect 12973 5956 12977 6012
rect 12977 5956 13033 6012
rect 13033 5956 13037 6012
rect 12973 5952 13037 5956
rect 13053 6012 13117 6016
rect 13053 5956 13057 6012
rect 13057 5956 13113 6012
rect 13113 5956 13117 6012
rect 13053 5952 13117 5956
rect 15332 5476 15396 5540
rect 3917 5468 3981 5472
rect 3917 5412 3921 5468
rect 3921 5412 3977 5468
rect 3977 5412 3981 5468
rect 3917 5408 3981 5412
rect 3997 5468 4061 5472
rect 3997 5412 4001 5468
rect 4001 5412 4057 5468
rect 4057 5412 4061 5468
rect 3997 5408 4061 5412
rect 4077 5468 4141 5472
rect 4077 5412 4081 5468
rect 4081 5412 4137 5468
rect 4137 5412 4141 5468
rect 4077 5408 4141 5412
rect 4157 5468 4221 5472
rect 4157 5412 4161 5468
rect 4161 5412 4217 5468
rect 4217 5412 4221 5468
rect 4157 5408 4221 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 15778 5468 15842 5472
rect 15778 5412 15782 5468
rect 15782 5412 15838 5468
rect 15838 5412 15842 5468
rect 15778 5408 15842 5412
rect 15858 5468 15922 5472
rect 15858 5412 15862 5468
rect 15862 5412 15918 5468
rect 15918 5412 15922 5468
rect 15858 5408 15922 5412
rect 15938 5468 16002 5472
rect 15938 5412 15942 5468
rect 15942 5412 15998 5468
rect 15998 5412 16002 5468
rect 15938 5408 16002 5412
rect 16018 5468 16082 5472
rect 16018 5412 16022 5468
rect 16022 5412 16078 5468
rect 16078 5412 16082 5468
rect 16018 5408 16082 5412
rect 12388 5204 12452 5268
rect 6882 4924 6946 4928
rect 6882 4868 6886 4924
rect 6886 4868 6942 4924
rect 6942 4868 6946 4924
rect 6882 4864 6946 4868
rect 6962 4924 7026 4928
rect 6962 4868 6966 4924
rect 6966 4868 7022 4924
rect 7022 4868 7026 4924
rect 6962 4864 7026 4868
rect 7042 4924 7106 4928
rect 7042 4868 7046 4924
rect 7046 4868 7102 4924
rect 7102 4868 7106 4924
rect 7042 4864 7106 4868
rect 7122 4924 7186 4928
rect 7122 4868 7126 4924
rect 7126 4868 7182 4924
rect 7182 4868 7186 4924
rect 7122 4864 7186 4868
rect 12813 4924 12877 4928
rect 12813 4868 12817 4924
rect 12817 4868 12873 4924
rect 12873 4868 12877 4924
rect 12813 4864 12877 4868
rect 12893 4924 12957 4928
rect 12893 4868 12897 4924
rect 12897 4868 12953 4924
rect 12953 4868 12957 4924
rect 12893 4864 12957 4868
rect 12973 4924 13037 4928
rect 12973 4868 12977 4924
rect 12977 4868 13033 4924
rect 13033 4868 13037 4924
rect 12973 4864 13037 4868
rect 13053 4924 13117 4928
rect 13053 4868 13057 4924
rect 13057 4868 13113 4924
rect 13113 4868 13117 4924
rect 13053 4864 13117 4868
rect 3917 4380 3981 4384
rect 3917 4324 3921 4380
rect 3921 4324 3977 4380
rect 3977 4324 3981 4380
rect 3917 4320 3981 4324
rect 3997 4380 4061 4384
rect 3997 4324 4001 4380
rect 4001 4324 4057 4380
rect 4057 4324 4061 4380
rect 3997 4320 4061 4324
rect 4077 4380 4141 4384
rect 4077 4324 4081 4380
rect 4081 4324 4137 4380
rect 4137 4324 4141 4380
rect 4077 4320 4141 4324
rect 4157 4380 4221 4384
rect 4157 4324 4161 4380
rect 4161 4324 4217 4380
rect 4217 4324 4221 4380
rect 4157 4320 4221 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 15778 4380 15842 4384
rect 15778 4324 15782 4380
rect 15782 4324 15838 4380
rect 15838 4324 15842 4380
rect 15778 4320 15842 4324
rect 15858 4380 15922 4384
rect 15858 4324 15862 4380
rect 15862 4324 15918 4380
rect 15918 4324 15922 4380
rect 15858 4320 15922 4324
rect 15938 4380 16002 4384
rect 15938 4324 15942 4380
rect 15942 4324 15998 4380
rect 15998 4324 16002 4380
rect 15938 4320 16002 4324
rect 16018 4380 16082 4384
rect 16018 4324 16022 4380
rect 16022 4324 16078 4380
rect 16078 4324 16082 4380
rect 16018 4320 16082 4324
rect 6882 3836 6946 3840
rect 6882 3780 6886 3836
rect 6886 3780 6942 3836
rect 6942 3780 6946 3836
rect 6882 3776 6946 3780
rect 6962 3836 7026 3840
rect 6962 3780 6966 3836
rect 6966 3780 7022 3836
rect 7022 3780 7026 3836
rect 6962 3776 7026 3780
rect 7042 3836 7106 3840
rect 7042 3780 7046 3836
rect 7046 3780 7102 3836
rect 7102 3780 7106 3836
rect 7042 3776 7106 3780
rect 7122 3836 7186 3840
rect 7122 3780 7126 3836
rect 7126 3780 7182 3836
rect 7182 3780 7186 3836
rect 7122 3776 7186 3780
rect 12813 3836 12877 3840
rect 12813 3780 12817 3836
rect 12817 3780 12873 3836
rect 12873 3780 12877 3836
rect 12813 3776 12877 3780
rect 12893 3836 12957 3840
rect 12893 3780 12897 3836
rect 12897 3780 12953 3836
rect 12953 3780 12957 3836
rect 12893 3776 12957 3780
rect 12973 3836 13037 3840
rect 12973 3780 12977 3836
rect 12977 3780 13033 3836
rect 13033 3780 13037 3836
rect 12973 3776 13037 3780
rect 13053 3836 13117 3840
rect 13053 3780 13057 3836
rect 13057 3780 13113 3836
rect 13113 3780 13117 3836
rect 13053 3776 13117 3780
rect 3917 3292 3981 3296
rect 3917 3236 3921 3292
rect 3921 3236 3977 3292
rect 3977 3236 3981 3292
rect 3917 3232 3981 3236
rect 3997 3292 4061 3296
rect 3997 3236 4001 3292
rect 4001 3236 4057 3292
rect 4057 3236 4061 3292
rect 3997 3232 4061 3236
rect 4077 3292 4141 3296
rect 4077 3236 4081 3292
rect 4081 3236 4137 3292
rect 4137 3236 4141 3292
rect 4077 3232 4141 3236
rect 4157 3292 4221 3296
rect 4157 3236 4161 3292
rect 4161 3236 4217 3292
rect 4217 3236 4221 3292
rect 4157 3232 4221 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 15778 3292 15842 3296
rect 15778 3236 15782 3292
rect 15782 3236 15838 3292
rect 15838 3236 15842 3292
rect 15778 3232 15842 3236
rect 15858 3292 15922 3296
rect 15858 3236 15862 3292
rect 15862 3236 15918 3292
rect 15918 3236 15922 3292
rect 15858 3232 15922 3236
rect 15938 3292 16002 3296
rect 15938 3236 15942 3292
rect 15942 3236 15998 3292
rect 15998 3236 16002 3292
rect 15938 3232 16002 3236
rect 16018 3292 16082 3296
rect 16018 3236 16022 3292
rect 16022 3236 16078 3292
rect 16078 3236 16082 3292
rect 16018 3232 16082 3236
rect 4292 2892 4356 2956
rect 6882 2748 6946 2752
rect 6882 2692 6886 2748
rect 6886 2692 6942 2748
rect 6942 2692 6946 2748
rect 6882 2688 6946 2692
rect 6962 2748 7026 2752
rect 6962 2692 6966 2748
rect 6966 2692 7022 2748
rect 7022 2692 7026 2748
rect 6962 2688 7026 2692
rect 7042 2748 7106 2752
rect 7042 2692 7046 2748
rect 7046 2692 7102 2748
rect 7102 2692 7106 2748
rect 7042 2688 7106 2692
rect 7122 2748 7186 2752
rect 7122 2692 7126 2748
rect 7126 2692 7182 2748
rect 7182 2692 7186 2748
rect 7122 2688 7186 2692
rect 12813 2748 12877 2752
rect 12813 2692 12817 2748
rect 12817 2692 12873 2748
rect 12873 2692 12877 2748
rect 12813 2688 12877 2692
rect 12893 2748 12957 2752
rect 12893 2692 12897 2748
rect 12897 2692 12953 2748
rect 12953 2692 12957 2748
rect 12893 2688 12957 2692
rect 12973 2748 13037 2752
rect 12973 2692 12977 2748
rect 12977 2692 13033 2748
rect 13033 2692 13037 2748
rect 12973 2688 13037 2692
rect 13053 2748 13117 2752
rect 13053 2692 13057 2748
rect 13057 2692 13113 2748
rect 13113 2692 13117 2748
rect 13053 2688 13117 2692
rect 13308 2544 13372 2548
rect 13308 2488 13322 2544
rect 13322 2488 13372 2544
rect 13308 2484 13372 2488
rect 3917 2204 3981 2208
rect 3917 2148 3921 2204
rect 3921 2148 3977 2204
rect 3977 2148 3981 2204
rect 3917 2144 3981 2148
rect 3997 2204 4061 2208
rect 3997 2148 4001 2204
rect 4001 2148 4057 2204
rect 4057 2148 4061 2204
rect 3997 2144 4061 2148
rect 4077 2204 4141 2208
rect 4077 2148 4081 2204
rect 4081 2148 4137 2204
rect 4137 2148 4141 2204
rect 4077 2144 4141 2148
rect 4157 2204 4221 2208
rect 4157 2148 4161 2204
rect 4161 2148 4217 2204
rect 4217 2148 4221 2204
rect 4157 2144 4221 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 15778 2204 15842 2208
rect 15778 2148 15782 2204
rect 15782 2148 15838 2204
rect 15838 2148 15842 2204
rect 15778 2144 15842 2148
rect 15858 2204 15922 2208
rect 15858 2148 15862 2204
rect 15862 2148 15918 2204
rect 15918 2148 15922 2204
rect 15858 2144 15922 2148
rect 15938 2204 16002 2208
rect 15938 2148 15942 2204
rect 15942 2148 15998 2204
rect 15998 2148 16002 2204
rect 15938 2144 16002 2148
rect 16018 2204 16082 2208
rect 16018 2148 16022 2204
rect 16022 2148 16078 2204
rect 16078 2148 16082 2204
rect 16018 2144 16082 2148
<< metal4 >>
rect 3909 14176 4229 14736
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 13088 4229 14112
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 12000 4229 13024
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 10912 4229 11936
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 9824 4229 10848
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 8736 4229 9760
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 7648 4229 8672
rect 6874 14720 7195 14736
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7195 14720
rect 6874 13632 7195 14656
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7195 13632
rect 6874 12544 7195 13568
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7195 12544
rect 6874 11456 7195 12480
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7195 11456
rect 6874 10368 7195 11392
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7195 10368
rect 6874 9280 7195 10304
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7195 9280
rect 4291 8532 4357 8533
rect 4291 8468 4292 8532
rect 4356 8468 4357 8532
rect 4291 8467 4357 8468
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 6560 4229 7584
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 5472 4229 6496
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 4384 4229 5408
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 3296 4229 4320
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 2208 4229 3232
rect 4294 2957 4354 8467
rect 6874 8192 7195 9216
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7195 8192
rect 6874 7104 7195 8128
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7195 7104
rect 6874 6016 7195 7040
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7195 6016
rect 6874 4928 7195 5952
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7195 4928
rect 6874 3840 7195 4864
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7195 3840
rect 4291 2956 4357 2957
rect 4291 2892 4292 2956
rect 4356 2892 4357 2956
rect 4291 2891 4357 2892
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2128 4229 2144
rect 6874 2752 7195 3776
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7195 2752
rect 6874 2128 7195 2688
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 12805 14720 13125 14736
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 13632 13125 14656
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 12544 13125 13568
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 11456 13125 12480
rect 15770 14176 16090 14736
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 15770 13088 16090 14112
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15770 12000 16090 13024
rect 16251 12476 16317 12477
rect 16251 12412 16252 12476
rect 16316 12412 16317 12476
rect 16251 12411 16317 12412
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15331 11932 15397 11933
rect 15331 11868 15332 11932
rect 15396 11868 15397 11932
rect 15331 11867 15397 11868
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 10368 13125 11392
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 12805 9280 13125 10304
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 8192 13125 9216
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 7104 13125 8128
rect 13307 7580 13373 7581
rect 13307 7516 13308 7580
rect 13372 7516 13373 7580
rect 13307 7515 13373 7516
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12387 7036 12453 7037
rect 12387 6972 12388 7036
rect 12452 6972 12453 7036
rect 12387 6971 12453 6972
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 12390 5269 12450 6971
rect 12805 6016 13125 7040
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12387 5268 12453 5269
rect 12387 5204 12388 5268
rect 12452 5204 12453 5268
rect 12387 5203 12453 5204
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12805 4928 13125 5952
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 3840 13125 4864
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 2752 13125 3776
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2128 13125 2688
rect 13310 2549 13370 7515
rect 15334 5541 15394 11867
rect 15770 10912 16090 11936
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 9824 16090 10848
rect 16254 10573 16314 12411
rect 16251 10572 16317 10573
rect 16251 10508 16252 10572
rect 16316 10508 16317 10572
rect 16251 10507 16317 10508
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 15770 8736 16090 9760
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 15770 7648 16090 8672
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 6560 16090 7584
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 15331 5540 15397 5541
rect 15331 5476 15332 5540
rect 15396 5476 15397 5540
rect 15331 5475 15397 5476
rect 15770 5472 16090 6496
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15770 4384 16090 5408
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 15770 3296 16090 4320
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 13307 2548 13373 2549
rect 13307 2484 13308 2548
rect 13372 2484 13373 2548
rect 13307 2483 13373 2484
rect 15770 2208 16090 3232
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 15770 2128 16090 2144
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608763979
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608763979
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_174
timestamp 1608763979
transform 1 0 17112 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_187
timestamp 1608763979
transform 1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608763979
transform 1 0 15456 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608763979
transform 1 0 15916 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608763979
transform 1 0 15364 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_153
timestamp 1608763979
transform 1 0 15180 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_159
timestamp 1608763979
transform 1 0 15732 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1608763979
transform 1 0 14352 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1608763979
transform 1 0 13340 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_142
timestamp 1608763979
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1608763979
transform 1 0 11132 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608763979
transform 1 0 12512 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_107
timestamp 1608763979
transform 1 0 10948 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_118
timestamp 1608763979
transform 1 0 11960 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_125
timestamp 1608763979
transform 1 0 12604 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1608763979
transform 1 0 10120 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608763979
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_91
timestamp 1608763979
transform 1 0 9476 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_94
timestamp 1608763979
transform 1 0 9752 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1608763979
transform 1 0 8648 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1608763979
transform 1 0 7636 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_63
timestamp 1608763979
transform 1 0 6900 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_80
timestamp 1608763979
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1608763979
transform 1 0 5796 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608763979
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_44
timestamp 1608763979
transform 1 0 5152 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_50
timestamp 1608763979
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_60
timestamp 1608763979
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608763979
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1608763979
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1608763979
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608763979
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1608763979
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1608763979
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608763979
transform -1 0 18860 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_188
timestamp 1608763979
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1608763979
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1608763979
transform 1 0 17388 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608763979
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1608763979
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1608763979
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608763979
transform 1 0 16008 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1608763979
transform 1 0 14996 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_160
timestamp 1608763979
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608763979
transform 1 0 13064 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_129
timestamp 1608763979
transform 1 0 12972 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_139
timestamp 1608763979
transform 1 0 13892 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763979
transform 1 0 11592 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608763979
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_112
timestamp 1608763979
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1608763979
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_123
timestamp 1608763979
transform 1 0 12420 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1608763979
transform 1 0 10580 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1608763979
transform 1 0 9568 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_90
timestamp 1608763979
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_101
timestamp 1608763979
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1608763979
transform 1 0 8556 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_71
timestamp 1608763979
transform 1 0 7636 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_79
timestamp 1608763979
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1608763979
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1608763979
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608763979
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_43
timestamp 1608763979
transform 1 0 5060 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_53
timestamp 1608763979
transform 1 0 5980 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1608763979
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_39
timestamp 1608763979
transform 1 0 4692 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608763979
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1608763979
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1608763979
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608763979
transform -1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608763979
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1608763979
transform 1 0 17480 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1608763979
transform 1 0 16836 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1608763979
transform 1 0 16468 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608763979
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_170
timestamp 1608763979
transform 1 0 16744 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_180
timestamp 1608763979
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_184
timestamp 1608763979
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_176
timestamp 1608763979
transform 1 0 17296 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_187
timestamp 1608763979
transform 1 0 18308 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763979
transform 1 0 14904 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1608763979
transform 1 0 15456 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608763979
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_147
timestamp 1608763979
transform 1 0 14628 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_166
timestamp 1608763979
transform 1 0 16376 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1608763979
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_154
timestamp 1608763979
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_165
timestamp 1608763979
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1608763979
transform 1 0 14168 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1608763979
transform 1 0 13156 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_19_139
timestamp 1608763979
transform 1 0 13892 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_129
timestamp 1608763979
transform 1 0 12972 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_140
timestamp 1608763979
transform 1 0 13984 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763979
transform 1 0 12420 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1608763979
transform 1 0 12144 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1608763979
transform 1 0 11316 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608763979
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_109
timestamp 1608763979
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1608763979
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_111
timestamp 1608763979
transform 1 0 11316 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_119
timestamp 1608763979
transform 1 0 12052 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1608763979
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1608763979
transform 1 0 10304 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1608763979
transform 1 0 10488 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608763979
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_97
timestamp 1608763979
transform 1 0 10028 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1608763979
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_96
timestamp 1608763979
transform 1 0 9936 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763979
transform 1 0 6900 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763979
transform 1 0 8556 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1608763979
transform 1 0 8556 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_79
timestamp 1608763979
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_76
timestamp 1608763979
transform 1 0 8096 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_80
timestamp 1608763979
transform 1 0 8464 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763979
transform 1 0 6624 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608763979
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1608763979
transform 1 0 6348 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_62
timestamp 1608763979
transform 1 0 6808 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_58
timestamp 1608763979
transform 1 0 6440 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1608763979
transform 1 0 5060 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1608763979
transform 1 0 5520 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1608763979
transform 1 0 5612 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_42
timestamp 1608763979
transform 1 0 4968 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_46
timestamp 1608763979
transform 1 0 5336 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_44
timestamp 1608763979
transform 1 0 5152 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_48
timestamp 1608763979
transform 1 0 5520 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763979
transform 1 0 3128 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608763979
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_38
timestamp 1608763979
transform 1 0 4600 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1608763979
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1608763979
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1608763979
transform 1 0 2484 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608763979
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608763979
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1608763979
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_18
timestamp 1608763979
transform 1 0 2760 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1608763979
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1608763979
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608763979
transform -1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763979
transform 1 0 16744 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_168
timestamp 1608763979
transform 1 0 16560 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_186
timestamp 1608763979
transform 1 0 18216 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1608763979
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1608763979
transform 1 0 15732 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608763979
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_148
timestamp 1608763979
transform 1 0 14720 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1608763979
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_157
timestamp 1608763979
transform 1 0 15548 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763979
transform 1 0 13248 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_130
timestamp 1608763979
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1608763979
transform 1 0 12236 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_116
timestamp 1608763979
transform 1 0 11776 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_120
timestamp 1608763979
transform 1 0 12144 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763979
transform 1 0 10304 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608763979
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1608763979
transform 1 0 8924 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1608763979
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_93
timestamp 1608763979
transform 1 0 9660 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_99
timestamp 1608763979
transform 1 0 10212 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1608763979
transform 1 0 7084 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1608763979
transform 1 0 8096 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_63
timestamp 1608763979
transform 1 0 6900 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_74
timestamp 1608763979
transform 1 0 7912 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1608763979
transform 1 0 6072 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_18_48
timestamp 1608763979
transform 1 0 5520 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763979
transform 1 0 4048 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608763979
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1608763979
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1608763979
transform 1 0 2944 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1608763979
transform 1 0 1840 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608763979
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1608763979
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1608763979
transform 1 0 1748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_17
timestamp 1608763979
transform 1 0 2668 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608763979
transform -1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608763979
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_173
timestamp 1608763979
transform 1 0 17020 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1608763979
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_184
timestamp 1608763979
transform 1 0 18032 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1608763979
transform 1 0 16192 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1608763979
transform 1 0 15180 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_150
timestamp 1608763979
transform 1 0 14904 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_162
timestamp 1608763979
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1608763979
transform 1 0 14076 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1608763979
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763979
transform 1 0 12420 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1608763979
transform 1 0 11316 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608763979
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_109
timestamp 1608763979
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1608763979
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1608763979
transform 1 0 9568 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_90
timestamp 1608763979
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_101
timestamp 1608763979
transform 1 0 10396 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763979
transform 1 0 7912 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_71
timestamp 1608763979
transform 1 0 7636 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1608763979
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1608763979
transform 1 0 5704 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608763979
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_45
timestamp 1608763979
transform 1 0 5244 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_49
timestamp 1608763979
transform 1 0 5612 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1608763979
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1608763979
transform 1 0 3220 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763979
transform 1 0 3772 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_21
timestamp 1608763979
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_27
timestamp 1608763979
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1608763979
transform 1 0 1656 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1608763979
transform 1 0 2208 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608763979
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1608763979
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_10
timestamp 1608763979
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608763979
transform -1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1608763979
transform 1 0 17388 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_173
timestamp 1608763979
transform 1 0 17020 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_186
timestamp 1608763979
transform 1 0 18216 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1608763979
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1608763979
transform 1 0 16192 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608763979
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1608763979
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_157
timestamp 1608763979
transform 1 0 15548 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_163
timestamp 1608763979
transform 1 0 16100 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1608763979
transform 1 0 13984 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1608763979
transform 1 0 13800 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763979
transform 1 0 12328 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1608763979
transform 1 0 11316 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763979
transform 1 0 11040 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_120
timestamp 1608763979
transform 1 0 12144 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1608763979
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608763979
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1608763979
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_102
timestamp 1608763979
transform 1 0 10488 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1608763979
transform 1 0 7544 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1608763979
transform 1 0 8556 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_68
timestamp 1608763979
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_79
timestamp 1608763979
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_0_
timestamp 1608763979
transform 1 0 6532 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_48
timestamp 1608763979
transform 1 0 5520 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_56
timestamp 1608763979
transform 1 0 6256 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763979
transform 1 0 4048 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608763979
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_28
timestamp 1608763979
transform 1 0 3680 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1608763979
transform 1 0 1656 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763979
transform 1 0 2208 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608763979
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1608763979
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_10
timestamp 1608763979
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608763979
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608763979
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1608763979
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_184
timestamp 1608763979
transform 1 0 18032 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763979
transform 1 0 14628 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763979
transform 1 0 16284 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_163
timestamp 1608763979
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1608763979
transform 1 0 13616 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_132
timestamp 1608763979
transform 1 0 13248 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_145
timestamp 1608763979
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1608763979
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1608763979
transform 1 0 11316 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608763979
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_110
timestamp 1608763979
transform 1 0 11224 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1608763979
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763979
transform 1 0 9016 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_84
timestamp 1608763979
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_102
timestamp 1608763979
transform 1 0 10488 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763979
transform 1 0 7360 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763979
transform 1 0 7084 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1608763979
transform 1 0 5428 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608763979
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_45
timestamp 1608763979
transform 1 0 5244 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_56
timestamp 1608763979
transform 1 0 6256 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1608763979
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_62
timestamp 1608763979
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1608763979
transform 1 0 4416 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1608763979
transform 1 0 3404 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_21
timestamp 1608763979
transform 1 0 3036 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_34
timestamp 1608763979
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1608763979
transform 1 0 1656 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1608763979
transform 1 0 2208 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608763979
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1608763979
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_10
timestamp 1608763979
transform 1 0 2024 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608763979
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608763979
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_189
timestamp 1608763979
transform 1 0 18492 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1608763979
transform 1 0 17848 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1608763979
transform 1 0 16744 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608763979
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_179
timestamp 1608763979
transform 1 0 17572 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_184
timestamp 1608763979
transform 1 0 18032 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_179
timestamp 1608763979
transform 1 0 17572 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_185
timestamp 1608763979
transform 1 0 18124 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763979
transform 1 0 16100 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608763979
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763979
transform 1 0 15456 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_158
timestamp 1608763979
transform 1 0 15640 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_147
timestamp 1608763979
transform 1 0 14628 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1608763979
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_159
timestamp 1608763979
transform 1 0 15732 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763979
transform 1 0 13156 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763979
transform 1 0 14168 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763979
transform 1 0 13432 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1608763979
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_137
timestamp 1608763979
transform 1 0 13708 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_141
timestamp 1608763979
transform 1 0 14076 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_129
timestamp 1608763979
transform 1 0 12972 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1608763979
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1608763979
transform 1 0 12144 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608763979
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_111
timestamp 1608763979
transform 1 0 11316 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_119
timestamp 1608763979
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_109
timestamp 1608763979
transform 1 0 11132 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_117
timestamp 1608763979
transform 1 0 11868 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1608763979
transform 1 0 9200 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763979
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763979
transform 1 0 9844 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608763979
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_86
timestamp 1608763979
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_91
timestamp 1608763979
transform 1 0 9476 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_89
timestamp 1608763979
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1608763979
transform 1 0 7176 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1608763979
transform 1 0 8188 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1608763979
transform 1 0 7452 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1608763979
transform 1 0 8464 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_75
timestamp 1608763979
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_67
timestamp 1608763979
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_78
timestamp 1608763979
transform 1 0 8280 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763979
transform 1 0 5796 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1608763979
transform 1 0 5704 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608763979
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763979
transform 1 0 5520 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_45
timestamp 1608763979
transform 1 0 5244 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_49
timestamp 1608763979
transform 1 0 5612 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1608763979
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1608763979
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_45
timestamp 1608763979
transform 1 0 5244 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1608763979
transform 1 0 4416 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1608763979
transform 1 0 4416 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608763979
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_33
timestamp 1608763979
transform 1 0 4140 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1608763979
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1608763979
transform 1 0 3036 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1608763979
transform 1 0 3772 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763979
transform 1 0 3588 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_27
timestamp 1608763979
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_25
timestamp 1608763979
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1608763979
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1608763979
transform 1 0 1564 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763979
transform 1 0 1380 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763979
transform 1 0 2116 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608763979
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608763979
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1608763979
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_9
timestamp 1608763979
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_19
timestamp 1608763979
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608763979
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763979
transform 1 0 16836 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_12_187
timestamp 1608763979
transform 1 0 18308 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1608763979
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608763979
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_146
timestamp 1608763979
transform 1 0 14536 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1608763979
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_163
timestamp 1608763979
transform 1 0 16100 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763979
transform 1 0 13064 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_128
timestamp 1608763979
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1608763979
transform 1 0 12052 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1608763979
transform 1 0 11040 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_117
timestamp 1608763979
transform 1 0 11868 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1608763979
transform 1 0 9016 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1608763979
transform 1 0 9844 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608763979
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_84
timestamp 1608763979
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_89
timestamp 1608763979
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1608763979
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_104
timestamp 1608763979
transform 1 0 10672 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763979
transform 1 0 7360 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_66
timestamp 1608763979
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763979
transform 1 0 5704 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_48
timestamp 1608763979
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763979
transform 1 0 4048 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608763979
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1608763979
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1608763979
transform 1 0 2944 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1608763979
transform 1 0 1840 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608763979
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1608763979
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1608763979
transform 1 0 1748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_17
timestamp 1608763979
transform 1 0 2668 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608763979
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_188
timestamp 1608763979
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1608763979
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608763979
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_178
timestamp 1608763979
transform 1 0 17480 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1608763979
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763979
transform 1 0 16008 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_11_153
timestamp 1608763979
transform 1 0 15180 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_161
timestamp 1608763979
transform 1 0 15916 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1608763979
transform 1 0 14352 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_139
timestamp 1608763979
transform 1 0 13892 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_143
timestamp 1608763979
transform 1 0 14260 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763979
transform 1 0 12420 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1608763979
transform 1 0 10948 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608763979
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763979
transform 1 0 11960 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_116
timestamp 1608763979
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1608763979
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763979
transform 1 0 9108 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_11_85
timestamp 1608763979
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763979
transform 1 0 7452 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_11_66
timestamp 1608763979
transform 1 0 7176 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1608763979
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1608763979
transform 1 0 5888 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608763979
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763979
transform 1 0 5612 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_44
timestamp 1608763979
transform 1 0 5152 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_48
timestamp 1608763979
transform 1 0 5520 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1608763979
transform 1 0 3312 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1608763979
transform 1 0 4324 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_23
timestamp 1608763979
transform 1 0 3220 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_33
timestamp 1608763979
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763979
transform 1 0 1380 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608763979
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_19
timestamp 1608763979
transform 1 0 2852 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608763979
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1608763979
transform 1 0 17848 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_178
timestamp 1608763979
transform 1 0 17480 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_186
timestamp 1608763979
transform 1 0 18216 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763979
transform 1 0 16008 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608763979
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1608763979
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_154
timestamp 1608763979
transform 1 0 15272 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1608763979
transform 1 0 14168 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1608763979
transform 1 0 13156 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_129
timestamp 1608763979
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_140
timestamp 1608763979
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1608763979
transform 1 0 12144 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_118
timestamp 1608763979
transform 1 0 11960 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1608763979
transform 1 0 9108 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763979
transform 1 0 10488 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1608763979
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608763979
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1608763979
transform 1 0 8924 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1608763979
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1608763979
transform 1 0 7084 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1608763979
transform 1 0 8096 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_74
timestamp 1608763979
transform 1 0 7912 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1608763979
transform 1 0 6256 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1608763979
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763979
transform 1 0 4784 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608763979
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1608763979
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_36
timestamp 1608763979
transform 1 0 4416 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1608763979
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1608763979
transform 1 0 2944 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1608763979
transform 1 0 1932 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608763979
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_7
timestamp 1608763979
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_18
timestamp 1608763979
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608763979
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1608763979
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1608763979
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1608763979
transform 1 0 17388 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608763979
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_172
timestamp 1608763979
transform 1 0 16928 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_176
timestamp 1608763979
transform 1 0 17296 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1608763979
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1608763979
transform 1 0 14720 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763979
transform 1 0 15456 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_151
timestamp 1608763979
transform 1 0 14996 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_155
timestamp 1608763979
transform 1 0 15364 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1608763979
transform 1 0 13616 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_134
timestamp 1608763979
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_145
timestamp 1608763979
transform 1 0 14444 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1608763979
transform 1 0 12604 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1608763979
transform 1 0 11316 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608763979
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_109
timestamp 1608763979
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1608763979
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1608763979
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1608763979
transform 1 0 10304 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_97
timestamp 1608763979
transform 1 0 10028 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763979
transform 1 0 8556 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1608763979
transform 1 0 7452 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_66
timestamp 1608763979
transform 1 0 7176 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_78
timestamp 1608763979
transform 1 0 8280 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1608763979
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763979
transform 1 0 4968 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608763979
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1608763979
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1608763979
transform 1 0 4232 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1608763979
transform 1 0 3220 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_21
timestamp 1608763979
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_32
timestamp 1608763979
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_38
timestamp 1608763979
transform 1 0 4600 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763979
transform 1 0 1564 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608763979
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1608763979
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608763979
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1608763979
transform 1 0 17848 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_174
timestamp 1608763979
transform 1 0 17112 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_186
timestamp 1608763979
transform 1 0 18216 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1608763979
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1608763979
transform 1 0 16284 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608763979
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763979
transform 1 0 14628 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_150
timestamp 1608763979
transform 1 0 14904 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1608763979
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1608763979
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_134
timestamp 1608763979
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_145
timestamp 1608763979
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1608763979
transform 1 0 12604 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1608763979
transform 1 0 11592 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_111
timestamp 1608763979
transform 1 0 11316 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_123
timestamp 1608763979
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1608763979
transform 1 0 9016 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763979
transform 1 0 9844 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608763979
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1608763979
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1608763979
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1608763979
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763979
transform 1 0 7360 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_66
timestamp 1608763979
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1608763979
transform 1 0 6348 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1608763979
transform 1 0 5336 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763979
transform 1 0 5060 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_55
timestamp 1608763979
transform 1 0 6164 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1608763979
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608763979
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1608763979
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_41
timestamp 1608763979
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1608763979
transform 1 0 1656 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763979
transform 1 0 2300 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608763979
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1608763979
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_10
timestamp 1608763979
transform 1 0 2024 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608763979
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608763979
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_188
timestamp 1608763979
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1608763979
transform 1 0 17848 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1608763979
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608763979
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_186
timestamp 1608763979
transform 1 0 18216 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1608763979
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1608763979
transform 1 0 17296 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1608763979
transform 1 0 17388 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_175
timestamp 1608763979
transform 1 0 17204 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_180
timestamp 1608763979
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_176
timestamp 1608763979
transform 1 0 17296 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_170
timestamp 1608763979
transform 1 0 16744 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1608763979
transform 1 0 14904 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1608763979
transform 1 0 15916 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1608763979
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608763979
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1608763979
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_163
timestamp 1608763979
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_148
timestamp 1608763979
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_159
timestamp 1608763979
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763979
transform 1 0 13248 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1608763979
transform 1 0 14168 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1608763979
transform 1 0 13156 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763979
transform 1 0 12972 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_129
timestamp 1608763979
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_140
timestamp 1608763979
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_127
timestamp 1608763979
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1608763979
transform 1 0 12512 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763979
transform 1 0 11500 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1608763979
transform 1 0 11316 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608763979
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_111
timestamp 1608763979
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_107
timestamp 1608763979
transform 1 0 10948 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1608763979
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_123
timestamp 1608763979
transform 1 0 12420 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1608763979
transform 1 0 10672 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763979
transform 1 0 9016 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763979
transform 1 0 9844 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608763979
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1608763979
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1608763979
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_84
timestamp 1608763979
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_102
timestamp 1608763979
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1608763979
transform 1 0 7084 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1608763979
transform 1 0 8464 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763979
transform 1 0 7912 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763979
transform 1 0 7636 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_63
timestamp 1608763979
transform 1 0 6900 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_69
timestamp 1608763979
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_78
timestamp 1608763979
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763979
transform 1 0 5428 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763979
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1608763979
transform 1 0 5520 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608763979
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763979
transform 1 0 5060 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_46
timestamp 1608763979
transform 1 0 5336 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_46
timestamp 1608763979
transform 1 0 5336 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1608763979
transform 1 0 6348 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1608763979
transform 1 0 3220 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763979
transform 1 0 3864 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1608763979
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608763979
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_21
timestamp 1608763979
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1608763979
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_41
timestamp 1608763979
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_28
timestamp 1608763979
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1608763979
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763979
transform 1 0 1564 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1608763979
transform 1 0 2852 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1608763979
transform 1 0 1840 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608763979
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608763979
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1608763979
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_6
timestamp 1608763979
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_17
timestamp 1608763979
transform 1 0 2668 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608763979
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1608763979
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1608763979
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608763979
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_178
timestamp 1608763979
transform 1 0 17480 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1608763979
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1608763979
transform 1 0 15548 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_155
timestamp 1608763979
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_166
timestamp 1608763979
transform 1 0 16376 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763979
transform 1 0 13892 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1608763979
transform 1 0 12880 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_127
timestamp 1608763979
transform 1 0 12788 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_137
timestamp 1608763979
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1608763979
transform 1 0 11684 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1608763979
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1608763979
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1608763979
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_123
timestamp 1608763979
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1608763979
transform 1 0 9660 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1608763979
transform 1 0 10672 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_91
timestamp 1608763979
transform 1 0 9476 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_102
timestamp 1608763979
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1608763979
transform 1 0 7636 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1608763979
transform 1 0 8648 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763979
transform 1 0 6900 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_69
timestamp 1608763979
transform 1 0 7452 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_80
timestamp 1608763979
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763979
transform 1 0 5796 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1608763979
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_49
timestamp 1608763979
transform 1 0 5612 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1608763979
transform 1 0 6348 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_62
timestamp 1608763979
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1608763979
transform 1 0 3772 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1608763979
transform 1 0 4784 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01
timestamp 1608763979
transform 1 0 3036 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_27
timestamp 1608763979
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_38
timestamp 1608763979
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763979
transform 1 0 1380 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608763979
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_19
timestamp 1608763979
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608763979
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1608763979
transform 1 0 17848 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1608763979
transform 1 0 17296 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_175
timestamp 1608763979
transform 1 0 17204 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_180
timestamp 1608763979
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_186
timestamp 1608763979
transform 1 0 18216 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1608763979
transform 1 0 14628 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1608763979
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1608763979
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_150
timestamp 1608763979
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_163
timestamp 1608763979
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1608763979
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_134
timestamp 1608763979
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_145
timestamp 1608763979
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763979
transform 1 0 11960 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1608763979
transform 1 0 10948 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_116
timestamp 1608763979
transform 1 0 11776 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1608763979
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1608763979
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763979
transform 1 0 10672 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1608763979
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_102
timestamp 1608763979
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1608763979
transform 1 0 7728 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763979
transform 1 0 8740 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_70
timestamp 1608763979
transform 1 0 7544 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_81
timestamp 1608763979
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1608763979
transform 1 0 5704 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1608763979
transform 1 0 6716 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_48
timestamp 1608763979
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_59
timestamp 1608763979
transform 1 0 6532 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763979
transform 1 0 4048 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1608763979
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1608763979
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1608763979
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1608763979
transform 1 0 2944 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1608763979
transform 1 0 1932 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608763979
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_7
timestamp 1608763979
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_18
timestamp 1608763979
transform 1 0 2760 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608763979
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_188
timestamp 1608763979
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1608763979
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1608763979
transform 1 0 17388 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1608763979
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1608763979
transform 1 0 16928 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_176
timestamp 1608763979
transform 1 0 17296 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1608763979
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1608763979
transform 1 0 14996 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_149
timestamp 1608763979
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_160
timestamp 1608763979
transform 1 0 15824 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763979
transform 1 0 13340 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_129
timestamp 1608763979
transform 1 0 12972 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763979
transform 1 0 12420 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1608763979
transform 1 0 11316 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1608763979
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_109
timestamp 1608763979
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1608763979
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763979
transform 1 0 9660 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_88
timestamp 1608763979
transform 1 0 9200 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_92
timestamp 1608763979
transform 1 0 9568 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763979
transform 1 0 7728 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_68
timestamp 1608763979
transform 1 0 7360 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1608763979
transform 1 0 5336 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763979
transform 1 0 6808 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1608763979
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_44
timestamp 1608763979
transform 1 0 5152 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_55
timestamp 1608763979
transform 1 0 6164 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763979
transform 1 0 3680 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_26
timestamp 1608763979
transform 1 0 3496 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1608763979
transform 1 0 1472 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763979
transform 1 0 2024 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608763979
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1608763979
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_8
timestamp 1608763979
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608763979
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1608763979
transform 1 0 17664 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1608763979
transform 1 0 17112 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_171
timestamp 1608763979
transform 1 0 16836 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_178
timestamp 1608763979
transform 1 0 17480 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_184
timestamp 1608763979
transform 1 0 18032 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1608763979
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1608763979
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_146
timestamp 1608763979
transform 1 0 14536 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1608763979
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_163
timestamp 1608763979
transform 1 0 16100 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1608763979
transform 1 0 13708 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_135
timestamp 1608763979
transform 1 0 13524 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763979
transform 1 0 12052 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_117
timestamp 1608763979
transform 1 0 11868 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763979
transform 1 0 10396 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763979
transform 1 0 9660 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1608763979
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1608763979
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_99
timestamp 1608763979
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763979
transform 1 0 7084 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763979
transform 1 0 8740 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_63
timestamp 1608763979
transform 1 0 6900 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_81
timestamp 1608763979
transform 1 0 8556 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763979
transform 1 0 5428 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1608763979
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1608763979
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_26
timestamp 1608763979
transform 1 0 3496 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_30
timestamp 1608763979
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_41
timestamp 1608763979
transform 1 0 4876 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1608763979
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1608763979
transform 1 0 2668 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763979
transform 1 0 1932 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608763979
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_7
timestamp 1608763979
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_15
timestamp 1608763979
transform 1 0 2484 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608763979
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608763979
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1608763979
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1608763979
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1608763979
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1608763979
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1608763979
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1608763979
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1608763979
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1608763979
transform 1 0 17664 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_176
timestamp 1608763979
transform 1 0 17296 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_176
timestamp 1608763979
transform 1 0 17296 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1608763979
transform 1 0 16928 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1608763979
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_170
timestamp 1608763979
transform 1 0 16744 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_170
timestamp 1608763979
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1608763979
transform 1 0 16376 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763979
transform 1 0 16192 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_162
timestamp 1608763979
transform 1 0 16008 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_162
timestamp 1608763979
transform 1 0 16008 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763979
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763979
transform 1 0 15456 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1608763979
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1608763979
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_154
timestamp 1608763979
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763979
transform 1 0 14628 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1608763979
transform 1 0 13432 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1608763979
transform 1 0 14444 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1608763979
transform 1 0 13616 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1608763979
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_145
timestamp 1608763979
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1608763979
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_143
timestamp 1608763979
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1608763979
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1608763979
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763979
transform 1 0 11776 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1608763979
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1608763979
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1608763979
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1608763979
transform 1 0 11868 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1608763979
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1608763979
transform 1 0 11040 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1608763979
transform 1 0 10764 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1608763979
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_106
timestamp 1608763979
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1608763979
transform 1 0 10028 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1608763979
transform 1 0 8832 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1608763979
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1608763979
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1608763979
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1608763979
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_93
timestamp 1608763979
transform 1 0 9660 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763979
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1608763979
transform 1 0 7820 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1608763979
transform 1 0 8648 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1608763979
transform 1 0 7636 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69
timestamp 1608763979
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80
timestamp 1608763979
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_71
timestamp 1608763979
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_82
timestamp 1608763979
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00
timestamp 1608763979
transform 1 0 5520 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1608763979
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1608763979
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1608763979
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1608763979
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_56
timestamp 1608763979
transform 1 0 6256 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp 1608763979
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1608763979
transform 1 0 5428 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46
timestamp 1608763979
transform 1 0 5336 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_45
timestamp 1608763979
transform 1 0 5244 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1608763979
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1608763979
transform 1 0 3128 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1608763979
transform 1 0 4416 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1608763979
transform 1 0 4508 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1608763979
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1608763979
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35
timestamp 1608763979
transform 1 0 4324 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_31
timestamp 1608763979
transform 1 0 3956 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_35
timestamp 1608763979
transform 1 0 4324 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1608763979
transform 1 0 2944 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_20
timestamp 1608763979
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1608763979
transform 1 0 2392 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1608763979
transform 1 0 2116 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11
timestamp 1608763979
transform 1 0 2116 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18
timestamp 1608763979
transform 1 0 2760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763979
transform 1 0 1564 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763979
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608763979
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608763979
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3
timestamp 1608763979
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_9
timestamp 1608763979
transform 1 0 1932 0 1 2720
box -38 -48 222 592
<< labels >>
rlabel metal2 s 1122 16200 1178 17000 4 IO_ISOL_N
port 1 nsew
rlabel metal2 s 17590 0 17646 800 4 SC_IN_BOT
port 2 nsew
rlabel metal2 s 3330 16200 3386 17000 4 SC_IN_TOP
port 3 nsew
rlabel metal2 s 18510 0 18566 800 4 SC_OUT_BOT
port 4 nsew
rlabel metal2 s 5538 16200 5594 17000 4 SC_OUT_TOP
port 5 nsew
rlabel metal2 s 1214 0 1270 800 4 bottom_grid_pin_0_
port 6 nsew
rlabel metal2 s 10322 0 10378 800 4 bottom_grid_pin_10_
port 7 nsew
rlabel metal2 s 11242 0 11298 800 4 bottom_grid_pin_11_
port 8 nsew
rlabel metal2 s 12162 0 12218 800 4 bottom_grid_pin_12_
port 9 nsew
rlabel metal2 s 13082 0 13138 800 4 bottom_grid_pin_13_
port 10 nsew
rlabel metal2 s 13910 0 13966 800 4 bottom_grid_pin_14_
port 11 nsew
rlabel metal2 s 14830 0 14886 800 4 bottom_grid_pin_15_
port 12 nsew
rlabel metal2 s 2134 0 2190 800 4 bottom_grid_pin_1_
port 13 nsew
rlabel metal2 s 3054 0 3110 800 4 bottom_grid_pin_2_
port 14 nsew
rlabel metal2 s 3974 0 4030 800 4 bottom_grid_pin_3_
port 15 nsew
rlabel metal2 s 4894 0 4950 800 4 bottom_grid_pin_4_
port 16 nsew
rlabel metal2 s 5814 0 5870 800 4 bottom_grid_pin_5_
port 17 nsew
rlabel metal2 s 6734 0 6790 800 4 bottom_grid_pin_6_
port 18 nsew
rlabel metal2 s 7562 0 7618 800 4 bottom_grid_pin_7_
port 19 nsew
rlabel metal2 s 8482 0 8538 800 4 bottom_grid_pin_8_
port 20 nsew
rlabel metal2 s 9402 0 9458 800 4 bottom_grid_pin_9_
port 21 nsew
rlabel metal2 s 15750 0 15806 800 4 bottom_width_0_height_0__pin_0_
port 22 nsew
rlabel metal2 s 16670 0 16726 800 4 bottom_width_0_height_0__pin_1_lower
port 23 nsew
rlabel metal2 s 386 0 442 800 4 bottom_width_0_height_0__pin_1_upper
port 24 nsew
rlabel metal2 s 7746 16200 7802 17000 4 ccff_head
port 25 nsew
rlabel metal2 s 9954 16200 10010 17000 4 ccff_tail
port 26 nsew
rlabel metal3 s 0 8848 800 8968 4 chanx_left_in[0]
port 27 nsew
rlabel metal3 s 0 12928 800 13048 4 chanx_left_in[10]
port 28 nsew
rlabel metal3 s 0 13336 800 13456 4 chanx_left_in[11]
port 29 nsew
rlabel metal3 s 0 13744 800 13864 4 chanx_left_in[12]
port 30 nsew
rlabel metal3 s 0 14152 800 14272 4 chanx_left_in[13]
port 31 nsew
rlabel metal3 s 0 14560 800 14680 4 chanx_left_in[14]
port 32 nsew
rlabel metal3 s 0 14968 800 15088 4 chanx_left_in[15]
port 33 nsew
rlabel metal3 s 0 15376 800 15496 4 chanx_left_in[16]
port 34 nsew
rlabel metal3 s 0 15784 800 15904 4 chanx_left_in[17]
port 35 nsew
rlabel metal3 s 0 16192 800 16312 4 chanx_left_in[18]
port 36 nsew
rlabel metal3 s 0 16600 800 16720 4 chanx_left_in[19]
port 37 nsew
rlabel metal3 s 0 9256 800 9376 4 chanx_left_in[1]
port 38 nsew
rlabel metal3 s 0 9664 800 9784 4 chanx_left_in[2]
port 39 nsew
rlabel metal3 s 0 10072 800 10192 4 chanx_left_in[3]
port 40 nsew
rlabel metal3 s 0 10480 800 10600 4 chanx_left_in[4]
port 41 nsew
rlabel metal3 s 0 10888 800 11008 4 chanx_left_in[5]
port 42 nsew
rlabel metal3 s 0 11296 800 11416 4 chanx_left_in[6]
port 43 nsew
rlabel metal3 s 0 11704 800 11824 4 chanx_left_in[7]
port 44 nsew
rlabel metal3 s 0 12112 800 12232 4 chanx_left_in[8]
port 45 nsew
rlabel metal3 s 0 12520 800 12640 4 chanx_left_in[9]
port 46 nsew
rlabel metal3 s 0 552 800 672 4 chanx_left_out[0]
port 47 nsew
rlabel metal3 s 0 4632 800 4752 4 chanx_left_out[10]
port 48 nsew
rlabel metal3 s 0 5040 800 5160 4 chanx_left_out[11]
port 49 nsew
rlabel metal3 s 0 5448 800 5568 4 chanx_left_out[12]
port 50 nsew
rlabel metal3 s 0 5856 800 5976 4 chanx_left_out[13]
port 51 nsew
rlabel metal3 s 0 6264 800 6384 4 chanx_left_out[14]
port 52 nsew
rlabel metal3 s 0 6672 800 6792 4 chanx_left_out[15]
port 53 nsew
rlabel metal3 s 0 7080 800 7200 4 chanx_left_out[16]
port 54 nsew
rlabel metal3 s 0 7488 800 7608 4 chanx_left_out[17]
port 55 nsew
rlabel metal3 s 0 7896 800 8016 4 chanx_left_out[18]
port 56 nsew
rlabel metal3 s 0 8304 800 8424 4 chanx_left_out[19]
port 57 nsew
rlabel metal3 s 0 960 800 1080 4 chanx_left_out[1]
port 58 nsew
rlabel metal3 s 0 1368 800 1488 4 chanx_left_out[2]
port 59 nsew
rlabel metal3 s 0 1776 800 1896 4 chanx_left_out[3]
port 60 nsew
rlabel metal3 s 0 2184 800 2304 4 chanx_left_out[4]
port 61 nsew
rlabel metal3 s 0 2592 800 2712 4 chanx_left_out[5]
port 62 nsew
rlabel metal3 s 0 3000 800 3120 4 chanx_left_out[6]
port 63 nsew
rlabel metal3 s 0 3408 800 3528 4 chanx_left_out[7]
port 64 nsew
rlabel metal3 s 0 3816 800 3936 4 chanx_left_out[8]
port 65 nsew
rlabel metal3 s 0 4224 800 4344 4 chanx_left_out[9]
port 66 nsew
rlabel metal3 s 19200 8576 20000 8696 4 chanx_right_in[0]
port 67 nsew
rlabel metal3 s 19200 12792 20000 12912 4 chanx_right_in[10]
port 68 nsew
rlabel metal3 s 19200 13200 20000 13320 4 chanx_right_in[11]
port 69 nsew
rlabel metal3 s 19200 13744 20000 13864 4 chanx_right_in[12]
port 70 nsew
rlabel metal3 s 19200 14152 20000 14272 4 chanx_right_in[13]
port 71 nsew
rlabel metal3 s 19200 14560 20000 14680 4 chanx_right_in[14]
port 72 nsew
rlabel metal3 s 19200 14968 20000 15088 4 chanx_right_in[15]
port 73 nsew
rlabel metal3 s 19200 15376 20000 15496 4 chanx_right_in[16]
port 74 nsew
rlabel metal3 s 19200 15784 20000 15904 4 chanx_right_in[17]
port 75 nsew
rlabel metal3 s 19200 16192 20000 16312 4 chanx_right_in[18]
port 76 nsew
rlabel metal3 s 19200 16600 20000 16720 4 chanx_right_in[19]
port 77 nsew
rlabel metal3 s 19200 8984 20000 9104 4 chanx_right_in[1]
port 78 nsew
rlabel metal3 s 19200 9392 20000 9512 4 chanx_right_in[2]
port 79 nsew
rlabel metal3 s 19200 9800 20000 9920 4 chanx_right_in[3]
port 80 nsew
rlabel metal3 s 19200 10344 20000 10464 4 chanx_right_in[4]
port 81 nsew
rlabel metal3 s 19200 10752 20000 10872 4 chanx_right_in[5]
port 82 nsew
rlabel metal3 s 19200 11160 20000 11280 4 chanx_right_in[6]
port 83 nsew
rlabel metal3 s 19200 11568 20000 11688 4 chanx_right_in[7]
port 84 nsew
rlabel metal3 s 19200 11976 20000 12096 4 chanx_right_in[8]
port 85 nsew
rlabel metal3 s 19200 12384 20000 12504 4 chanx_right_in[9]
port 86 nsew
rlabel metal3 s 19200 144 20000 264 4 chanx_right_out[0]
port 87 nsew
rlabel metal3 s 19200 4360 20000 4480 4 chanx_right_out[10]
port 88 nsew
rlabel metal3 s 19200 4768 20000 4888 4 chanx_right_out[11]
port 89 nsew
rlabel metal3 s 19200 5176 20000 5296 4 chanx_right_out[12]
port 90 nsew
rlabel metal3 s 19200 5584 20000 5704 4 chanx_right_out[13]
port 91 nsew
rlabel metal3 s 19200 5992 20000 6112 4 chanx_right_out[14]
port 92 nsew
rlabel metal3 s 19200 6400 20000 6520 4 chanx_right_out[15]
port 93 nsew
rlabel metal3 s 19200 6944 20000 7064 4 chanx_right_out[16]
port 94 nsew
rlabel metal3 s 19200 7352 20000 7472 4 chanx_right_out[17]
port 95 nsew
rlabel metal3 s 19200 7760 20000 7880 4 chanx_right_out[18]
port 96 nsew
rlabel metal3 s 19200 8168 20000 8288 4 chanx_right_out[19]
port 97 nsew
rlabel metal3 s 19200 552 20000 672 4 chanx_right_out[1]
port 98 nsew
rlabel metal3 s 19200 960 20000 1080 4 chanx_right_out[2]
port 99 nsew
rlabel metal3 s 19200 1368 20000 1488 4 chanx_right_out[3]
port 100 nsew
rlabel metal3 s 19200 1776 20000 1896 4 chanx_right_out[4]
port 101 nsew
rlabel metal3 s 19200 2184 20000 2304 4 chanx_right_out[5]
port 102 nsew
rlabel metal3 s 19200 2592 20000 2712 4 chanx_right_out[6]
port 103 nsew
rlabel metal3 s 19200 3000 20000 3120 4 chanx_right_out[7]
port 104 nsew
rlabel metal3 s 19200 3544 20000 3664 4 chanx_right_out[8]
port 105 nsew
rlabel metal3 s 19200 3952 20000 4072 4 chanx_right_out[9]
port 106 nsew
rlabel metal2 s 14370 16200 14426 17000 4 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 107 nsew
rlabel metal2 s 16578 16200 16634 17000 4 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 108 nsew
rlabel metal2 s 18786 16200 18842 17000 4 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 109 nsew
rlabel metal2 s 19430 0 19486 800 4 prog_clk_0_S_in
port 110 nsew
rlabel metal3 s 0 144 800 264 4 prog_clk_0_W_out
port 111 nsew
rlabel metal2 s 12162 16200 12218 17000 4 top_grid_pin_0_
port 112 nsew
rlabel metal4 s 3909 2128 4229 14736 4 VPWR
port 113 nsew
rlabel metal4 s 6875 2128 7195 14736 4 VGND
port 114 nsew
<< properties >>
string FIXED_BBOX 0 0 20000 17000
string GDS_FILE /ef/openfpga/openlane/runs/cbx_1__2_/results/magic/cbx_1__2_.gds
string GDS_END 1030846
string GDS_START 98316
<< end >>
